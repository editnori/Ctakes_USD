 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|43,52|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|43,52|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|43,57|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|77,86|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|77,86|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|77,91|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|133,136|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|144,151|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|144,151|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|153,161|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|SIMPLE_SEGMENT|164,173|false|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|164,173|false|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|164,173|false|false|false|C0020517|Hypersensitivity|Allergies
Attribute|Clinical Attribute|SIMPLE_SEGMENT|185,194|false|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|185,194|false|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|185,194|false|false|false|C0020517|Hypersensitivity|Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|197,219|true|false|false|C0041755|Adverse reaction to drug|Adverse Drug Reactions
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|205,209|false|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|Drug
Finding|Finding|SIMPLE_SEGMENT|205,209|false|false|false|C0740721|Drug problem|Drug
Finding|Pathologic Function|SIMPLE_SEGMENT|205,219|true|false|false|C0041755|Adverse reaction to drug|Drug Reactions
Event|Event|SIMPLE_SEGMENT|210,219|false|false|false|||Reactions
Event|Event|SIMPLE_SEGMENT|222,231|false|false|false|||Attending
Finding|Functional Concept|SIMPLE_SEGMENT|222,231|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|SIMPLE_SEGMENT|239,254|false|false|false|C0277786|Chief complaint (finding)|Chief Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|245,254|false|false|false|C3864418||Complaint
Event|Event|SIMPLE_SEGMENT|245,254|false|false|false|||Complaint
Finding|Finding|SIMPLE_SEGMENT|245,254|false|false|false|C5441521|Complaint (finding)|Complaint
Event|Event|SIMPLE_SEGMENT|257,264|false|false|false|||dyspnea
Finding|Finding|SIMPLE_SEGMENT|257,264|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|257,264|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|257,276|false|false|false|C0231807|Dyspnea on exertion|dyspnea on exertion
Event|Event|SIMPLE_SEGMENT|268,276|false|false|false|||exertion
Finding|Organism Function|SIMPLE_SEGMENT|268,276|false|false|false|C0015264|Exertion|exertion
Finding|Classification|SIMPLE_SEGMENT|280,285|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|SIMPLE_SEGMENT|286,294|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|286,294|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|298,316|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|307,316|false|false|false|C0945766||Procedure
Event|Event|SIMPLE_SEGMENT|307,316|false|false|false|||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|307,316|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|307,316|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|307,316|false|false|false|C0184661|Interventional procedure|Procedure
Event|Event|SIMPLE_SEGMENT|326,333|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|326,333|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|326,333|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|326,333|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|326,336|false|false|false|C0262926|Medical History|History of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|326,352|false|false|false|C0488508||History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|326,352|false|false|false|C0262512|History of present illness (finding)|History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|337,344|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Idea or Concept|SIMPLE_SEGMENT|337,344|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Finding|SIMPLE_SEGMENT|337,352|false|false|false|C4264312|Present illness|Present Illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|345,352|false|false|false|C0221423|Illness (finding)|Illness
Finding|Body Substance|SIMPLE_SEGMENT|354,361|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|354,361|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|354,361|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|371,375|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|SIMPLE_SEGMENT|371,375|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Event|Event|SIMPLE_SEGMENT|376,379|false|false|false|||old
Drug|Chemical Viewed Structurally|SIMPLE_SEGMENT|398,405|false|false|false|C0302912|Radicals (chemistry)|radical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|398,416|false|false|false|C0194401|Complete cystectomy|radical cystectomy
Event|Event|SIMPLE_SEGMENT|406,416|false|false|false|||cystectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|406,416|false|false|false|C0010651|Cystectomy|cystectomy
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|428,433|false|false|false|C0020885|ileum|ileal
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|428,441|false|false|false|C0441253|Structure of ileal conduit|ileal conduit
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|428,441|false|false|false|C0348002|Ileal conduit procedure|ileal conduit
Event|Activity|SIMPLE_SEGMENT|442,450|false|false|false|C1706214|Creation|creation
Event|Event|SIMPLE_SEGMENT|442,450|false|false|false|||creation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|442,450|false|false|false|C0441513|Surgical construction|creation
Event|Event|SIMPLE_SEGMENT|464,470|false|false|false|||course
Event|Event|SIMPLE_SEGMENT|472,483|false|false|false|||complicated
Event|Event|SIMPLE_SEGMENT|487,497|false|false|false|||bacteremia
Finding|Finding|SIMPLE_SEGMENT|487,497|false|false|false|C0004610|Bacteremia|bacteremia
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|502,509|false|false|false|C0000833|Abscess|abscess
Event|Event|SIMPLE_SEGMENT|502,509|false|false|false|||abscess
Finding|Intellectual Product|SIMPLE_SEGMENT|502,509|false|false|false|C1546533||abscess
Event|Event|SIMPLE_SEGMENT|511,514|false|false|false|||LLE
Anatomy|Body Location or Region|SIMPLE_SEGMENT|515,518|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|515,518|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|515,518|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Event|Event|SIMPLE_SEGMENT|515,518|false|false|false|||DVT
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|523,535|false|false|false|C0355642|Drugs used in migraine prophylaxis|prophylactic
Event|Event|SIMPLE_SEGMENT|523,535|false|false|false|||prophylactic
Finding|Functional Concept|SIMPLE_SEGMENT|523,535|false|false|false|C0445202|Prophylactic behavior|prophylactic
Drug|Organic Chemical|SIMPLE_SEGMENT|544,551|false|false|false|C0728963|Lovenox|lovenox
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|544,551|false|false|false|C0728963|Lovenox|lovenox
Event|Event|SIMPLE_SEGMENT|544,551|false|false|false|||lovenox
Event|Event|SIMPLE_SEGMENT|557,565|false|false|false|||presents
Event|Event|SIMPLE_SEGMENT|571,578|false|false|false|||dyspnea
Finding|Finding|SIMPLE_SEGMENT|571,578|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|571,578|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|571,590|false|false|false|C0231807|Dyspnea on exertion|dyspnea on exertion
Event|Event|SIMPLE_SEGMENT|582,590|false|false|false|||exertion
Finding|Organism Function|SIMPLE_SEGMENT|582,590|false|false|false|C0015264|Exertion|exertion
Finding|Body Substance|SIMPLE_SEGMENT|620,627|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|620,627|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|620,627|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|642,650|false|false|false|||admitted
Event|Occupational Activity|SIMPLE_SEGMENT|666,673|false|false|false|C0557854|Services|service
Finding|Idea or Concept|SIMPLE_SEGMENT|666,673|false|false|false|C3245478|ActInformationPrivacyReason - service|service
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|696,704|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Event|Event|SIMPLE_SEGMENT|705,717|false|false|false|||exenteration
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|705,717|false|false|false|C0015258||exenteration
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|723,728|false|false|false|C0020885|ileum|ileal
Event|Event|SIMPLE_SEGMENT|730,737|false|false|false|||conduit
Event|Event|SIMPLE_SEGMENT|747,757|false|false|false|||discharged
Event|Event|SIMPLE_SEGMENT|761,766|false|false|false|||rehab
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|761,766|false|false|false|C0034991|Rehabilitation therapy|rehab
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|770,782|false|false|false|C0355642|Drugs used in migraine prophylaxis|prophylactic
Event|Event|SIMPLE_SEGMENT|770,782|false|false|false|||prophylactic
Finding|Functional Concept|SIMPLE_SEGMENT|770,782|false|false|false|C0445202|Prophylactic behavior|prophylactic
Event|Event|SIMPLE_SEGMENT|783,789|false|false|false|||dosing
Drug|Organic Chemical|SIMPLE_SEGMENT|791,798|false|false|false|C0728963|Lovenox|lovenox
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|791,798|false|false|false|C0728963|Lovenox|lovenox
Event|Event|SIMPLE_SEGMENT|791,798|false|false|false|||lovenox
Finding|Idea or Concept|SIMPLE_SEGMENT|805,810|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Intellectual Product|SIMPLE_SEGMENT|805,810|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Intellectual Product|SIMPLE_SEGMENT|820,824|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|SIMPLE_SEGMENT|825,835|false|false|false|||readmitted
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|850,855|false|false|false|C1258215;C4019039|Ileus;Intestinal obstruction co-occurrent and due to decreased peristalsis|ileus
Event|Event|SIMPLE_SEGMENT|850,855|false|false|false|||ileus
Event|Event|SIMPLE_SEGMENT|870,883|false|false|false|||decompression
Finding|Functional Concept|SIMPLE_SEGMENT|870,883|false|false|false|C1965697|Decompression - action (qualifier value)|decompression
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|870,883|false|false|false|C0011117|external decompression|decompression
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|870,883|false|false|false|C0021153;C1829459|Decompression;Decompressive incision|decompression
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|885,888|false|false|false|C0027303;C1313790|NADP;TAPBP protein, human|TPN
Drug|Biologically Active Substance|SIMPLE_SEGMENT|885,888|false|false|false|C0027303;C1313790|NADP;TAPBP protein, human|TPN
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|885,888|false|false|false|C0027303;C1313790|NADP;TAPBP protein, human|TPN
Event|Event|SIMPLE_SEGMENT|885,888|false|false|false|||TPN
Finding|Gene or Genome|SIMPLE_SEGMENT|885,888|false|false|false|C1420583;C3813711|TAPBP gene;TAPBP wt Allele|TPN
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|885,888|false|false|false|C0030548|Parenteral Nutrition, Total|TPN
Event|Event|SIMPLE_SEGMENT|894,898|false|false|false|||grew
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|923,926|false|false|false|C0238052|Xanthomatosis, Cerebrotendinous|CTX
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|923,926|false|false|false|C0010377;C0010583;C5574748|C-Terminal Telopeptide Type 1 Collagen, human;Crotoxin;cyclophosphamide|CTX
Drug|Biologically Active Substance|SIMPLE_SEGMENT|923,926|false|false|false|C0010377;C0010583;C5574748|C-Terminal Telopeptide Type 1 Collagen, human;Crotoxin;cyclophosphamide|CTX
Drug|Enzyme|SIMPLE_SEGMENT|923,926|false|false|false|C0010377;C0010583;C5574748|C-Terminal Telopeptide Type 1 Collagen, human;Crotoxin;cyclophosphamide|CTX
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|923,926|false|false|false|C0010377;C0010583;C5574748|C-Terminal Telopeptide Type 1 Collagen, human;Crotoxin;cyclophosphamide|CTX
Drug|Organic Chemical|SIMPLE_SEGMENT|923,926|false|false|false|C0010377;C0010583;C5574748|C-Terminal Telopeptide Type 1 Collagen, human;Crotoxin;cyclophosphamide|CTX
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|923,926|false|false|false|C0010377;C0010583;C5574748|C-Terminal Telopeptide Type 1 Collagen, human;Crotoxin;cyclophosphamide|CTX
Event|Event|SIMPLE_SEGMENT|923,926|false|false|false|||CTX
Finding|Gene or Genome|SIMPLE_SEGMENT|923,926|false|false|false|C1413864;C3539598|CYP27A1 gene;CYP27A1 wt Allele|CTX
Event|Event|SIMPLE_SEGMENT|931,938|false|false|false|||started
Event|Event|SIMPLE_SEGMENT|940,942|false|false|false|||CT
Event|Event|SIMPLE_SEGMENT|943,949|false|false|false|||showed
Event|Event|SIMPLE_SEGMENT|950,965|false|false|false|||intra-abdominal
Finding|Functional Concept|SIMPLE_SEGMENT|950,965|false|false|false|C1512911|Intraabdominal Route of Administration|intra-abdominal
Event|Event|SIMPLE_SEGMENT|967,976|false|false|false|||interloop
Finding|Gene or Genome|SIMPLE_SEGMENT|979,985|false|false|false|C1424587|LITAF gene|simple
Drug|Substance|SIMPLE_SEGMENT|986,991|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|986,991|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|986,991|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|992,1002|false|false|false|||collection
Finding|Conceptual Entity|SIMPLE_SEGMENT|992,1002|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|SIMPLE_SEGMENT|992,1002|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|SIMPLE_SEGMENT|992,1002|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|SIMPLE_SEGMENT|992,1002|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1007,1010|false|false|false|C0230180|Structure of left lower quadrant of abdomen|LLQ
Drug|Substance|SIMPLE_SEGMENT|1011,1016|false|false|false|C1550628|Drain - SpecimenType|drain
Event|Event|SIMPLE_SEGMENT|1011,1016|false|false|false|||drain
Finding|Intellectual Product|SIMPLE_SEGMENT|1011,1016|false|false|false|C1546604|Drain Specimen Code|drain
Event|Event|SIMPLE_SEGMENT|1021,1027|false|false|false|||placed
Finding|Body Substance|SIMPLE_SEGMENT|1036,1043|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1036,1043|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1036,1043|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|1045,1053|false|false|false|||improved
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1063,1066|false|false|false|C0006430|Burning Mouth Syndrome|BMs
Event|Event|SIMPLE_SEGMENT|1063,1066|false|false|false|||BMs
Event|Event|SIMPLE_SEGMENT|1094,1104|false|false|false|||discharged
Drug|Organic Chemical|SIMPLE_SEGMENT|1109,1114|false|false|false|C0701042|Cipro|cipro
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1109,1114|false|false|false|C0701042|Cipro|cipro
Event|Event|SIMPLE_SEGMENT|1109,1114|false|false|false|||cipro
Drug|Organic Chemical|SIMPLE_SEGMENT|1115,1121|false|false|false|C0699678|Flagyl|flagyl
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1115,1121|false|false|false|C0699678|Flagyl|flagyl
Event|Event|SIMPLE_SEGMENT|1115,1121|false|false|false|||flagyl
Event|Event|SIMPLE_SEGMENT|1136,1146|false|false|false|||discharged
Drug|Organic Chemical|SIMPLE_SEGMENT|1153,1160|false|false|false|C0591139|Bactrim|Bactrim
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1153,1160|false|false|false|C0591139|Bactrim|Bactrim
Event|Event|SIMPLE_SEGMENT|1153,1160|false|false|false|||Bactrim
Event|Event|SIMPLE_SEGMENT|1165,1173|false|false|false|||presumed
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1175,1178|false|false|false|C0042029|Urinary tract infection|UTI
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1175,1178|false|false|false|C0077906|urinastatin|UTI
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1175,1178|false|false|false|C0077906|urinastatin|UTI
Event|Event|SIMPLE_SEGMENT|1175,1178|false|false|false|||UTI
Finding|Gene or Genome|SIMPLE_SEGMENT|1175,1178|false|false|false|C1412376;C5780748|AMBP gene;AMBP wt Allele|UTI
Event|Event|SIMPLE_SEGMENT|1211,1215|false|false|false|||took
Event|Event|SIMPLE_SEGMENT|1235,1244|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|1235,1244|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|SIMPLE_SEGMENT|1254,1259|false|false|false|||noted
Finding|Finding|SIMPLE_SEGMENT|1268,1271|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|1268,1271|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1286,1291|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|1286,1291|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|1286,1291|false|false|false|C0013604|Edema|edema
Finding|Finding|SIMPLE_SEGMENT|1307,1311|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|1307,1311|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|1307,1311|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|SIMPLE_SEGMENT|1312,1318|false|false|false|||showed
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1324,1328|false|false|false|C4318566|Deep Resection Margin|deep
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1324,1333|false|false|false|C0226514|Structure of deep vein|deep vein
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1324,1344|false|false|false|C0149871;C0340708|Deep Vein Thrombosis;Deep vein thrombosis of lower limb|deep vein thrombosis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1329,1333|false|false|false|C0042449|Veins|vein
Finding|Pathologic Function|SIMPLE_SEGMENT|1329,1344|false|false|false|C0042487|Venous Thrombosis|vein thrombosis
Event|Event|SIMPLE_SEGMENT|1334,1344|false|false|false|||thrombosis
Finding|Pathologic Function|SIMPLE_SEGMENT|1334,1344|false|false|false|C0040053|Thrombosis|thrombosis
Event|Event|SIMPLE_SEGMENT|1352,1362|false|false|false|||duplicated
Finding|Finding|SIMPLE_SEGMENT|1352,1362|false|false|false|C0332597|Duplication (finding)|duplicated
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1372,1378|false|false|false|C4522154|Distal Resection Margin|distal
Finding|Functional Concept|SIMPLE_SEGMENT|1379,1383|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1384,1391|false|false|false|C0015811|Femur|femoral
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1384,1397|false|false|false|C0015809|Femoral vein|femoral veins
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1392,1397|false|false|false|C0042449|Veins|veins
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1392,1397|false|false|false|C0398102|Procedure on vein|veins
Event|Event|SIMPLE_SEGMENT|1407,1417|false|false|false|||discharged
Drug|Organic Chemical|SIMPLE_SEGMENT|1423,1433|false|false|false|C0206460|enoxaparin|Enoxaparin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1423,1433|false|false|false|C0206460|enoxaparin|Enoxaparin
Event|Event|SIMPLE_SEGMENT|1423,1433|false|false|false|||Enoxaparin
Drug|Organic Chemical|SIMPLE_SEGMENT|1423,1440|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1423,1440|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1434,1440|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|1434,1440|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1434,1440|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|SIMPLE_SEGMENT|1434,1440|false|false|false|||Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|1434,1440|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1434,1440|false|false|false|C0337443|Sodium measurement|Sodium
Event|Event|SIMPLE_SEGMENT|1461,1468|false|false|false|||reports
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1478,1481|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|1478,1481|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1478,1481|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1478,1481|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|SIMPLE_SEGMENT|1478,1481|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|1478,1481|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|SIMPLE_SEGMENT|1478,1481|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1478,1481|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|SIMPLE_SEGMENT|1478,1481|false|false|false|||PCP
Finding|Gene or Genome|SIMPLE_SEGMENT|1478,1481|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|SIMPLE_SEGMENT|1478,1481|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Event|SIMPLE_SEGMENT|1483,1490|false|false|false|||started
Finding|Intellectual Product|SIMPLE_SEGMENT|1519,1523|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|SIMPLE_SEGMENT|1540,1551|false|false|false|||improvement
Finding|Conceptual Entity|SIMPLE_SEGMENT|1540,1551|false|false|false|C2986411|Improvement|improvement
Event|Event|SIMPLE_SEGMENT|1559,1567|false|false|false|||swelling
Finding|Finding|SIMPLE_SEGMENT|1559,1567|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|SIMPLE_SEGMENT|1559,1567|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1577,1583|false|false|false|C4255046||report
Event|Event|SIMPLE_SEGMENT|1577,1583|false|false|false|||report
Finding|Intellectual Product|SIMPLE_SEGMENT|1577,1583|false|false|false|C0684224|Report (document)|report
Procedure|Health Care Activity|SIMPLE_SEGMENT|1577,1583|false|false|false|C0700287|Reporting|report
Finding|Functional Concept|SIMPLE_SEGMENT|1587,1593|false|false|false|C0205341;C1705914|Repeat;Repeat Object|repeat
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1606,1611|false|false|false|C0034991|Rehabilitation therapy|rehab
Event|Event|SIMPLE_SEGMENT|1612,1620|false|false|false|||facility
Finding|Intellectual Product|SIMPLE_SEGMENT|1612,1620|false|false|false|C4695111|ADMIN.FACILITY|facility
Event|Event|SIMPLE_SEGMENT|1631,1639|false|false|false|||negative
Finding|Classification|SIMPLE_SEGMENT|1631,1639|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|1631,1639|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1631,1639|false|false|false|C5237010|Expression Negative|negative
Finding|Finding|SIMPLE_SEGMENT|1631,1643|false|false|false|C0205160|Negative|negative for
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1644,1647|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1644,1647|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1644,1647|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Event|Event|SIMPLE_SEGMENT|1644,1647|false|false|false|||DVT
Finding|Body Substance|SIMPLE_SEGMENT|1650,1657|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1650,1657|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1650,1657|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|1658,1665|false|false|false|||reports
Event|Event|SIMPLE_SEGMENT|1675,1684|false|false|false|||recovered
Finding|Finding|SIMPLE_SEGMENT|1685,1689|false|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|1722,1726|false|false|false|||well
Finding|Finding|SIMPLE_SEGMENT|1722,1726|false|false|false|C5575035|Well (answer to question)|well
Procedure|Health Care Activity|SIMPLE_SEGMENT|1734,1749|false|false|false|C1456630|Assisted Living|assisted living
Event|Event|SIMPLE_SEGMENT|1743,1749|false|false|false|||living
Finding|Conceptual Entity|SIMPLE_SEGMENT|1743,1749|false|false|false|C0595998;C4520849;C4551704|Alive;Household composition;Living|living
Finding|Finding|SIMPLE_SEGMENT|1743,1749|false|false|false|C0595998;C4520849;C4551704|Alive;Household composition;Living|living
Finding|Intellectual Product|SIMPLE_SEGMENT|1750,1758|false|false|false|C4695111|ADMIN.FACILITY|facility
Finding|Intellectual Product|SIMPLE_SEGMENT|1770,1774|false|false|false|C1561540|Transaction counts and value totals - week|week
Finding|Gene or Genome|SIMPLE_SEGMENT|1775,1778|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Event|Event|SIMPLE_SEGMENT|1789,1794|false|false|false|||began
Event|Event|SIMPLE_SEGMENT|1808,1815|false|false|false|||dyspnea
Finding|Finding|SIMPLE_SEGMENT|1808,1815|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|1808,1815|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|1808,1827|false|false|false|C0231807|Dyspnea on exertion|dyspnea on exertion
Event|Event|SIMPLE_SEGMENT|1819,1827|false|false|false|||exertion
Finding|Organism Function|SIMPLE_SEGMENT|1819,1827|false|false|false|C0015264|Exertion|exertion
Event|Event|SIMPLE_SEGMENT|1833,1839|false|false|false|||states
Event|Event|SIMPLE_SEGMENT|1863,1867|false|false|false|||able
Finding|Finding|SIMPLE_SEGMENT|1863,1867|false|false|false|C1299581|Able (qualifier value)|able
Event|Event|SIMPLE_SEGMENT|1871,1879|false|false|false|||ambulate
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|1882,1887|false|false|false|C1706085|Block Dosage Form|block
Event|Event|SIMPLE_SEGMENT|1882,1887|false|false|false|||block
Finding|Body Substance|SIMPLE_SEGMENT|1882,1887|false|false|false|C0028778;C0332206;C1533157|Blocking;Fixed Block;Obstruction|block
Finding|Finding|SIMPLE_SEGMENT|1882,1887|false|false|false|C0028778;C0332206;C1533157|Blocking;Fixed Block;Obstruction|block
Finding|Functional Concept|SIMPLE_SEGMENT|1882,1887|false|false|false|C0028778;C0332206;C1533157|Blocking;Fixed Block;Obstruction|block
Event|Event|SIMPLE_SEGMENT|1895,1903|false|false|false|||stopping
Event|Event|SIMPLE_SEGMENT|1908,1913|false|false|false|||catch
Finding|Sign or Symptom|SIMPLE_SEGMENT|1908,1913|false|false|false|C0231617|Catch - Finding of sensory dimension of pain|catch
Event|Event|SIMPLE_SEGMENT|1918,1924|false|false|false|||breath
Finding|Body Substance|SIMPLE_SEGMENT|1918,1924|false|false|false|C0225386|Breath|breath
Finding|Intellectual Product|SIMPLE_SEGMENT|1946,1950|false|false|false|C1561540|Transaction counts and value totals - week|week
Event|Event|SIMPLE_SEGMENT|1964,1970|false|false|false|||unable
Finding|Finding|SIMPLE_SEGMENT|1964,1970|false|false|false|C1299582|Unable|unable
Event|Event|SIMPLE_SEGMENT|1996,2001|false|false|false|||steps
Finding|Conceptual Entity|SIMPLE_SEGMENT|1996,2001|false|false|false|C1261552|Step (specific stage)|steps
Procedure|Health Care Activity|SIMPLE_SEGMENT|1996,2001|false|false|false|C4722257|STEPS to Enhance Physical Activity|steps
Event|Event|SIMPLE_SEGMENT|2007,2013|false|false|false|||states
Event|Event|SIMPLE_SEGMENT|2026,2032|false|false|false|||become
Event|Event|SIMPLE_SEGMENT|2052,2061|false|false|false|||difficult
Finding|Finding|SIMPLE_SEGMENT|2052,2061|false|false|false|C0332218|Difficult (qualifier value)|difficult
Event|Event|SIMPLE_SEGMENT|2065,2073|false|false|false|||ambulate
Event|Event|SIMPLE_SEGMENT|2083,2090|false|false|false|||bedroom
Event|Event|SIMPLE_SEGMENT|2099,2107|false|false|false|||bathroom
Event|Event|SIMPLE_SEGMENT|2114,2121|false|false|false|||visited
Finding|Functional Concept|SIMPLE_SEGMENT|2136,2146|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|ambulatory
Finding|Idea or Concept|SIMPLE_SEGMENT|2136,2146|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|ambulatory
Finding|Intellectual Product|SIMPLE_SEGMENT|2136,2146|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|ambulatory
Procedure|Health Care Activity|SIMPLE_SEGMENT|2136,2146|false|false|false|C1561560|ambulatory encounter|ambulatory
Event|Event|SIMPLE_SEGMENT|2147,2157|false|false|false|||saturation
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|2147,2157|false|false|false|C0522534|Saturated|saturation
Event|Event|SIMPLE_SEGMENT|2163,2168|false|false|false|||noted
Event|Event|SIMPLE_SEGMENT|2202,2213|false|false|false|||tachycardia
Finding|Finding|SIMPLE_SEGMENT|2202,2213|false|false|false|C0039231;C3827868|Tachycardia;Tachycardia by ECG Finding|tachycardia
Event|Event|SIMPLE_SEGMENT|2223,2229|false|false|false|||pallor
Finding|Finding|SIMPLE_SEGMENT|2223,2229|false|false|false|C0241137|Pallor of skin|pallor
Event|Event|SIMPLE_SEGMENT|2234,2245|false|false|false|||diaphoresis
Finding|Finding|SIMPLE_SEGMENT|2234,2245|false|false|false|C0700590|Increased sweating|diaphoresis
Event|Event|SIMPLE_SEGMENT|2251,2259|false|false|false|||endorses
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2271,2274|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Finding|Pathologic Function|SIMPLE_SEGMENT|2271,2283|false|true|false|C0581394|Swelling of lower limb|leg swelling
Event|Event|SIMPLE_SEGMENT|2275,2283|false|false|false|||swelling
Finding|Finding|SIMPLE_SEGMENT|2275,2283|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|SIMPLE_SEGMENT|2275,2283|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Functional Concept|SIMPLE_SEGMENT|2285,2289|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Event|Event|SIMPLE_SEGMENT|2290,2295|false|false|false|||worse
Finding|Finding|SIMPLE_SEGMENT|2290,2295|false|false|false|C1457868;C1550463|Observation Interpretation - worse;Worse|worse
Finding|Idea or Concept|SIMPLE_SEGMENT|2290,2295|false|false|false|C1457868;C1550463|Observation Interpretation - worse;Worse|worse
Event|Event|SIMPLE_SEGMENT|2301,2306|false|false|false|||right
Finding|Functional Concept|SIMPLE_SEGMENT|2301,2306|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Event|Event|SIMPLE_SEGMENT|2316,2322|false|false|false|||states
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2332,2338|false|false|false|C0039866|Thigh structure|thighs
Event|Event|SIMPLE_SEGMENT|2340,2344|false|false|false|||feel
Finding|Mental Process|SIMPLE_SEGMENT|2340,2344|false|false|false|C1527305|Feelings|feel
Event|Event|SIMPLE_SEGMENT|2358,2364|false|false|false|||denies
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2380,2385|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|2380,2385|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2380,2390|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|2380,2390|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2386,2390|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|2386,2390|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|2386,2390|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|2386,2390|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|2392,2397|false|false|false|||fever
Finding|Finding|SIMPLE_SEGMENT|2392,2397|true|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|2392,2397|true|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Event|Event|SIMPLE_SEGMENT|2399,2405|false|false|false|||chills
Finding|Sign or Symptom|SIMPLE_SEGMENT|2399,2405|true|false|false|C0085593|Chills|chills
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2408,2412|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|2408,2412|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|2408,2412|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|2408,2412|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2418,2422|false|false|false|C4318566|Deep Resection Margin|deep
Event|Event|SIMPLE_SEGMENT|2423,2434|false|false|false|||inspiration
Finding|Organism Function|SIMPLE_SEGMENT|2423,2434|false|false|false|C0004048|Inspiration (function)|inspiration
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2436,2445|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|SIMPLE_SEGMENT|2436,2450|false|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2446,2450|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|2446,2450|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|2446,2450|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|2446,2450|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|2452,2458|false|false|false|||rashes
Finding|Sign or Symptom|SIMPLE_SEGMENT|2452,2458|false|false|false|C0015230;C5779628|Exanthema;Skin rash|rashes
Event|Event|SIMPLE_SEGMENT|2460,2469|false|false|false|||dizziness
Finding|Sign or Symptom|SIMPLE_SEGMENT|2460,2469|false|false|false|C0012833;C0042571|Dizziness;Vertigo|dizziness
Event|Event|SIMPLE_SEGMENT|2472,2487|false|false|false|||lightheadedness
Finding|Sign or Symptom|SIMPLE_SEGMENT|2472,2487|false|false|false|C0220870|Lightheadedness|lightheadedness
Finding|Idea or Concept|SIMPLE_SEGMENT|2503,2510|false|false|false|C1555582|Initial (abbreviation)|initial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2543,2548|false|false|false|C0028429||Nasal
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|2543,2548|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Organic Chemical|SIMPLE_SEGMENT|2543,2548|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2543,2548|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Finding|Finding|SIMPLE_SEGMENT|2543,2548|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Finding|Functional Concept|SIMPLE_SEGMENT|2543,2548|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2549,2556|false|false|false|C1550232|Body Parts - Cannula|Cannula
Finding|Body Substance|SIMPLE_SEGMENT|2549,2556|false|false|false|C1546577;C1550622|Specimen Type - Cannula|Cannula
Finding|Intellectual Product|SIMPLE_SEGMENT|2549,2556|false|false|false|C1546577;C1550622|Specimen Type - Cannula|Cannula
Event|Event|SIMPLE_SEGMENT|2562,2570|false|false|false|||physical
Finding|Finding|SIMPLE_SEGMENT|2562,2570|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Finding|Functional Concept|SIMPLE_SEGMENT|2562,2570|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|2562,2570|false|false|false|C0031809|Physical Examination|physical
Finding|Finding|SIMPLE_SEGMENT|2562,2575|false|false|false|C1509143|physical examination (physical finding)|physical exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2562,2575|false|false|false|C0031809|Physical Examination|physical exam
Event|Event|SIMPLE_SEGMENT|2571,2575|false|false|false|||exam
Finding|Functional Concept|SIMPLE_SEGMENT|2571,2575|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2571,2575|false|false|false|C0582103|Medical Examination|exam
Event|Event|SIMPLE_SEGMENT|2580,2588|false|false|false|||recorded
Finding|Body Substance|SIMPLE_SEGMENT|2592,2599|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|2592,2599|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|2592,2599|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2637,2640|false|false|false|C0023759|Lip structure|lip
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2637,2640|false|false|false|C0153932;C0264511|Benign neoplasm of the lip;Lymphoid interstitial pneumonia|lip
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2637,2640|false|false|false|C0153932;C0264511|Benign neoplasm of the lip;Lymphoid interstitial pneumonia|lip
Finding|Gene or Genome|SIMPLE_SEGMENT|2637,2640|false|false|false|C1846919;C3889123|SMG1 gene;SMG1 wt Allele|lip
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2641,2650|false|false|false|C5885990||breathing
Event|Event|SIMPLE_SEGMENT|2641,2650|false|false|false|||breathing
Finding|Finding|SIMPLE_SEGMENT|2641,2650|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|SIMPLE_SEGMENT|2641,2650|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|SIMPLE_SEGMENT|2641,2650|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|SIMPLE_SEGMENT|2641,2650|false|false|false|C1160636|respiratory system process|breathing
Event|Event|SIMPLE_SEGMENT|2652,2658|false|false|false|||unable
Finding|Finding|SIMPLE_SEGMENT|2652,2658|false|false|false|C1299582|Unable|unable
Finding|Finding|SIMPLE_SEGMENT|2652,2667|false|false|false|C0564216;C4722246|Unable to Speak at All;Unable to speak (finding)|unable to speak
Event|Event|SIMPLE_SEGMENT|2662,2667|false|false|false|||speak
Finding|Finding|SIMPLE_SEGMENT|2662,2667|false|false|false|C0234856;C0600116;C1547187|Does speak;Speak - language ability;Speaking (function)|speak
Finding|Idea or Concept|SIMPLE_SEGMENT|2662,2667|false|false|false|C0234856;C0600116;C1547187|Does speak;Speak - language ability;Speaking (function)|speak
Finding|Individual Behavior|SIMPLE_SEGMENT|2662,2667|false|false|false|C0234856;C0600116;C1547187|Does speak;Speak - language ability;Speaking (function)|speak
Event|Event|SIMPLE_SEGMENT|2676,2685|false|false|false|||sentences
Finding|Intellectual Product|SIMPLE_SEGMENT|2676,2685|false|false|false|C0876929|Sentence|sentences
Event|Event|SIMPLE_SEGMENT|2694,2702|false|false|false|||becoming
Finding|Sign or Symptom|SIMPLE_SEGMENT|2703,2718|false|false|false|C0013404|Dyspnea|short of breath
Finding|Body Substance|SIMPLE_SEGMENT|2712,2718|false|false|false|C0225386|Breath|breath
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|2720,2728|false|false|false|C0559495|Urological stoma|urostomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2720,2728|false|false|false|C0856443|Urostomy procedure|urostomy
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2729,2734|false|false|false|C0222017|Abdominal skin pouch|pouch
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2738,2741|false|false|false|C0230178|Structure of right lower quadrant of abdomen|RLQ
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|2743,2748|false|false|false|C1955856|Surgical Stoma|stoma
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2759,2764|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|2759,2764|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|2759,2764|false|false|false|C0013604|Edema|edema
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2778,2783|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|2778,2783|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2778,2795|false|false|false|C0023216|Lower Extremity|lower extremities
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2784,2795|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Event|Event|SIMPLE_SEGMENT|2806,2810|false|false|false|||labs
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2806,2810|false|false|false|C0587081|Laboratory test finding|labs
Event|Event|SIMPLE_SEGMENT|2816,2823|false|false|false|||notable
Event|Event|SIMPLE_SEGMENT|2835,2838|false|false|false|||Hct
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2835,2838|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2835,2838|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Event|Event|SIMPLE_SEGMENT|2843,2846|false|false|false|||plt
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2843,2846|false|false|false|C0201617|Primed lymphocyte test|plt
Finding|Gene or Genome|SIMPLE_SEGMENT|2856,2861|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Anatomy|Cell|SIMPLE_SEGMENT|2873,2876|false|false|false|C0023516|Leukocytes|WBC
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2890,2893|false|false|false|C0267963|Exocrine pancreatic insufficiency|epi
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2890,2893|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|epi
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2890,2893|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|epi
Drug|Hormone|SIMPLE_SEGMENT|2890,2893|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|epi
Drug|Organic Chemical|SIMPLE_SEGMENT|2890,2893|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|epi
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2890,2893|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|epi
Event|Event|SIMPLE_SEGMENT|2890,2893|false|false|false|||epi
Finding|Gene or Genome|SIMPLE_SEGMENT|2890,2893|false|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|epi
Finding|Intellectual Product|SIMPLE_SEGMENT|2890,2893|false|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|epi
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2890,2893|false|false|false|C0162734;C3641909|Echo-Planar Imaging;Electronic Portal Imaging|epi
Finding|Finding|SIMPLE_SEGMENT|2900,2903|false|false|false|C5848551|Neg - answer|neg
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2908,2914|false|false|false|C5574646|Natriuretic Peptides B, human|proBNP
Drug|Hormone|SIMPLE_SEGMENT|2908,2914|false|false|false|C5574646|Natriuretic Peptides B, human|proBNP
Event|Event|SIMPLE_SEGMENT|2915,2921|false|false|false|||normal
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2923,2926|false|false|false|C3813556|Cancer/Testis Antigen|CTA
Event|Event|SIMPLE_SEGMENT|2923,2926|false|false|false|||CTA
Finding|Gene or Genome|SIMPLE_SEGMENT|2923,2926|false|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2923,2926|false|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2927,2932|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|2927,2932|false|false|false|C0741025|Chest problem|chest
Event|Event|SIMPLE_SEGMENT|2933,2939|false|false|false|||showed
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2954,2963|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2954,2963|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|2954,2963|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|SIMPLE_SEGMENT|2954,2972|false|false|false|C0034065|Pulmonary Embolism|pulmonary embolism
Event|Event|SIMPLE_SEGMENT|2964,2972|false|false|false|||embolism
Finding|Finding|SIMPLE_SEGMENT|2964,2972|false|false|false|C0013922;C1704212|Embolism;Embolus|embolism
Finding|Pathologic Function|SIMPLE_SEGMENT|2964,2972|false|false|false|C0013922;C1704212|Embolism;Embolus|embolism
Event|Event|SIMPLE_SEGMENT|2978,2986|false|false|false|||thrombus
Finding|Pathologic Function|SIMPLE_SEGMENT|2978,2986|false|false|false|C0087086;C0302148|Blood Clot;Thrombus|thrombus
Event|Event|SIMPLE_SEGMENT|2987,2991|false|false|false|||seen
Event|Event|SIMPLE_SEGMENT|2992,3001|false|false|false|||extending
Finding|Functional Concept|SIMPLE_SEGMENT|3012,3017|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3012,3039|false|false|false|C0226054;C0923924|Right pulmonary arterial tree;Right pulmonary artery|right main pulmonary artery
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3023,3032|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3023,3032|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|3023,3032|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3023,3039|false|false|false|C0034052|Pulmonary artery structure|pulmonary artery
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3033,3039|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|SIMPLE_SEGMENT|3033,3039|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Finding|Functional Concept|SIMPLE_SEGMENT|3077,3082|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Event|Event|SIMPLE_SEGMENT|3090,3096|false|false|false|||middle
Finding|Intellectual Product|SIMPLE_SEGMENT|3090,3096|false|false|false|C1552826|Table Cell Vertical Align - middle|middle
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3102,3107|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|3102,3107|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3102,3112|false|false|false|C0225758|Structure of lower lobe of lung|lower lobe
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3108,3112|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|SIMPLE_SEGMENT|3108,3112|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3108,3122|false|false|false|C0225752|Structure of lobe of lung|lobe pulmonary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3113,3122|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3113,3122|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|3113,3122|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3124,3132|false|false|false|C0003842;C0226004|Arterial system;Arteries|arteries
Anatomy|Body System|SIMPLE_SEGMENT|3124,3132|false|false|false|C0003842;C0226004|Arterial system;Arteries|arteries
Event|Event|SIMPLE_SEGMENT|3124,3132|false|false|false|||arteries
Procedure|Health Care Activity|SIMPLE_SEGMENT|3124,3132|false|false|false|C0397581|Procedure on artery|arteries
Finding|Functional Concept|SIMPLE_SEGMENT|3137,3142|true|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3137,3148|false|false|false|C0225808|Right side of heart|right heart
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3143,3148|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3143,3148|true|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|3143,3148|true|false|false|C0795691|HEART PROBLEM|heart
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|3149,3155|true|false|false|C0080194|Muscle strain|strain
Event|Event|SIMPLE_SEGMENT|3149,3155|false|false|false|||strain
Finding|Idea or Concept|SIMPLE_SEGMENT|3149,3155|true|false|false|C0442694;C1510453;C1548152;C2987481|Emotional Strain;Nature of Abnormal Testing - Strain;Straining (finding);strain symptom|strain
Finding|Mental Process|SIMPLE_SEGMENT|3149,3155|true|false|false|C0442694;C1510453;C1548152;C2987481|Emotional Strain;Nature of Abnormal Testing - Strain;Straining (finding);strain symptom|strain
Finding|Physiologic Function|SIMPLE_SEGMENT|3149,3155|true|false|false|C0442694;C1510453;C1548152;C2987481|Emotional Strain;Nature of Abnormal Testing - Strain;Straining (finding);strain symptom|strain
Finding|Sign or Symptom|SIMPLE_SEGMENT|3149,3155|true|false|false|C0442694;C1510453;C1548152;C2987481|Emotional Strain;Nature of Abnormal Testing - Strain;Straining (finding);strain symptom|strain
Event|Event|SIMPLE_SEGMENT|3156,3166|false|false|false|||identified
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3204,3213|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3204,3213|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|3204,3213|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|SIMPLE_SEGMENT|3204,3220|false|false|false|C0034065|Pulmonary Embolism|pulmonary emboli
Event|Event|SIMPLE_SEGMENT|3214,3220|false|false|false|||emboli
Finding|Finding|SIMPLE_SEGMENT|3214,3220|false|false|false|C1704212|Embolus|emboli
Event|Event|SIMPLE_SEGMENT|3221,3225|false|false|false|||seen
Event|Event|SIMPLE_SEGMENT|3261,3269|false|false|false|||branches
Finding|Functional Concept|SIMPLE_SEGMENT|3277,3281|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3292,3297|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|3292,3297|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3298,3303|false|false|false|C0796494|lobe|lobes
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3317,3326|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3317,3326|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|3317,3326|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Finding|SIMPLE_SEGMENT|3317,3334|false|false|false|C0748164|Multiple Pulmonary Nodules|pulmonary nodules
Event|Event|SIMPLE_SEGMENT|3327,3334|false|false|false|||nodules
Event|Event|SIMPLE_SEGMENT|3339,3344|false|false|false|||noted
Event|Event|SIMPLE_SEGMENT|3349,3354|false|false|false|||noted
Event|Event|SIMPLE_SEGMENT|3395,3405|false|false|false|||spiculated
Event|Event|SIMPLE_SEGMENT|3410,3419|false|false|false|||measuring
Finding|Functional Concept|SIMPLE_SEGMENT|3439,3444|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3439,3456|false|false|false|C4281590|Structure of middle lobe of right lung|right middle lobe
Finding|Intellectual Product|SIMPLE_SEGMENT|3445,3451|false|false|false|C1552826|Table Cell Vertical Align - middle|middle
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3445,3456|false|false|false|C4281590|Structure of middle lobe of right lung|middle lobe
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3452,3456|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|SIMPLE_SEGMENT|3452,3456|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Event|Event|SIMPLE_SEGMENT|3458,3468|false|false|false|||suspicious
Finding|Finding|SIMPLE_SEGMENT|3458,3483|false|false|false|C4050405|Suspicious for Malignancy|suspicious for malignancy
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3473,3483|false|true|false|C0006826;C1306459|Malignant Neoplasms;Primary malignant neoplasm|malignancy
Event|Event|SIMPLE_SEGMENT|3473,3483|false|false|false|||malignancy
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3501,3504|false|false|false|C0032743;C0040398|Positron-Emission Tomography;Tomography, Emission-Computed|PET
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3501,3507|false|false|false|C1699633|PET/CT scan|PET-CT
Event|Event|SIMPLE_SEGMENT|3505,3507|false|false|false|||CT
Event|Event|SIMPLE_SEGMENT|3516,3529|false|false|false|||demonstration
Finding|Functional Concept|SIMPLE_SEGMENT|3535,3539|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3535,3546|false|false|false|C0222601|Left breast|left breast
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3540,3546|false|false|false|C0006141|Breast|breast
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3540,3546|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|breast
Finding|Finding|SIMPLE_SEGMENT|3540,3546|false|false|false|C0567499|Breast problem|breast
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3540,3546|false|false|false|C0191838|Procedures on breast|breast
Finding|Finding|SIMPLE_SEGMENT|3540,3554|false|false|false|C0024103|Mass in breast|breast nodules
Event|Event|SIMPLE_SEGMENT|3547,3554|false|false|false|||nodules
Event|Event|SIMPLE_SEGMENT|3566,3577|false|false|false|||correlation
Event|Event|SIMPLE_SEGMENT|3583,3594|false|false|false|||mammography
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3583,3594|false|false|false|C0024671;C0848600|Mammography;Mammography, Female|mammography
Event|Event|SIMPLE_SEGMENT|3599,3609|false|false|false|||ultrasound
Finding|Functional Concept|SIMPLE_SEGMENT|3599,3609|false|false|false|C0220934|Ultrasonic|ultrasound
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3599,3609|false|false|false|C0041621;C1456803|Ultrasonic Shockwave;Ultrasonics (sound)|ultrasound
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3599,3609|false|false|false|C0041618;C1315081|Ultrasonography;Urological ultrasound|ultrasound
Event|Event|SIMPLE_SEGMENT|3613,3622|false|false|false|||suggested
Event|Event|SIMPLE_SEGMENT|3625,3628|false|false|false|||EKG
Finding|Intellectual Product|SIMPLE_SEGMENT|3625,3628|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3625,3628|false|false|false|C1623258|Electrocardiography|EKG
Event|Event|SIMPLE_SEGMENT|3629,3635|false|false|false|||showed
Event|Event|SIMPLE_SEGMENT|3636,3639|false|false|false|||NSR
Finding|Molecular Function|SIMPLE_SEGMENT|3636,3639|false|false|false|C1704493;C2700623|Neutral Sidebent Rotated|NSR
Finding|Pathologic Function|SIMPLE_SEGMENT|3636,3639|false|false|false|C1704493;C2700623|Neutral Sidebent Rotated|NSR
Anatomy|Cell Component|SIMPLE_SEGMENT|3654,3657|false|false|false|C5239889|protein aggregate center|PAC
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3654,3657|false|false|false|C0033036|Atrial Premature Complexes|PAC
Event|Event|SIMPLE_SEGMENT|3654,3657|false|false|false|||PAC
Finding|Finding|SIMPLE_SEGMENT|3654,3657|false|false|false|C1823219;C4082832|Atrial Premature Complex by ECG Finding;PACC1 gene|PAC
Finding|Gene or Genome|SIMPLE_SEGMENT|3654,3657|false|false|false|C1823219;C4082832|Atrial Premature Complex by ECG Finding;PACC1 gene|PAC
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3654,3657|false|false|false|C0280547;C1879916|CAP Regimen;cisplatin/cyclophosphamide/doxorubicin protocol|PAC
Finding|Body Substance|SIMPLE_SEGMENT|3659,3666|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|3659,3666|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|3659,3666|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Organic Chemical|SIMPLE_SEGMENT|3694,3707|false|false|false|C0008809|ciprofloxacin|Ciprofloxacin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3694,3707|false|false|false|C0008809|ciprofloxacin|Ciprofloxacin
Drug|Antibiotic|SIMPLE_SEGMENT|3694,3711|false|false|false|C0282104|ciprofloxacin hydrochloride|Ciprofloxacin HCl
Drug|Organic Chemical|SIMPLE_SEGMENT|3694,3711|false|false|false|C0282104|ciprofloxacin hydrochloride|Ciprofloxacin HCl
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3708,3711|false|false|false|C0023443|Hairy Cell Leukemia|HCl
Drug|Immunologic Factor|SIMPLE_SEGMENT|3708,3711|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Inorganic Chemical|SIMPLE_SEGMENT|3708,3711|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3708,3711|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Event|Event|SIMPLE_SEGMENT|3708,3711|false|false|false|||HCl
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3733,3740|false|false|false|C0019134;C0770546|heparin;heparin, porcine|Heparin
Drug|Organic Chemical|SIMPLE_SEGMENT|3733,3740|false|false|false|C0019134;C0770546|heparin;heparin, porcine|Heparin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3733,3740|false|false|false|C0019134;C0770546|heparin;heparin, porcine|Heparin
Event|Event|SIMPLE_SEGMENT|3733,3740|false|false|false|||Heparin
Event|Event|SIMPLE_SEGMENT|3746,3750|false|false|false|||UNIT
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3765,3772|false|false|false|C0019134;C0770546|heparin;heparin, porcine|Heparin
Drug|Organic Chemical|SIMPLE_SEGMENT|3765,3772|false|false|false|C0019134;C0770546|heparin;heparin, porcine|Heparin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3765,3772|false|false|false|C0019134;C0770546|heparin;heparin, porcine|Heparin
Event|Event|SIMPLE_SEGMENT|3765,3772|false|false|false|||Heparin
Event|Event|SIMPLE_SEGMENT|3776,3784|false|false|false|||Transfer
Finding|Functional Concept|SIMPLE_SEGMENT|3776,3784|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|Transfer
Finding|Idea or Concept|SIMPLE_SEGMENT|3776,3784|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|Transfer
Procedure|Health Care Activity|SIMPLE_SEGMENT|3776,3784|false|false|false|C4706767|Transfer (immobility management)|Transfer
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3816,3821|false|false|false|C0028429||Nasal
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3816,3821|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Organic Chemical|SIMPLE_SEGMENT|3816,3821|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3816,3821|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Finding|Finding|SIMPLE_SEGMENT|3816,3821|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Finding|Functional Concept|SIMPLE_SEGMENT|3816,3821|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3822,3829|false|false|false|C1550232|Body Parts - Cannula|Cannula
Finding|Body Substance|SIMPLE_SEGMENT|3822,3829|false|false|false|C1546577;C1550622|Specimen Type - Cannula|Cannula
Finding|Intellectual Product|SIMPLE_SEGMENT|3822,3829|false|false|false|C1546577;C1550622|Specimen Type - Cannula|Cannula
Event|Event|SIMPLE_SEGMENT|3837,3841|false|false|false|||seen
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|3849,3854|false|false|false|C3714591|Floor (anatomic)|floor
Event|Event|SIMPLE_SEGMENT|3860,3867|false|false|false|||reports
Finding|Idea or Concept|SIMPLE_SEGMENT|3868,3879|false|false|false|C0750502|Significant|significant
Event|Event|SIMPLE_SEGMENT|3880,3887|false|false|false|||dyspnea
Finding|Finding|SIMPLE_SEGMENT|3880,3887|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|3880,3887|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Event|Event|SIMPLE_SEGMENT|3902,3910|false|false|false|||exertion
Finding|Organism Function|SIMPLE_SEGMENT|3902,3910|false|false|false|C0015264|Exertion|exertion
Event|Event|SIMPLE_SEGMENT|3912,3918|false|false|false|||Denies
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3919,3924|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|3919,3924|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3919,3929|true|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|3919,3929|true|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3925,3929|true|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|3925,3929|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|3925,3929|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|3925,3929|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|3931,3943|false|false|false|||palpitations
Finding|Finding|SIMPLE_SEGMENT|3931,3943|true|false|false|C0030252|Palpitations|palpitations
Event|Event|SIMPLE_SEGMENT|3946,3961|false|false|false|||lightheadedness
Finding|Sign or Symptom|SIMPLE_SEGMENT|3946,3961|false|false|false|C0220870|Lightheadedness|lightheadedness
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|3975,3978|false|false|false|C0262327|rostral sulcus|ROS
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3975,3978|false|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|3975,3978|false|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Drug|Organic Chemical|SIMPLE_SEGMENT|3975,3978|false|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3975,3978|false|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Event|Event|SIMPLE_SEGMENT|3975,3978|false|false|false|||ROS
Finding|Gene or Genome|SIMPLE_SEGMENT|3975,3978|false|false|false|C0812281;C1709820|ROS1 gene;ROS1 wt Allele|ROS
Procedure|Health Care Activity|SIMPLE_SEGMENT|3975,3978|false|false|false|C0489633|Review of systems (procedure)|ROS
Event|Event|SIMPLE_SEGMENT|3983,3992|false|false|false|||conducted
Event|Event|SIMPLE_SEGMENT|4001,4009|false|false|false|||negative
Finding|Classification|SIMPLE_SEGMENT|4001,4009|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|4001,4009|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4001,4009|false|false|false|C5237010|Expression Negative|negative
Finding|Idea or Concept|SIMPLE_SEGMENT|4020,4025|false|false|false|C1552828|Table Frame - above|above
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4034,4037|false|false|false|C0268529|Proline dehydrogenase deficiency|HPI
Event|Event|SIMPLE_SEGMENT|4034,4037|false|false|false|||HPI
Finding|Finding|SIMPLE_SEGMENT|4034,4037|false|false|false|C0262512;C1323983|History of present illness (finding);allene oxide synthase activity|HPI
Finding|Molecular Function|SIMPLE_SEGMENT|4034,4037|false|false|false|C0262512;C1323983|History of present illness (finding);allene oxide synthase activity|HPI
Finding|Finding|SIMPLE_SEGMENT|4041,4061|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Event|Event|SIMPLE_SEGMENT|4046,4053|false|false|false|||Medical
Finding|Functional Concept|SIMPLE_SEGMENT|4046,4053|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|4046,4053|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|4046,4053|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|4046,4053|false|false|false|C0199168|Medical service|Medical
Finding|Finding|SIMPLE_SEGMENT|4046,4061|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|4054,4061|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|4054,4061|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|4054,4061|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4063,4075|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|SIMPLE_SEGMENT|4063,4075|false|false|false|||Hypertension
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4077,4089|false|false|false|C0031150|Laparoscopy|laparoscopic
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4077,4105|false|false|false|C0162522|Cholecystectomy, Laparoscopic|laparoscopic cholecystectomy
Event|Event|SIMPLE_SEGMENT|4090,4105|false|false|false|||cholecystectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4090,4105|false|false|false|C0008320|Cholecystectomy procedure|cholecystectomy
Finding|Functional Concept|SIMPLE_SEGMENT|4107,4111|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4107,4116|false|false|false|C0230432;C4281599|Structure of left knee;Structure of left knee region|left knee
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4107,4116|false|false|false|C0230432;C4281599|Structure of left knee;Structure of left knee region|left knee
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4112,4116|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4112,4116|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4112,4116|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4112,4116|false|false|false|C0562271|Examination of knee joint|knee
Event|Event|SIMPLE_SEGMENT|4118,4129|false|false|false|||replacement
Finding|Functional Concept|SIMPLE_SEGMENT|4118,4129|false|false|false|C0559956|Replacement|replacement
Procedure|Health Care Activity|SIMPLE_SEGMENT|4118,4129|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|replacement
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4118,4129|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|replacement
Finding|Gene or Genome|SIMPLE_SEGMENT|4147,4150|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Event|Event|SIMPLE_SEGMENT|4152,4163|false|false|false|||laminectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4152,4163|false|false|false|C0022983|Laminectomy|laminectomy
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4176,4179|false|false|false|C1114365||age
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4176,4179|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|SIMPLE_SEGMENT|4176,4179|false|false|false|C0162574|Glycation End Products, Advanced|age
Event|Event|SIMPLE_SEGMENT|4176,4179|false|false|false|||age
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4190,4197|false|false|false|C0042232|Vagina|vaginal
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4190,4197|false|false|false|C1272941|Vaginal Dosage Form|vaginal
Finding|Finding|SIMPLE_SEGMENT|4190,4197|false|false|false|C1522570;C4521343|Vaginal (intended site);Vaginal Route of Administration|vaginal
Finding|Functional Concept|SIMPLE_SEGMENT|4190,4197|false|false|false|C1522570;C4521343|Vaginal (intended site);Vaginal Route of Administration|vaginal
Event|Event|SIMPLE_SEGMENT|4198,4208|false|false|false|||deliveries
Event|Event|SIMPLE_SEGMENT|4240,4252|false|false|false|||laparoscopic
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4240,4252|false|false|false|C0031150|Laparoscopy|laparoscopic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4263,4269|false|false|false|C0030797|Pelvis|pelvic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4263,4280|false|false|false|C0729595|Pelvic lymph node group|pelvic lymph node
Finding|Body Substance|SIMPLE_SEGMENT|4270,4275|false|false|false|C0024202|Lymph|lymph
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4270,4280|false|false|false|C0024204|lymph nodes|lymph node
Event|Event|SIMPLE_SEGMENT|4282,4292|false|false|false|||dissection
Finding|Pathologic Function|SIMPLE_SEGMENT|4282,4292|false|false|false|C0333288|Dissecting hemorrhage|dissection
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4282,4292|false|false|false|C0012737|Tissue Dissection|dissection
Event|Event|SIMPLE_SEGMENT|4312,4324|false|false|false|||hysterectomy
Finding|Finding|SIMPLE_SEGMENT|4312,4324|false|false|false|C1548863|Consent Type - Hysterectomy|hysterectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4312,4324|false|false|false|C0020699|Hysterectomy|hysterectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4329,4351|false|false|false|C0278321|Bilateral oophorectomy|bilateral oophorectomy
Event|Event|SIMPLE_SEGMENT|4339,4351|false|false|false|||oophorectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4339,4351|false|false|false|C0029936|Ovariectomy|oophorectomy
Finding|Gene or Genome|SIMPLE_SEGMENT|4357,4362|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Finding|Finding|SIMPLE_SEGMENT|4357,4369|false|false|false|C0151994|Enlarged uterus|large uterus
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4363,4369|false|false|false|C0042149;C1519876;C4266525|Mouse Uterus;Pelvis>Uterus;Uterus|uterus
Anatomy|Tissue|SIMPLE_SEGMENT|4363,4369|false|false|false|C0042149;C1519876;C4266525|Mouse Uterus;Pelvis>Uterus;Uterus|uterus
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4363,4369|false|false|false|C0042131;C0496919|Neoplasm of uncertain or unknown behavior of uterus;Uterine Diseases|uterus
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4363,4369|false|false|false|C0042131;C0496919|Neoplasm of uncertain or unknown behavior of uterus;Uterine Diseases|uterus
Event|Event|SIMPLE_SEGMENT|4363,4369|false|false|false|||uterus
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4363,4369|false|false|false|C0869889|examination of uterus|uterus
Finding|Gene or Genome|SIMPLE_SEGMENT|4400,4405|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4406,4413|false|false|false|C0023267|Fibroid Tumor|fibroid
Event|Event|SIMPLE_SEGMENT|4406,4413|false|false|false|||fibroid
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4418,4430|false|false|false|C0031150|Laparoscopy|Laparoscopic
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4418,4449|false|false|false|C5879917|Laparoscopic radical cystectomy|Laparoscopic radical cystectomy
Drug|Chemical Viewed Structurally|SIMPLE_SEGMENT|4431,4438|false|false|false|C0302912|Radicals (chemistry)|radical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4431,4449|false|false|false|C0194401|Complete cystectomy|radical cystectomy
Event|Event|SIMPLE_SEGMENT|4439,4449|false|false|false|||cystectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4439,4449|false|false|false|C0010651|Cystectomy|cystectomy
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4454,4462|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Event|Event|SIMPLE_SEGMENT|4463,4474|false|false|false|||vaginectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4463,4474|false|false|false|C0195130|Vaginectomy|vaginectomy
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4481,4488|false|false|false|C0042232|Vagina|vaginal
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4481,4488|false|false|false|C1272941|Vaginal Dosage Form|vaginal
Finding|Finding|SIMPLE_SEGMENT|4481,4488|false|false|false|C1522570;C4521343|Vaginal (intended site);Vaginal Route of Administration|vaginal
Finding|Functional Concept|SIMPLE_SEGMENT|4481,4488|false|false|false|C1522570;C4521343|Vaginal (intended site);Vaginal Route of Administration|vaginal
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4481,4503|false|false|false|C0195196|Reconstruction of vagina|vaginal reconstruction
Event|Event|SIMPLE_SEGMENT|4489,4503|false|false|false|||reconstruction
Procedure|Machine Activity|SIMPLE_SEGMENT|4489,4503|false|false|false|C0020912;C0524865|Optical Image Reconstruction;Reconstructive Surgical Procedures|reconstruction
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4489,4503|false|false|false|C0020912;C0524865|Optical Image Reconstruction;Reconstructive Surgical Procedures|reconstruction
Finding|Functional Concept|SIMPLE_SEGMENT|4508,4514|false|false|false|C0728831|Social|Social
Finding|Finding|SIMPLE_SEGMENT|4508,4522|false|false|false|C0424945;C3714536|Social History;Social and personal history|Social History
Event|Event|SIMPLE_SEGMENT|4515,4522|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|4515,4522|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|4515,4522|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|4515,4522|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Classification|SIMPLE_SEGMENT|4528,4534|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|SIMPLE_SEGMENT|4528,4534|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|SIMPLE_SEGMENT|4528,4534|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|SIMPLE_SEGMENT|4528,4534|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Finding|SIMPLE_SEGMENT|4528,4542|false|false|false|C0241889|Family Medical History|Family History
Event|Event|SIMPLE_SEGMENT|4535,4542|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|4535,4542|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|4535,4542|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|4535,4542|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Event|Event|SIMPLE_SEGMENT|4544,4552|false|false|false|||Negative
Finding|Classification|SIMPLE_SEGMENT|4544,4552|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|Negative
Finding|Finding|SIMPLE_SEGMENT|4544,4552|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|Negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4544,4552|false|false|false|C5237010|Expression Negative|Negative
Finding|Finding|SIMPLE_SEGMENT|4544,4556|false|false|false|C0205160|Negative|Negative for
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4557,4564|false|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4557,4564|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Event|Event|SIMPLE_SEGMENT|4557,4564|false|false|false|||bladder
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4557,4564|false|false|false|C0872388|Procedures on bladder|bladder
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4557,4567|false|true|false|C0005684|Malignant neoplasm of urinary bladder|bladder CA
Event|Event|SIMPLE_SEGMENT|4572,4580|false|false|false|||Physical
Finding|Finding|SIMPLE_SEGMENT|4572,4580|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|4572,4580|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|4572,4580|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|4572,4585|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|4572,4585|false|false|false|C0031809|Physical Examination|Physical Exam
Event|Event|SIMPLE_SEGMENT|4581,4585|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|4581,4585|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|4581,4585|false|false|false|C0582103|Medical Examination|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|4587,4596|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|SIMPLE_SEGMENT|4597,4601|false|false|false|||EXAM
Finding|Functional Concept|SIMPLE_SEGMENT|4597,4601|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|SIMPLE_SEGMENT|4597,4601|false|false|false|C0582103|Medical Examination|EXAM
Finding|Classification|SIMPLE_SEGMENT|4604,4607|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Finding|Gene or Genome|SIMPLE_SEGMENT|4604,4607|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4609,4612|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4609,4612|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4609,4612|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|4609,4612|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4609,4612|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|SIMPLE_SEGMENT|4609,4612|false|false|false|||NAD
Finding|Finding|SIMPLE_SEGMENT|4609,4612|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Event|Event|SIMPLE_SEGMENT|4614,4622|false|false|false|||speaking
Finding|Idea or Concept|SIMPLE_SEGMENT|4628,4632|false|false|false|C1705313|Term (lexical)|word
Event|Event|SIMPLE_SEGMENT|4633,4642|false|false|false|||sentences
Finding|Intellectual Product|SIMPLE_SEGMENT|4633,4642|false|false|false|C0876929|Sentence|sentences
Event|Event|SIMPLE_SEGMENT|4644,4650|false|false|false|||pursed
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4651,4654|false|false|false|C0023759|Lip structure|lip
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4651,4654|false|false|false|C0153932;C0264511|Benign neoplasm of the lip;Lymphoid interstitial pneumonia|lip
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4651,4654|false|false|false|C0153932;C0264511|Benign neoplasm of the lip;Lymphoid interstitial pneumonia|lip
Finding|Gene or Genome|SIMPLE_SEGMENT|4651,4654|false|false|false|C1846919;C3889123|SMG1 gene;SMG1 wt Allele|lip
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4655,4664|false|false|false|C5885990||breathing
Event|Event|SIMPLE_SEGMENT|4655,4664|false|false|false|||breathing
Finding|Finding|SIMPLE_SEGMENT|4655,4664|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|SIMPLE_SEGMENT|4655,4664|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|SIMPLE_SEGMENT|4655,4664|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|SIMPLE_SEGMENT|4655,4664|false|false|false|C1160636|respiratory system process|breathing
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|4670,4686|true|false|false|C0158784|Accessory skeletal muscle|accessory muscle
Finding|Finding|SIMPLE_SEGMENT|4670,4690|true|false|false|C1821466|Use of accessory muscles|accessory muscle use
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4680,4686|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Anatomy|Tissue|SIMPLE_SEGMENT|4680,4686|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Event|Event|SIMPLE_SEGMENT|4687,4690|false|false|false|||use
Finding|Functional Concept|SIMPLE_SEGMENT|4687,4690|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|SIMPLE_SEGMENT|4687,4690|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Event|Event|SIMPLE_SEGMENT|4692,4697|false|false|false|||lying
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4701,4704|false|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Event|Event|SIMPLE_SEGMENT|4701,4704|false|false|false|||bed
Finding|Intellectual Product|SIMPLE_SEGMENT|4701,4704|false|false|false|C2346952|Bachelor of Education|bed
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4706,4710|false|false|false|C0015392|Eye|Eyes
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4706,4710|false|false|false|C5848506||Eyes
Event|Event|SIMPLE_SEGMENT|4712,4716|false|false|false|||EOMI
Event|Event|SIMPLE_SEGMENT|4726,4735|false|false|false|||anicteric
Finding|Finding|SIMPLE_SEGMENT|4726,4735|false|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4739,4742|false|false|false|C0150934;C0175196|Ear, nose and throat;Structure of entorhinal cortex|ENT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4739,4742|false|false|false|C0150934;C0175196|Ear, nose and throat;Structure of entorhinal cortex|ENT
Finding|Gene or Genome|SIMPLE_SEGMENT|4739,4742|false|false|false|C0262471;C1417861;C3889152|ENT problem;NT5E gene;NT5E wt Allele|ENT
Finding|Sign or Symptom|SIMPLE_SEGMENT|4739,4742|false|false|false|C0262471;C1417861;C3889152|ENT problem;NT5E gene;NT5E wt Allele|ENT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4744,4747|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4744,4747|false|false|false|C0026987|Myelofibrosis|MMM
Event|Event|SIMPLE_SEGMENT|4744,4747|false|false|false|||MMM
Event|Event|SIMPLE_SEGMENT|4752,4757|false|false|false|||clear
Finding|Idea or Concept|SIMPLE_SEGMENT|4752,4757|false|false|false|C1550016|Remote control command - Clear|clear
Event|Event|SIMPLE_SEGMENT|4771,4774|false|false|false|||RRR
Event|Event|SIMPLE_SEGMENT|4779,4782|false|false|false|||MRG
Finding|Gene or Genome|SIMPLE_SEGMENT|4779,4782|true|false|false|C1422304|MAS1L gene|MRG
Drug|Food|SIMPLE_SEGMENT|4789,4795|false|false|false|C5890763||pulses
Event|Event|SIMPLE_SEGMENT|4789,4795|false|false|false|||pulses
Finding|Physiologic Function|SIMPLE_SEGMENT|4789,4795|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|SIMPLE_SEGMENT|4789,4795|false|false|false|C0034107|Pulse taking|pulses
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4800,4805|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|4800,4805|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|4800,4805|false|false|false|C0013604|Edema|edema
Event|Event|SIMPLE_SEGMENT|4824,4835|false|false|false|||compression
Finding|Functional Concept|SIMPLE_SEGMENT|4824,4835|false|false|false|C0332459;C4551657|Compressed structure|compression
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|4824,4835|false|false|false|C0728907|Compression|compression
Procedure|Machine Activity|SIMPLE_SEGMENT|4824,4835|false|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4824,4835|false|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Event|Event|SIMPLE_SEGMENT|4836,4845|false|false|false|||stockings
Event|Activity|SIMPLE_SEGMENT|4849,4854|false|false|false|C1882509|put - instruction imperative|place
Event|Event|SIMPLE_SEGMENT|4849,4854|false|false|false|||place
Finding|Functional Concept|SIMPLE_SEGMENT|4849,4854|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|SIMPLE_SEGMENT|4849,4854|false|false|false|C1533810||place
Event|Event|SIMPLE_SEGMENT|4859,4862|false|false|false|||JVD
Finding|Finding|SIMPLE_SEGMENT|4859,4862|true|false|false|C0425687|Jugular venous engorgement|JVD
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4865,4869|false|false|false|C0231832|Respiratory rate|Resp
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4865,4869|false|false|false|C0851355|Respiratory, thoracic and mediastinal disorders|Resp
Event|Event|SIMPLE_SEGMENT|4865,4869|false|false|false|||Resp
Event|Event|SIMPLE_SEGMENT|4878,4884|false|false|false|||effort
Finding|Organism Function|SIMPLE_SEGMENT|4878,4884|false|false|false|C0015264|Exertion|effort
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|4889,4905|true|false|false|C0158784|Accessory skeletal muscle|accessory muscle
Finding|Finding|SIMPLE_SEGMENT|4889,4909|true|false|false|C1821466|Use of accessory muscles|accessory muscle use
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4899,4905|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Anatomy|Tissue|SIMPLE_SEGMENT|4899,4905|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Event|Event|SIMPLE_SEGMENT|4906,4909|false|false|false|||use
Finding|Functional Concept|SIMPLE_SEGMENT|4906,4909|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|SIMPLE_SEGMENT|4906,4909|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4911,4916|false|false|false|C0024109|Lung|lungs
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4917,4920|false|false|false|C3813556|Cancer/Testis Antigen|CTA
Event|Event|SIMPLE_SEGMENT|4917,4920|false|false|false|||CTA
Finding|Gene or Genome|SIMPLE_SEGMENT|4917,4920|false|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4917,4920|false|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4929,4937|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Event|Event|SIMPLE_SEGMENT|4938,4950|false|false|false|||auscultation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4938,4950|false|false|false|C0004339|Auscultation|auscultation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4957,4961|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|SIMPLE_SEGMENT|4957,4961|false|false|false|||soft
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|4976,4984|false|false|false|C0559495|Urological stoma|Urostomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4976,4984|false|false|false|C0856443|Urostomy procedure|Urostomy
Finding|Finding|SIMPLE_SEGMENT|4976,4989|false|false|false|C4053891|Urostomy Site|Urostomy site
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4985,4989|false|false|false|C1515974|Anatomic Site|site
Finding|Intellectual Product|SIMPLE_SEGMENT|4985,4989|false|false|false|C1546778||site
Event|Event|SIMPLE_SEGMENT|4999,5005|false|false|false|||appear
Event|Event|SIMPLE_SEGMENT|5006,5014|false|false|false|||infected
Finding|Finding|SIMPLE_SEGMENT|5006,5014|false|true|false|C0439663|Infected|infected
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|5016,5019|false|false|false|C0022681|Medullary sponge kidney|MSK
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5016,5019|false|false|false|C0022681|Medullary sponge kidney|MSK
Event|Event|SIMPLE_SEGMENT|5016,5019|false|false|false|||MSK
Finding|Gene or Genome|SIMPLE_SEGMENT|5016,5019|false|false|false|C1420279|SIK1 gene|MSK
Finding|Idea or Concept|SIMPLE_SEGMENT|5024,5035|false|false|false|C0750502|Significant|significant
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|5036,5044|true|false|false|C0022821;C0022822;C0265673|Acquired kyphosis;Congenital kyphosis;Kyphosis deformity of spine|kyphosis
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|5036,5044|true|false|false|C0022821;C0022822;C0265673|Acquired kyphosis;Congenital kyphosis;Kyphosis deformity of spine|kyphosis
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|5036,5044|true|false|false|C0022821;C0022822;C0265673|Acquired kyphosis;Congenital kyphosis;Kyphosis deformity of spine|kyphosis
Event|Event|SIMPLE_SEGMENT|5036,5044|false|false|false|||kyphosis
Finding|Finding|SIMPLE_SEGMENT|5036,5044|true|false|false|C2115817|kyphosis|kyphosis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5058,5067|true|false|false|C0039103|Synovitis|synovitis
Event|Event|SIMPLE_SEGMENT|5058,5067|false|false|false|||synovitis
Anatomy|Body System|SIMPLE_SEGMENT|5070,5074|false|false|false|C1123023;C4520765|Skin;Skin, Human|Skin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5070,5074|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|Skin
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5070,5074|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|Skin
Finding|Body Substance|SIMPLE_SEGMENT|5070,5074|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|Skin
Finding|Intellectual Product|SIMPLE_SEGMENT|5070,5074|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|Skin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5087,5091|true|false|false|C5779629|Eruption of skin (disorder)|rash
Event|Event|SIMPLE_SEGMENT|5087,5091|false|false|false|||rash
Finding|Pathologic Function|SIMPLE_SEGMENT|5087,5091|true|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Sign or Symptom|SIMPLE_SEGMENT|5087,5091|true|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Event|Event|SIMPLE_SEGMENT|5096,5104|false|false|false|||jaundice
Finding|Finding|SIMPLE_SEGMENT|5096,5104|true|false|false|C0022346;C2010848;C2203646|Icterus;jaundice;yellow skin or eyes (symptom)|jaundice
Finding|Sign or Symptom|SIMPLE_SEGMENT|5096,5104|true|false|false|C0022346;C2010848;C2203646|Icterus;jaundice;yellow skin or eyes (symptom)|jaundice
Event|Event|SIMPLE_SEGMENT|5114,5119|false|false|false|||AAOx3
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5124,5130|false|false|false|C0015450|Face|facial
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5124,5136|true|false|false|C0427055|Facial Paresis|facial droop
Finding|Finding|SIMPLE_SEGMENT|5124,5136|true|false|false|C4022719|Unilateral facial palsy|facial droop
Event|Event|SIMPLE_SEGMENT|5131,5136|false|false|false|||droop
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|5139,5144|false|false|false|C0004936;C1306597|Mental disorders;Psychiatric problem|Psych
Event|Event|SIMPLE_SEGMENT|5139,5144|false|false|false|||Psych
Event|Event|SIMPLE_SEGMENT|5151,5156|false|false|false|||range
Finding|Intellectual Product|SIMPLE_SEGMENT|5151,5156|false|false|false|C3542016|Concept model range (foundation metadata concept)|range
Event|Event|SIMPLE_SEGMENT|5160,5166|false|false|false|||affect
Finding|Mental Process|SIMPLE_SEGMENT|5160,5166|false|false|false|C0001721|Affect (mental function)|affect
Procedure|Health Care Activity|SIMPLE_SEGMENT|5160,5166|false|false|false|C2237113|assessment of affect|affect
Finding|Body Substance|SIMPLE_SEGMENT|5169,5178|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|5169,5178|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|5169,5178|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|5169,5178|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|SIMPLE_SEGMENT|5179,5183|false|false|false|||EXAM
Finding|Functional Concept|SIMPLE_SEGMENT|5179,5183|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|SIMPLE_SEGMENT|5179,5183|false|false|false|C0582103|Medical Examination|EXAM
Event|Event|SIMPLE_SEGMENT|5185,5191|false|false|false|||vitals
Finding|Classification|SIMPLE_SEGMENT|5218,5221|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Finding|Gene or Genome|SIMPLE_SEGMENT|5218,5221|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Event|Event|SIMPLE_SEGMENT|5223,5228|false|false|false|||Lying
Finding|Individual Behavior|SIMPLE_SEGMENT|5223,5228|false|false|false|C0600261|Telling untruths|Lying
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5232,5235|false|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Finding|Intellectual Product|SIMPLE_SEGMENT|5232,5235|false|false|false|C2346952|Bachelor of Education|bed
Finding|Idea or Concept|SIMPLE_SEGMENT|5242,5250|true|false|false|C0750489|apparent|apparent
Event|Event|SIMPLE_SEGMENT|5251,5259|false|false|false|||distress
Finding|Finding|SIMPLE_SEGMENT|5251,5259|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|SIMPLE_SEGMENT|5251,5259|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5260,5265|false|false|false|C1512338|HEENT|HEENT
Event|Event|SIMPLE_SEGMENT|5267,5276|false|false|false|||Anicteric
Finding|Finding|SIMPLE_SEGMENT|5267,5276|false|false|false|C0205180|Anicteric|Anicteric
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5278,5281|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5278,5281|false|false|false|C0026987|Myelofibrosis|MMM
Anatomy|Body System|SIMPLE_SEGMENT|5282,5296|false|false|false|C0007226;C3887460|Cardiovascular;Cardiovascular system|Cardiovascular
Event|Event|SIMPLE_SEGMENT|5298,5301|false|false|false|||RRR
Finding|Functional Concept|SIMPLE_SEGMENT|5320,5325|true|false|false|C1552823|Table Cell Horizontal Align - right|right
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5332,5337|true|false|false|C3714496|Chronic obstructive pulmonary disease of horses|heave
Event|Event|SIMPLE_SEGMENT|5332,5337|false|false|false|||heave
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|5344,5352|false|false|false|C0039155|Systole|systolic
Finding|Finding|SIMPLE_SEGMENT|5344,5359|false|false|false|C0232257|Systolic Murmurs|systolic murmur
Event|Event|SIMPLE_SEGMENT|5353,5359|false|false|false|||murmur
Finding|Finding|SIMPLE_SEGMENT|5353,5359|false|false|false|C0018808|Heart murmur|murmur
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5361,5370|false|false|false|C0024109|Lung|Pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5361,5370|false|false|false|C2707265||Pulmonary
Finding|Finding|SIMPLE_SEGMENT|5361,5370|false|false|false|C4522268|Pulmonary (intended site)|Pulmonary
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5372,5376|false|false|false|C0024109;C4037972|Chest>Lung;Lung|Lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5372,5376|false|false|false|C0024109;C4037972|Chest>Lung;Lung|Lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5372,5376|false|false|false|C0024115|Lung diseases|Lung
Finding|Finding|SIMPLE_SEGMENT|5372,5376|false|false|false|C0740941|Lung Problem|Lung
Event|Event|SIMPLE_SEGMENT|5377,5383|false|false|false|||fields
Event|Event|SIMPLE_SEGMENT|5384,5389|false|false|false|||clear
Finding|Idea or Concept|SIMPLE_SEGMENT|5384,5389|false|false|false|C1550016|Remote control command - Clear|clear
Event|Event|SIMPLE_SEGMENT|5393,5405|false|false|false|||auscultation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5393,5405|false|false|false|C0004339|Auscultation|auscultation
Event|Event|SIMPLE_SEGMENT|5422,5430|false|false|false|||crackles
Finding|Finding|SIMPLE_SEGMENT|5422,5430|false|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Event|Event|SIMPLE_SEGMENT|5434,5442|false|false|false|||wheezing
Finding|Sign or Symptom|SIMPLE_SEGMENT|5434,5442|false|false|false|C0043144|Wheezing|wheezing
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5449,5453|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Event|Event|SIMPLE_SEGMENT|5449,5453|false|false|false|||Soft
Event|Event|SIMPLE_SEGMENT|5455,5464|false|false|false|||distended
Finding|Finding|SIMPLE_SEGMENT|5455,5464|false|false|false|C0700124|Dilated|distended
Event|Event|SIMPLE_SEGMENT|5466,5475|false|false|false|||nontender
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5477,5482|false|false|false|C0021853|Intestines|bowel
Finding|Finding|SIMPLE_SEGMENT|5477,5489|false|false|false|C0232693|Bowel sounds|bowel sounds
Event|Event|SIMPLE_SEGMENT|5483,5489|false|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|5483,5489|false|false|false|C0037709||sounds
Finding|Finding|SIMPLE_SEGMENT|5490,5497|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|SIMPLE_SEGMENT|5490,5497|false|false|false|C0150312;C0449450|Present;Presentation|present
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|5499,5507|false|false|false|C0559495|Urological stoma|urostomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5499,5507|false|false|false|C0856443|Urostomy procedure|urostomy
Event|Activity|SIMPLE_SEGMENT|5512,5517|false|false|false|C1882509|put - instruction imperative|place
Event|Event|SIMPLE_SEGMENT|5512,5517|false|false|false|||place
Finding|Functional Concept|SIMPLE_SEGMENT|5512,5517|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|SIMPLE_SEGMENT|5512,5517|false|false|false|C1533810||place
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5519,5530|false|false|false|C0015385;C0278454|All extremities;Limb structure|Extremities
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5535,5540|true|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|5535,5540|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|5535,5540|true|false|false|C0013604|Edema|edema
Finding|Functional Concept|SIMPLE_SEGMENT|5549,5553|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5549,5557|false|false|false|C0230416;C0230443|Left lower extremity;Structure of left lower leg|left leg
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5554,5557|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Event|Event|SIMPLE_SEGMENT|5566,5572|false|false|false|||larger
Event|Event|SIMPLE_SEGMENT|5578,5583|false|false|false|||right
Finding|Functional Concept|SIMPLE_SEGMENT|5578,5583|false|true|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5585,5588|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Event|Event|SIMPLE_SEGMENT|5590,5594|false|false|false|||warm
Finding|Finding|SIMPLE_SEGMENT|5590,5594|false|false|false|C0582051|Feels warm|warm
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|5590,5594|false|false|false|C0687712|warming process|warm
Finding|Finding|SIMPLE_SEGMENT|5596,5600|false|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|5601,5609|false|false|false|||perfused
Finding|Functional Concept|SIMPLE_SEGMENT|5615,5620|false|false|false|C1513492|motor movement|motor
Finding|Finding|SIMPLE_SEGMENT|5615,5629|false|false|false|C5551447|Motor function (finding)|motor function
Phenomenon|Biologic Function|SIMPLE_SEGMENT|5615,5629|false|false|false|C0234130|Motor function (observable entity)|motor function
Event|Event|SIMPLE_SEGMENT|5621,5629|false|false|false|||function
Finding|Finding|SIMPLE_SEGMENT|5621,5629|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|SIMPLE_SEGMENT|5621,5629|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|SIMPLE_SEGMENT|5621,5629|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|SIMPLE_SEGMENT|5621,5629|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Event|Event|SIMPLE_SEGMENT|5630,5636|false|false|false|||intact
Finding|Finding|SIMPLE_SEGMENT|5630,5636|false|false|false|C1554187|Gender Status - Intact|intact
Finding|Functional Concept|SIMPLE_SEGMENT|5642,5646|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5648,5653|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|5648,5653|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5648,5657|false|false|false|C1140621;C4299093|Leg;Lower extremity>Lower leg|lower leg
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5654,5657|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Event|Event|SIMPLE_SEGMENT|5661,5668|false|false|false|||wrapped
Event|Event|SIMPLE_SEGMENT|5693,5697|false|false|false|||LABS
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5693,5697|false|false|false|C0587081|Laboratory test finding|LABS
Procedure|Health Care Activity|SIMPLE_SEGMENT|5726,5735|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5736,5740|false|false|false|C0587081|Laboratory test finding|labs
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5756,5763|false|false|false|C0017725|glucose|GLUCOSE
Drug|Organic Chemical|SIMPLE_SEGMENT|5756,5763|false|false|false|C0017725|glucose|GLUCOSE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5756,5763|false|false|false|C0017725|glucose|GLUCOSE
Event|Event|SIMPLE_SEGMENT|5756,5763|false|false|false|||GLUCOSE
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5756,5763|false|false|false|C5781949|Glucose^1.5H post dose glucagon|GLUCOSE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5756,5763|false|false|false|C0337438|Glucose measurement|GLUCOSE
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5769,5773|false|false|false|C0041942|urea|UREA
Drug|Organic Chemical|SIMPLE_SEGMENT|5769,5773|false|false|false|C0041942|urea|UREA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5769,5773|false|false|false|C0041942|urea|UREA
Event|Event|SIMPLE_SEGMENT|5769,5773|false|false|false|||UREA
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5769,5773|false|false|false|C0523961|Urea measurement|UREA
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5790,5796|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|5790,5796|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5790,5796|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Event|Event|SIMPLE_SEGMENT|5790,5796|false|false|false|||SODIUM
Finding|Physiologic Function|SIMPLE_SEGMENT|5790,5796|false|false|false|C4553025|Sodium metabolic function|SODIUM
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5790,5796|false|false|false|C0337443|Sodium measurement|SODIUM
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5802,5811|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|5802,5811|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Food|SIMPLE_SEGMENT|5802,5811|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5802,5811|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5802,5811|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Event|Event|SIMPLE_SEGMENT|5802,5811|false|false|false|||POTASSIUM
Finding|Physiologic Function|SIMPLE_SEGMENT|5802,5811|false|false|false|C4553027|Potassium metabolic function|POTASSIUM
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5802,5811|false|false|false|C0202194|Potassium measurement|POTASSIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|5816,5824|false|false|false|C0008203;C0596019|Chlorides;chloride ion|CHLORIDE
Event|Event|SIMPLE_SEGMENT|5816,5824|false|false|false|||CHLORIDE
Finding|Physiologic Function|SIMPLE_SEGMENT|5816,5824|false|false|false|C4553021|Chloride metabolic function|CHLORIDE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5816,5824|false|false|false|C0201952|Chloride measurement|CHLORIDE
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5834,5837|false|false|false|C0007012|carbon dioxide|CO2
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5834,5837|false|false|false|C0007012|carbon dioxide|CO2
Event|Event|SIMPLE_SEGMENT|5834,5837|false|false|false|||CO2
Finding|Finding|SIMPLE_SEGMENT|5834,5837|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Finding|Gene or Genome|SIMPLE_SEGMENT|5834,5837|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|5841,5846|false|false|false|C0003075|Anions|ANION
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5841,5850|false|false|false|C0003074|Anion Gap|ANION GAP
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5841,5850|false|false|false|C1509129|Anion gap result|ANION GAP
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5841,5850|false|false|false|C0201889;C2189246|Anion gap measurement;blood anion gap (lab test)|ANION GAP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5847,5850|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5847,5850|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Event|Event|SIMPLE_SEGMENT|5847,5850|false|false|false|||GAP
Finding|Gene or Genome|SIMPLE_SEGMENT|5847,5850|false|false|false|C1419277;C2984552|RASA1 gene;RASA1 wt Allele|GAP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5896,5902|false|false|false|C5574646|Natriuretic Peptides B, human|proBNP
Drug|Hormone|SIMPLE_SEGMENT|5896,5902|false|false|false|C5574646|Natriuretic Peptides B, human|proBNP
Event|Event|SIMPLE_SEGMENT|5896,5902|false|false|false|||proBNP
Anatomy|Cell|SIMPLE_SEGMENT|5921,5924|false|false|false|C0023516|Leukocytes|WBC
Event|Event|SIMPLE_SEGMENT|5921,5924|false|false|false|||WBC
Anatomy|Cell|SIMPLE_SEGMENT|5929,5932|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5929,5932|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5929,5932|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5939,5942|false|false|false|C0019046|Hemoglobin|HGB
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5939,5942|false|false|false|C0019046|Hemoglobin|HGB
Event|Event|SIMPLE_SEGMENT|5939,5942|false|false|false|||HGB
Finding|Gene or Genome|SIMPLE_SEGMENT|5939,5942|false|false|false|C1424337|CYGB gene|HGB
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5939,5942|false|false|false|C0019029|Hemoglobin concentration|HGB
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5948,5951|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5948,5951|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Disorder|Virus|SIMPLE_SEGMENT|5958,5961|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|5958,5961|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5958,5961|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5958,5961|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5958,5961|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|5966,5969|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5966,5969|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|5966,5969|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|5966,5969|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|5966,5969|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5966,5969|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|SIMPLE_SEGMENT|5975,5979|false|false|false|||MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5975,5979|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Event|Event|SIMPLE_SEGMENT|6021,6024|false|false|false|||PLT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6021,6024|false|false|false|C0201617|Primed lymphocyte test|PLT
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6054,6057|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|SIMPLE_SEGMENT|6054,6057|false|false|false|||PTT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6054,6057|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Finding|Body Substance|SIMPLE_SEGMENT|6068,6077|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|6068,6077|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|6068,6077|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|6068,6077|false|false|false|C0030685|Patient Discharge|Discharge
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6078,6082|false|false|false|C0587081|Laboratory test finding|labs
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6096,6101|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|6096,6101|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|6096,6101|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|6102,6105|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|6112,6115|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6112,6115|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6112,6115|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6122,6125|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6122,6125|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|6122,6125|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6122,6125|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6131,6134|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6131,6134|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|6142,6145|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|6142,6145|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6142,6145|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6142,6145|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6142,6145|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|6149,6152|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6149,6152|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|6149,6152|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|6149,6152|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|6149,6152|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6149,6152|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|SIMPLE_SEGMENT|6158,6162|false|false|false|||MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6158,6162|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6190,6193|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6210,6215|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|6210,6215|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|6210,6215|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|6210,6223|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6210,6223|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6210,6223|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6216,6223|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|6216,6223|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6216,6223|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|6216,6223|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6216,6223|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6216,6223|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|SIMPLE_SEGMENT|6267,6271|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6267,6271|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6267,6271|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6296,6301|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|6296,6301|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|6296,6301|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6296,6309|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6302,6309|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|6302,6309|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|6302,6309|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6302,6309|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|6302,6309|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|SIMPLE_SEGMENT|6302,6309|false|false|false|||Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|6302,6309|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6302,6309|false|false|false|C0201925|Calcium measurement|Calcium
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6343,6348|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|6343,6348|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|6343,6348|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6375,6378|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6375,6378|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Drug|Hormone|SIMPLE_SEGMENT|6375,6378|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6375,6378|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Finding|Gene or Genome|SIMPLE_SEGMENT|6375,6378|false|false|false|C1334121;C1336604;C1705002|IL5 gene;TERF1 gene;TERF1 wt Allele|TRF
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6396,6401|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|6396,6401|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|6396,6401|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6396,6406|false|false|false|C0853169|Blood iron measurement|BLOOD Iron
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6402,6406|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|6402,6406|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6402,6406|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Event|Event|SIMPLE_SEGMENT|6402,6406|false|false|false|||Iron
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6402,6406|false|false|false|C0337439|Iron measurement|Iron
Event|Event|SIMPLE_SEGMENT|6412,6424|false|false|false|||MICROBIOLOGY
Finding|Functional Concept|SIMPLE_SEGMENT|6412,6424|false|false|false|C0025953;C1571921;C4049106|Microbiological;Microbiology - Laboratory Class;Microbiology Diagnostic Service Section ID|MICROBIOLOGY
Finding|Intellectual Product|SIMPLE_SEGMENT|6412,6424|false|false|false|C0025953;C1571921;C4049106|Microbiological;Microbiology - Laboratory Class;Microbiology Diagnostic Service Section ID|MICROBIOLOGY
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6412,6424|false|false|false|C0085672|Microbiology procedure|MICROBIOLOGY
Finding|Body Substance|SIMPLE_SEGMENT|6464,6469|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|6464,6469|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|6464,6469|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Idea or Concept|SIMPLE_SEGMENT|6501,6506|false|false|false|C1546485|Diagnosis Type - Final|FINAL
Finding|Intellectual Product|SIMPLE_SEGMENT|6501,6513|false|false|false|C0460114|Final report|FINAL REPORT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6507,6513|false|false|false|C4255046||REPORT
Event|Event|SIMPLE_SEGMENT|6507,6513|false|false|false|||REPORT
Finding|Intellectual Product|SIMPLE_SEGMENT|6507,6513|false|false|false|C0684224|Report (document)|REPORT
Procedure|Health Care Activity|SIMPLE_SEGMENT|6507,6513|false|false|false|C0700287|Reporting|REPORT
Finding|Body Substance|SIMPLE_SEGMENT|6522,6527|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|6522,6527|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|6522,6527|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6522,6535|false|false|false|C0430404|Urine culture|URINE CULTURE
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6528,6535|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|SIMPLE_SEGMENT|6528,6535|false|false|false|||CULTURE
Finding|Functional Concept|SIMPLE_SEGMENT|6528,6535|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|SIMPLE_SEGMENT|6528,6535|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6528,6535|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Event|Event|SIMPLE_SEGMENT|6537,6542|false|false|false|||Final
Finding|Idea or Concept|SIMPLE_SEGMENT|6537,6542|false|false|false|C1546485|Diagnosis Type - Final|Final
Event|Event|SIMPLE_SEGMENT|6555,6560|false|false|false|||MIXED
Anatomy|Cell|SIMPLE_SEGMENT|6584,6590|false|false|false|C1947989|Colony (cells or organisms)|COLONY
Event|Event|SIMPLE_SEGMENT|6599,6609|false|false|false|||CONSISTENT
Finding|Idea or Concept|SIMPLE_SEGMENT|6599,6609|false|false|false|C0332290|Consistent with|CONSISTENT
Anatomy|Body System|SIMPLE_SEGMENT|6616,6620|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6616,6620|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6616,6620|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Event|Event|SIMPLE_SEGMENT|6616,6620|false|false|false|||SKIN
Finding|Body Substance|SIMPLE_SEGMENT|6616,6620|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|SIMPLE_SEGMENT|6616,6620|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Event|Event|SIMPLE_SEGMENT|6630,6631|false|false|false|||/
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6634,6641|false|false|false|C0017420;C0559522|Genital system;Genitalia|GENITAL
Anatomy|Body System|SIMPLE_SEGMENT|6634,6641|false|false|false|C0017420;C0559522|Genital system;Genitalia|GENITAL
Finding|Body Substance|SIMPLE_SEGMENT|6634,6641|false|false|false|C1546649;C1550642|Specimen Type - Genital|GENITAL
Finding|Intellectual Product|SIMPLE_SEGMENT|6634,6641|false|false|false|C1546649;C1550642|Specimen Type - Genital|GENITAL
Event|Event|SIMPLE_SEGMENT|6642,6655|false|false|false|||CONTAMINATION
Finding|Idea or Concept|SIMPLE_SEGMENT|6642,6655|false|false|false|C2349974|Contamination|CONTAMINATION
Phenomenon|Human-caused Phenomenon or Process|SIMPLE_SEGMENT|6642,6655|false|false|false|C0259846|adulteration|CONTAMINATION
Event|Event|SIMPLE_SEGMENT|6677,6679|false|false|false|||SP
Finding|Functional Concept|SIMPLE_SEGMENT|6735,6744|false|false|false|C1285553|Interprets|INTERPRET
Event|Event|SIMPLE_SEGMENT|6745,6752|false|false|false|||RESULTS
Event|Event|SIMPLE_SEGMENT|6758,6765|false|false|false|||CAUTION
Event|Event|SIMPLE_SEGMENT|6799,6812|false|false|false|||SENSITIVITIES
Finding|Finding|SIMPLE_SEGMENT|6799,6812|false|false|false|C0427965|Antimicrobial susceptibility|SENSITIVITIES
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6814,6817|false|false|false|C2732473|Ductal Carcinoma In Situ with Microinvasion|MIC
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|6814,6817|false|false|false|C0066256|methyl isocyanate|MIC
Drug|Organic Chemical|SIMPLE_SEGMENT|6814,6817|false|false|false|C0066256|methyl isocyanate|MIC
Event|Event|SIMPLE_SEGMENT|6814,6817|false|false|false|||MIC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6814,6817|false|false|false|C0281162;C0427978|Minimum Inhibitory Concentration Test;cisplatin/ifosfamide/mitomycin protocol|MIC
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6814,6817|false|false|false|C0281162;C0427978|Minimum Inhibitory Concentration Test;cisplatin/ifosfamide/mitomycin protocol|MIC
Event|Event|SIMPLE_SEGMENT|6832,6835|false|false|false|||MCG
Event|Event|SIMPLE_SEGMENT|6962,6964|false|false|false|||SP
Drug|Antibiotic|SIMPLE_SEGMENT|7000,7010|false|false|false|C0002680;C2095775|ampicillin;ampicillins|AMPICILLIN
Drug|Organic Chemical|SIMPLE_SEGMENT|7000,7010|false|false|false|C0002680;C2095775|ampicillin;ampicillins|AMPICILLIN
Drug|Organic Chemical|SIMPLE_SEGMENT|7031,7045|false|false|false|C0028156|nitrofurantoin|NITROFURANTOIN
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7031,7045|false|false|false|C0028156|nitrofurantoin|NITROFURANTOIN
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|7062,7074|false|false|false|C0481114|Tetracyclines causing adverse effects in therapeutic use|TETRACYCLINE
Drug|Antibiotic|SIMPLE_SEGMENT|7062,7074|false|false|false|C0039644;C1744619|Tetracycline Antibiotics;tetracycline|TETRACYCLINE
Drug|Organic Chemical|SIMPLE_SEGMENT|7062,7074|false|false|false|C0039644;C1744619|Tetracycline Antibiotics;tetracycline|TETRACYCLINE
Event|Event|SIMPLE_SEGMENT|7062,7074|false|false|false|||TETRACYCLINE
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7093,7103|false|false|false|C0042313|vancomycin|VANCOMYCIN
Drug|Antibiotic|SIMPLE_SEGMENT|7093,7103|false|false|false|C0042313|vancomycin|VANCOMYCIN
Event|Event|SIMPLE_SEGMENT|7093,7103|false|false|false|||VANCOMYCIN
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7093,7103|false|false|false|C0489941|Vancomycin measurement|VANCOMYCIN
Event|Event|SIMPLE_SEGMENT|7125,7132|false|false|false|||IMAGING
Finding|Finding|SIMPLE_SEGMENT|7125,7132|false|false|false|C0740845|Imaging problem|IMAGING
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7125,7132|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|IMAGING
Event|Event|SIMPLE_SEGMENT|7164,7167|false|false|false|||CXR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7164,7167|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|SIMPLE_SEGMENT|7168,7178|false|false|false|||IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|7168,7178|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|7168,7178|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Event|Event|SIMPLE_SEGMENT|7186,7196|false|false|false|||congestion
Finding|Pathologic Function|SIMPLE_SEGMENT|7186,7196|false|false|false|C0700148|Congestion|congestion
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7205,7210|false|false|false|C0398650|Immune thrombocytopenic purpura|frank
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7211,7216|true|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|7211,7216|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|7211,7216|true|false|false|C0013604|Edema|edema
Event|Event|SIMPLE_SEGMENT|7234,7239|false|false|false|||signs
Finding|Finding|SIMPLE_SEGMENT|7234,7239|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|SIMPLE_SEGMENT|7234,7239|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7243,7252|false|false|false|C0032285|Pneumonia|pneumonia
Event|Event|SIMPLE_SEGMENT|7243,7252|false|false|false|||pneumonia
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7259,7262|false|false|false|C3813556|Cancer/Testis Antigen|CTA
Event|Event|SIMPLE_SEGMENT|7259,7262|false|false|false|||CTA
Finding|Gene or Genome|SIMPLE_SEGMENT|7259,7262|false|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7259,7262|false|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7263,7268|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|7263,7268|false|false|false|C0741025|Chest problem|chest
Event|Event|SIMPLE_SEGMENT|7269,7275|false|false|false|||showed
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7290,7299|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7290,7299|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|7290,7299|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|SIMPLE_SEGMENT|7290,7308|false|false|false|C0034065|Pulmonary Embolism|pulmonary embolism
Event|Event|SIMPLE_SEGMENT|7300,7308|false|false|false|||embolism
Finding|Finding|SIMPLE_SEGMENT|7300,7308|false|false|false|C0013922;C1704212|Embolism;Embolus|embolism
Finding|Pathologic Function|SIMPLE_SEGMENT|7300,7308|false|false|false|C0013922;C1704212|Embolism;Embolus|embolism
Event|Event|SIMPLE_SEGMENT|7314,7322|false|false|false|||thrombus
Finding|Pathologic Function|SIMPLE_SEGMENT|7314,7322|false|false|false|C0087086;C0302148|Blood Clot;Thrombus|thrombus
Event|Event|SIMPLE_SEGMENT|7323,7327|false|false|false|||seen
Event|Event|SIMPLE_SEGMENT|7328,7337|false|false|false|||extending
Finding|Functional Concept|SIMPLE_SEGMENT|7348,7353|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7348,7375|false|false|false|C0226054;C0923924|Right pulmonary arterial tree;Right pulmonary artery|right main pulmonary artery
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7359,7368|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7359,7368|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|7359,7368|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7359,7375|false|false|false|C0034052|Pulmonary artery structure|pulmonary artery
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7369,7375|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|SIMPLE_SEGMENT|7369,7375|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Finding|Functional Concept|SIMPLE_SEGMENT|7413,7418|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Event|Event|SIMPLE_SEGMENT|7426,7432|false|false|false|||middle
Finding|Intellectual Product|SIMPLE_SEGMENT|7426,7432|false|false|false|C1552826|Table Cell Vertical Align - middle|middle
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7438,7443|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|7438,7443|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7438,7448|false|false|false|C0225758|Structure of lower lobe of lung|lower lobe
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7444,7448|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|SIMPLE_SEGMENT|7444,7448|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7444,7458|false|false|false|C0225752|Structure of lobe of lung|lobe pulmonary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7449,7458|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7449,7458|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|7449,7458|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7460,7468|false|false|false|C0003842;C0226004|Arterial system;Arteries|arteries
Anatomy|Body System|SIMPLE_SEGMENT|7460,7468|false|false|false|C0003842;C0226004|Arterial system;Arteries|arteries
Event|Event|SIMPLE_SEGMENT|7460,7468|false|false|false|||arteries
Procedure|Health Care Activity|SIMPLE_SEGMENT|7460,7468|false|false|false|C0397581|Procedure on artery|arteries
Finding|Functional Concept|SIMPLE_SEGMENT|7473,7478|true|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7473,7484|false|false|false|C0225808|Right side of heart|right heart
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7479,7484|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7479,7484|true|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|7479,7484|true|false|false|C0795691|HEART PROBLEM|heart
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|7485,7491|true|false|false|C0080194|Muscle strain|strain
Event|Event|SIMPLE_SEGMENT|7485,7491|false|false|false|||strain
Finding|Idea or Concept|SIMPLE_SEGMENT|7485,7491|true|false|false|C0442694;C1510453;C1548152;C2987481|Emotional Strain;Nature of Abnormal Testing - Strain;Straining (finding);strain symptom|strain
Finding|Mental Process|SIMPLE_SEGMENT|7485,7491|true|false|false|C0442694;C1510453;C1548152;C2987481|Emotional Strain;Nature of Abnormal Testing - Strain;Straining (finding);strain symptom|strain
Finding|Physiologic Function|SIMPLE_SEGMENT|7485,7491|true|false|false|C0442694;C1510453;C1548152;C2987481|Emotional Strain;Nature of Abnormal Testing - Strain;Straining (finding);strain symptom|strain
Finding|Sign or Symptom|SIMPLE_SEGMENT|7485,7491|true|false|false|C0442694;C1510453;C1548152;C2987481|Emotional Strain;Nature of Abnormal Testing - Strain;Straining (finding);strain symptom|strain
Event|Event|SIMPLE_SEGMENT|7492,7502|false|false|false|||identified
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7540,7549|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7540,7549|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|7540,7549|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|SIMPLE_SEGMENT|7540,7556|false|false|false|C0034065|Pulmonary Embolism|pulmonary emboli
Event|Event|SIMPLE_SEGMENT|7550,7556|false|false|false|||emboli
Finding|Finding|SIMPLE_SEGMENT|7550,7556|false|false|false|C1704212|Embolus|emboli
Event|Event|SIMPLE_SEGMENT|7557,7561|false|false|false|||seen
Event|Event|SIMPLE_SEGMENT|7597,7605|false|false|false|||branches
Finding|Functional Concept|SIMPLE_SEGMENT|7613,7617|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7628,7633|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|7628,7633|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7634,7639|false|false|false|C0796494|lobe|lobes
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7653,7662|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7653,7662|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|7653,7662|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Finding|SIMPLE_SEGMENT|7653,7670|false|false|false|C0748164|Multiple Pulmonary Nodules|pulmonary nodules
Event|Event|SIMPLE_SEGMENT|7663,7670|false|false|false|||nodules
Event|Event|SIMPLE_SEGMENT|7675,7680|false|false|false|||noted
Event|Event|SIMPLE_SEGMENT|7685,7690|false|false|false|||noted
Event|Event|SIMPLE_SEGMENT|7731,7741|false|false|false|||spiculated
Event|Event|SIMPLE_SEGMENT|7746,7755|false|false|false|||measuring
Finding|Functional Concept|SIMPLE_SEGMENT|7775,7780|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7775,7792|false|false|false|C4281590|Structure of middle lobe of right lung|right middle lobe
Finding|Intellectual Product|SIMPLE_SEGMENT|7781,7787|false|false|false|C1552826|Table Cell Vertical Align - middle|middle
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7781,7792|false|false|false|C4281590|Structure of middle lobe of right lung|middle lobe
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7788,7792|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|SIMPLE_SEGMENT|7788,7792|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Event|Event|SIMPLE_SEGMENT|7794,7804|false|false|false|||suspicious
Finding|Finding|SIMPLE_SEGMENT|7794,7819|false|false|false|C4050405|Suspicious for Malignancy|suspicious for malignancy
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7809,7819|false|true|false|C0006826;C1306459|Malignant Neoplasms;Primary malignant neoplasm|malignancy
Event|Event|SIMPLE_SEGMENT|7809,7819|false|false|false|||malignancy
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7837,7840|false|false|false|C0032743;C0040398|Positron-Emission Tomography;Tomography, Emission-Computed|PET
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7837,7843|false|false|false|C1699633|PET/CT scan|PET-CT
Event|Event|SIMPLE_SEGMENT|7841,7843|false|false|false|||CT
Event|Event|SIMPLE_SEGMENT|7852,7865|false|false|false|||demonstration
Finding|Functional Concept|SIMPLE_SEGMENT|7871,7875|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7871,7882|false|false|false|C0222601|Left breast|left breast
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7876,7882|false|false|false|C0006141|Breast|breast
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7876,7882|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|breast
Finding|Finding|SIMPLE_SEGMENT|7876,7882|false|false|false|C0567499|Breast problem|breast
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7876,7882|false|false|false|C0191838|Procedures on breast|breast
Finding|Finding|SIMPLE_SEGMENT|7876,7890|false|false|false|C0024103|Mass in breast|breast nodules
Event|Event|SIMPLE_SEGMENT|7883,7890|false|false|false|||nodules
Event|Event|SIMPLE_SEGMENT|7902,7913|false|false|false|||correlation
Event|Event|SIMPLE_SEGMENT|7919,7930|false|false|false|||mammography
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7919,7930|false|false|false|C0024671;C0848600|Mammography;Mammography, Female|mammography
Event|Event|SIMPLE_SEGMENT|7935,7945|false|false|false|||ultrasound
Finding|Functional Concept|SIMPLE_SEGMENT|7935,7945|false|false|false|C0220934|Ultrasonic|ultrasound
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|7935,7945|false|false|false|C0041621;C1456803|Ultrasonic Shockwave;Ultrasonics (sound)|ultrasound
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7935,7945|false|false|false|C0041618;C1315081|Ultrasonography;Urological ultrasound|ultrasound
Event|Event|SIMPLE_SEGMENT|7949,7958|false|false|false|||suggested
Event|Event|SIMPLE_SEGMENT|7970,7980|false|false|false|||IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|7970,7980|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|7970,7980|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|7985,7993|false|false|false|C1552654|Parameterized Data Type - Interval|Interval
Event|Event|SIMPLE_SEGMENT|7994,8005|false|false|false|||progression
Finding|Functional Concept|SIMPLE_SEGMENT|7994,8005|false|false|false|C0242656;C0449258|Disease Progression;Progression|progression
Finding|Pathologic Function|SIMPLE_SEGMENT|7994,8005|false|false|false|C0242656;C0449258|Disease Progression;Progression|progression
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8009,8013|false|false|false|C4318566|Deep Resection Margin|deep
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8009,8018|false|false|false|C0226514|Structure of deep vein|deep vein
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8009,8029|false|false|false|C0149871;C0340708|Deep Vein Thrombosis;Deep vein thrombosis of lower limb|deep vein thrombosis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8014,8018|false|false|false|C0042449|Veins|vein
Finding|Pathologic Function|SIMPLE_SEGMENT|8014,8029|false|false|false|C0042487|Venous Thrombosis|vein thrombosis
Event|Event|SIMPLE_SEGMENT|8019,8029|false|false|false|||thrombosis
Finding|Pathologic Function|SIMPLE_SEGMENT|8019,8029|false|false|false|C0040053|Thrombosis|thrombosis
Finding|Functional Concept|SIMPLE_SEGMENT|8037,8041|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|SIMPLE_SEGMENT|8043,8048|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|8043,8048|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8043,8058|false|false|false|C0023216|Lower Extremity|lower extremity
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8049,8058|false|false|false|C0015385|Limb structure|extremity
Finding|Functional Concept|SIMPLE_SEGMENT|8065,8074|false|false|false|C1947917|Occluded|occlusive
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|8065,8083|false|false|false|C0333203|Occlusive thrombus|occlusive thrombus
Event|Event|SIMPLE_SEGMENT|8075,8083|false|false|false|||thrombus
Finding|Pathologic Function|SIMPLE_SEGMENT|8075,8083|false|false|false|C0087086;C0302148|Blood Clot;Thrombus|thrombus
Event|Event|SIMPLE_SEGMENT|8084,8093|false|false|false|||involving
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8106,8113|false|false|false|C0015811|Femur|femoral
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8106,8118|false|false|false|C0015809|Femoral vein|femoral vein
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8114,8118|false|false|false|C0042449|Veins|vein
Event|Event|SIMPLE_SEGMENT|8136,8145|false|false|false|||involving
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8158,8164|false|false|false|C4522154|Distal Resection Margin|distal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8166,8173|false|false|false|C0015811|Femur|femoral
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8166,8178|false|false|false|C0015809|Femoral vein|femoral vein
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8174,8178|false|false|false|C0042449|Veins|vein
Finding|Functional Concept|SIMPLE_SEGMENT|8190,8200|false|false|false|C1524062|Additional|additional
Event|Event|SIMPLE_SEGMENT|8214,8222|false|false|false|||thrombus
Finding|Pathologic Function|SIMPLE_SEGMENT|8214,8222|false|false|false|C0087086;C0302148|Blood Clot;Thrombus|thrombus
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8231,8235|false|false|false|C4318566|Deep Resection Margin|deep
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8231,8248|false|false|false|C0226841|Structure of profunda femoris vein|deep femoral vein
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8236,8243|false|false|false|C0015811|Femur|femoral
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8236,8248|false|false|false|C0015809|Femoral vein|femoral vein
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8244,8248|false|false|false|C0042449|Veins|vein
Finding|Functional Concept|SIMPLE_SEGMENT|8255,8259|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Finding|Functional Concept|SIMPLE_SEGMENT|8260,8266|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Finding|Intellectual Product|SIMPLE_SEGMENT|8260,8266|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8267,8274|false|false|false|C0015811|Femur|femoral
Anatomy|Body Location or Region|SIMPLE_SEGMENT|8279,8288|false|false|false|C0442037|popliteal|popliteal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8279,8294|false|false|false|C0032652|Structure of popliteal vein|popliteal veins
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8289,8294|false|false|false|C0042449|Veins|veins
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8289,8294|false|false|false|C0398102|Procedure on vein|veins
Event|Event|SIMPLE_SEGMENT|8300,8306|false|false|false|||patent
Finding|Intellectual Product|SIMPLE_SEGMENT|8300,8306|false|false|false|C0030650|Legal patent|patent
Anatomy|Body Location or Region|SIMPLE_SEGMENT|8325,8329|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8325,8329|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8330,8335|false|false|false|C0042449|Veins|veins
Event|Event|SIMPLE_SEGMENT|8330,8335|false|false|false|||veins
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8330,8335|true|false|false|C0398102|Procedure on vein|veins
Event|Event|SIMPLE_SEGMENT|8345,8355|false|false|false|||visualized
Event|Event|SIMPLE_SEGMENT|8367,8376|false|false|false|||overlying
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8377,8385|false|false|false|C1705365|Dressing Dosage Form|dressing
Event|Event|SIMPLE_SEGMENT|8377,8385|false|false|false|||dressing
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|8377,8385|false|false|false|C0518459;C1305428|Ability to dress|dressing
Finding|Finding|SIMPLE_SEGMENT|8377,8385|false|false|false|C0518459;C1305428|Ability to dress|dressing
Procedure|Health Care Activity|SIMPLE_SEGMENT|8377,8385|false|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|dressing
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8377,8385|false|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|dressing
Event|Event|SIMPLE_SEGMENT|8400,8408|false|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|8400,8408|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|8400,8411|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8412,8416|true|false|false|C4318566|Deep Resection Margin|deep
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8417,8423|false|false|false|C0042449|Veins|venous
Event|Event|SIMPLE_SEGMENT|8425,8435|false|false|false|||thrombosis
Finding|Pathologic Function|SIMPLE_SEGMENT|8425,8435|false|false|false|C0040053|Thrombosis|thrombosis
Finding|Functional Concept|SIMPLE_SEGMENT|8443,8448|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8443,8464|false|false|false|C0230415|Right lower extremity|right lower extremity
Anatomy|Body Location or Region|SIMPLE_SEGMENT|8449,8454|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|8449,8454|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8449,8464|false|false|false|C0023216|Lower Extremity|lower extremity
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8455,8464|false|false|false|C0015385|Limb structure|extremity
Event|Event|SIMPLE_SEGMENT|8471,8474|false|false|false|||TTE
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8471,8474|false|false|false|C0430462|Transthoracic echocardiography|TTE
Event|Event|SIMPLE_SEGMENT|8476,8487|false|false|false|||Conclusions
Finding|Idea or Concept|SIMPLE_SEGMENT|8476,8487|false|false|false|C1707478|Conclusion|Conclusions
Finding|Functional Concept|SIMPLE_SEGMENT|8492,8496|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8492,8503|false|false|false|C0225860|Left atrial structure|left atrium
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8497,8503|false|false|false|C0018792|Heart Atrium|atrium
Event|Event|SIMPLE_SEGMENT|8507,8513|false|false|false|||normal
Finding|Functional Concept|SIMPLE_SEGMENT|8537,8542|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8543,8549|false|false|false|C0018792|Heart Atrium|atrial
Event|Event|SIMPLE_SEGMENT|8551,8559|false|false|false|||pressure
Finding|Finding|SIMPLE_SEGMENT|8551,8559|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|SIMPLE_SEGMENT|8551,8559|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|8551,8559|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|8551,8559|false|false|false|C0033095||pressure
Finding|Functional Concept|SIMPLE_SEGMENT|8573,8577|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8573,8594|false|false|false|C0504053|Wall of left ventricle|Left ventricular wall
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8578,8589|false|false|false|C0018827|Heart Ventricle|ventricular
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8578,8594|false|false|false|C0507618|Wall of ventricle|ventricular wall
Finding|Finding|SIMPLE_SEGMENT|8578,8604|false|false|false|C2024242|cardiac evaluation of ventricular wall thickness|ventricular wall thickness
Event|Event|SIMPLE_SEGMENT|8595,8604|false|false|false|||thickness
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|8606,8612|false|false|false|C0333343|Body cavities|cavity
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|8606,8612|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8606,8612|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|8631,8639|false|false|false|C0039155|Systole|systolic
Event|Event|SIMPLE_SEGMENT|8640,8648|false|false|false|||function
Finding|Finding|SIMPLE_SEGMENT|8640,8648|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|SIMPLE_SEGMENT|8640,8648|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|SIMPLE_SEGMENT|8640,8648|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|SIMPLE_SEGMENT|8640,8648|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Event|Event|SIMPLE_SEGMENT|8653,8659|false|false|false|||normal
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8661,8665|false|false|false|C0428772|Left ventricular ejection fraction|LVEF
Event|Event|SIMPLE_SEGMENT|8661,8665|false|false|false|||LVEF
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8661,8665|false|false|false|C3837267|LVEF (procedure)|LVEF
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8673,8680|false|false|false|C0554756|Doppler studies|Doppler
Event|Event|SIMPLE_SEGMENT|8681,8691|false|false|false|||parameters
Finding|Finding|SIMPLE_SEGMENT|8681,8691|false|false|false|C0449381|Observation parameter|parameters
Event|Event|SIMPLE_SEGMENT|8701,8711|false|false|false|||consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|8701,8711|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|8701,8716|false|false|false|C0332290|Consistent with|consistent with
Finding|Classification|SIMPLE_SEGMENT|8712,8722|false|false|false|C0441800|Grade|with Grade
Finding|Classification|SIMPLE_SEGMENT|8717,8722|false|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|Grade
Finding|Finding|SIMPLE_SEGMENT|8717,8722|false|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|Grade
Finding|Finding|SIMPLE_SEGMENT|8717,8724|false|false|false|C0475269;C0687695;C4049998|Clavien-Dindo Grade I;Grade 1 (qualifier value);Tumor grade G1|Grade I
Finding|Intellectual Product|SIMPLE_SEGMENT|8717,8724|false|false|false|C0475269;C0687695;C4049998|Clavien-Dindo Grade I;Grade 1 (qualifier value);Tumor grade G1|Grade I
Finding|Intellectual Product|SIMPLE_SEGMENT|8726,8730|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Functional Concept|SIMPLE_SEGMENT|8732,8736|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8738,8749|false|false|false|C0018827|Heart Ventricle|ventricular
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8750,8759|false|false|false|C0012000|Diastole|diastolic
Finding|Pathologic Function|SIMPLE_SEGMENT|8750,8771|false|false|false|C0520863|Diastolic dysfunction|diastolic dysfunction
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8760,8771|false|false|false|C3887505|DYSFUNCTION - SKIN DISORDERS|dysfunction
Event|Event|SIMPLE_SEGMENT|8760,8771|false|false|false|||dysfunction
Finding|Conceptual Entity|SIMPLE_SEGMENT|8760,8771|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Functional Concept|SIMPLE_SEGMENT|8760,8771|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Pathologic Function|SIMPLE_SEGMENT|8760,8771|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Functional Concept|SIMPLE_SEGMENT|8773,8778|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8779,8790|false|false|false|C0018827|Heart Ventricle|ventricular
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8791,8798|false|false|false|C0935616|chamber [body part]|chamber
Event|Event|SIMPLE_SEGMENT|8809,8813|false|false|false|||free
Finding|Functional Concept|SIMPLE_SEGMENT|8809,8813|false|false|false|C0332296|Free of (attribute)|free
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8814,8825|false|false|false|C1980023|Wall motion|wall motion
Event|Event|SIMPLE_SEGMENT|8819,8825|false|false|false|||motion
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|8819,8825|false|false|false|C0026597|Motion|motion
Event|Event|SIMPLE_SEGMENT|8830,8836|false|false|false|||normal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8842,8848|false|false|false|C0003483|Aorta|aortic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8842,8854|false|false|false|C0003501;C4533215|Aortic valve structure;Chest>Aortic valve|aortic valve
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8849,8854|false|false|false|C1186983|Anatomical valve|valve
Event|Event|SIMPLE_SEGMENT|8876,8885|false|false|false|||thickened
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8904,8910|false|false|false|C0003483|Aorta|aortic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8904,8916|false|false|false|C0003501;C4533215|Aortic valve structure;Chest>Aortic valve|aortic valve
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|8904,8925|true|false|false|C5193127;C5700069|AORTIC VALVE DISEASE 3;Stenosis of aorta|aortic valve stenosis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8904,8925|true|false|false|C5193127;C5700069|AORTIC VALVE DISEASE 3;Stenosis of aorta|aortic valve stenosis
Finding|Pathologic Function|SIMPLE_SEGMENT|8904,8925|true|false|false|C0003507|Aortic Valve Stenosis|aortic valve stenosis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8911,8916|false|false|false|C1186983|Anatomical valve|valve
Event|Event|SIMPLE_SEGMENT|8917,8925|false|false|false|||stenosis
Finding|Pathologic Function|SIMPLE_SEGMENT|8917,8925|true|false|false|C1261287|Stenosis|stenosis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8936,8956|false|false|false|C0026266|Mitral Valve Insufficiency|mitral regurgitation
Event|Event|SIMPLE_SEGMENT|8943,8956|false|false|false|||regurgitation
Finding|Finding|SIMPLE_SEGMENT|8943,8956|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|SIMPLE_SEGMENT|8943,8956|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|SIMPLE_SEGMENT|8943,8956|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Event|Event|SIMPLE_SEGMENT|8960,8964|false|false|false|||seen
Finding|Intellectual Product|SIMPLE_SEGMENT|8975,8979|false|false|false|C1547225|Mild Severity of Illness Code|mild
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8980,8989|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8980,8989|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|8980,8989|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8991,8997|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|SIMPLE_SEGMENT|8991,8997|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|8998,9006|false|false|false|C0039155|Systole|systolic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8998,9019|false|false|false|C0221155|Systolic Hypertension|systolic hypertension
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9007,9019|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|SIMPLE_SEGMENT|9007,9019|false|false|false|||hypertension
Event|Event|SIMPLE_SEGMENT|9027,9030|false|false|false|||CXR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|9027,9030|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|SIMPLE_SEGMENT|9031,9041|false|false|false|||IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|9031,9041|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|9031,9041|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Event|Event|SIMPLE_SEGMENT|9044,9052|false|false|false|||Compared
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9056,9061|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|9056,9061|false|false|false|C0741025|Chest problem|chest
Event|Event|SIMPLE_SEGMENT|9062,9073|false|false|false|||radiographs
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|9062,9073|false|false|false|C1306645|Plain x-ray|radiographs
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9092,9097|false|false|false|C0018787;C4037974|Chest>Heart;Heart|Heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|9092,9097|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|Heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|9092,9097|false|false|false|C0795691|HEART PROBLEM|Heart
Finding|Finding|SIMPLE_SEGMENT|9092,9102|false|false|false|C0744689|heart size|Heart size
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9116,9121|false|false|false|C0024109|Lung|Lungs
Event|Event|SIMPLE_SEGMENT|9130,9135|false|false|false|||clear
Finding|Idea or Concept|SIMPLE_SEGMENT|9130,9135|false|false|false|C1550016|Remote control command - Clear|clear
Anatomy|Tissue|SIMPLE_SEGMENT|9141,9148|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9141,9148|true|false|false|C0032226|Pleural Diseases|pleural
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|9150,9161|false|false|false|C0000768|Congenital Abnormality|abnormality
Event|Event|SIMPLE_SEGMENT|9150,9161|false|false|false|||abnormality
Finding|Finding|SIMPLE_SEGMENT|9150,9161|false|false|false|C1704258|Abnormality|abnormality
Event|Event|SIMPLE_SEGMENT|9165,9173|false|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|9165,9173|false|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|9165,9176|false|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9177,9184|false|false|false|C0719205|Central brand of multivitamin with minerals|central
Drug|Vitamin|SIMPLE_SEGMENT|9177,9184|false|false|false|C0719205|Central brand of multivitamin with minerals|central
Event|Event|SIMPLE_SEGMENT|9177,9184|false|false|false|||central
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9177,9184|false|false|false|C1879652|Central Minus|central
Finding|Body Substance|SIMPLE_SEGMENT|9177,9190|false|false|false|C1179479|Central lymph|central lymph
Finding|Body Substance|SIMPLE_SEGMENT|9185,9190|false|false|false|C0024202|Lymph|lymph
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9185,9195|false|false|false|C0024204|lymph nodes|lymph node
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9185,9207|false|false|false|C0497156|Lymphadenopathy|lymph node enlargement
Finding|Sign or Symptom|SIMPLE_SEGMENT|9185,9207|false|false|false|C4282165|Swollen Lymph Node|lymph node enlargement
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|9196,9207|false|false|false|C2711450|Enlargement (morphologic abnormality)|enlargement
Event|Event|SIMPLE_SEGMENT|9196,9207|false|false|false|||enlargement
Finding|Pathologic Function|SIMPLE_SEGMENT|9196,9207|false|false|false|C0020564|Hypertrophy|enlargement
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9196,9207|false|false|false|C1293134|Enlargement procedure|enlargement
Finding|Intellectual Product|SIMPLE_SEGMENT|9212,9217|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|Brief
Finding|Idea or Concept|SIMPLE_SEGMENT|9218,9226|false|false|false|C1547192|Organization unit type - Hospital|Hospital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9218,9233|false|false|false|C0488549||Hospital Course
Finding|Finding|SIMPLE_SEGMENT|9218,9233|false|false|false|C0489547|Hospital course|Hospital Course
Drug|Chemical Viewed Structurally|SIMPLE_SEGMENT|9270,9277|false|false|false|C0302912|Radicals (chemistry)|radical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9270,9288|false|false|false|C0194401|Complete cystectomy|radical cystectomy
Event|Event|SIMPLE_SEGMENT|9278,9288|false|false|false|||cystectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9278,9288|false|false|false|C0010651|Cystectomy|cystectomy
Event|Event|SIMPLE_SEGMENT|9293,9303|false|false|false|||omplicated
Finding|Finding|SIMPLE_SEGMENT|9307,9317|false|false|false|C0004610|Bacteremia|bacteremia
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9323,9330|false|false|false|C0000833|Abscess|abscess
Event|Event|SIMPLE_SEGMENT|9323,9330|false|false|false|||abscess
Finding|Intellectual Product|SIMPLE_SEGMENT|9323,9330|false|false|false|C1546533||abscess
Event|Event|SIMPLE_SEGMENT|9332,9335|false|false|false|||LLE
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9336,9339|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9336,9339|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9336,9339|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Event|Event|SIMPLE_SEGMENT|9336,9339|false|false|false|||DVT
Drug|Organic Chemical|SIMPLE_SEGMENT|9360,9367|false|false|false|C0728963|Lovenox|lovenox
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9360,9367|false|false|false|C0728963|Lovenox|lovenox
Event|Event|SIMPLE_SEGMENT|9360,9367|false|false|false|||lovenox
Event|Event|SIMPLE_SEGMENT|9372,9380|false|false|false|||presents
Event|Event|SIMPLE_SEGMENT|9387,9394|false|false|false|||dyspnea
Finding|Finding|SIMPLE_SEGMENT|9387,9394|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|9387,9394|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|9387,9406|false|false|false|C0231807|Dyspnea on exertion|dyspnea on exertion
Event|Event|SIMPLE_SEGMENT|9398,9406|false|false|false|||exertion
Finding|Organism Function|SIMPLE_SEGMENT|9398,9406|false|false|false|C0015264|Exertion|exertion
Event|Event|SIMPLE_SEGMENT|9411,9418|false|false|false|||dyspnea
Finding|Finding|SIMPLE_SEGMENT|9411,9418|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|9411,9418|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|9411,9430|false|false|false|C0231807|Dyspnea on exertion|dyspnea on exertion
Event|Event|SIMPLE_SEGMENT|9422,9430|false|false|false|||exertion
Finding|Organism Function|SIMPLE_SEGMENT|9422,9430|false|false|false|C0015264|Exertion|exertion
Event|Event|SIMPLE_SEGMENT|9435,9440|false|false|false|||found
Finding|Gene or Genome|SIMPLE_SEGMENT|9450,9455|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Event|Event|SIMPLE_SEGMENT|9463,9474|false|false|false|||progression
Finding|Functional Concept|SIMPLE_SEGMENT|9463,9474|false|false|false|C0242656;C0449258|Disease Progression;Progression|progression
Finding|Pathologic Function|SIMPLE_SEGMENT|9463,9474|false|false|false|C0242656;C0449258|Disease Progression;Progression|progression
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9478,9481|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9478,9481|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9478,9481|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Event|Event|SIMPLE_SEGMENT|9478,9481|false|false|false|||DVT
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9489,9492|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9489,9492|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9489,9492|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Finding|Finding|SIMPLE_SEGMENT|9494,9500|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Finding|Idea or Concept|SIMPLE_SEGMENT|9494,9500|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Event|Event|SIMPLE_SEGMENT|9501,9504|false|false|false|||due
Finding|Functional Concept|SIMPLE_SEGMENT|9501,9504|false|true|false|C0678226;C3146286|Due;Due to|due
Finding|Idea or Concept|SIMPLE_SEGMENT|9501,9504|false|true|false|C0678226;C3146286|Due;Due to|due
Finding|Functional Concept|SIMPLE_SEGMENT|9501,9507|false|true|false|C0678226|Due to|due to
Event|Event|SIMPLE_SEGMENT|9508,9522|false|false|false|||undertreatment
Procedure|Health Care Activity|SIMPLE_SEGMENT|9508,9522|false|true|false|C5828474|Undertreatment|undertreatment
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9536,9539|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9536,9539|false|true|false|C2926618||DVT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9536,9539|false|true|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Event|Event|SIMPLE_SEGMENT|9536,9539|false|false|false|||DVT
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9546,9558|false|false|false|C0355642|Drugs used in migraine prophylaxis|prophylactic
Event|Event|SIMPLE_SEGMENT|9546,9558|false|false|false|||prophylactic
Finding|Functional Concept|SIMPLE_SEGMENT|9546,9558|false|false|false|C0445202|Prophylactic behavior|prophylactic
Event|Event|SIMPLE_SEGMENT|9559,9565|false|false|false|||dosing
Drug|Organic Chemical|SIMPLE_SEGMENT|9569,9576|false|false|false|C0728963|Lovenox|lovenox
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9569,9576|false|false|false|C0728963|Lovenox|lovenox
Event|Event|SIMPLE_SEGMENT|9569,9576|false|false|false|||lovenox
Event|Event|SIMPLE_SEGMENT|9584,9595|false|false|false|||underdosing
Drug|Organic Chemical|SIMPLE_SEGMENT|9599,9606|false|false|false|C0728963|Lovenox|lovenox
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9599,9606|false|false|false|C0728963|Lovenox|lovenox
Event|Event|SIMPLE_SEGMENT|9599,9606|false|false|false|||lovenox
Event|Event|SIMPLE_SEGMENT|9622,9629|false|false|false|||thought
Event|Event|SIMPLE_SEGMENT|9636,9645|false|false|false|||treatment
Finding|Conceptual Entity|SIMPLE_SEGMENT|9636,9645|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|SIMPLE_SEGMENT|9636,9645|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|SIMPLE_SEGMENT|9636,9645|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9636,9645|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Finding|Finding|SIMPLE_SEGMENT|9636,9653|false|false|false|C0162643;C0438286;C1547544|Absent response to treatment;Charge Type Reason - Treatment Failure;treatment failure|treatment failure
Finding|Idea or Concept|SIMPLE_SEGMENT|9636,9653|false|false|false|C0162643;C0438286;C1547544|Absent response to treatment;Charge Type Reason - Treatment Failure;treatment failure|treatment failure
Event|Event|SIMPLE_SEGMENT|9646,9653|false|false|false|||failure
Finding|Functional Concept|SIMPLE_SEGMENT|9646,9653|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|SIMPLE_SEGMENT|9646,9653|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|SIMPLE_SEGMENT|9646,9653|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9658,9661|false|false|false|C3498924|lamina IVC|IVC
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|9658,9661|false|false|false|C4085887|Inspiratory Vital Capacity Test|IVC
Event|Event|SIMPLE_SEGMENT|9662,9668|false|false|false|||filter
Finding|Body Substance|SIMPLE_SEGMENT|9662,9668|false|false|false|C1522664;C1546637;C1550638;C1704449|Filter (function);Specimen Type - Filter;filter information process|filter
Finding|Conceptual Entity|SIMPLE_SEGMENT|9662,9668|false|false|false|C1522664;C1546637;C1550638;C1704449|Filter (function);Specimen Type - Filter;filter information process|filter
Finding|Intellectual Product|SIMPLE_SEGMENT|9662,9668|false|false|false|C1522664;C1546637;C1550638;C1704449|Filter (function);Specimen Type - Filter;filter information process|filter
Event|Event|SIMPLE_SEGMENT|9674,9682|false|false|false|||deferred
Event|Event|SIMPLE_SEGMENT|9695,9700|false|false|false|||signs
Finding|Finding|SIMPLE_SEGMENT|9695,9700|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|SIMPLE_SEGMENT|9695,9700|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|SIMPLE_SEGMENT|9704,9709|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9704,9715|false|false|false|C0225808|Right side of heart|right heart
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9710,9715|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|9710,9715|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|9710,9715|false|false|false|C0795691|HEART PROBLEM|heart
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|9716,9722|true|false|false|C0080194|Muscle strain|strain
Event|Event|SIMPLE_SEGMENT|9716,9722|false|false|false|||strain
Finding|Idea or Concept|SIMPLE_SEGMENT|9716,9722|true|false|false|C0442694;C1510453;C1548152;C2987481|Emotional Strain;Nature of Abnormal Testing - Strain;Straining (finding);strain symptom|strain
Finding|Mental Process|SIMPLE_SEGMENT|9716,9722|true|false|false|C0442694;C1510453;C1548152;C2987481|Emotional Strain;Nature of Abnormal Testing - Strain;Straining (finding);strain symptom|strain
Finding|Physiologic Function|SIMPLE_SEGMENT|9716,9722|true|false|false|C0442694;C1510453;C1548152;C2987481|Emotional Strain;Nature of Abnormal Testing - Strain;Straining (finding);strain symptom|strain
Finding|Sign or Symptom|SIMPLE_SEGMENT|9716,9722|true|false|false|C0442694;C1510453;C1548152;C2987481|Emotional Strain;Nature of Abnormal Testing - Strain;Straining (finding);strain symptom|strain
Event|Event|SIMPLE_SEGMENT|9726,9733|false|false|false|||imaging
Finding|Finding|SIMPLE_SEGMENT|9726,9733|false|false|false|C0740845|Imaging problem|imaging
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|9726,9733|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|imaging
Event|Event|SIMPLE_SEGMENT|9736,9739|false|false|false|||EKG
Finding|Intellectual Product|SIMPLE_SEGMENT|9736,9739|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|9736,9739|false|false|false|C1623258|Electrocardiography|EKG
Event|Event|SIMPLE_SEGMENT|9741,9745|false|false|false|||exam
Finding|Functional Concept|SIMPLE_SEGMENT|9741,9745|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|9741,9745|false|false|false|C0582103|Medical Examination|exam
Event|Event|SIMPLE_SEGMENT|9747,9750|false|false|false|||TTE
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|9747,9750|false|false|false|C0430462|Transthoracic echocardiography|TTE
Event|Event|SIMPLE_SEGMENT|9751,9757|false|false|false|||showed
Event|Event|SIMPLE_SEGMENT|9761,9769|false|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|9761,9769|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|9761,9772|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Finding|Functional Concept|SIMPLE_SEGMENT|9773,9778|true|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9773,9784|false|false|false|C0225808|Right side of heart|right heart
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9779,9784|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|9779,9784|true|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|9779,9784|true|false|false|C0795691|HEART PROBLEM|heart
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|9785,9791|true|false|false|C0080194|Muscle strain|strain
Event|Event|SIMPLE_SEGMENT|9785,9791|false|false|false|||strain
Finding|Idea or Concept|SIMPLE_SEGMENT|9785,9791|true|false|false|C0442694;C1510453;C1548152;C2987481|Emotional Strain;Nature of Abnormal Testing - Strain;Straining (finding);strain symptom|strain
Finding|Mental Process|SIMPLE_SEGMENT|9785,9791|true|false|false|C0442694;C1510453;C1548152;C2987481|Emotional Strain;Nature of Abnormal Testing - Strain;Straining (finding);strain symptom|strain
Finding|Physiologic Function|SIMPLE_SEGMENT|9785,9791|true|false|false|C0442694;C1510453;C1548152;C2987481|Emotional Strain;Nature of Abnormal Testing - Strain;Straining (finding);strain symptom|strain
Finding|Sign or Symptom|SIMPLE_SEGMENT|9785,9791|true|false|false|C0442694;C1510453;C1548152;C2987481|Emotional Strain;Nature of Abnormal Testing - Strain;Straining (finding);strain symptom|strain
Event|Event|SIMPLE_SEGMENT|9802,9809|false|false|false|||treated
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9817,9824|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Organic Chemical|SIMPLE_SEGMENT|9817,9824|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9817,9824|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Event|Event|SIMPLE_SEGMENT|9817,9824|false|false|false|||heparin
Disorder|Neoplastic Process|SIMPLE_SEGMENT|9825,9828|false|false|false|C1135868|Gestational Trophoblastic Neoplasms|gtt
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9825,9828|false|false|false|C0991568|Drops - Drug Form|gtt
Event|Event|SIMPLE_SEGMENT|9825,9828|false|false|false|||gtt
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9825,9828|false|false|false|C0017741|Glucose tolerance test|gtt
Finding|Intellectual Product|SIMPLE_SEGMENT|9830,9834|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|SIMPLE_SEGMENT|9835,9847|false|false|false|||transitioned
Event|Event|SIMPLE_SEGMENT|9851,9860|false|false|false|||treatment
Finding|Conceptual Entity|SIMPLE_SEGMENT|9851,9860|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|SIMPLE_SEGMENT|9851,9860|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|SIMPLE_SEGMENT|9851,9860|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9851,9860|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Event|Event|SIMPLE_SEGMENT|9861,9865|false|false|false|||dose
Drug|Organic Chemical|SIMPLE_SEGMENT|9867,9874|false|false|false|C0728963|Lovenox|lovenox
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9867,9874|false|false|false|C0728963|Lovenox|lovenox
Disorder|Neoplastic Process|SIMPLE_SEGMENT|9881,9891|false|false|false|C0006826;C1306459|Malignant Neoplasms;Primary malignant neoplasm|malignancy
Event|Event|SIMPLE_SEGMENT|9881,9891|false|false|false|||malignancy
Event|Event|SIMPLE_SEGMENT|9903,9913|false|false|false|||thrombosis
Finding|Pathologic Function|SIMPLE_SEGMENT|9903,9913|false|false|false|C0040053|Thrombosis|thrombosis
Event|Event|SIMPLE_SEGMENT|9917,9922|false|false|false|||noted
Drug|Organic Chemical|SIMPLE_SEGMENT|9926,9930|false|false|false|C0009074|clotrimazole|CLOT
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9926,9930|false|false|false|C0009074|clotrimazole|CLOT
Event|Event|SIMPLE_SEGMENT|9926,9930|false|false|false|||CLOT
Finding|Pathologic Function|SIMPLE_SEGMENT|9926,9930|false|false|false|C0302148|Blood Clot|CLOT
Event|Event|SIMPLE_SEGMENT|9932,9937|false|false|false|||trial
Procedure|Research Activity|SIMPLE_SEGMENT|9932,9937|false|false|false|C0008976|Clinical Trials|trial
Event|Event|SIMPLE_SEGMENT|9952,9963|false|false|false|||symptomatic
Finding|Functional Concept|SIMPLE_SEGMENT|9952,9963|false|false|false|C0231220|Symptomatic|symptomatic
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9977,9983|false|false|false|C0030054|oxygen|oxygen
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|9977,9983|false|false|false|C0030054|oxygen|oxygen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9977,9983|false|false|false|C0030054|oxygen|oxygen
Event|Event|SIMPLE_SEGMENT|9977,9983|false|false|false|||oxygen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9977,9983|false|false|false|C0184633|Oxygen Therapy Care|oxygen
Event|Event|SIMPLE_SEGMENT|9985,10000|false|false|false|||supplementation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9985,10000|false|false|false|C0242297|Dietary Supplementation|supplementation
Event|Event|SIMPLE_SEGMENT|10009,10017|false|false|false|||improved
Event|Event|SIMPLE_SEGMENT|10025,10040|false|false|false|||hospitalization
Procedure|Health Care Activity|SIMPLE_SEGMENT|10025,10040|false|false|false|C0019993|Hospitalization|hospitalization
Drug|Biologically Active Substance|SIMPLE_SEGMENT|10055,10061|false|false|false|C0030054|oxygen|oxygen
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|10055,10061|false|false|false|C0030054|oxygen|oxygen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10055,10061|false|false|false|C0030054|oxygen|oxygen
Event|Event|SIMPLE_SEGMENT|10055,10061|false|false|false|||oxygen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10055,10061|false|false|false|C0184633|Oxygen Therapy Care|oxygen
Event|Event|SIMPLE_SEGMENT|10065,10074|false|false|false|||tolerated
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10079,10088|false|false|false|C0024109|Lung|Pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10079,10088|false|false|false|C2707265||Pulmonary
Finding|Finding|SIMPLE_SEGMENT|10079,10088|false|false|false|C4522268|Pulmonary (intended site)|Pulmonary
Finding|Finding|SIMPLE_SEGMENT|10079,10096|false|false|false|C0748164|Multiple Pulmonary Nodules|Pulmonary nodules
Event|Event|SIMPLE_SEGMENT|10089,10096|false|false|false|||nodules
Event|Event|SIMPLE_SEGMENT|10115,10121|false|false|false|||masses
Event|Event|SIMPLE_SEGMENT|10132,10137|false|false|false|||noted
Event|Event|SIMPLE_SEGMENT|10142,10144|false|false|false|||CT
Anatomy|Body Location or Region|SIMPLE_SEGMENT|10176,10180|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10176,10180|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10176,10180|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|SIMPLE_SEGMENT|10176,10180|false|false|false|C0740941|Lung Problem|lung
Disorder|Neoplastic Process|SIMPLE_SEGMENT|10176,10191|false|true|false|C0242379|Malignant neoplasm of lung|lung malignancy
Disorder|Neoplastic Process|SIMPLE_SEGMENT|10181,10191|false|true|false|C0006826;C1306459|Malignant Neoplasms;Primary malignant neoplasm|malignancy
Event|Event|SIMPLE_SEGMENT|10181,10191|false|false|false|||malignancy
Event|Event|SIMPLE_SEGMENT|10195,10199|false|false|false|||mets
Finding|Gene or Genome|SIMPLE_SEGMENT|10195,10199|false|false|false|C0812270;C1705694|ETV3 gene;ETV3 wt Allele|mets
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|10202,10209|false|false|false|C1705970|Electrical Current|Current
Event|Event|SIMPLE_SEGMENT|10210,10212|false|false|false|||CT
Event|Event|SIMPLE_SEGMENT|10213,10219|false|false|false|||showed
Finding|Intellectual Product|SIMPLE_SEGMENT|10220,10226|false|false|false|C1547311|Patient Condition Code - Stable|stable
Event|Event|SIMPLE_SEGMENT|10227,10234|false|false|false|||nodules
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10235,10240|false|false|false|C1410088|Still|still
Disorder|Neoplastic Process|SIMPLE_SEGMENT|10257,10267|false|false|false|C0006826;C1306459|Malignant Neoplasms;Primary malignant neoplasm|malignancy
Event|Event|SIMPLE_SEGMENT|10257,10267|false|false|false|||malignancy
Event|Event|SIMPLE_SEGMENT|10277,10286|false|false|false|||evaluated
Anatomy|Body Location or Region|SIMPLE_SEGMENT|10294,10302|false|false|false|C0817096|Chest|thoracic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10294,10302|false|false|false|C5779551|Dissecting Thoracic Aortic Aneurysm|thoracic
Event|Event|SIMPLE_SEGMENT|10313,10324|false|false|false|||recommended
Event|Event|SIMPLE_SEGMENT|10328,10334|false|false|false|||biopsy
Finding|Finding|SIMPLE_SEGMENT|10328,10334|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Finding|Intellectual Product|SIMPLE_SEGMENT|10328,10334|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10328,10334|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Procedure|Health Care Activity|SIMPLE_SEGMENT|10328,10334|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Event|Event|SIMPLE_SEGMENT|10339,10351|false|false|false|||surveillance
Event|Occupational Activity|SIMPLE_SEGMENT|10339,10351|false|false|false|C0684245|legal surveillance|surveillance
Finding|Functional Concept|SIMPLE_SEGMENT|10339,10351|false|false|false|C0220920|surveillance aspects|surveillance
Procedure|Health Care Activity|SIMPLE_SEGMENT|10339,10351|false|false|false|C0733511|Medical Surveillance|surveillance
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|10363,10370|false|false|false|C1705970|Electrical Current|current
Anatomy|Body Location or Region|SIMPLE_SEGMENT|10375,10378|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10375,10378|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10375,10378|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Finding|Classification|SIMPLE_SEGMENT|10384,10390|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|10384,10390|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|10384,10390|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|10384,10390|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Body Substance|SIMPLE_SEGMENT|10399,10406|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|10399,10406|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|10399,10406|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|10407,10414|false|false|false|||decided
Event|Event|SIMPLE_SEGMENT|10419,10431|false|false|false|||surveillance
Event|Occupational Activity|SIMPLE_SEGMENT|10419,10431|false|false|false|C0684245|legal surveillance|surveillance
Finding|Functional Concept|SIMPLE_SEGMENT|10419,10431|false|false|false|C0220920|surveillance aspects|surveillance
Procedure|Health Care Activity|SIMPLE_SEGMENT|10419,10431|false|false|false|C0733511|Medical Surveillance|surveillance
Finding|Finding|SIMPLE_SEGMENT|10441,10445|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|10441,10445|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|10441,10445|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|SIMPLE_SEGMENT|10457,10463|false|false|false|||follow
Finding|Intellectual Product|SIMPLE_SEGMENT|10476,10488|false|false|false|C1547426|Location Service Code - Primary Care|primary care
Procedure|Health Care Activity|SIMPLE_SEGMENT|10476,10488|false|false|false|C0033137|Primary Health Care|primary care
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10476,10497|false|false|false|C2735025||primary care provider
Finding|Idea or Concept|SIMPLE_SEGMENT|10476,10497|false|false|false|C1547431|Primary Care Provider - Provider role|primary care provider
Event|Activity|SIMPLE_SEGMENT|10484,10488|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|10484,10488|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|10484,10488|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|10484,10488|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Functional Concept|SIMPLE_SEGMENT|10489,10497|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|provider
Finding|Intellectual Product|SIMPLE_SEGMENT|10489,10497|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|provider
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10516,10519|false|false|false|C0042029|Urinary tract infection|UTI
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10516,10519|false|false|false|C0077906|urinastatin|UTI
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10516,10519|false|false|false|C0077906|urinastatin|UTI
Event|Event|SIMPLE_SEGMENT|10516,10519|false|false|false|||UTI
Finding|Gene or Genome|SIMPLE_SEGMENT|10516,10519|false|false|false|C1412376;C5780748|AMBP gene;AMBP wt Allele|UTI
Event|Event|SIMPLE_SEGMENT|10528,10533|false|false|false|||noted
Anatomy|Cell|SIMPLE_SEGMENT|10549,10552|false|false|false|C0023516|Leukocytes|WBC
Event|Event|SIMPLE_SEGMENT|10549,10552|false|false|false|||WBC
Finding|Mental Process|SIMPLE_SEGMENT|10560,10567|false|false|false|C0542559|contextual factors|setting
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|10581,10589|false|false|false|C0559495|Urological stoma|urostomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10581,10589|false|false|false|C0856443|Urostomy procedure|urostomy
Event|Event|SIMPLE_SEGMENT|10590,10597|false|false|false|||growing
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10629,10641|false|false|false|C0023518|Leukocytosis|leukocytosis
Event|Event|SIMPLE_SEGMENT|10629,10641|false|false|false|||leukocytosis
Finding|Finding|SIMPLE_SEGMENT|10629,10641|false|false|false|C0750426|Blood leukocyte number above reference range|leukocytosis
Event|Event|SIMPLE_SEGMENT|10647,10656|false|false|false|||proceeded
Event|Event|SIMPLE_SEGMENT|10662,10671|false|false|false|||treatment
Finding|Conceptual Entity|SIMPLE_SEGMENT|10662,10671|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|SIMPLE_SEGMENT|10662,10671|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|SIMPLE_SEGMENT|10662,10671|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10662,10671|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Event|Event|SIMPLE_SEGMENT|10681,10688|false|false|false|||started
Finding|Finding|SIMPLE_SEGMENT|10689,10694|false|false|false|C3714655|On IV|on IV
Drug|Antibiotic|SIMPLE_SEGMENT|10695,10705|false|false|false|C0002680;C2095775|ampicillin;ampicillins|Ampicillin
Drug|Organic Chemical|SIMPLE_SEGMENT|10695,10705|false|false|false|C0002680;C2095775|ampicillin;ampicillins|Ampicillin
Event|Event|SIMPLE_SEGMENT|10695,10705|false|false|false|||Ampicillin
Event|Event|SIMPLE_SEGMENT|10711,10723|false|false|false|||transitioned
Drug|Organic Chemical|SIMPLE_SEGMENT|10727,10735|false|false|false|C0591750|Macrobid|macrobid
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10727,10735|false|false|false|C0591750|Macrobid|macrobid
Event|Event|SIMPLE_SEGMENT|10746,10757|false|false|false|||sensitivies
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10759,10771|false|false|false|C0023518|Leukocytosis|Leukocytosis
Event|Event|SIMPLE_SEGMENT|10759,10771|false|false|false|||Leukocytosis
Finding|Finding|SIMPLE_SEGMENT|10759,10771|false|false|false|C0750426|Blood leukocyte number above reference range|Leukocytosis
Event|Event|SIMPLE_SEGMENT|10773,10781|false|false|false|||improved
Drug|Antibiotic|SIMPLE_SEGMENT|10785,10796|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|SIMPLE_SEGMENT|10785,10796|false|false|false|||antibiotics
Event|Event|SIMPLE_SEGMENT|10809,10817|false|false|false|||complete
Finding|Idea or Concept|SIMPLE_SEGMENT|10822,10825|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|10822,10825|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|10826,10832|false|false|false|||course
Finding|Idea or Concept|SIMPLE_SEGMENT|10834,10837|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|10834,10837|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Idea or Concept|SIMPLE_SEGMENT|10847,10850|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|10847,10850|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Finding|SIMPLE_SEGMENT|10847,10852|false|false|false|C3842672|Day 7|day 7
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10874,10880|false|false|false|C0002871|Anemia|Anemia
Event|Event|SIMPLE_SEGMENT|10874,10880|false|false|false|||Anemia
Event|Event|SIMPLE_SEGMENT|10885,10890|false|false|false|||signs
Finding|Finding|SIMPLE_SEGMENT|10885,10890|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|SIMPLE_SEGMENT|10885,10890|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Event|Event|SIMPLE_SEGMENT|10894,10902|false|false|false|||bleeding
Finding|Pathologic Function|SIMPLE_SEGMENT|10894,10902|true|false|false|C0019080|Hemorrhage|bleeding
Event|Event|SIMPLE_SEGMENT|10907,10916|false|false|false|||hemolysis
Finding|Cell Function|SIMPLE_SEGMENT|10907,10916|true|false|false|C0019054;C1553188;C2937287;C2945560|Hemolysis (biological function);Hemolysis (disorder);Hemolysis (finding)|hemolysis
Finding|Finding|SIMPLE_SEGMENT|10907,10916|true|false|false|C0019054;C1553188;C2937287;C2945560|Hemolysis (biological function);Hemolysis (disorder);Hemolysis (finding)|hemolysis
Finding|Pathologic Function|SIMPLE_SEGMENT|10907,10916|true|false|false|C0019054;C1553188;C2937287;C2945560|Hemolysis (biological function);Hemolysis (disorder);Hemolysis (finding)|hemolysis
Event|Event|SIMPLE_SEGMENT|10922,10929|false|false|false|||dropped
Event|Event|SIMPLE_SEGMENT|10933,10938|false|false|false|||nadir
Event|Event|SIMPLE_SEGMENT|10947,10953|false|false|false|||stable
Finding|Intellectual Product|SIMPLE_SEGMENT|10947,10953|false|false|false|C1547311|Patient Condition Code - Stable|stable
Event|Event|SIMPLE_SEGMENT|10957,10966|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|10957,10966|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|10957,10966|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|10957,10966|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|10957,10966|false|false|false|C0030685|Patient Discharge|discharge
Drug|Biologically Active Substance|SIMPLE_SEGMENT|10975,10979|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|10975,10979|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10975,10979|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Event|Event|SIMPLE_SEGMENT|10975,10979|false|false|false|||Iron
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10975,10979|false|false|false|C0337439|Iron measurement|Iron
Event|Event|SIMPLE_SEGMENT|10981,10988|false|false|false|||studies
Procedure|Research Activity|SIMPLE_SEGMENT|10981,10988|false|false|false|C0947630|Scientific Study|studies
Event|Event|SIMPLE_SEGMENT|10989,10999|false|false|false|||consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|10989,10999|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|10989,11004|false|false|false|C0332290|Consistent with|consistent with
Finding|Finding|SIMPLE_SEGMENT|11005,11011|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|11005,11011|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Finding|SIMPLE_SEGMENT|11012,11023|false|true|false|C3811910|combination - answer to question|combination
Drug|Biologically Active Substance|SIMPLE_SEGMENT|11024,11028|false|true|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|11024,11028|false|true|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11024,11028|false|true|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|11024,11028|false|true|false|C0337439|Iron measurement|iron
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11024,11039|false|true|false|C0162316;C0240066|Iron deficiency;Iron deficiency anemia|iron deficiency
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11029,11039|false|true|false|C0162429|Malnutrition|deficiency
Event|Event|SIMPLE_SEGMENT|11029,11039|false|false|false|||deficiency
Finding|Functional Concept|SIMPLE_SEGMENT|11029,11039|false|true|false|C0011155|Deficiency|deficiency
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11041,11047|false|false|false|C0002871|Anemia|anemia
Event|Event|SIMPLE_SEGMENT|11041,11047|false|false|false|||anemia
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11052,11058|false|false|false|C0002871|Anemia|anemia
Event|Event|SIMPLE_SEGMENT|11052,11058|false|false|false|||anemia
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11052,11077|false|false|false|C0002873|Anemia of chronic disease|anemia of chronic disease
Finding|Intellectual Product|SIMPLE_SEGMENT|11062,11069|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|11062,11069|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11062,11077|false|false|false|C0008679|Chronic disease|chronic disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11070,11077|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|11070,11077|false|false|false|||disease
Finding|Finding|SIMPLE_SEGMENT|11083,11086|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|SIMPLE_SEGMENT|11083,11086|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Finding|SIMPLE_SEGMENT|11083,11091|false|false|false|C0860975|Iron low|low iron
Drug|Biologically Active Substance|SIMPLE_SEGMENT|11087,11091|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|11087,11091|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11087,11091|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Event|Event|SIMPLE_SEGMENT|11087,11091|false|false|false|||iron
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|11087,11091|false|false|false|C0337439|Iron measurement|iron
Event|Event|SIMPLE_SEGMENT|11096,11104|false|false|false|||elevated
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|11106,11114|false|false|false|C0015879|Ferritin|ferritin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|11106,11114|false|false|false|C0015879|Ferritin|ferritin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11106,11114|false|false|false|C0015879|Ferritin|ferritin
Event|Event|SIMPLE_SEGMENT|11106,11114|false|false|false|||ferritin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|11106,11114|false|false|false|C0373607|Ferritin measurement|ferritin
Finding|Finding|SIMPLE_SEGMENT|11119,11122|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|SIMPLE_SEGMENT|11119,11122|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Event|Event|SIMPLE_SEGMENT|11123,11127|false|false|false|||TIBC
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|11123,11127|false|false|false|C0036835|Total Iron-Binding Capacity result|TIBC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|11123,11127|false|false|false|C1283048|Total iron binding capacity measurement|TIBC
Event|Event|SIMPLE_SEGMENT|11135,11144|false|false|false|||recommend
Event|Event|SIMPLE_SEGMENT|11145,11153|false|false|false|||checking
Event|Event|SIMPLE_SEGMENT|11164,11174|false|false|false|||outpatient
Finding|Classification|SIMPLE_SEGMENT|11164,11174|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|11164,11174|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|SIMPLE_SEGMENT|11179,11183|false|false|false|||work
Event|Occupational Activity|SIMPLE_SEGMENT|11179,11183|false|false|false|C0043227|Work|work
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|11179,11186|false|false|false|C0750430|Work-up|work-up
Event|Event|SIMPLE_SEGMENT|11190,11196|false|false|false|||needed
Event|Event|SIMPLE_SEGMENT|11205,11213|false|false|false|||swelling
Finding|Finding|SIMPLE_SEGMENT|11205,11213|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|SIMPLE_SEGMENT|11205,11213|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Event|Event|SIMPLE_SEGMENT|11222,11236|false|false|false|||multifactorial
Finding|Finding|SIMPLE_SEGMENT|11222,11236|false|false|false|C1837655|Multifactorial|multifactorial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11247,11253|false|false|false|C0042449|Veins|venous
Event|Event|SIMPLE_SEGMENT|11255,11268|false|false|false|||insufficiency
Finding|Functional Concept|SIMPLE_SEGMENT|11255,11268|false|false|false|C0231179|Insufficiency|insufficiency
Finding|Finding|SIMPLE_SEGMENT|11273,11277|false|false|false|C5575035|Well (answer to question)|well
Anatomy|Body Location or Region|SIMPLE_SEGMENT|11291,11294|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11291,11294|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11291,11294|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Event|Event|SIMPLE_SEGMENT|11291,11294|false|false|false|||DVT
Event|Event|SIMPLE_SEGMENT|11300,11309|false|false|false|||responded
Event|Event|SIMPLE_SEGMENT|11317,11321|false|false|false|||well
Finding|Finding|SIMPLE_SEGMENT|11317,11321|false|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|11327,11338|false|false|false|||compression
Finding|Functional Concept|SIMPLE_SEGMENT|11327,11338|false|false|false|C0332459;C4551657|Compressed structure|compression
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|11327,11338|false|false|false|C0728907|Compression|compression
Procedure|Machine Activity|SIMPLE_SEGMENT|11327,11338|false|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11327,11338|false|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Event|Event|SIMPLE_SEGMENT|11339,11348|false|false|false|||stockings
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11359,11366|false|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|SIMPLE_SEGMENT|11359,11366|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11359,11366|false|false|false|C0872388|Procedures on bladder|bladder
Disorder|Neoplastic Process|SIMPLE_SEGMENT|11359,11373|false|false|false|C0005684;C0005695;C0699885|Bladder Neoplasm;Carcinoma of bladder;Malignant neoplasm of urinary bladder|bladder cancer
Disorder|Neoplastic Process|SIMPLE_SEGMENT|11367,11373|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|SIMPLE_SEGMENT|11367,11373|false|false|false|||cancer
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11383,11388|false|false|false|C0401496|Transurethral resection of neoplasm of bladder|TURBT
Finding|Finding|SIMPLE_SEGMENT|11390,11394|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|SIMPLE_SEGMENT|11390,11394|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|SIMPLE_SEGMENT|11390,11394|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Classification|SIMPLE_SEGMENT|11395,11400|false|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|grade
Finding|Finding|SIMPLE_SEGMENT|11395,11400|false|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|grade
Anatomy|Cell Component|SIMPLE_SEGMENT|11401,11404|false|false|false|C1167383|membrane attack complex location|TCC
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11401,11404|false|false|false|C1861305|TARSAL-CARPAL COALITION SYNDROME|TCC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|11401,11404|false|false|false|C0077072;C5552697|Membrane Attack Complex;triclocarban|TCC
Drug|Biologically Active Substance|SIMPLE_SEGMENT|11401,11404|false|false|false|C0077072;C5552697|Membrane Attack Complex;triclocarban|TCC
Drug|Organic Chemical|SIMPLE_SEGMENT|11401,11404|false|false|false|C0077072;C5552697|Membrane Attack Complex;triclocarban|TCC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11401,11404|false|false|false|C0077072;C5552697|Membrane Attack Complex;triclocarban|TCC
Event|Event|SIMPLE_SEGMENT|11401,11404|false|false|false|||TCC
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11414,11420|true|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Anatomy|Tissue|SIMPLE_SEGMENT|11414,11420|true|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Event|Event|SIMPLE_SEGMENT|11421,11431|false|false|false|||identified
Finding|Intellectual Product|SIMPLE_SEGMENT|11434,11438|false|false|false|C1720594|Then - dosing instruction fragment|Then
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11447,11453|false|false|false|C0030797|Pelvis|pelvic
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|11447,11457|false|false|false|C0203201|Magnetic Resonance Imaging (MRI) of Pelvis|pelvic MRI
Event|Event|SIMPLE_SEGMENT|11454,11457|false|false|false|||MRI
Finding|Gene or Genome|SIMPLE_SEGMENT|11454,11457|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|11454,11457|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|SIMPLE_SEGMENT|11454,11457|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Event|Event|SIMPLE_SEGMENT|11458,11464|false|false|false|||showed
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11466,11473|false|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|SIMPLE_SEGMENT|11466,11473|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11466,11473|false|false|false|C0872388|Procedures on bladder|bladder
Finding|Finding|SIMPLE_SEGMENT|11466,11478|false|false|false|C0238775|Mass of urinary bladder|bladder mass
Finding|Finding|SIMPLE_SEGMENT|11474,11478|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|SIMPLE_SEGMENT|11474,11478|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|SIMPLE_SEGMENT|11474,11478|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Disorder|Neoplastic Process|SIMPLE_SEGMENT|11479,11487|false|false|false|C1269955|Tumor Cell Invasion|invasion
Event|Event|SIMPLE_SEGMENT|11479,11487|false|false|false|||invasion
Finding|Pathologic Function|SIMPLE_SEGMENT|11479,11487|false|false|false|C2699153|Cell Invasion|invasion
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11501,11505|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Anatomy|Body Location or Region|SIMPLE_SEGMENT|11501,11512|false|false|false|C0225317;C4532079|Neck+Chest>Soft tissue;soft tissue|soft tissue
Anatomy|Tissue|SIMPLE_SEGMENT|11501,11512|false|false|false|C0225317;C4532079|Neck+Chest>Soft tissue;soft tissue|soft tissue
Anatomy|Tissue|SIMPLE_SEGMENT|11506,11512|false|false|false|C0040300|Body tissue|tissue
Finding|Intellectual Product|SIMPLE_SEGMENT|11506,11512|false|false|false|C1547928|Tissue Specimen Code|tissue
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11514,11522|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11523,11530|false|false|false|C0042232|Vagina|vaginal
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|11523,11530|false|false|false|C1272941|Vaginal Dosage Form|vaginal
Finding|Finding|SIMPLE_SEGMENT|11523,11530|false|false|false|C1522570;C4521343|Vaginal (intended site);Vaginal Route of Administration|vaginal
Finding|Functional Concept|SIMPLE_SEGMENT|11523,11530|false|false|false|C1522570;C4521343|Vaginal (intended site);Vaginal Route of Administration|vaginal
Event|Event|SIMPLE_SEGMENT|11540,11545|false|false|false|||right
Finding|Functional Concept|SIMPLE_SEGMENT|11540,11545|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Event|Event|SIMPLE_SEGMENT|11554,11560|false|false|false|||lesion
Finding|Finding|SIMPLE_SEGMENT|11554,11560|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|SIMPLE_SEGMENT|11554,11560|false|false|false|C0221198;C1546698|Lesion|lesion
Event|Event|SIMPLE_SEGMENT|11581,11588|false|false|false|||robotic
Event|Event|SIMPLE_SEGMENT|11590,11593|false|false|false|||TAH
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11590,11593|false|false|false|C0404079|Total abdominal hysterectomy|TAH
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|11594,11597|false|false|false|C0054252|Buthionine Sulfoximine|BSO
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|11594,11597|false|false|false|C0054252|Buthionine Sulfoximine|BSO
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11594,11597|false|false|false|C0054252|Buthionine Sulfoximine|BSO
Event|Event|SIMPLE_SEGMENT|11594,11597|false|false|false|||BSO
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11599,11602|false|false|false|C0396060|Congenital laryngeal adductor palsy|lap
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|11599,11602|false|false|false|C1870042|ACP2 protein, human|lap
Drug|Enzyme|SIMPLE_SEGMENT|11599,11602|false|false|false|C1870042|ACP2 protein, human|lap
Event|Event|SIMPLE_SEGMENT|11599,11602|false|false|false|||lap
Finding|Finding|SIMPLE_SEGMENT|11599,11602|false|false|false|C0456170;C1412132;C1413323;C1423544;C1424863;C1425522;C2827449;C3540509;C5575443;C5890955|ACP2 gene;ACP2 wt Allele;CEBPB gene;CEBPB wt Allele;CENPJ gene;LAP3 gene;LAP3 wt Allele;Left atrial pressure;PICALM gene;PICALM wt Allele|lap
Finding|Gene or Genome|SIMPLE_SEGMENT|11599,11602|false|false|false|C0456170;C1412132;C1413323;C1423544;C1424863;C1425522;C2827449;C3540509;C5575443;C5890955|ACP2 gene;ACP2 wt Allele;CEBPB gene;CEBPB wt Allele;CENPJ gene;LAP3 gene;LAP3 wt Allele;Left atrial pressure;PICALM gene;PICALM wt Allele|lap
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|11599,11602|false|false|false|C0031150|Laparoscopy|lap
Drug|Chemical Viewed Structurally|SIMPLE_SEGMENT|11603,11610|false|false|false|C0302912|Radicals (chemistry)|radical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11603,11621|false|false|false|C0194401|Complete cystectomy|radical cystectomy
Event|Event|SIMPLE_SEGMENT|11611,11621|false|false|false|||cystectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11611,11621|false|false|false|C0010651|Cystectomy|cystectomy
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11626,11634|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Event|Event|SIMPLE_SEGMENT|11635,11646|false|false|false|||vaginectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11635,11646|false|false|false|C0195130|Vaginectomy|vaginectomy
Event|Event|SIMPLE_SEGMENT|11653,11662|false|false|false|||pathology
Finding|Functional Concept|SIMPLE_SEGMENT|11653,11662|false|false|false|C0205469;C0677042|Pathological aspects;Pathology processes|pathology
Finding|Pathologic Function|SIMPLE_SEGMENT|11653,11662|false|false|false|C0205469;C0677042|Pathological aspects;Pathology processes|pathology
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|11653,11662|false|false|false|C0919386|Pathology procedure|pathology
Event|Event|SIMPLE_SEGMENT|11663,11670|false|false|false|||showing
Finding|Finding|SIMPLE_SEGMENT|11671,11675|false|false|false|C1711132|pT2b TNM Finding|pT2b
Event|Event|SIMPLE_SEGMENT|11686,11693|false|false|false|||margins
Event|Event|SIMPLE_SEGMENT|11694,11702|false|false|false|||negative
Finding|Classification|SIMPLE_SEGMENT|11694,11702|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|11694,11702|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|11694,11702|false|false|false|C5237010|Expression Negative|negative
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11707,11711|true|false|false|C0270724|Infantile Neuroaxonal Dystrophy|plan
Event|Event|SIMPLE_SEGMENT|11707,11711|false|false|false|||plan
Finding|Functional Concept|SIMPLE_SEGMENT|11707,11711|true|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Intellectual Product|SIMPLE_SEGMENT|11707,11711|true|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Mental Process|SIMPLE_SEGMENT|11707,11711|true|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Event|Event|SIMPLE_SEGMENT|11729,11736|false|false|false|||therapy
Finding|Finding|SIMPLE_SEGMENT|11729,11736|true|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|SIMPLE_SEGMENT|11729,11736|true|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11729,11736|true|false|false|C0087111|Therapeutic procedure|therapy
Finding|Finding|SIMPLE_SEGMENT|11745,11749|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|11745,11749|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|11745,11749|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Body Substance|SIMPLE_SEGMENT|11767,11774|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|11767,11774|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|11767,11774|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|11778,11782|false|false|false|||safe
Finding|Intellectual Product|SIMPLE_SEGMENT|11778,11782|false|false|false|C4684764|SAFE-Biopharma Standard|safe
Event|Event|SIMPLE_SEGMENT|11786,11795|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|11786,11795|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|11786,11795|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|11786,11795|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|11786,11795|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|SIMPLE_SEGMENT|11819,11824|false|false|false|||spent
Event|Event|SIMPLE_SEGMENT|11829,11838|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|11829,11838|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|11829,11838|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|11829,11838|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|11829,11838|false|false|false|C0030685|Patient Discharge|discharge
Finding|Idea or Concept|SIMPLE_SEGMENT|11839,11842|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|11839,11842|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Occupational Activity|SIMPLE_SEGMENT|11843,11853|false|false|false|C0001554;C1273870|Administration occupational activities;Management procedure|management
Procedure|Health Care Activity|SIMPLE_SEGMENT|11843,11853|false|false|false|C0376636|Disease Management|management
Event|Event|SIMPLE_SEGMENT|11854,11862|false|false|false|||services
Event|Occupational Activity|SIMPLE_SEGMENT|11854,11862|false|false|false|C0557854|Services|services
Procedure|Health Care Activity|SIMPLE_SEGMENT|11854,11862|false|false|false|C1704289|Clinical Service|services
Finding|Idea or Concept|SIMPLE_SEGMENT|11865,11877|false|false|false|C1548597|Marketing basis - Transitional|Transitional
Event|Event|SIMPLE_SEGMENT|11878,11884|false|false|false|||issues
Event|Event|SIMPLE_SEGMENT|11897,11901|false|false|false|||need
Event|Event|SIMPLE_SEGMENT|11902,11908|false|false|false|||follow
Anatomy|Body Location or Region|SIMPLE_SEGMENT|11912,11917|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|11912,11917|false|false|false|C0741025|Chest problem|chest
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|11912,11920|false|false|false|C0202823|Chest CT|chest CT
Event|Event|SIMPLE_SEGMENT|11918,11920|false|false|false|||CT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11925,11934|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11925,11934|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|11925,11934|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Finding|SIMPLE_SEGMENT|11925,11942|false|false|false|C0748164|Multiple Pulmonary Nodules|pulmonary nodules
Event|Event|SIMPLE_SEGMENT|11935,11942|false|false|false|||nodules
Drug|Organic Chemical|SIMPLE_SEGMENT|11967,11975|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11967,11975|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|SIMPLE_SEGMENT|11967,11975|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Finding|Functional Concept|SIMPLE_SEGMENT|11967,11975|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|SIMPLE_SEGMENT|11967,11975|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|SIMPLE_SEGMENT|11978,11981|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|11978,11981|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|11982,11988|false|false|false|||course
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11993,11996|false|false|false|C0042029|Urinary tract infection|UTI
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|11993,11996|false|false|false|C0077906|urinastatin|UTI
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11993,11996|false|false|false|C0077906|urinastatin|UTI
Event|Event|SIMPLE_SEGMENT|11993,11996|false|false|false|||UTI
Finding|Gene or Genome|SIMPLE_SEGMENT|11993,11996|false|false|false|C1412376;C5780748|AMBP gene;AMBP wt Allele|UTI
Drug|Organic Chemical|SIMPLE_SEGMENT|12002,12010|false|false|false|C0591750|Macrobid|macrobid
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12002,12010|false|false|false|C0591750|Macrobid|macrobid
Event|Event|SIMPLE_SEGMENT|12002,12010|false|false|false|||macrobid
Event|Event|SIMPLE_SEGMENT|12012,12015|false|false|false|||day
Finding|Idea or Concept|SIMPLE_SEGMENT|12012,12015|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|12012,12015|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Finding|SIMPLE_SEGMENT|12012,12017|false|false|false|C3842672|Day 7|day 7
Drug|Biologically Active Substance|SIMPLE_SEGMENT|12034,12040|false|false|false|C0030054|oxygen|oxygen
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|12034,12040|false|false|false|C0030054|oxygen|oxygen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12034,12040|false|false|false|C0030054|oxygen|oxygen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|12034,12040|false|false|false|C0184633|Oxygen Therapy Care|oxygen
Finding|Finding|SIMPLE_SEGMENT|12034,12048|false|false|false|C1546419|Ambulatory Status - Oxygen therapy|oxygen therapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|12034,12048|false|false|false|C0184633;C3665674|Oxygen Therapy Care;Warburg Therapy|oxygen therapy
Event|Event|SIMPLE_SEGMENT|12041,12048|false|false|false|||therapy
Finding|Finding|SIMPLE_SEGMENT|12041,12048|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|SIMPLE_SEGMENT|12041,12048|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|12041,12048|false|false|false|C0087111|Therapeutic procedure|therapy
Finding|Finding|SIMPLE_SEGMENT|12053,12057|false|false|false|C0043084|Weaning|wean
Event|Event|SIMPLE_SEGMENT|12061,12070|false|false|false|||tolerated
Drug|Substance|SIMPLE_SEGMENT|12074,12082|false|false|false|C0721534|Maintain brand of benzocaine|maintain
Event|Activity|SIMPLE_SEGMENT|12074,12082|false|false|false|C0024501|Maintenance|maintain
Event|Event|SIMPLE_SEGMENT|12087,12090|false|false|false|||sat
Event|Event|SIMPLE_SEGMENT|12107,12112|false|false|false|||check
Anatomy|Cell Component|SIMPLE_SEGMENT|12113,12116|false|false|false|C2263086|Nuclear cap binding complex location|CBC
Event|Event|SIMPLE_SEGMENT|12113,12116|false|false|false|||CBC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|12113,12116|false|false|false|C0009555|Complete Blood Count|CBC
Event|Event|SIMPLE_SEGMENT|12127,12133|false|false|false|||ensure
Event|Event|SIMPLE_SEGMENT|12134,12143|false|false|false|||stability
Event|Event|SIMPLE_SEGMENT|12156,12167|false|false|false|||demonstrate
Event|Event|SIMPLE_SEGMENT|12168,12178|false|false|false|||resolution
Finding|Conceptual Entity|SIMPLE_SEGMENT|12168,12178|false|false|false|C1514893;C2699488|Resolution;physiologic resolution|resolution
Finding|Pathologic Function|SIMPLE_SEGMENT|12168,12178|false|false|false|C1514893;C2699488|Resolution;physiologic resolution|resolution
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12182,12194|false|false|false|C0023518|Leukocytosis|leukocytosis
Event|Event|SIMPLE_SEGMENT|12182,12194|false|false|false|||leukocytosis
Finding|Finding|SIMPLE_SEGMENT|12182,12194|false|false|false|C0750426|Blood leukocyte number above reference range|leukocytosis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12197,12200|false|false|false|C0162531|Hereditary Coproporphyria|HCP
Event|Event|SIMPLE_SEGMENT|12197,12200|false|false|false|||HCP
Finding|Gene or Genome|SIMPLE_SEGMENT|12197,12200|false|false|false|C1335283;C1412376;C1413681;C1705637;C5780748|AMBP gene;AMBP wt Allele;CPOX gene;PTPN6 gene;PTPN6 wt Allele|HCP
Finding|Gene or Genome|SIMPLE_SEGMENT|12202,12205|false|false|false|C1420310|SON gene|son
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12222,12233|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12222,12233|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|12222,12233|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|12222,12233|false|false|false|C4284232|Medications|Medications
Finding|Finding|SIMPLE_SEGMENT|12222,12246|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|SIMPLE_SEGMENT|12237,12246|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|12237,12246|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12265,12275|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|12265,12275|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|12265,12280|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|SIMPLE_SEGMENT|12276,12280|false|false|false|||list
Finding|Intellectual Product|SIMPLE_SEGMENT|12276,12280|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|SIMPLE_SEGMENT|12288,12298|false|false|false|||inaccurate
Event|Event|SIMPLE_SEGMENT|12303,12311|false|false|false|||requires
Event|Event|SIMPLE_SEGMENT|12320,12333|false|false|false|||investigation
Finding|Intellectual Product|SIMPLE_SEGMENT|12320,12333|false|false|false|C1552578|Act Class - investigation|investigation
Procedure|Health Care Activity|SIMPLE_SEGMENT|12320,12333|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|investigation
Drug|Organic Chemical|SIMPLE_SEGMENT|12338,12351|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12338,12351|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|SIMPLE_SEGMENT|12338,12351|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|12338,12351|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Drug|Organic Chemical|SIMPLE_SEGMENT|12370,12378|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12370,12378|false|false|false|C1692318|docusate|Docusate
Event|Event|SIMPLE_SEGMENT|12370,12378|false|false|false|||Docusate
Drug|Organic Chemical|SIMPLE_SEGMENT|12370,12385|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12370,12385|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|12379,12385|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|12379,12385|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12379,12385|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|SIMPLE_SEGMENT|12379,12385|false|false|false|||Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|12379,12385|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|12379,12385|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|12396,12399|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|12396,12399|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|12396,12399|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|12396,12399|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|12396,12399|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|12404,12414|false|false|false|C0206460|enoxaparin|Enoxaparin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12404,12414|false|false|false|C0206460|enoxaparin|Enoxaparin
Event|Event|SIMPLE_SEGMENT|12404,12414|false|false|false|||Enoxaparin
Drug|Organic Chemical|SIMPLE_SEGMENT|12404,12421|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12404,12421|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|12415,12421|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|12415,12421|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12415,12421|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|SIMPLE_SEGMENT|12415,12421|false|false|false|||Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|12415,12421|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|12415,12421|false|false|false|C0337443|Sodium measurement|Sodium
Event|Event|SIMPLE_SEGMENT|12438,12443|false|false|false|||Start
Finding|Idea or Concept|SIMPLE_SEGMENT|12462,12466|false|false|false|C1552851|next - HtmlLinkType|Next
Event|Event|SIMPLE_SEGMENT|12467,12474|false|false|false|||Routine
Finding|Idea or Concept|SIMPLE_SEGMENT|12467,12474|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|Routine
Finding|Intellectual Product|SIMPLE_SEGMENT|12467,12474|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|Routine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|12467,12474|false|false|false|C1979801|Routine coag|Routine
Event|Occupational Activity|SIMPLE_SEGMENT|12475,12489|false|false|false|C0001554|Administration occupational activities|Administration
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|12475,12489|false|false|false|C1533734|Administration (procedure)|Administration
Finding|Finding|SIMPLE_SEGMENT|12490,12494|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Finding|Idea or Concept|SIMPLE_SEGMENT|12490,12494|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Finding|Intellectual Product|SIMPLE_SEGMENT|12490,12494|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|12499,12512|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Hormone|SIMPLE_SEGMENT|12499,12512|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Organic Chemical|SIMPLE_SEGMENT|12499,12512|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12499,12512|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Event|Event|SIMPLE_SEGMENT|12499,12512|false|false|false|||Levothyroxine
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|12499,12519|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Hormone|SIMPLE_SEGMENT|12499,12519|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12499,12519|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|12513,12519|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|12513,12519|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12513,12519|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|SIMPLE_SEGMENT|12513,12519|false|false|false|||Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|12513,12519|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|12513,12519|false|false|false|C0337443|Sodium measurement|Sodium
Drug|Organic Chemical|SIMPLE_SEGMENT|12541,12553|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12541,12553|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|SIMPLE_SEGMENT|12571,12579|false|false|false|C0126174|losartan|Losartan
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12571,12579|false|false|false|C0126174|losartan|Losartan
Event|Event|SIMPLE_SEGMENT|12571,12579|false|false|false|||Losartan
Drug|Organic Chemical|SIMPLE_SEGMENT|12571,12589|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12571,12589|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|12580,12589|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|12580,12589|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Food|SIMPLE_SEGMENT|12580,12589|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|12580,12589|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12580,12589|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Event|Event|SIMPLE_SEGMENT|12580,12589|false|false|false|||Potassium
Finding|Physiologic Function|SIMPLE_SEGMENT|12580,12589|false|false|false|C4553027|Potassium metabolic function|Potassium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|12580,12589|false|false|false|C0202194|Potassium measurement|Potassium
Drug|Organic Chemical|SIMPLE_SEGMENT|12609,12618|false|false|false|C0030049|oxycodone|OxyCODONE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12609,12618|false|false|false|C0030049|oxycodone|OxyCODONE
Event|Event|SIMPLE_SEGMENT|12609,12618|false|false|false|||OxyCODONE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|12609,12618|false|false|false|C0524222|Oxycodone measurement|OxyCODONE
Finding|Idea or Concept|SIMPLE_SEGMENT|12620,12629|false|false|false|C1548167;C1697779|Query Priority - Immediate;immediate - ResponseCode|Immediate
Finding|Intellectual Product|SIMPLE_SEGMENT|12620,12629|false|false|false|C1548167;C1697779|Query Priority - Immediate;immediate - ResponseCode|Immediate
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|12620,12637|false|false|false|C1708470|Immediate Release Dosage Form|Immediate Release
Event|Event|SIMPLE_SEGMENT|12630,12637|false|false|false|||Release
Finding|Functional Concept|SIMPLE_SEGMENT|12630,12637|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|12630,12637|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|12630,12637|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Finding|Gene or Genome|SIMPLE_SEGMENT|12651,12654|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12655,12659|false|false|false|C2598155||Pain
Event|Event|SIMPLE_SEGMENT|12655,12659|false|false|false|||Pain
Finding|Functional Concept|SIMPLE_SEGMENT|12655,12659|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|12655,12659|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Finding|SIMPLE_SEGMENT|12662,12670|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Intellectual Product|SIMPLE_SEGMENT|12662,12670|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Drug|Organic Chemical|SIMPLE_SEGMENT|12676,12685|false|false|false|C0024002|lorazepam|LORazepam
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12676,12685|false|false|false|C0024002|lorazepam|LORazepam
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|12697,12700|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|12697,12700|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|12697,12700|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|12697,12700|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|12697,12700|false|false|false|C1332410|BID gene|BID
Finding|Gene or Genome|SIMPLE_SEGMENT|12701,12704|false|false|false|C1422467|CIAO3 gene|PRN
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|12705,12712|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Event|Event|SIMPLE_SEGMENT|12705,12712|false|false|false|||anxiety
Finding|Sign or Symptom|SIMPLE_SEGMENT|12705,12712|false|false|false|C0860603|Anxiety symptoms|anxiety
Drug|Organic Chemical|SIMPLE_SEGMENT|12717,12722|false|false|false|C3489575|sennosides, USP|Senna
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12717,12722|false|false|false|C3489575|sennosides, USP|Senna
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|12733,12736|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|12733,12736|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|12733,12736|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|12733,12736|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|12733,12736|false|false|false|C1332410|BID gene|BID
Event|Event|SIMPLE_SEGMENT|12741,12750|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|12741,12750|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|12741,12750|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|12741,12750|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|12741,12750|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|12741,12762|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12751,12762|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12751,12762|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|12751,12762|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|12751,12762|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|SIMPLE_SEGMENT|12768,12782|false|false|false|C0028156|nitrofurantoin|Nitrofurantoin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12768,12782|false|false|false|C0028156|nitrofurantoin|Nitrofurantoin
Drug|Organic Chemical|SIMPLE_SEGMENT|12792,12800|false|false|false|C0591750|Macrobid|MacroBID
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12792,12800|false|false|false|C0591750|Macrobid|MacroBID
Finding|Idea or Concept|SIMPLE_SEGMENT|12823,12826|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|12823,12826|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|SIMPLE_SEGMENT|12834,12844|false|false|false|C0206460|enoxaparin|Enoxaparin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12834,12844|false|false|false|C0206460|enoxaparin|Enoxaparin
Drug|Organic Chemical|SIMPLE_SEGMENT|12834,12851|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12834,12851|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|12845,12851|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|12845,12851|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12845,12851|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|SIMPLE_SEGMENT|12845,12851|false|false|false|||Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|12845,12851|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|12845,12851|false|false|false|C0337443|Sodium measurement|Sodium
Event|Event|SIMPLE_SEGMENT|12867,12872|false|false|false|||Start
Finding|Idea or Concept|SIMPLE_SEGMENT|12899,12903|false|false|false|C1552851|next - HtmlLinkType|Next
Finding|Idea or Concept|SIMPLE_SEGMENT|12904,12911|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|Routine
Finding|Intellectual Product|SIMPLE_SEGMENT|12904,12911|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|Routine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|12904,12911|false|false|false|C1979801|Routine coag|Routine
Event|Event|SIMPLE_SEGMENT|12912,12926|false|false|false|||Administration
Event|Occupational Activity|SIMPLE_SEGMENT|12912,12926|false|false|false|C0001554|Administration occupational activities|Administration
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|12912,12926|false|false|false|C1533734|Administration (procedure)|Administration
Finding|Finding|SIMPLE_SEGMENT|12928,12932|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Finding|Idea or Concept|SIMPLE_SEGMENT|12928,12932|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Finding|Intellectual Product|SIMPLE_SEGMENT|12928,12932|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Drug|Organic Chemical|SIMPLE_SEGMENT|12939,12948|false|false|false|C0024002|lorazepam|LORazepam
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12939,12948|false|false|false|C0024002|lorazepam|LORazepam
Finding|Gene or Genome|SIMPLE_SEGMENT|12964,12967|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12968,12976|false|false|false|C1950154|Insomnia homeopathic medication|insomnia
Event|Event|SIMPLE_SEGMENT|12968,12976|false|false|false|||insomnia
Finding|Sign or Symptom|SIMPLE_SEGMENT|12968,12976|false|false|false|C0917801|Sleeplessness|insomnia
Event|Event|SIMPLE_SEGMENT|12978,12980|false|false|false|||RX
Drug|Organic Chemical|SIMPLE_SEGMENT|12982,12991|false|false|false|C0024002|lorazepam|lorazepam
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12982,12991|false|false|false|C0024002|lorazepam|lorazepam
Event|Event|SIMPLE_SEGMENT|12982,12991|false|false|false|||lorazepam
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|13014,13017|false|false|false|C0039225|Tablet Dosage Form|tab
Event|Event|SIMPLE_SEGMENT|13014,13017|false|false|false|||tab
Finding|Functional Concept|SIMPLE_SEGMENT|13018,13026|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|13021,13026|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|13021,13026|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Gene or Genome|SIMPLE_SEGMENT|13031,13034|false|false|false|C1422467|CIAO3 gene|prn
Event|Activity|SIMPLE_SEGMENT|13035,13039|false|false|false|C1880359|Dispense (activity)|Disp
Event|Event|SIMPLE_SEGMENT|13035,13039|false|false|false|||Disp
Finding|Gene or Genome|SIMPLE_SEGMENT|13035,13039|false|false|false|C2828567|PRSS30P gene|Disp
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|13045,13051|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|13052,13059|false|false|false|||Refills
Finding|Idea or Concept|SIMPLE_SEGMENT|13052,13059|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|13068,13081|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13068,13081|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|SIMPLE_SEGMENT|13068,13081|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|13068,13081|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Drug|Organic Chemical|SIMPLE_SEGMENT|13102,13114|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13102,13114|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|SIMPLE_SEGMENT|13134,13142|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13134,13142|false|false|false|C1692318|docusate|Docusate
Event|Event|SIMPLE_SEGMENT|13134,13142|false|false|false|||Docusate
Drug|Organic Chemical|SIMPLE_SEGMENT|13134,13149|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13134,13149|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|13143,13149|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|13143,13149|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13143,13149|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|SIMPLE_SEGMENT|13143,13149|false|false|false|||Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|13143,13149|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|13143,13149|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|13160,13163|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|13160,13163|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|13160,13163|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|13160,13163|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|13160,13163|false|false|false|C1332410|BID gene|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|13170,13183|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Hormone|SIMPLE_SEGMENT|13170,13183|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Organic Chemical|SIMPLE_SEGMENT|13170,13183|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13170,13183|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|13170,13190|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Hormone|SIMPLE_SEGMENT|13170,13190|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13170,13190|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|13184,13190|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|13184,13190|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13184,13190|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|SIMPLE_SEGMENT|13184,13190|false|false|false|||Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|13184,13190|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|13184,13190|false|false|false|C0337443|Sodium measurement|Sodium
Drug|Organic Chemical|SIMPLE_SEGMENT|13214,13223|false|false|false|C0030049|oxycodone|OxyCODONE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13214,13223|false|false|false|C0030049|oxycodone|OxyCODONE
Event|Event|SIMPLE_SEGMENT|13214,13223|false|false|false|||OxyCODONE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|13214,13223|false|false|false|C0524222|Oxycodone measurement|OxyCODONE
Finding|Idea or Concept|SIMPLE_SEGMENT|13225,13234|false|false|false|C1548167;C1697779|Query Priority - Immediate;immediate - ResponseCode|Immediate
Finding|Intellectual Product|SIMPLE_SEGMENT|13225,13234|false|false|false|C1548167;C1697779|Query Priority - Immediate;immediate - ResponseCode|Immediate
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|13225,13242|false|false|false|C1708470|Immediate Release Dosage Form|Immediate Release
Event|Event|SIMPLE_SEGMENT|13235,13242|false|false|false|||Release
Finding|Functional Concept|SIMPLE_SEGMENT|13235,13242|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|13235,13242|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|13235,13242|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Finding|Gene or Genome|SIMPLE_SEGMENT|13256,13259|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13260,13264|false|false|false|C2598155||Pain
Finding|Functional Concept|SIMPLE_SEGMENT|13260,13264|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|13260,13264|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Finding|SIMPLE_SEGMENT|13268,13276|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Intellectual Product|SIMPLE_SEGMENT|13268,13276|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Event|Event|SIMPLE_SEGMENT|13278,13280|false|false|false|||RX
Drug|Organic Chemical|SIMPLE_SEGMENT|13282,13291|false|false|false|C0030049|oxycodone|oxycodone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13282,13291|false|false|false|C0030049|oxycodone|oxycodone
Event|Event|SIMPLE_SEGMENT|13282,13291|false|false|false|||oxycodone
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|13282,13291|false|false|false|C0524222|Oxycodone measurement|oxycodone
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|13299,13305|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|SIMPLE_SEGMENT|13309,13317|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|13312,13317|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|13312,13317|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Gene or Genome|SIMPLE_SEGMENT|13322,13325|false|false|false|C1422467|CIAO3 gene|prn
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|13335,13341|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|13335,13341|false|false|false|||Tablet
Event|Event|SIMPLE_SEGMENT|13343,13350|false|false|false|||Refills
Finding|Idea or Concept|SIMPLE_SEGMENT|13343,13350|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|13359,13364|false|false|false|C3489575|sennosides, USP|Senna
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13359,13364|false|false|false|C3489575|sennosides, USP|Senna
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|13375,13378|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|13375,13378|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|13375,13378|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|13375,13378|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|13375,13378|false|false|false|C1332410|BID gene|BID
Event|Event|SIMPLE_SEGMENT|13384,13393|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|13384,13393|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|13384,13393|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|13384,13393|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|13384,13393|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13384,13405|false|false|false|C4019243||Discharge Disposition
Finding|Finding|SIMPLE_SEGMENT|13384,13405|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13394,13405|false|false|false|C2926604||Disposition
Event|Event|SIMPLE_SEGMENT|13394,13405|false|false|false|||Disposition
Procedure|Health Care Activity|SIMPLE_SEGMENT|13394,13405|false|false|false|C0184758|Patient disposition|Disposition
Finding|Finding|SIMPLE_SEGMENT|13407,13415|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|SIMPLE_SEGMENT|13407,13415|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Procedure|Health Care Activity|SIMPLE_SEGMENT|13407,13420|false|false|false|C0023977|long-term care|Extended Care
Event|Activity|SIMPLE_SEGMENT|13416,13420|false|false|false|C1947933|care activity|Care
Event|Event|SIMPLE_SEGMENT|13416,13420|false|false|false|||Care
Finding|Finding|SIMPLE_SEGMENT|13416,13420|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|SIMPLE_SEGMENT|13416,13420|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Event|Event|SIMPLE_SEGMENT|13423,13431|false|false|false|||Facility
Finding|Intellectual Product|SIMPLE_SEGMENT|13423,13431|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|SIMPLE_SEGMENT|13439,13448|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|13439,13448|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|13439,13448|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|13439,13448|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|13439,13448|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|13439,13458|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13449,13458|false|false|false|C0945731||Diagnosis
Event|Event|SIMPLE_SEGMENT|13449,13458|false|false|false|||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|13449,13458|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|13449,13458|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|13449,13458|false|false|false|C0011900|Diagnosis|Diagnosis
Event|Event|SIMPLE_SEGMENT|13465,13474|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|13465,13474|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|13465,13474|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|13465,13474|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|13465,13474|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13475,13484|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13475,13484|false|false|false|C0012634|Disease|Condition
Event|Event|SIMPLE_SEGMENT|13475,13484|false|false|false|||Condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|13475,13484|false|false|false|C1705253|Logical Condition|Condition
Finding|Mental Process|SIMPLE_SEGMENT|13486,13492|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13486,13499|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|SIMPLE_SEGMENT|13486,13499|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13493,13499|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|13493,13499|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|13501,13506|false|false|false|||Clear
Finding|Idea or Concept|SIMPLE_SEGMENT|13501,13506|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|SIMPLE_SEGMENT|13511,13519|false|false|false|||coherent
Finding|Finding|SIMPLE_SEGMENT|13511,13519|false|false|false|C4068804|Coherent|coherent
Event|Event|SIMPLE_SEGMENT|13521,13526|false|false|false|||Level
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13521,13543|false|false|false|C4050479||Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|13521,13543|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|SIMPLE_SEGMENT|13530,13543|false|false|false|||Consciousness
Finding|Finding|SIMPLE_SEGMENT|13530,13543|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|SIMPLE_SEGMENT|13530,13543|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13545,13550|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|13545,13550|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13545,13550|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|SIMPLE_SEGMENT|13545,13550|false|false|false|||Alert
Finding|Finding|SIMPLE_SEGMENT|13545,13550|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|13545,13550|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|13545,13550|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|SIMPLE_SEGMENT|13555,13566|false|false|false|||interactive
Finding|Functional Concept|SIMPLE_SEGMENT|13555,13566|false|false|false|C1704675|Interaction|interactive
Event|Activity|SIMPLE_SEGMENT|13568,13576|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|13568,13576|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|SIMPLE_SEGMENT|13568,13576|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13577,13583|false|false|false|C5889824||Status
Event|Event|SIMPLE_SEGMENT|13577,13583|false|false|false|||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|13577,13583|false|false|false|C1546481|What subject filter - Status|Status
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13592,13595|false|false|false|C3159311|BORNHOLM EYE DISEASE|Bed
Event|Event|SIMPLE_SEGMENT|13592,13595|false|false|false|||Bed
Finding|Intellectual Product|SIMPLE_SEGMENT|13592,13595|false|false|false|C2346952|Bachelor of Education|Bed
Event|Event|SIMPLE_SEGMENT|13601,13611|false|false|false|||assistance
Finding|Social Behavior|SIMPLE_SEGMENT|13601,13611|false|false|false|C0018896|Helping Behavior|assistance
Event|Event|SIMPLE_SEGMENT|13625,13635|false|false|false|||wheelchair
Finding|Finding|SIMPLE_SEGMENT|13625,13635|false|false|false|C2135586;C4321408|Wheelchair Usually Used;has wheelchair at home (history)|wheelchair
Event|Event|SIMPLE_SEGMENT|13640,13649|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|13640,13649|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|13640,13649|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|13640,13649|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|13640,13649|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13640,13662|false|false|false|C3669312||Discharge Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|13640,13662|false|false|false|C4282220|Discharge instructions|Discharge Instructions
Procedure|Health Care Activity|SIMPLE_SEGMENT|13640,13662|false|false|false|C2266673|hospital discharge instructions (treatment)|Discharge Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13650,13662|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|13650,13662|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|13650,13662|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Event|Event|SIMPLE_SEGMENT|13681,13689|false|false|false|||pleasure
Finding|Intellectual Product|SIMPLE_SEGMENT|13681,13689|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|SIMPLE_SEGMENT|13681,13689|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|SIMPLE_SEGMENT|13697,13701|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|13697,13701|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|13697,13701|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|13697,13701|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Event|Event|SIMPLE_SEGMENT|13719,13728|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|13719,13728|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|SIMPLE_SEGMENT|13746,13754|false|false|false|||admitted
Drug|Organic Chemical|SIMPLE_SEGMENT|13761,13765|false|false|false|C0009074|clotrimazole|clot
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13761,13765|false|false|false|C0009074|clotrimazole|clot
Event|Event|SIMPLE_SEGMENT|13761,13765|false|false|false|||clot
Finding|Pathologic Function|SIMPLE_SEGMENT|13761,13765|false|false|false|C0302148|Blood Clot|clot
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|13774,13779|false|false|false|C0024109|Lung|lungs
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|13785,13788|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Event|Event|SIMPLE_SEGMENT|13799,13806|false|false|false|||treated
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13814,13819|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|13814,13819|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|13814,13819|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Event|Event|SIMPLE_SEGMENT|13820,13827|false|false|false|||thinner
Event|Event|SIMPLE_SEGMENT|13838,13842|false|false|false|||need
Event|Event|SIMPLE_SEGMENT|13847,13855|false|false|false|||continue
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13860,13865|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|13860,13865|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|13860,13865|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Event|Event|SIMPLE_SEGMENT|13866,13873|false|false|false|||thinner
Event|Event|SIMPLE_SEGMENT|13889,13896|false|false|false|||treated
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|13903,13910|false|false|false|C0042027|Urinary tract|urinary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|13912,13917|false|false|false|C1185740|Tract|tract
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13918,13927|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|SIMPLE_SEGMENT|13918,13927|false|false|false|||infection
Finding|Pathologic Function|SIMPLE_SEGMENT|13918,13927|false|false|false|C3714514|Infection|infection
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|13938,13947|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13938,13947|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|13938,13947|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Finding|SIMPLE_SEGMENT|13938,13955|false|false|false|C0748164|Multiple Pulmonary Nodules|pulmonary nodules
Event|Event|SIMPLE_SEGMENT|13948,13955|false|false|false|||nodules
Event|Event|SIMPLE_SEGMENT|13968,13974|false|false|false|||follow
Finding|Intellectual Product|SIMPLE_SEGMENT|13989,14001|false|false|false|C1547426|Location Service Code - Primary Care|primary care
Procedure|Health Care Activity|SIMPLE_SEGMENT|13989,14001|false|false|false|C0033137|Primary Health Care|primary care
Event|Activity|SIMPLE_SEGMENT|13997,14001|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|13997,14001|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|13997,14001|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|13997,14001|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|14002,14008|false|false|false|C2348314|Doctor - Title|doctor
Procedure|Health Care Activity|SIMPLE_SEGMENT|14013,14021|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14022,14034|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|14022,14034|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|14022,14034|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

