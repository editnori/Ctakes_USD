CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|true|false||Unit
null|Unit device|Device|true|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|true|false||Unit
null|Unit of Measure|LabModifier|true|false||Unit
null|Unit|LabModifier|true|false||Unit
null|Enzyme Unit|LabModifier|true|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Pharmaceutical Preparations|Drug|false|false||MEDICINEnull|Medicine|Title|false|false||MEDICINEnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|lisinopril|Drug|false|false||lisinopril
null|lisinopril|Drug|false|false||lisinoprilnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Chief complaint (finding)|Finding|false|false||Chief Complaintnull|Complaint (finding)|Finding|false|false||Complaintnull|null|Attribute|false|false||Complaintnull|Chest Pain|Finding|false|false||chest painnull|null|Attribute|false|false||chest painnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Cardiac catheterisation as the cause of abnormal reaction of the patient, or of later complication, without mention of misadventure at the time of the procedure|Disorder|false|false||cardiac catheterizationnull|Diagnostic Service Section ID - Cardiac Catheterization|Finding|false|false||cardiac catheterizationnull|Consent Type - Cardiac Catheterization|Procedure|false|false||cardiac catheterization
null|Cardiac Catheterization Procedures|Procedure|false|false||cardiac catheterizationnull|Cardiac attachment|Finding|false|false||cardiacnull|Heart|Anatomy|false|false||cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||cardiacnull|Catheterization|Procedure|false|false||catheterizationnull|History of present illness (finding)|Finding|false|false||History of Present Illnessnull|null|Attribute|false|false||History of Present Illnessnull|Medical History|Finding|false|false||History ofnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Present illness|Finding|false|false||Present Illnessnull|Present|Finding|false|false||Present
null|Presentation|Finding|false|false||Presentnull|Illness (finding)|Finding|false|false||Illnessnull|PMH - past medical history|Finding|false|false||PMH
null|Medical History|Finding|false|false||PMHnull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|SERPINA5 protein, human|Drug|false|false||PCI
null|SERPINA5 protein, human|Drug|false|false||PCInull|Peritoneal Cancer Index|Finding|false|false||PCI
null|SERPINA5 wt Allele|Finding|false|false||PCI
null|SERPINA5 gene|Finding|false|false||PCInull|Percutaneous Coronary Intervention|Procedure|false|false||PCI
null|photochemical internalization|Procedure|false|false||PCI
null|Prophylactic Cranial Irradiation|Procedure|false|false||PCInull|Picocurie|LabModifier|false|false||PCInull|matrix metalloproteinase 7 activity|Finding|false|false||pumpnull|null|Device|false|false||pumpnull|Pump Dosing Unit|LabModifier|false|false||pumpnull|Coronary Artery Bypass Surgery|Procedure|false|false||CABGnull|Leukocyte adhesion deficiency type 1|Disorder|false|false||LAD
null|Leukocyte adhesion deficiency|Disorder|false|false||LADnull|ITGB2 wt Allele|Finding|false|false||LAD
null|DLD gene|Finding|false|false||LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false||LADnull|Ladino Language|Entity|false|false||LADnull|Scalable Vector Graphics|Entity|false|false||SVGnull|diagnosis aspects|Finding|false|false||diagnull|Diagnosis|Procedure|false|false||diagnull|Type 2|Finding|false|false||type 2null|Type - ParameterizedDataType|Finding|false|false||type
null|SGCG gene|Finding|false|false||typenull|null|Modifier|false|false||typenull|insulin, regular, human|Drug|false|false||insulin
null|Insulin [EPC]|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulinnull|INS gene|Finding|false|false||insulinnull|Insulin measurement|Procedure|false|false||insulinnull|Hypertensive disease|Disorder|false|false||HTNnull|Hyperlipidemia|Disorder|false|false||hyperlipidemia
null|Hyperlipoproteinemias|Disorder|false|false||hyperlipidemianull|Serum lipids high (finding)|Finding|false|false||hyperlipidemianull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Sharp sensation quality|Finding|false|false||sharp
null|SPEN wt Allele|Finding|false|false||sharp
null|SPEN gene|Finding|false|false||sharpnull|Left sided|Modifier|false|false||left-sidednull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Chest Pain|Finding|false|false||chest painnull|null|Attribute|false|false||chest painnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Dyspnea|Finding|false|false||SOBnull|Chest Pain|Finding|false|false||chest painnull|null|Attribute|false|false||chest painnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pinched|Disorder|false|false||pinchingnull|Specimen Type - Bone|Finding|false|false||bone
null|null|Finding|false|false||bonenull|Skeletal bone|Anatomy|false|false||bone
null|XXX bone|Anatomy|false|false||bonenull|Episode of|Time|false|false||episodesnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|per day|Time|false|false||/daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Always - AcknowledgementCondition|Finding|false|false||always
null|All of the Time|Finding|false|false||alwaysnull|Always (frequency)|Time|false|false||alwaysnull|At rest (qualifier value)|Finding|false|false||at restnull|REST protein, human|Drug|false|false||rest
null|REST protein, human|Drug|false|false||restnull|REST gene|Finding|false|false||rest
null|site-specific telomere resolvase activity|Finding|false|false||rest
null|Rest|Finding|false|false||restnull|Episode of|Time|false|false||episodesnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Last|Modifier|false|false||lastnull|Approximate|Modifier|false|false||approximatelynull|5 minutes Office visit|Procedure|false|false||5 minutesnull|5 minutes|Time|false|false||5 minutesnull|Minute of time|Time|false|false||minutesnull|Minute Unit of Plane Angle|LabModifier|false|false||minutes
null|Minute (diminutive)|LabModifier|false|false||minutes
null|Small|LabModifier|false|false||minutesnull|nitroglycerin|Drug|false|false||nitroglycerin
null|nitroglycerin|Drug|false|false||nitroglycerinnull|Administration Method - Pain|Finding|true|false||pain
null|Pain|Finding|true|false||painnull|null|Attribute|true|false||painnull|Exertion|Finding|true|false||exertionnull|Eating|Finding|true|false||eatingnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|Authorization Mode - Phone|Finding|false|false||phone
null|Visit User Code - Phone|Finding|false|false||phone
null|Telephone Number|Finding|false|false||phone
null|MDFAttributeType - Phone|Finding|false|false||phonenull|Telephone|Device|false|false||phonenull|Person location type - Phone|Modifier|false|false||phonenull|Similarity|Modifier|false|false||similarnull|Vomiting|Finding|false|false||vomitingnull|Last|Modifier|false|false||lastnull|Night time|Time|false|false||nightnull|Increased sweating|Finding|true|false||diaphoresisnull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|Has patient|Finding|false|false||patient hasnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Increasing breathlessness|Finding|false|false||increased shortness of breathnull|Dyspnea|Finding|false|false||shortness of breathnull|null|Attribute|false|false||shortness of breathnull|Breath|Finding|false|false||breathnull|day|Time|false|false||daysnull|sleeping upright or using specific number of extra pillows (orthopnea)|Finding|false|false||orthopnea
null|Orthopnea|Finding|false|false||orthopneanull|year|Time|false|false||yearsnull|Paroxysmal nocturnal dyspnea|Disorder|true|false||PNDnull|NPPA wt Allele|Finding|true|false||PND
null|NPPA gene|Finding|true|false||PNDnull|Edema of lower extremity|Finding|true|false||lower extremity edemanull|Lower Extremity|Anatomy|true|false||lower extremitynull|Body Site Modifier - Lower|Anatomy|true|false||lowernull|Lower (action)|Event|true|false||lowernull|Lower - spatial qualifier|Modifier|true|false||lowernull|Peripheral edema|Finding|true|false||extremity edemanull|Limb structure|Anatomy|true|false||extremitynull|Edema|Finding|true|false||edemanull|null|Attribute|true|false||edemanull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Regular|Modifier|false|false||regularnull|Rhythm|Finding|false|false||rhythm
null|rhythmic process (biological)|Finding|false|false||rhythmnull|Lung|Anatomy|false|false||Lungsnull|cetrimonium bromide|Drug|false|false||CTABnull|Sequence Chromatogram|Finding|false|false||tracenull|Trace Dosing Unit|LabModifier|false|false||trace
null|trace amount|LabModifier|false|false||trace
null|unknown - trace|LabModifier|false|false||tracenull|Edema|Finding|true|false||edemanull|null|Attribute|true|false||edemanull|Left lower extremity|Anatomy|true|false||left lower extremitynull|Table Cell Horizontal Align - left|Finding|true|false||leftnull|Left sided|Modifier|true|false||left
null|Left|Modifier|true|false||leftnull|Lower Extremity|Anatomy|true|false||lower extremitynull|Body Site Modifier - Lower|Anatomy|true|false||lowernull|Lower (action)|Event|true|false||lowernull|Lower - spatial qualifier|Modifier|true|false||lowernull|Limb structure|Anatomy|true|false||extremitynull|Structure of right lower leg|Anatomy|true|false||right leg
null|Right lower extremity|Anatomy|true|false||right legnull|Table Cell Horizontal Align - right|Finding|true|false||rightnull|Right sided|Modifier|true|false||right
null|Right|Modifier|true|false||rightnull|Leg|Anatomy|true|false||leg
null|Lower Extremity|Anatomy|true|false||legnull|Initial (abbreviation)|Finding|false|false||initialnull|Initially|Time|false|false||initialnull|Firstly|Modifier|false|false||initialnull|Laboratory test finding|Lab|false|false||Labsnull|Imaging problem|Finding|false|false||imagingnull|Diagnostic Imaging|Procedure|false|false||imaging
null|Imaging Techniques|Procedure|false|false||imagingnull|Imaging Technology|Title|false|false||imagingnull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|Plain chest X-ray|Procedure|false|false||CXRnull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|Moderate - Severity of Illness Code|Finding|false|false||moderate
null|Moderate|Finding|false|false||moderatenull|Moderate (severity modifier)|Modifier|false|false||moderate
null|Moderate - Allergy Severity|Modifier|false|false||moderate
null|Moderation|Modifier|false|false||moderatenull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Pleural Diseases|Disorder|false|false||pleuralnull|Pleura|Anatomy|false|false||pleuralnull|Pleural|Modifier|false|false||pleuralnull|Effusion (substance)|Finding|false|false||effusion
null|null|Finding|false|false||effusion
null|effusion|Finding|false|false||effusionnull|Adjacent|Modifier|false|false||adjacentnull|Atelectasis|Finding|false|false||atelectasisnull|Structure of base of left lung|Anatomy|false|false||left lung basenull|Left lung|Anatomy|false|false||left lungnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Basal segment of lung|Anatomy|false|false||lung basenull|Lung diseases|Disorder|false|false||lungnull|Lung Problem|Finding|false|false||lungnull|Chest>Lung|Anatomy|false|false||lung
null|Lung|Anatomy|false|false||lungnull|nitrogenous base|Drug|false|false||base
null|Base|Drug|false|false||base
null|Dental Base|Drug|false|false||base
null|base - RoleClass|Drug|false|false||basenull|Base - General Qualifier|Finding|false|false||base
null|BPIFA4P gene|Finding|false|false||base
null|Base - RX Component Type|Finding|false|false||basenull|Anatomical base|Anatomy|false|false||basenull|Base - unit of product usage|LabModifier|false|false||basenull|Complete Blood Count|Procedure|false|false||CBCnull|Nuclear cap binding complex location|Anatomy|false|false||CBCnull|null|Finding|false|false||within normal limitsnull|Limited (extensiveness)|Finding|false|false||limitsnull|Electrolytes|Drug|false|false||electrolytes
null|Electrolytes|Drug|false|false||electrolytes
null|Electrolyte [EPC]|Drug|false|false||electrolytesnull|null|Finding|false|false||within normal limitsnull|Limited (extensiveness)|Finding|false|false||limitsnull|Troponin|Drug|false|false||troponin
null|Troponin|Drug|false|false||troponinnull|Troponin measurement|Procedure|false|false||troponinnull|Fibrin fragment D|Drug|false|false||D-dimer
null|Fibrin fragment D|Drug|false|false||D-dimernull|dimer|Drug|false|false||dimernull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Evidence of (contextual qualifier)|Finding|true|false||evidence fornull|Evidence|Finding|true|false||evidencenull|Pulmonary Embolism|Finding|true|false||pulmonary embolusnull|Pulmonary (intended site)|Finding|true|false||pulmonarynull|Lung|Anatomy|true|false||pulmonarynull|null|Attribute|true|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|true|false||pulmonarynull|null|Finding|true|false||embolus
null|Embolus|Finding|true|false||embolusnull|Small|LabModifier|false|false||smallnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Pleural effusion (disorder)|Finding|false|false||pleural effusion
null|Pleural effusion fluid|Finding|false|false||pleural effusion
null|null|Finding|false|false||pleural effusionnull|Pleural Diseases|Disorder|false|false||pleuralnull|Pleura|Anatomy|false|false||pleuralnull|Pleural|Modifier|false|false||pleuralnull|Effusion (substance)|Finding|false|false||effusion
null|null|Finding|false|false||effusion
null|effusion|Finding|false|false||effusionnull|Adjacent|Modifier|false|false||adjacentnull|Atelectasis|Finding|false|false||atelectasisnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|aspirin|Drug|false|false||aspirin
null|aspirin|Drug|false|false||aspirinnull|nitroglycerin|Drug|false|false||nitroglycerin
null|nitroglycerin|Drug|false|false||nitroglycerinnull|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparinnull|Response Modality - Bolus|Finding|false|false||bolus
null|Bolus of ingested food|Finding|false|false||bolusnull|bolus infusion|Procedure|false|false||bolusnull|Bolus Dosing Unit|LabModifier|false|false||bolusnull|Transfer - product ownership|Finding|false|false||transfer
null|Transfer Technique|Finding|false|false||transfer
null|ActClass - transfer|Finding|false|false||transfer
null|null|Finding|false|false||transfernull|Transfer (immobility management)|Procedure|false|false||transfernull|arrival - ActRelationshipType|Finding|false|false||arrivalnull|null|Event|false|false||arrivalnull|Floor (anatomic)|Anatomy|false|false||floornull|floor (object)|Device|false|false||floornull|Floor - story of building|Entity|false|false||floornull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Feeling comfortable|Finding|false|false||comfortablenull|Review of systems (procedure)|Procedure|false|false||REVIEW OF SYSTEMSnull|null|Attribute|false|false||REVIEW OF SYSTEMS
null|null|Attribute|false|false||REVIEW OF SYSTEMSnull|Review of|Finding|false|false||REVIEW OFnull|Review (Publication Type)|Finding|false|false||REVIEW
null|Act Class - review|Finding|false|false||REVIEWnull|System|Finding|false|false||SYSTEMSnull|Review of systems (procedure)|Procedure|false|false||review of systemsnull|null|Attribute|false|false||review of systems
null|null|Attribute|false|false||review of systemsnull|Review of|Finding|false|false||review ofnull|Review (Publication Type)|Finding|false|false||review
null|Act Class - review|Finding|false|false||reviewnull|System|Finding|false|false||systemsnull|null|Time|true|false||priornull|Medical History|Finding|true|false||history ofnull|History of present illness (finding)|Finding|true|false||history
null|History of previous events|Finding|true|false||history
null|Historical aspects qualifier|Finding|true|false||history
null|Medical History|Finding|true|false||history
null|Concept History|Finding|true|false||historynull|History|Subject|true|false||historynull|Cerebrovascular accident|Disorder|true|false||strokenull|Stroke (heart beat)|Finding|true|false||strokenull|Transient Cerebral Ischemia|Disorder|true|false||TIA
null|Transient Ischemic Attack|Disorder|true|false||TIAnull|Tacca leontopetaloides|Entity|true|false||TIAnull|Deep Vein Thrombosis|Disorder|false|false||deep venous thrombosisnull|Deep Resection Margin|Attribute|false|false||deepnull|Deep (qualifier value)|Modifier|false|false||deepnull|Venous thrombosis after immobility|Finding|false|false||venous thrombosis
null|Venous Thrombosis|Finding|false|false||venous thrombosisnull|Veins|Anatomy|false|false||venousnull|Venous|Modifier|false|false||venousnull|Thrombosis|Finding|false|false||thrombosisnull|Pulmonary Embolism|Finding|false|false||pulmonary embolismnull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Embolism|Finding|false|false||embolism
null|Embolus|Finding|false|false||embolismnull|Hemorrhage|Finding|false|false||bleedingnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Myalgia|Finding|false|false||myalgiasnull|Arthralgia|Finding|false|false||joint painsnull|Joint problem|Finding|false|false||jointnull|null|Anatomy|false|false||joint
null|Joints|Anatomy|false|false||joint
null|Articular system|Anatomy|false|false||jointnull|Joint Device|Device|false|false||jointnull|Pain|Finding|false|false||painsnull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|Hemoptysis|Finding|false|false||hemoptysisnull|Black - ethnic group (ethnic group)|Subject|false|false||black
null|Black race|Subject|false|false||black
null|African|Subject|false|false||blacknull|Black - Structured Product Labeling Color|Modifier|false|false||black
null|Black color|Modifier|false|false||blacknull|Feces|Finding|false|false||stoolsnull|null|Attribute|false|false||stoolsnull|Stool seat|Device|false|false||stoolsnull|Red stools|Finding|false|false||red stoolsnull|DYRK3 gene|Finding|false|false||red
null|Redness|Finding|false|false||red
null|IK gene|Finding|false|false||rednull|Radiological Exposure Device|Device|false|false||rednull|Red color|Modifier|false|false||rednull|Feces|Finding|false|false||stoolsnull|null|Attribute|false|false||stoolsnull|Stool seat|Device|false|false||stoolsnull|Recent|Time|true|false||recentnull|Fever|Finding|true|false||feversnull|Chills|Finding|true|false||chillsnull|Rigor - Temperature-associated observation|Finding|true|false||rigorsnull|exercise induced|Finding|true|false||exertionalnull|Buttocks|Anatomy|true|false||buttocknull|Pain in calf|Finding|true|false||calf painnull|Structure of calf of leg|Anatomy|true|false||calf
null|null|Anatomy|true|false||calfnull|Cattle calf (organism)|Entity|true|false||calfnull|Administration Method - Pain|Finding|true|false||pain
null|Pain|Finding|true|false||painnull|null|Attribute|true|false||painnull|Review of systems (procedure)|Procedure|false|false||review of systemsnull|null|Attribute|false|false||review of systems
null|null|Attribute|false|false||review of systemsnull|Review of|Finding|false|false||review ofnull|Review (Publication Type)|Finding|false|false||review
null|Act Class - review|Finding|false|false||reviewnull|System|Finding|false|false||systemsnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|PMH - past medical history|Finding|false|false||Past Medical History
null|Medical History|Finding|false|false||Past Medical Historynull|Medical History|Finding|false|false||Medical Historynull|Medical referral type|Finding|false|false||Medical
null|Medical|Finding|false|false||Medical
null|Medical school type|Finding|false|false||Medicalnull|Medical service|Procedure|false|false||Medicalnull|Medical History|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|History of present illness (finding)|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|cardiac risk factors|Finding|false|false||CARDIAC RISK FACTORSnull|CARD.RISK|Finding|false|false||CARDIAC RISKnull|Cardiac attachment|Finding|false|false||CARDIACnull|Heart|Anatomy|false|false||CARDIACnull|Cardiac - anatomy qualifier|Modifier|false|false||CARDIACnull|risk factors - observation list|Finding|false|false||RISK FACTORS
null|risk factors|Finding|false|false||RISK FACTORS
null|History of - risk factor|Finding|false|false||RISK FACTORSnull|null|Attribute|false|false||RISK FACTORSnull|Risk|Finding|false|false||RISKnull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||Diabetes
null|Diabetes|Disorder|false|false||Diabetes
null|Diabetes Mellitus|Disorder|false|false||Diabetesnull|Dyslipidemias|Disorder|false|false||Dyslipidemianull|Hypertensive disease|Disorder|false|false||HTNnull|Cardiac attachment|Finding|true|false||CARDIACnull|Heart|Anatomy|false|false||CARDIACnull|Cardiac - anatomy qualifier|Modifier|false|false||CARDIACnull|History of present illness (finding)|Finding|false|false||HISTORY
null|History of previous events|Finding|false|false||HISTORY
null|Historical aspects qualifier|Finding|false|false||HISTORY
null|Medical History|Finding|false|false||HISTORY
null|Concept History|Finding|false|false||HISTORYnull|History|Subject|false|false||HISTORYnull|Coronary Artery Disease|Disorder|false|false||Coronary artery disease
null|Coronary Arteriosclerosis|Disorder|false|false||Coronary artery diseasenull|Coronary artery|Anatomy|false|false||Coronary arterynull|Heart|Anatomy|false|false||Coronarynull|Coronary|Modifier|false|false||Coronarynull|Arteriopathic disease|Disorder|false|false||artery diseasenull|Arterial system|Anatomy|false|false||artery
null|Arteries|Anatomy|false|false||arterynull|Disease|Disorder|false|false||diseasenull|diastolic congestive heart failure|Disorder|false|false||Diastolic congestive heart failurenull|Diastole|Attribute|false|false||Diastolicnull|Congestive heart failure|Disorder|false|false||congestive heart failurenull|Congestive|Modifier|false|false||congestivenull|Congestive heart failure|Disorder|false|false||heart failure
null|Heart failure|Disorder|false|false||heart failurenull|Malignant neoplasm of heart|Disorder|false|false||heart
null|benign neoplasm of heart|Disorder|false|false||heartnull|HEART PROBLEM|Finding|false|false||heartnull|Chest>Heart|Anatomy|false|false||heart
null|Heart|Anatomy|false|false||heartnull|Failure (biologic function)|Finding|false|false||failure
null|Failure|Finding|false|false||failure
null|Personal failure|Finding|false|false||failurenull|Coronary Artery Bypass Surgery|Procedure|false|false||CABGnull|Coronary Artery Bypass Surgery|Procedure|false|false||CABGnull|Coronary Artery Bypass, Off-Pump|Procedure|false|false||Off pump coronary artery bypassnull|matrix metalloproteinase 7 activity|Finding|false|false||pumpnull|null|Device|false|false||pumpnull|Pump Dosing Unit|LabModifier|false|false||pumpnull|Coronary Artery Bypass Surgery|Procedure|false|false||coronary artery bypass graftnull|coronary artery graft device|Device|false|false||coronary artery bypass graftnull|Coronary Artery Bypass Surgery|Procedure|false|false||coronary artery bypassnull|Coronary artery|Anatomy|false|false||coronary arterynull|Heart|Anatomy|false|false||coronarynull|Coronary|Modifier|false|false||coronarynull|Arterial bypass graft|Procedure|false|false||artery bypass graftnull|Arterial system|Anatomy|false|false||artery
null|Arteries|Anatomy|false|false||arterynull|Bypass graft|Procedure|false|false||bypass graftnull|Creation of shunt|Procedure|false|false||bypassnull|Graft Dosage Form|Drug|false|false||graft
null|Graft material|Drug|false|false||graftnull|Graft - Specimen Source Codes|Finding|false|false||graftnull|Graft Procedures on the Head|Procedure|false|false||graft
null|Grafting procedure|Procedure|false|false||graftnull|Transplanted tissue|Anatomy|false|false||graftnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Structure of internal thoracic artery|Anatomy|false|false||internal mammary arterynull|Code System Type - Internal|Modifier|false|false||internal
null|Internal Surface|Modifier|false|false||internal
null|Internal|Modifier|false|false||internalnull|Mammary Arteries|Anatomy|false|false||mammary arterynull|Mammary gland|Anatomy|false|false||mammary
null|Breast|Anatomy|false|false||mammarynull|Arterial system|Anatomy|false|false||artery
null|Arteries|Anatomy|false|false||arterynull|Anterior descending branch of left coronary artery|Anatomy|false|false||left anterior descending artery
null|null|Anatomy|false|false||left anterior descending arterynull|Left anterior|Modifier|false|false||left anteriornull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Adenohypophyseal Diseases|Disorder|false|false||anteriornull|Anterior|Modifier|false|false||anteriornull|Sequencing - Descending|Finding|false|false||descendingnull|Descending|Modifier|false|false||descendingnull|Arterial system|Anatomy|false|false||artery
null|Arteries|Anatomy|false|false||arterynull|Great saphenous vein structure|Anatomy|false|false||saphenous vein
null|Saphenous Vein|Anatomy|false|false||saphenous veinnull|Veins|Anatomy|false|false||veinnull|Graft material|Drug|false|false||graftsnull|Transplanted tissue|Anatomy|false|false||graftsnull|grafting qualifier|Modifier|false|false||graftsnull|Diagonal|Modifier|false|false||diagonalnull|Obtuse|Modifier|false|false||obtusenull|Target Awareness - marginal|Finding|false|false||marginalnull|Marginal (quality)|Modifier|false|false||marginal
null|Marginal|Modifier|false|false||marginalnull|Procedure on artery|Procedure|false|false||arteriesnull|Arteries|Anatomy|false|false||arteries
null|Arterial system|Anatomy|false|false||arteriesnull|Percutaneous Coronary Intervention|Procedure|false|false||PERCUTANEOUS CORONARY INTERVENTIONSnull|Percutaneous Route of Drug Administration|Finding|false|false||PERCUTANEOUSnull|Percutaneous|Modifier|false|false||PERCUTANEOUSnull|Heart|Anatomy|false|false||CORONARYnull|Coronary|Modifier|false|false||CORONARYnull|Nursing interventions|Procedure|false|false||INTERVENTIONS
null|Intervention regimes|Procedure|false|false||INTERVENTIONSnull|null|Attribute|false|false||INTERVENTIONSnull|Burning Mouth Syndrome|Disorder|false|false||BMSnull|Proximal Resection Margin|Attribute|false|false||proximalnull|Proximal|Modifier|false|false||proximalnull|Leukocyte adhesion deficiency type 1|Disorder|false|false||LAD
null|Leukocyte adhesion deficiency|Disorder|false|false||LADnull|ITGB2 wt Allele|Finding|false|false||LAD
null|DLD gene|Finding|false|false||LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false||LADnull|Ladino Language|Entity|false|false||LADnull|DES protein, human|Drug|false|false||DES
null|Desmosine|Drug|false|false||DES
null|Desmosine|Drug|false|false||DES
null|DES protein, human|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DESnull|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|Disorder|false|false||DESnull|DES gene|Finding|false|false||DESnull|Middle|Modifier|false|false||midnull|Leukocyte adhesion deficiency type 1|Disorder|false|false||LAD
null|Leukocyte adhesion deficiency|Disorder|false|false||LADnull|ITGB2 wt Allele|Finding|false|false||LAD
null|DLD gene|Finding|false|false||LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false||LADnull|Ladino Language|Entity|false|false||LADnull|DES protein, human|Drug|false|false||DES
null|Desmosine|Drug|false|false||DES
null|Desmosine|Drug|false|false||DES
null|DES protein, human|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DESnull|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|Disorder|false|false||DESnull|DES gene|Finding|false|false||DESnull|Graph Edge|Finding|false|false||edgenull|Along edge (qualifier value)|Modifier|false|false||edgenull|Middle|Modifier|false|false||midnull|Leukocyte adhesion deficiency type 1|Disorder|false|false||LAD
null|Leukocyte adhesion deficiency|Disorder|false|false||LADnull|ITGB2 wt Allele|Finding|false|false||LAD
null|DLD gene|Finding|false|false||LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false||LADnull|Ladino Language|Entity|false|false||LADnull|DES protein, human|Drug|false|false||DES
null|Desmosine|Drug|false|false||DES
null|Desmosine|Drug|false|false||DES
null|DES protein, human|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DESnull|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|Disorder|false|false||DESnull|DES gene|Finding|false|false||DESnull|Stenosis|Finding|false|false||stenosisnull|Stenosis <Pimeliinae>|Entity|false|false||stenosisnull|Stenosis Morphology|Modifier|false|false||stenosisnull|Distal Resection Margin|Attribute|false|false||distalnull|Distal (qualifier value)|Modifier|false|false||distalnull|null|Device|false|false||stentnull|DES protein, human|Drug|false|false||DES
null|Desmosine|Drug|false|false||DES
null|Desmosine|Drug|false|false||DES
null|DES protein, human|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DESnull|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|Disorder|false|false||DESnull|DES gene|Finding|false|false||DESnull|Pacing up and down|Finding|false|false||PACINGnull|Disruptive, Impulse Control, and Conduct Disorders|Disorder|false|false||ICD
null|Type II Mucolipidosis|Disorder|false|false||ICDnull|International Classification of Diseases|Finding|false|false||ICD
null|GNPTAB wt Allele|Finding|false|false||ICDnull|Icd Regimen|Procedure|false|false||ICDnull|between lunch and dinner|Time|false|false||ICDnull|Morbid obesity|Disorder|true|false||Morbid obesitynull|Obesity|Disorder|true|false||obesitynull|BODY MASS INDEX QUANTITATIVE TRAIT LOCUS 20|Finding|true|false||obesitynull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|Gastroesophageal reflux disease|Disorder|false|false||GERDnull|Right tendinous cuff|Anatomy|false|false||Right rotator cuffnull|Table Cell Horizontal Align - right|Finding|false|false||Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|Rotator Cuff Injuries|Disorder|false|false||rotator cuff injurynull|Rotator Cuff|Anatomy|false|false||rotator cuffnull|null|Device|false|false||rotatornull|Cuffing (morphologic abnormality)|Finding|false|false||cuffnull|Cuff - body part|Anatomy|false|false||cuffnull|Cuff Device|Device|false|false||cuffnull|Traumatic AND/OR non-traumatic injury|Disorder|false|false||injury
null|Traumatic injury|Disorder|false|false||injurynull|Bursitis|Disorder|false|false||bursitisnull|Migraine Disorders|Disorder|false|false||Migrainesnull|Cancer patients and suicide and depression|Disorder|false|false||Depression
null|Mental Depression|Disorder|false|false||Depression
null|Depressive disorder|Disorder|false|false||Depression
null|Depressed mood|Disorder|false|false||Depressionnull|Depression - motion|Finding|false|false||Depression
null|null|Finding|false|false||Depressionnull|Depression - recess|Modifier|false|false||Depressionnull|Degenerative polyarthritis|Disorder|false|false||DJDnull|Hemorrhoids|Disorder|false|false||Hemorrhoidsnull|Rosacea|Disorder|false|false||Rosaceanull|Rosacea <Prayinae>|Entity|false|false||Rosaceanull|Social and personal history|Finding|false|false||Social History
null|Social History|Finding|false|false||Social Historynull|Social|Finding|false|false||Socialnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Family Medical History|Finding|false|false||Family Historynull|Entity Name Part Type - family|Finding|false|false||Family
null|Last Name|Finding|false|false||Family
null|Living Arrangement - Family|Finding|false|false||Family
null|Family (taxonomic)|Finding|false|false||Family
null|Family Collection|Finding|false|false||Familynull|Family|Subject|false|false||Familynull|History of present illness (finding)|Finding|false|true||History
null|History of previous events|Finding|false|true||History
null|Historical aspects qualifier|Finding|false|true||History
null|Medical History|Finding|false|true||History
null|Concept History|Finding|false|true||Historynull|History|Subject|false|false||Historynull|Ward (environment)|Device|false|false||wardnull|Ward (person)|Subject|false|false||wardnull|Ward (environment)|Entity|false|false||wardnull|ErbB Receptors|Drug|true|false||her family
null|ErbB Receptors|Drug|true|false||her familynull|ErbB Receptors|Finding|true|false||her familynull|Entity Name Part Type - family|Finding|true|false||family
null|Last Name|Finding|true|false||family
null|Living Arrangement - Family|Finding|true|false||family
null|Family (taxonomic)|Finding|true|false||family
null|Family Collection|Finding|true|false||familynull|Family|Subject|true|false||familynull|physical examination (physical finding)|Finding|false|false||Physical Examnull|Physical Examination|Procedure|false|false||Physical Examnull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||GENERALnull|General medical service|Procedure|false|false||GENERALnull|Generalized|Modifier|false|false||GENERALnull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|Oriented to place|Finding|false|false||Orientednull|Orientation, Spatial|Modifier|false|false||Orientednull|Mood (psychological function)|Finding|false|false||Mood
null|mood (physical finding)|Finding|false|false||Mood
null|Mood (attribute)|Finding|false|false||Moodnull|null|Attribute|false|false||Moodnull|Appropriate|Modifier|false|false||appropriatenull|HEENT|Anatomy|false|false||HEENTnull|Scleral Diseases|Disorder|false|false||Scleranull|examination of sclera|Procedure|false|false||Scleranull|Sclera|Anatomy|false|false||Scleranull|Anicteric|Finding|false|false||anictericnull|Pupil equal round and reacting to light|Finding|false|false||PERRLnull|Malignant neoplasm of conjunctiva|Disorder|true|false||Conjunctiva
null|Benign neoplasm of conjunctiva|Disorder|true|false||Conjunctiva
null|Conjunctival Diseases|Disorder|true|false||Conjunctivanull|Specimen Type - Conjunctiva|Finding|true|false||Conjunctiva
null|null|Finding|true|false||Conjunctivanull|examination of conjunctiva|Procedure|true|false||Conjunctiva
null|Procedure on conjunctiva|Procedure|true|false||Conjunctivanull|Structure of palpebral conjunctiva|Anatomy|true|false||Conjunctiva
null|conjunctiva|Anatomy|true|false||Conjunctivanull|Pink color|Modifier|true|false||pinknull|Pallor of skin|Finding|true|false||pallornull|Cyanosis|Finding|true|false||cyanosisnull|Oral mucous membrane structure|Anatomy|true|false||oral mucosanull|Oral Dosage Form|Drug|true|false||oralnull|Oral Route of Administration|Finding|true|false||oral
null|Oral (intended site)|Finding|true|false||oralnull|Oral cavity|Anatomy|true|false||oralnull|Oral|Modifier|true|false||oralnull|null|Finding|true|false||mucosanull|Mucous Membrane|Anatomy|true|false||mucosanull|Passive joint movement of neck (finding)|Finding|true|false||NECK
null|Neck problem|Finding|true|false||NECKnull|dendritic spine neck|Anatomy|true|false||NECK
null|Neck|Anatomy|true|false||NECKnull|Supple|Finding|true|false||Supplenull|Jugular venous pressure|Finding|true|false||JVPnull|Cardiac attachment|Finding|true|false||CARDIACnull|Heart|Anatomy|true|false||CARDIACnull|Cardiac - anatomy qualifier|Modifier|true|false||CARDIACnull|Point of Maximum Impulse|Finding|true|false||PMI
null|TMEM11 gene|Finding|true|false||PMI
null|PMM2 wt Allele|Finding|true|false||PMI
null|PMM2 gene|Finding|true|false||PMI
null|MPI gene|Finding|true|false||PMInull|Prostate Mechanical Imager|Device|true|false||PMInull|Space of intercostal compartment|Anatomy|false|false||intercostal space
null|Structure of intercostal space|Anatomy|false|false||intercostal spacenull|Intercostal|Modifier|false|false||intercostalnull|Space (Astronomy)|Phenomenon|false|false||spacenull|Space - property|Modifier|false|false||spacenull|Midclavicular|Modifier|false|false||midclavicularnull|Line Specimen|Drug|false|false||line
null|Long Interspersed Elements|Drug|false|false||line
null|Long Interspersed Elements|Drug|false|false||linenull|line source specimen code|Finding|false|false||linenull|Intravascular line|Device|false|false||linenull|Linear|Modifier|false|false||linenull|Line Unit of Length|LabModifier|false|false||linenull|midline cell component|Anatomy|false|false||Midlinenull|Midline (qualifier value)|Modifier|false|false||Midlinenull|Scar Tissue|Finding|false|false||scar
null|Cicatrix|Finding|false|false||scar
null|RPS4X gene|Finding|false|false||scarnull|recent surgery|Finding|false|false||recent surgerynull|Recent|Time|false|false||recentnull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Lung|Anatomy|true|false||LUNGSnull|Deformity of chest wall|Disorder|true|false||chest wall deformitiesnull|Chest wall structure|Anatomy|true|false||chest wall
null|Chest>Chest wall|Anatomy|true|false||chest wallnull|Chest problem|Finding|true|false||chestnull|Chest|Anatomy|true|false||chest
null|Anterior thoracic region|Anatomy|true|false||chestnull|Walls of a building|Device|true|false||wallnull|Congenital Abnormality|Disorder|true|false||deformitiesnull|deformities qualifier|Modifier|true|false||deformitiesnull|Congenital scoliosis|Disorder|true|false||scoliosis
null|null|Disorder|true|false||scoliosis
null|Acquired scoliosis|Disorder|true|false||scoliosisnull|Kyphosis deformity of spine|Disorder|true|false||kyphosis
null|Acquired kyphosis|Disorder|true|false||kyphosis
null|Congenital kyphosis|Disorder|true|false||kyphosisnull|kyphosis|Finding|true|false||kyphosisnull|Respiratory, thoracic and mediastinal disorders|Disorder|true|false||Respnull|Respiratory rate|Attribute|true|false||Respnull|Unlabored|Finding|true|false||unlaborednull|Use of accessory muscles|Finding|true|false||accessory muscle usenull|Accessory skeletal muscle|Disorder|true|false||accessory musclenull|Accessory|Device|true|false||accessorynull|Muscle (organ)|Anatomy|true|false||muscle
null|Muscle Tissue|Anatomy|true|false||musclenull|Use - dosing instruction imperative|Finding|true|false||use
null|utilization qualifier|Finding|true|false||use
null|Usage|Finding|true|false||usenull|cetrimonium bromide|Drug|true|false||CTABnull|Basilar Rales|Finding|true|false||crackles
null|Rales|Finding|true|false||cracklesnull|Wheezing|Finding|true|false||wheezesnull|Rhonchi|Finding|true|false||rhonchinull|Malignant neoplasm of abdomen|Disorder|false|false||ABDOMENnull|Abdomen problem|Finding|false|false||ABDOMENnull|Abdomen|Anatomy|false|false||ABDOMEN
null|Abdominal Cavity|Anatomy|false|false||ABDOMENnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||Softnull|Soft|Modifier|false|false||Softnull|LRRC4B gene|Finding|true|false||HSMnull|Emotional tenderness|Finding|true|false||tenderness
null|Sore to touch|Finding|true|false||tendernessnull|All extremities|Anatomy|true|false||EXTREMITIES
null|Limb structure|Anatomy|true|false||EXTREMITIESnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Intake|Finding|false|false||Intakenull|Measurement of fluid intake|Procedure|false|false||Intake
null|Intake (treatment)|Procedure|false|false||Intakenull|system output|Finding|false|false||Outputnull|Measurement of fluid output|Procedure|false|false||Outputnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||GENERALnull|General medical service|Procedure|false|false||GENERALnull|Generalized|Modifier|false|false||GENERALnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|HEENT|Anatomy|false|false||HEENTnull|PERRLA|Finding|false|false||PERRLAnull|Anicteric|Finding|false|false||anictericnull|dry mucous membranes|Finding|true|false||dry mucous membranesnull|moisture of mucous membranes (physical finding)|Finding|true|false||mucous membranesnull|Mucous Membrane|Anatomy|true|false||mucous membranesnull|Mucus (substance)|Finding|true|false||mucous
null|mucus layer|Finding|true|false||mucousnull|Mucous appearance|Modifier|true|false||mucousnull|Membrane Tissue|Anatomy|true|false||membranesnull|Remote control command - Clear|Finding|true|false||clearnull|Clear|Modifier|true|false||clear
null|Transparent (qualitative concept)|Modifier|true|false||clearnull|Jugular venous pressure|Finding|true|false||JVPnull|Malignant neoplasm of heart|Disorder|true|false||HEART
null|benign neoplasm of heart|Disorder|true|false||HEARTnull|HEART PROBLEM|Finding|true|false||HEARTnull|Chest>Heart|Anatomy|true|false||HEART
null|Heart|Anatomy|true|false||HEARTnull|MAS1L gene|Finding|true|false||MRGnull|Scar Tissue|Finding|false|false||Scar
null|Cicatrix|Finding|false|false||Scar
null|RPS4X gene|Finding|false|false||Scarnull|recent surgery|Finding|false|false||recent surgerynull|Recent|Time|false|false||recentnull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Present|Finding|false|false||present
null|Presentation|Finding|false|false||presentnull|midline cell component|Anatomy|false|false||midlinenull|Midline (qualifier value)|Modifier|false|false||midlinenull|Traumatic Wound|Disorder|true|false||Wound
null|Wounds and Injuries|Disorder|true|false||Wound
null|Traumatic injury|Disorder|true|false||Woundnull|Route of Administration - Wound|Finding|true|false||Wound
null|null|Finding|true|false||Wound
null|Specimen Type - Wound|Finding|true|false||Woundnull|Well (answer to question)|Finding|true|false||wellnull|Well (container)|Device|true|false||wellnull|Microplate Well|Modifier|true|false||well
null|Good|Modifier|true|false||well
null|Healthy|Modifier|true|false||wellnull|Emotional tenderness|Finding|true|false||tenderness
null|Sore to touch|Finding|true|false||tendernessnull|Scar Tissue|Finding|true|false||scar
null|Cicatrix|Finding|true|false||scar
null|RPS4X gene|Finding|true|false||scarnull|Intensity and Distress 1|Finding|false|false||Slightnull|Slight (qualifier value)|Modifier|false|false||Slight
null|Mild (qualifier value)|Modifier|false|false||Slightnull|Erythema|Disorder|false|false||erythemanull|nitrogenous base|Drug|false|false||base
null|Base|Drug|false|false||base
null|Dental Base|Drug|false|false||base
null|base - RoleClass|Drug|false|false||basenull|Base - General Qualifier|Finding|false|false||base
null|BPIFA4P gene|Finding|false|false||base
null|Base - RX Component Type|Finding|false|false||basenull|Anatomical base|Anatomy|false|false||basenull|Base - unit of product usage|LabModifier|false|false||basenull|Academic Research Enhancement Awards|Event|false|false||areanull|Geographic Locations|Entity|false|false||areanull|Area|Modifier|false|false||areanull|Scar Tissue|Finding|false|false||scar
null|Cicatrix|Finding|false|false||scar
null|RPS4X gene|Finding|false|false||scarnull|Present|Finding|false|false||present
null|Presentation|Finding|false|false||presentnull|Act Relationship Subset - previous|Time|false|false||previous
null|Previous|Time|false|false||previousnull|Sterile maggot wound debridement|Procedure|false|false||debridement
null|Debridement|Procedure|false|false||debridementnull|Lung|Anatomy|false|false||LUNGSnull|Basilar Rales|Finding|false|false||crackles
null|Rales|Finding|false|false||cracklesnull|Present|Finding|false|false||present
null|Presentation|Finding|false|false||presentnull|Base|Drug|false|false||basesnull|Base - unit of product usage|LabModifier|false|false||basesnull|Wheezing|Finding|true|false||wheezesnull|Respiration|Finding|false|false||Respirationsnull|Unlabored|Finding|false|false||unlaborednull|Malignant neoplasm of abdomen|Disorder|false|false||ABDOMENnull|Abdomen problem|Finding|false|false||ABDOMENnull|Abdomen|Anatomy|false|false||ABDOMEN
null|Abdominal Cavity|Anatomy|false|false||ABDOMENnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|true|false||softnull|Soft|Modifier|true|false||softnull|LRRC4B gene|Finding|true|false||HSMnull|All extremities|Anatomy|true|false||EXTREMITIES
null|Limb structure|Anatomy|true|false||EXTREMITIESnull|Peripheral pulse|Finding|false|false||peripheral pulsesnull|Peripheral|Modifier|false|false||peripheralnull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false||pulsesnull|Neurology speciality|Title|false|false||NEUROnull|Neurologic (qualifier value)|Modifier|false|false||NEUROnull|Awake (finding)|Finding|false|false||awakenull|Awakening (time frame)|Time|false|false||awakenull|Central Nervous System|Anatomy|false|false||CNsnull|Clinical Nurse Specialists|Subject|false|false||CNsnull|Certified Nurse Specialist|Title|false|false||CNsnull|Staphylococcus, coagulase negative (organism)|Entity|false|false||CNsnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|Laboratory test finding|Lab|false|false||labsnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||HGB
null|Hemoglobin|Drug|false|false||HGBnull|CYGB gene|Finding|false|false||HGBnull|Hemoglobin concentration|Lab|false|false||HGBnull|Hemopoietic stem cell transplant|Procedure|false|false||HCT
null|Hematocrit Measurement|Procedure|false|false||HCTnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Monos|Drug|false|false||MONOS
null|Mono-S|Drug|false|false||MONOS
null|Monos|Drug|false|false||MONOSnull|SARCOIDOSIS, EARLY-ONSET|Disorder|false|false||EOS
null|Familial eosinophilia|Disorder|false|false||EOSnull|PRSS33 gene|Finding|false|false||EOS
null|IKZF4 gene|Finding|false|false||EOSnull|Eos <Loriini>|Entity|false|false||EOSnull|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSEnull|Glucose measurement|Procedure|false|false||GLUCOSEnull|Glucose^1.5H post dose glucagon|Lab|false|false||GLUCOSEnull|urea|Drug|false|false||UREA
null|urea|Drug|false|false||UREA
null|urea|Drug|false|false||UREAnull|Urea measurement|Procedure|false|false||UREAnull|Sodium supplements|Drug|false|false||SODIUM
null|sodium|Drug|false|false||SODIUM
null|sodium|Drug|false|false||SODIUM
null|Sodium Drug Class|Drug|false|false||SODIUMnull|Sodium metabolic function|Finding|false|false||SODIUMnull|Sodium measurement|Procedure|false|false||SODIUMnull|Potassium Drug Class|Drug|false|false||POTASSIUM
null|Dietary Potassium|Drug|false|false||POTASSIUM
null|potassium|Drug|false|false||POTASSIUM
null|potassium|Drug|false|false||POTASSIUM
null|potassium|Drug|false|false||POTASSIUM
null|Potassium supplement|Drug|false|false||POTASSIUM
null|Potassium supplement|Drug|false|false||POTASSIUMnull|Potassium metabolic function|Finding|false|false||POTASSIUMnull|Potassium measurement|Procedure|false|false||POTASSIUMnull|chloride ion|Drug|false|false||CHLORIDE
null|Chlorides|Drug|false|false||CHLORIDEnull|Chloride metabolic function|Finding|false|false||CHLORIDEnull|Chloride measurement|Procedure|false|false||CHLORIDEnull|Total|Modifier|false|false||TOTALnull|carbon dioxide|Drug|false|false||CO2
null|carbon dioxide|Drug|false|false||CO2null|MT-CO2 gene|Finding|false|false||CO2
null|null|Finding|false|false||CO2
null|C2 wt Allele|Finding|false|false||CO2null|blood anion gap (lab test)|Procedure|false|false||ANION GAP
null|Anion gap measurement|Procedure|false|false||ANION GAPnull|Anion Gap|Attribute|false|false||ANION GAPnull|Anion gap result|Lab|false|false||ANION GAPnull|Anions|Drug|false|false||ANIONnull|Ras GTPase-Activating Protein 1, Human|Drug|false|false||GAP
null|Ras GTPase-Activating Protein 1, Human|Drug|false|false||GAP
null|GTPase-Activating Proteins|Drug|false|false||GAP
null|GTPase-Activating Proteins|Drug|false|false||GAPnull|RASA1 wt Allele|Finding|false|false||GAP
null|RASA1 gene|Finding|false|false||GAPnull|Gap (space)|Modifier|false|false||GAPnull|Mandibular right central incisor mesial prosthesis|Device|false|false||25PMnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Creatine Kinase|Drug|false|false||CPK
null|Creatine Kinase|Drug|false|false||CPKnull|PIK3C2A gene|Finding|false|false||CPKnull|Creatine kinase measurement|Procedure|false|false||CPKnull|Fibrin fragment D|Drug|false|false||D-DIMER
null|Fibrin fragment D|Drug|false|false||D-DIMERnull|dimer|Drug|false|false||DIMERnull|Laboratory test finding|Lab|false|false||labsnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MB
null|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MBnull|creatine kinase activity|Finding|false|false||CK-MBnull|Serum creatine phosphokinase MB isoenzyme measurement|Procedure|false|false||CK-MB
null|Creatine kinase MB measurement|Procedure|false|false||CK-MBnull|MB 3|Drug|false|false||MB-3null|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MB
null|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MBnull|creatine kinase activity|Finding|false|false||CK-MBnull|Serum creatine phosphokinase MB isoenzyme measurement|Procedure|false|false||CK-MB
null|Creatine kinase MB measurement|Procedure|false|false||CK-MBnull|MB 3|Drug|false|false||MB-3null|Imaging problem|Finding|false|false||Imagingnull|Diagnostic Imaging|Procedure|false|false||Imaging
null|Imaging Techniques|Procedure|false|false||Imagingnull|Imaging Technology|Title|false|false||Imagingnull|Scientific Study|Procedure|false|false||studiesnull|Electrocardiogram image|Finding|false|false||EKG
null|Electrocardiogram|Finding|false|false||EKGnull|Electrocardiography|Procedure|false|false||EKGnull|On admission|Time|false|false||on admissionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Sinus Tachycardia|Disorder|false|false||Sinus tachycardianull|continuous electrocardiogram sinus tachycardia|Finding|false|false||Sinus tachycardia
null|Sinus Tachycardia by ECG Finding|Finding|false|false||Sinus tachycardianull|Sinus brand of acetaminophen-pseudoephedrine|Drug|false|false||Sinus
null|Sinus brand of acetaminophen-pseudoephedrine|Drug|false|false||Sinusnull|pathologic fistula|Disorder|false|false||Sinusnull|Sinus - general anatomical term|Anatomy|false|false||Sinus
null|Nasal sinus|Anatomy|false|false||Sinusnull|Tachycardia by ECG Finding|Finding|false|false||tachycardia
null|Tachycardia|Finding|false|false||tachycardianull|Extensive|Modifier|false|false||Extensivenull|ST segment|Finding|false|false||ST segmentnull|Anatomical segmentation|Modifier|false|false||segmentnull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|Ischemia|Finding|false|false||ischemianull|Ischemia Procedure|Procedure|false|false||ischemianull|Act Relationship Subset - previous|Time|true|false||previous
null|Previous|Time|true|false||previousnull|Changing|Finding|true|false||changenull|Change - procedure|Procedure|true|false||changenull|Delta (difference)|LabModifier|true|false||change
null|Changed status|LabModifier|true|false||changenull|Plain chest X-ray|Procedure|false|false||CXRnull|Query Status Code - new|Finding|false|false||New
null|Act Status - new|Finding|false|false||Newnull|Newar Language|Entity|false|false||Newnull|New|Modifier|false|false||Newnull|Moderate - Severity of Illness Code|Finding|false|false||moderate
null|Moderate|Finding|false|false||moderatenull|Moderate (severity modifier)|Modifier|false|false||moderate
null|Moderate - Allergy Severity|Modifier|false|false||moderate
null|Moderation|Modifier|false|false||moderatenull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Pleural effusion (disorder)|Finding|false|false||pleural effusion
null|Pleural effusion fluid|Finding|false|false||pleural effusion
null|null|Finding|false|false||pleural effusionnull|Pleural Diseases|Disorder|false|false||pleuralnull|Pleura|Anatomy|false|false||pleuralnull|Pleural|Modifier|false|false||pleuralnull|Effusion (substance)|Finding|false|false||effusion
null|null|Finding|false|false||effusion
null|effusion|Finding|false|false||effusionnull|Adjacent|Modifier|false|false||adjacentnull|Atelectasis|Finding|false|false||atelectasisnull|Structure of base of left lung|Anatomy|false|false||left lung basenull|Left lung|Anatomy|false|false||left lungnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Basal segment of lung|Anatomy|false|false||lung basenull|Lung diseases|Disorder|false|false||lungnull|Lung Problem|Finding|false|false||lungnull|Chest>Lung|Anatomy|false|false||lung
null|Lung|Anatomy|false|false||lungnull|nitrogenous base|Drug|false|false||base
null|Base|Drug|false|false||base
null|Dental Base|Drug|false|false||base
null|base - RoleClass|Drug|false|false||basenull|Base - General Qualifier|Finding|false|false||base
null|BPIFA4P gene|Finding|false|false||base
null|Base - RX Component Type|Finding|false|false||basenull|Anatomical base|Anatomy|false|false||basenull|Base - unit of product usage|LabModifier|false|false||basenull|Cancer/Testis Antigen|Drug|false|false||CTAnull|PCYT1A wt Allele|Finding|false|false||CTA
null|CERNA3 gene|Finding|false|false||CTAnull|Cardiac Computerized Tomographic Angiography|Procedure|false|false||CTAnull|Chest problem|Finding|false|false||Chestnull|Chest|Anatomy|false|false||Chest
null|Anterior thoracic region|Anatomy|false|false||Chestnull|Evidence of (contextual qualifier)|Finding|true|false||evidence fornull|Evidence|Finding|true|false||evidencenull|Pulmonary Embolism|Finding|true|false||pulmonary embolusnull|Pulmonary (intended site)|Finding|true|false||pulmonarynull|Lung|Anatomy|true|false||pulmonarynull|null|Attribute|true|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|true|false||pulmonarynull|null|Finding|true|false||embolus
null|Embolus|Finding|true|false||embolusnull|Small|LabModifier|false|false||Smallnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Pleural effusion (disorder)|Finding|false|false||pleural effusion
null|Pleural effusion fluid|Finding|false|false||pleural effusion
null|null|Finding|false|false||pleural effusionnull|Pleural Diseases|Disorder|false|false||pleuralnull|Pleura|Anatomy|false|false||pleuralnull|Pleural|Modifier|false|false||pleuralnull|Effusion (substance)|Finding|false|false||effusion
null|null|Finding|false|false||effusion
null|effusion|Finding|false|false||effusionnull|Adjacent|Modifier|false|false||adjacentnull|Atelectasis|Finding|false|false||atelectasisnull|Possible|Finding|false|false||Possiblenull|Possible diagnosis|Modifier|false|false||Possible
null|Possibly Related to Intervention|Modifier|false|false||Possiblenull|Calcified (qualifier value)|Modifier|false|false||calcifiednull|Aneurysm of splenic artery|Disorder|false|false||splenic artery aneurysmnull|Structure of splenic artery|Anatomy|false|false||splenic artery
null|Abdomen>Splenic artery|Anatomy|false|false||splenic arterynull|Spleen|Anatomy|false|false||splenicnull|Arterial system|Anatomy|false|false||artery
null|Arteries|Anatomy|false|false||arterynull|Aneurysm|Finding|false|false||aneurysmnull|Protein Domain|Drug|false|false||regionnull|Geographic Locations|Entity|false|false||regionnull|regional|Modifier|false|false||regionnull|Hilum|Anatomy|false|false||hilumnull|Cardiac catheterisation as the cause of abnormal reaction of the patient, or of later complication, without mention of misadventure at the time of the procedure|Disorder|false|false||Cardiac catheterizationnull|Diagnostic Service Section ID - Cardiac Catheterization|Finding|false|false||Cardiac catheterizationnull|Consent Type - Cardiac Catheterization|Procedure|false|false||Cardiac catheterization
null|Cardiac Catheterization Procedures|Procedure|false|false||Cardiac catheterizationnull|Cardiac attachment|Finding|false|false||Cardiacnull|Heart|Anatomy|false|false||Cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||Cardiacnull|Catheterization|Procedure|false|false||catheterizationnull|Consent Type - Coronary Angiography|Procedure|false|false||coronary angiography
null|Coronary angiography|Procedure|false|false||coronary angiographynull|Heart|Anatomy|false|false||coronarynull|Coronary|Modifier|false|false||coronarynull|angiogram|Procedure|false|false||angiographynull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Dominant|Finding|false|false||dominantnull|System (basic dose form)|Drug|false|false||systemnull|System, LOINC Axis 4|Finding|false|false||system
null|System|Finding|false|false||systemnull|Device system|Device|false|false||system
null|System - kit|Device|false|false||systemnull|System (unit of presentation)|LabModifier|false|false||systemnull|Coronary Vessels|Anatomy|false|false||vessel coronarynull|Vessel Positions|Anatomy|false|false||vessel
null|Blood Vessel|Anatomy|false|false||vesselnull|Vessel (unit of presentation)|LabModifier|false|false||vesselnull|Coronary Artery Disease|Disorder|false|false||coronary disease
null|Coronary heart disease|Disorder|false|false||coronary diseasenull|Heart|Anatomy|false|false||coronarynull|Coronary|Modifier|false|false||coronarynull|Disease|Disorder|false|false||diseasenull|Native (qualifier value)|Finding|false|false||nativenull|Blood Vessel|Anatomy|false|false||vesselsnull|apparent|Finding|true|false||apparentnull|Disease|Disorder|true|false||diseasenull|Leukocyte adhesion deficiency type 1|Disorder|false|false||LAD
null|Leukocyte adhesion deficiency|Disorder|false|false||LADnull|ITGB2 wt Allele|Finding|false|false||LAD
null|DLD gene|Finding|false|false||LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false||LADnull|Ladino Language|Entity|false|false||LADnull|Lesion|Finding|false|false||lesion
null|null|Finding|false|false||lesionnull|null|Time|false|false||priornull|null|Device|false|false||stentnull|Small|LabModifier|false|false||smallnull|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group|Finding|false|false||poor
null|Patient Condition Code - Poor|Finding|false|false||poornull|Poverty|Subject|false|false||poornull|Language Proficiency - Poor|Modifier|false|false||poor
null|Specimen Quality - Poor|Modifier|false|false||poor
null|Poor - grade|Modifier|false|false||poor
null|Poor - qualifier|Modifier|false|false||poornull|Flow|Phenomenon|false|false||flownull|Methylcytosine Dioxygenase TET1|Drug|false|false||LCx
null|Methylcytosine Dioxygenase TET1|Drug|false|false||LCxnull|TET1 wt Allele|Finding|false|false||LCx
null|TET1 gene|Finding|false|false||LCxnull|Stenosis|Finding|false|false||stenosisnull|Stenosis <Pimeliinae>|Entity|false|false||stenosisnull|Stenosis Morphology|Modifier|false|false||stenosisnull|Participation Type - origin|Finding|false|false||origin
null|National origin|Finding|false|false||originnull|Beginning|Time|false|false||originnull|apparent|Finding|true|false||apparentnull|Disease|Disorder|true|false||diseasenull|Arteries|Anatomy|false|false||Arterialnull|Arterial|Modifier|false|false||Arterialnull|Conduit implant|Device|false|false||conduitnull|angiogram|Procedure|false|false||angiographynull|Lima|Entity|false|false||LIMAnull|Graft Dosage Form|Drug|false|false||graft
null|Graft material|Drug|false|false||graftnull|Graft - Specimen Source Codes|Finding|false|false||graftnull|Graft Procedures on the Head|Procedure|false|false||graft
null|Grafting procedure|Procedure|false|false||graftnull|Transplanted tissue|Anatomy|false|false||graftnull|Legal patent|Finding|false|false||patentnull|Open|Modifier|false|false||patentnull|Veins|Anatomy|false|false||Venousnull|Venous|Modifier|false|false||Venousnull|Conduit implant|Device|false|false||conduitnull|angiogram|Procedure|false|false||angiographynull|Legal patent|Finding|false|false||patentnull|Open|Modifier|false|false||patentnull|Scalable Vector Graphics|Entity|false|false||SVGnull|Retrograde direction|Modifier|false|false||retrograde
null|Retrograde approach|Modifier|false|false||retrogradenull|Stenosis|Finding|false|false||stenosisnull|Stenosis <Pimeliinae>|Entity|false|false||stenosisnull|Stenosis Morphology|Modifier|false|false||stenosisnull|Small|LabModifier|false|false||smallnull|Scalable Vector Graphics|Entity|false|false||SVGnull|Small|LabModifier|false|false||smallnull|Diagonal|Modifier|false|false||diagonalnull|Occluded|Finding|false|false||occluded
null|Obstruction|Finding|false|false||occludednull|Unable|Finding|false|false||unablenull|Limited component (foundation metadata concept)|Finding|false|false||Limited
null|Limited (extensiveness)|Finding|false|false||Limitednull|Hemodynamics|Finding|false|false||hemodynamicsnull|hemodynamics (procedure)|Procedure|false|false||hemodynamicsnull|Hypertensive disease|Disorder|false|false||systemic hypertensionnull|Systemic Route of Administration|Finding|false|false||systemic
null|Systemic|Finding|false|false||systemicnull|Hypertensive disease|Disorder|false|false||hypertensionnull|Aortic Pressure|Lab|false|false||aortic pressurenull|Aorta|Anatomy|false|false||aorticnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|mmHg|LabModifier|false|false||mm Hgnull|Final diagnosis (discharge)|Modifier|false|false||FINAL DIAGNOSISnull|Diagnosis Type - Final|Finding|false|false||FINALnull|Final|Time|false|false||FINALnull|End-stage|Modifier|false|false||FINALnull|Diagnosis Classification - Diagnosis|Finding|false|false||DIAGNOSIS
null|diagnosis aspects|Finding|false|false||DIAGNOSISnull|Diagnosis|Procedure|false|false||DIAGNOSISnull|null|Attribute|false|false||DIAGNOSISnull|Coronary Vessels|Anatomy|false|false||vessel coronarynull|Vessel Positions|Anatomy|false|false||vessel
null|Blood Vessel|Anatomy|false|false||vesselnull|Vessel (unit of presentation)|LabModifier|false|false||vesselnull|Coronary Artery Disease|Disorder|false|false||coronary artery disease
null|Coronary Arteriosclerosis|Disorder|false|false||coronary artery diseasenull|Coronary artery|Anatomy|false|false||coronary arterynull|Heart|Anatomy|false|false||coronarynull|Coronary|Modifier|false|false||coronarynull|Arteriopathic disease|Disorder|false|false||artery diseasenull|Arteries|Anatomy|false|false||artery
null|Arterial system|Anatomy|false|false||arterynull|Disease|Disorder|false|false||diseasenull|Native (qualifier value)|Finding|false|false||nativenull|Procedure on artery|Procedure|false|false||arteriesnull|Arteries|Anatomy|false|false||arteries
null|Arterial system|Anatomy|false|false||arteriesnull|Legal patent|Finding|false|false||Patentnull|Open|Modifier|false|false||Patentnull|Lima|Entity|false|false||LIMAnull|Leukocyte adhesion deficiency type 1|Disorder|false|false||LAD
null|Leukocyte adhesion deficiency|Disorder|false|false||LADnull|ITGB2 wt Allele|Finding|false|false||LAD
null|DLD gene|Finding|false|false||LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false||LADnull|Ladino Language|Entity|false|false||LADnull|Legal patent|Finding|false|false||patentnull|Open|Modifier|false|false||patentnull|Scalable Vector Graphics|Entity|false|false||SVGnull|Occluded|Finding|false|false||occluded
null|Obstruction|Finding|false|false||occludednull|Scalable Vector Graphics|Entity|false|false||SVGnull|Small|LabModifier|false|false||smallnull|Diagonal|Modifier|false|false||diagonalnull|Macromolecular Branch|Drug|false|false||branchnull|Branch of|Modifier|false|false||branchnull|BRIEF Health Literacy Screening Tool|Finding|false|false||Brief
null|Behavior Rating Inventory of Executive Function|Finding|false|false||Briefnull|Brief|Time|false|false||Briefnull|Shortened|Modifier|false|false||Briefnull|Hospital course|Finding|false|false||Hospital Coursenull|null|Attribute|false|false||Hospital Coursenull|Organization unit type - Hospital|Finding|false|false||Hospitalnull|Hospitals|Device|false|false||Hospitalnull|Hospitals|Entity|false|false||Hospitalnull|Hospital environment|Modifier|false|false||Hospitalnull|Course|Time|false|false||Coursenull|Transaction counts and value totals - year|Finding|false|false||year
null|Precision - year|Finding|false|false||yearnull|year|Time|false|false||yearnull|Old|Time|false|false||oldnull|Females|Subject|false|false||female
null|Woman|Subject|false|false||femalenull|Female, Self-Report|Modifier|false|false||female
null|Female Phenotype|Modifier|false|false||femalenull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|SERPINA5 protein, human|Drug|false|false||PCI
null|SERPINA5 protein, human|Drug|false|false||PCInull|Peritoneal Cancer Index|Finding|false|false||PCI
null|SERPINA5 wt Allele|Finding|false|false||PCI
null|SERPINA5 gene|Finding|false|false||PCInull|Percutaneous Coronary Intervention|Procedure|false|false||PCI
null|photochemical internalization|Procedure|false|false||PCI
null|Prophylactic Cranial Irradiation|Procedure|false|false||PCInull|Picocurie|LabModifier|false|false||PCInull|Coronary Artery Bypass Surgery|Procedure|false|false||CABGnull|Type 2|Finding|false|false||type 2null|Type - ParameterizedDataType|Finding|false|false||type
null|SGCG gene|Finding|false|false||typenull|null|Modifier|false|false||typenull|insulin, regular, human|Drug|false|false||insulin
null|Insulin [EPC]|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulinnull|INS gene|Finding|false|false||insulinnull|Insulin measurement|Procedure|false|false||insulinnull|Hypertensive disease|Disorder|false|false||HTNnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Left sided chest pain|Finding|false|false||left sided chest painnull|Left sided|Modifier|false|false||left sided
null|Left|Modifier|false|false||left sidednull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Chest Pain|Finding|false|false||chest painnull|null|Attribute|false|false||chest painnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Dyspnea|Finding|false|false||SOBnull|Chest Pain|Finding|false|false||Chest Painnull|null|Attribute|false|false||Chest Painnull|Chest problem|Finding|false|false||Chestnull|Chest|Anatomy|false|false||Chest
null|Anterior thoracic region|Anatomy|false|false||Chestnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Recent|Time|false|false||recentnull|Coronary Artery Bypass Surgery|Procedure|false|false||CABGnull|Chest Pain|Finding|false|false||chest painnull|null|Attribute|false|false||chest painnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Troponin|Drug|false|false||troponins
null|Troponin|Drug|false|false||troponinsnull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|Mental Depression|Disorder|false|false||depressionsnull|Consistent with|Finding|false|false||consistent withnull|Compatible|Modifier|false|false||consistent withnull|Consistent with|Finding|false|false||consistentnull|null|Disorder|false|false||NSTEMInull|null|Finding|false|false||NSTEMInull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Troponin|Drug|false|false||troponins
null|Troponin|Drug|false|false||troponinsnull|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparinnull|Drops - Drug Form|Drug|false|false||gttnull|Gestational Trophoblastic Neoplasms|Disorder|false|false||gttnull|Glucose tolerance test|Procedure|false|false||gttnull|Drop Dosing Unit|LabModifier|false|false||gtt
null|Medical Drop|LabModifier|false|false||gttnull|Cardiac Catheterization Procedures|Procedure|false|false||cardiac cathnull|Cardiac attachment|Finding|false|false||cardiacnull|Heart|Anatomy|false|false||cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||cardiacnull|Catheterization|Procedure|false|false||cathnull|Morning|Time|false|false||morningnull|Catheterization|Procedure|false|false||Catheterizationnull|Complete obstruction|Disorder|false|false||occlusionnull|Cardiovascular occlusion|Finding|false|false||occlusion
null|Occluded|Finding|false|false||occlusion
null|Dental Occlusion|Finding|false|false||occlusion
null|Obstruction|Finding|false|false||occlusion
null|null|Finding|false|false||occlusionnull|Scalable Vector Graphics|Entity|false|false||SVGnull|Diagonal|Modifier|false|false||diagonalnull|Possible|Finding|false|false||possiblynull|Possible diagnosis|Modifier|false|false||possiblynull|Electrical Current|Phenomenon|false|false||currentnull|Current (present time)|Time|false|false||currentnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Intervention regimes|Procedure|true|false||intervention
null|Nursing interventions|Procedure|true|false||intervention
null|Interventional procedure|Procedure|true|false||interventionnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|metoprolol|Drug|false|false||metoprolol
null|metoprolol|Drug|false|false||metoprololnull|Transcription Initiation|Finding|false|false||initiation
null|Initiation|Finding|false|false||initiation
null|null|Finding|false|false||initiationnull|AOD use initiation|Time|false|false||initiationnull|losartan|Drug|false|false||losartan
null|losartan|Drug|false|false||losartannull|Transcription Initiation|Finding|false|false||initiation
null|Initiation|Finding|false|false||initiation
null|null|Finding|false|false||initiationnull|AOD use initiation|Time|false|false||initiationnull|Imdur|Drug|false|false||imdur
null|Imdur|Drug|false|false||imdurnull|Potential|Modifier|false|false||potentialnull|Etiology aspects|Finding|false|false||causes
null|Etiology|Finding|false|false||causesnull|Chest Pain|Finding|false|false||chest painnull|null|Attribute|false|false||chest painnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Rh Negative Blood Group|Finding|true|false||negative
null|Negative|Finding|true|false||negative
null|Negative Finding|Finding|true|false||negativenull|Expression Negative|Lab|true|false||negativenull|Negative - qualifier|Modifier|true|false||negative
null|Negative Charge|Modifier|true|false||negativenull|Negative Number|LabModifier|true|false||negativenull|Cancer/Testis Antigen|Drug|true|false||CTAnull|PCYT1A wt Allele|Finding|true|false||CTA
null|CERNA3 gene|Finding|true|false||CTAnull|Cardiac Computerized Tomographic Angiography|Procedure|true|false||CTAnull|Pericarditis|Disorder|false|false||pericarditisnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Consistent with|Finding|false|false||consistentnull|Exam|Finding|true|false||examnull|Medical Examination|Procedure|true|false||examnull|Electrocardiogram image|Finding|true|false||EKG
null|Electrocardiogram|Finding|true|false||EKGnull|Electrocardiography|Procedure|true|false||EKGnull|Consistent with|Finding|true|false||consistentnull|Has patient|Finding|true|false||patient hasnull|Relationship modifier - Patient|Finding|true|false||patient
null|Specimen Type - Patient|Finding|true|false||patient
null|Mail Claim Party - Patient|Finding|true|false||patient
null|Report source - Patient|Finding|true|false||patient
null|null|Finding|true|false||patient
null|Disabled Person Code - Patient|Finding|true|false||patientnull|Patients|Subject|true|false||patientnull|Veterinary Patient|Entity|true|false||patientnull|Consistent with|Finding|false|false||consistentnull|Analgesics and non-steroidal anti-inflammatory drugs|Drug|false|false||NSAIDs
null|Anti-Inflammatory Agents, Non-Steroidal|Drug|false|false||NSAIDsnull|Tietze's Syndrome|Disorder|false|false||costochondritis
null|Costal chondritis|Disorder|false|false||costochondritisnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Pleurisy|Disorder|false|false||pleuritisnull|Secondary to|Modifier|false|false||secondary tonull|Neoplasm Metastasis|Disorder|false|false||secondarynull|metastatic qualifier|Finding|false|false||secondarynull|Secondary to|Modifier|false|false||secondarynull|second (number)|LabModifier|false|false||secondarynull|Pleural effusion (disorder)|Finding|false|false||pleural effusion
null|Pleural effusion fluid|Finding|false|false||pleural effusion
null|null|Finding|false|false||pleural effusionnull|Pleural Diseases|Disorder|false|false||pleuralnull|Pleura|Anatomy|false|false||pleuralnull|Pleural|Modifier|false|false||pleuralnull|Effusion (substance)|Finding|false|false||effusion
null|null|Finding|false|false||effusion
null|effusion|Finding|false|false||effusionnull|Very|Modifier|false|false||verynull|Small|LabModifier|false|false||smallnull|Effusion (substance)|Finding|false|false||effusion
null|null|Finding|false|false||effusion
null|effusion|Finding|false|false||effusionnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Coronary Artery Bypass Surgery|Procedure|false|false||CABGnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Cardiologists|Subject|false|false||cardiologistnull|Imdur|Drug|false|false||imdur
null|Imdur|Drug|false|false||imdurnull|Blood pressure finding|Finding|false|false||blood pressure
null|Systemic arterial pressure|Finding|false|false||blood pressure
null|Blood Pressure|Finding|false|false||blood pressurenull|Blood pressure determination|Procedure|false|false||blood pressurenull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|Acute Kidney Insufficiency|Disorder|false|false||Acute renal insufficiency
null|Kidney Failure, Acute|Disorder|false|false||Acute renal insufficiencynull|Admission Level of Care Code - Acute|Finding|false|false||Acute
null|Acute - Triage Code|Finding|false|false||Acutenull|acute|Time|false|false||Acutenull|Renal Insufficiency|Disorder|false|false||renal insufficiency
null|Kidney Failure|Disorder|false|false||renal insufficiencynull|Urologic Diseases|Disorder|false|false||renalnull|Kidney|Anatomy|false|false||renalnull|Insufficiency|Finding|false|false||insufficiencynull|On admission|Time|false|false||On admissionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Creatinine increased|Finding|false|false||creatinine elevatednull|creatinine|Drug|false|false||creatinine
null|creatinine|Drug|false|false||creatininenull|Creatinine metabolic function|Finding|false|false||creatininenull|Creatinine measurement|Procedure|false|false||creatininenull|Elevated|Modifier|false|false||elevated
null|High|Modifier|false|false||elevatednull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|dehydration (Na, H2O)|Disorder|false|false||dehydration
null|Dehydration|Disorder|false|false||dehydrationnull|Dehydration procedure|Procedure|false|false||dehydrationnull|creatinine|Drug|false|false||creatinine
null|creatinine|Drug|false|false||creatininenull|Creatinine metabolic function|Finding|false|false||creatininenull|Creatinine measurement|Procedure|false|false||creatininenull|Overnight|Time|false|false||overnightnull|Gentle|Drug|false|false||gentle
null|Gentle|Drug|false|false||gentlenull|Liquid substance|Drug|false|false||fluidsnull|Mouse Body Fluid or Substance|Finding|false|false||fluidsnull|Fluid Therapy|Procedure|false|false||fluidsnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Inhaler|Device|false|false||inhalersnull|albuterol|Drug|false|false||albuterol
null|albuterol|Drug|false|false||albuterolnull|fluticasone|Drug|false|false||fluticasone
null|fluticasone|Drug|false|false||fluticasonenull|insulin glargine|Drug|false|false||glargine
null|insulin glargine|Drug|false|false||glargine
null|insulin glargine|Drug|false|false||glarginenull|Unit - NCI Thesaurus Property|LabModifier|false|false||units
null|Unit of Measure|LabModifier|false|false||units
null|Unit|LabModifier|false|false||unitsnull|SHORT STATURE, IDIOPATHIC, X-LINKED|Disorder|false|false||ISSnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|atorvastatin|Drug|false|false||atorvastatin
null|atorvastatin|Drug|false|false||atorvastatinnull|Gastroesophageal reflux disease|Disorder|false|false||GERDnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|pantoprazole|Drug|false|false||pantoprazole
null|pantoprazole|Drug|false|false||pantoprazolenull|Marketing basis - Transitional|Finding|false|false||Transitionalnull|Transitional cell morphology|Modifier|false|false||Transitionalnull|New medications|Drug|false|false||NEW MEDICATIONSnull|Query Status Code - new|Finding|false|false||NEW
null|Act Status - new|Finding|false|false||NEWnull|Newar Language|Entity|false|false||NEWnull|New|Modifier|false|false||NEWnull|Pharmaceutical Preparations|Drug|false|false||MEDICATIONSnull|Medications|Finding|false|false||MEDICATIONSnull|null|Attribute|false|false||MEDICATIONS
null|null|Attribute|false|false||MEDICATIONSnull|losartan|Drug|false|false||losartan
null|losartan|Drug|false|false||losartannull|Imdur|Drug|false|false||imdur
null|Imdur|Drug|false|false||imdurnull|Pharmaceutical Preparations|Drug|false|false||MEDICATIONnull|medication - HL7 publishing domain|Finding|false|false||MEDICATION
null|Medications|Finding|false|false||MEDICATIONnull|Changing|Finding|false|false||CHANGESnull|Changed status|LabModifier|false|false||CHANGESnull|metoprolol|Drug|false|false||metoprolol
null|metoprolol|Drug|false|false||metoprololnull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|Continuous|Finding|false|false||ongoingnull|Chest Pain|Finding|false|false||chest painnull|null|Attribute|false|false||chest painnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Imdur|Drug|false|false||imdur
null|Imdur|Drug|false|false||imdurnull|Angina Pectoris|Finding|false|false||anginal painnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Tietze's Syndrome|Disorder|false|false||costochondritis
null|Costal chondritis|Disorder|false|false||costochondritisnull|Pericarditis|Disorder|false|false||pericarditisnull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|MEDICATION LIST|Finding|false|false||Medication listnull|Pharmaceutical Preparations|Drug|false|false||Medicationnull|medication - HL7 publishing domain|Finding|false|false||Medication
null|Medications|Finding|false|false||Medicationnull|List|Finding|false|false||list
null|Sequence Data Type|Finding|false|false||listnull|Accurate (qualifier value)|Modifier|false|false||accuratenull|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||completenull|Completion Status for valid values - Complete|Finding|false|false||complete
null|Data operation - complete|Finding|false|false||complete
null|Finish - dosing instruction imperative|Finding|false|false||completenull|Complete|Modifier|false|false||completenull|albuterol|Drug|false|false||Albuterol
null|albuterol|Drug|false|false||Albuterolnull|Inhaler (unit of presentation)|Finding|false|false||Inhalernull|Inhaler|Device|false|false||Inhalernull|Inhaler Dosing Unit|LabModifier|false|false||Inhalernull|Puff Dosing Unit|LabModifier|false|false||PUFF
null|Picofarad|LabModifier|false|false||PUFFnull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Dyspnea|Finding|false|false||SOBnull|atorvastatin|Drug|false|false||Atorvastatin
null|atorvastatin|Drug|false|false||Atorvastatinnull|Daily|Time|false|false||DAILYnull|clopidogrel|Drug|false|false||Clopidogrel
null|clopidogrel|Drug|false|false||Clopidogrelnull|Daily|Time|false|false||DAILYnull|fluticasone propionate|Drug|false|false||Fluticasone Propionate
null|fluticasone propionate|Drug|false|false||Fluticasone Propionatenull|fluticasone|Drug|false|false||Fluticasone
null|fluticasone|Drug|false|false||Fluticasonenull|propionate|Drug|false|false||Propionate
null|Propionates|Drug|false|false||Propionatenull|Puff Dosing Unit|LabModifier|false|false||PUFF
null|Picofarad|LabModifier|false|false||PUFFnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|insulin glargine|Drug|false|false||Glargine
null|insulin glargine|Drug|false|false||Glargine
null|insulin glargine|Drug|false|false||Glarginenull|Unit - NCI Thesaurus Property|LabModifier|false|false||Units
null|Unit of Measure|LabModifier|false|false||Units
null|Unit|LabModifier|false|false||Unitsnull|Bedtime (qualifier value)|Time|false|false||Bedtime
null|Once a day, at bedtime|Time|false|false||Bedtimenull|insulin, regular, human|Drug|false|false||Insulin
null|Insulin [EPC]|Drug|false|false||Insulin
null|INS protein, human|Drug|false|false||Insulin
null|INS protein, human|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Insulin Drug Class|Drug|false|false||Insulin
null|Insulin Drug Class|Drug|false|false||Insulin
null|insulin, regular, human|Drug|false|false||Insulin
null|insulin, regular, human|Drug|false|false||Insulinnull|INS gene|Finding|false|false||Insulinnull|Insulin measurement|Procedure|false|false||Insulinnull|sliding scale|Procedure|false|false||Sliding Scalenull|Sliding|Finding|false|false||Slidingnull|Scale, LOINC Axis 5|Finding|false|false||Scale
null|Base Number|Finding|false|false||Scale
null|Scale - rank|Finding|false|false||Scalenull|Integumentary scale|Anatomy|false|false||Scalenull|Weight measurement scales|Device|false|false||Scalenull|Scaling|Event|false|false||Scalenull|insulin, regular, human|Drug|false|false||Insulin
null|Insulin [EPC]|Drug|false|false||Insulin
null|INS protein, human|Drug|false|false||Insulin
null|INS protein, human|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Insulin Drug Class|Drug|false|false||Insulin
null|Insulin Drug Class|Drug|false|false||Insulin
null|insulin, regular, human|Drug|false|false||Insulin
null|insulin, regular, human|Drug|false|false||Insulinnull|INS gene|Finding|false|false||Insulinnull|Insulin measurement|Procedure|false|false||Insulinnull|metoprolol tartrate|Drug|false|false||Metoprolol Tartrate
null|metoprolol tartrate|Drug|false|false||Metoprolol Tartratenull|metoprolol|Drug|false|false||Metoprolol
null|metoprolol|Drug|false|false||Metoprololnull|tartrate|Drug|false|false||Tartrate
null|Tartrates|Drug|false|false||Tartrate
null|tartrate|Drug|false|false||Tartratenull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|Hold - dosing instruction fragment|Finding|false|false||Hold
null|hold - Data Operation|Finding|false|false||Holdnull|Hold (action)|Event|false|false||Holdnull|Androgen Binding Protein|Drug|false|false||SBP
null|Androgen Binding Protein|Drug|false|false||SBPnull|CCHCR1 wt Allele|Finding|false|false||SBP
null|SHBG wt Allele|Finding|false|false||SBPnull|Systolic blood pressure measurement|Procedure|false|false||SBPnull|Systolic Pressure|Attribute|false|false||SBPnull|MetroGel|Drug|false|false||Metrogel
null|MetroGel|Drug|false|false||Metrogelnull|metronidazole|Drug|false|false||metroNIDAZOLE
null|metronidazole|Drug|false|false||metroNIDAZOLEnull|Topical Dosage Form|Drug|false|false||Topicalnull|Topical Route of Administration|Finding|false|false||Topicalnull|Topical surface|Modifier|false|false||Topicalnull|Daily|Time|false|false||Dailynull|acetaminophen / oxycodone|Drug|false|false||Oxycodone-Acetaminophennull|oxycodone|Drug|false|false||Oxycodone
null|oxycodone|Drug|false|false||Oxycodonenull|Oxycodone measurement|Procedure|false|false||Oxycodonenull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Tablet Dosage Form|Drug|false|false||TABnull|Tablet Dosing Unit|LabModifier|false|false||TABnull|Every eight hours|Time|false|false||Q8Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|pantoprazole|Drug|false|false||Pantoprazole
null|pantoprazole|Drug|false|false||Pantoprazolenull|Every twenty four hours|Time|false|false||Q24Hnull|ropinirole|Drug|false|false||Ropinirole
null|ropinirole|Drug|false|false||Ropinirolenull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|aspirin|Drug|false|false||Aspirin
null|aspirin|Drug|false|false||Aspirinnull|Daily|Time|false|false||DAILYnull|Vitamin D Drug Class|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|D Vitamin|Drug|false|false||Vitamin D
null|Vitamin D [EPC]|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|Vitamin D Drug Class|Drug|false|false||Vitamin Dnull|Vitamin D measurement|Procedure|false|false||Vitamin Dnull|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitaminnull|Storage Unit|Device|false|false||UNIT
null|Unit device|Device|false|false||UNITnull|Unit - NCI Thesaurus Property|LabModifier|false|false||UNIT
null|Unit of Measure|LabModifier|false|false||UNIT
null|Unit|LabModifier|false|false||UNIT
null|Enzyme Unit|LabModifier|false|false||UNITnull|Daily|Time|false|false||DAILYnull|ibuprofen|Drug|false|false||Ibuprofen
null|ibuprofen|Drug|false|false||Ibuprofennull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|albuterol|Drug|false|false||Albuterol
null|albuterol|Drug|false|false||Albuterolnull|Inhaler (unit of presentation)|Finding|false|false||Inhalernull|Inhaler|Device|false|false||Inhalernull|Inhaler Dosing Unit|LabModifier|false|false||Inhalernull|Puff Dosing Unit|LabModifier|false|false||PUFF
null|Picofarad|LabModifier|false|false||PUFFnull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Dyspnea|Finding|false|false||SOBnull|aspirin|Drug|false|false||Aspirin
null|aspirin|Drug|false|false||Aspirinnull|Daily|Time|false|false||DAILYnull|aspirin|Drug|false|false||aspirin
null|aspirin|Drug|false|false||aspirinnull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Daily|Time|false|false||dailynull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|atorvastatin|Drug|false|false||Atorvastatin
null|atorvastatin|Drug|false|false||Atorvastatinnull|Daily|Time|false|false||DAILYnull|atorvastatin|Drug|false|false||atorvastatin
null|atorvastatin|Drug|false|false||atorvastatinnull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Daily|Time|false|false||dailynull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|insulin glargine|Drug|false|false||Glargine
null|insulin glargine|Drug|false|false||Glargine
null|insulin glargine|Drug|false|false||Glarginenull|Unit - NCI Thesaurus Property|LabModifier|false|false||Units
null|Unit of Measure|LabModifier|false|false||Units
null|Unit|LabModifier|false|false||Unitsnull|Bedtime (qualifier value)|Time|false|false||Bedtime
null|Once a day, at bedtime|Time|false|false||Bedtimenull|insulin, regular, human|Drug|false|false||Insulin
null|Insulin [EPC]|Drug|false|false||Insulin
null|INS protein, human|Drug|false|false||Insulin
null|INS protein, human|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Insulin Drug Class|Drug|false|false||Insulin
null|Insulin Drug Class|Drug|false|false||Insulin
null|insulin, regular, human|Drug|false|false||Insulin
null|insulin, regular, human|Drug|false|false||Insulinnull|INS gene|Finding|false|false||Insulinnull|Insulin measurement|Procedure|false|false||Insulinnull|sliding scale|Procedure|false|false||Sliding Scalenull|Sliding|Finding|false|false||Slidingnull|Scale, LOINC Axis 5|Finding|false|false||Scale
null|Base Number|Finding|false|false||Scale
null|Scale - rank|Finding|false|false||Scalenull|Integumentary scale|Anatomy|false|false||Scalenull|Weight measurement scales|Device|false|false||Scalenull|Scaling|Event|false|false||Scalenull|insulin, regular, human|Drug|false|false||Insulin
null|Insulin [EPC]|Drug|false|false||Insulin
null|INS protein, human|Drug|false|false||Insulin
null|INS protein, human|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Insulin Drug Class|Drug|false|false||Insulin
null|Insulin Drug Class|Drug|false|false||Insulin
null|insulin, regular, human|Drug|false|false||Insulin
null|insulin, regular, human|Drug|false|false||Insulinnull|INS gene|Finding|false|false||Insulinnull|Insulin measurement|Procedure|false|false||Insulinnull|metoprolol tartrate|Drug|false|false||Metoprolol Tartrate
null|metoprolol tartrate|Drug|false|false||Metoprolol Tartratenull|metoprolol|Drug|false|false||Metoprolol
null|metoprolol|Drug|false|false||Metoprololnull|tartrate|Drug|false|false||Tartrate
null|Tartrates|Drug|false|false||Tartrate
null|tartrate|Drug|false|false||Tartratenull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|metoprolol tartrate|Drug|false|false||metoprolol tartrate
null|metoprolol tartrate|Drug|false|false||metoprolol tartratenull|metoprolol|Drug|false|false||metoprolol
null|metoprolol|Drug|false|false||metoprololnull|tartrate|Drug|false|false||tartrate
null|Tartrates|Drug|false|false||tartrate
null|tartrate|Drug|false|false||tartratenull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Thrice|LabModifier|false|false||three timesnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|pantoprazole|Drug|false|false||Pantoprazole
null|pantoprazole|Drug|false|false||Pantoprazolenull|Every twenty four hours|Time|false|false||Q24Hnull|pantoprazole|Drug|false|false||pantoprazole
null|pantoprazole|Drug|false|false||pantoprazolenull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Daily|Time|false|false||dailynull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|ropinirole|Drug|false|false||Ropinirole
null|ropinirole|Drug|false|false||Ropinirolenull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|Vitamin D Drug Class|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|D Vitamin|Drug|false|false||Vitamin D
null|Vitamin D [EPC]|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|Vitamin D Drug Class|Drug|false|false||Vitamin Dnull|Vitamin D measurement|Procedure|false|false||Vitamin Dnull|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitaminnull|Storage Unit|Device|false|false||UNIT
null|Unit device|Device|false|false||UNITnull|Unit - NCI Thesaurus Property|LabModifier|false|false||UNIT
null|Unit of Measure|LabModifier|false|false||UNIT
null|Unit|LabModifier|false|false||UNIT
null|Enzyme Unit|LabModifier|false|false||UNITnull|Daily|Time|false|false||DAILYnull|isosorbide mononitrate|Drug|false|false||Isosorbide Mononitrate
null|isosorbide mononitrate|Drug|false|false||Isosorbide Mononitratenull|isosorbide|Drug|false|false||Isosorbide
null|isosorbide|Drug|false|false||Isosorbidenull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Daily|Time|false|false||DAILYnull|isosorbide mononitrate|Drug|false|false||isosorbide mononitrate
null|isosorbide mononitrate|Drug|false|false||isosorbide mononitratenull|isosorbide|Drug|false|false||isosorbide
null|isosorbide|Drug|false|false||isosorbidenull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Daily|Time|false|false||dailynull|PRSS30P gene|Finding|false|false||Dispnull|Dispense (activity)|Event|false|false||Dispnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|MetroGel|Drug|false|false||Metrogel
null|MetroGel|Drug|false|false||Metrogelnull|metronidazole|Drug|false|false||metroNIDAZOLE
null|metronidazole|Drug|false|false||metroNIDAZOLEnull|Topical Dosage Form|Drug|false|false||Topicalnull|Topical Route of Administration|Finding|false|false||Topicalnull|Topical surface|Modifier|false|false||Topicalnull|Daily|Time|false|false||Dailynull|acetaminophen / oxycodone|Drug|false|false||Oxycodone-Acetaminophennull|oxycodone|Drug|false|false||Oxycodone
null|oxycodone|Drug|false|false||Oxycodonenull|Oxycodone measurement|Procedure|false|false||Oxycodonenull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Tablet Dosage Form|Drug|false|false||TABnull|Tablet Dosing Unit|LabModifier|false|false||TABnull|Every eight hours|Time|false|false||Q8Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|losartan potassium|Drug|false|false||Losartan Potassium
null|losartan potassium|Drug|false|false||Losartan Potassiumnull|losartan|Drug|false|false||Losartan
null|losartan|Drug|false|false||Losartannull|Potassium Drug Class|Drug|false|false||Potassium
null|Dietary Potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassiumnull|Potassium metabolic function|Finding|false|false||Potassiumnull|Potassium measurement|Procedure|false|false||Potassiumnull|Daily|Time|false|false||DAILYnull|losartan|Drug|false|false||losartan
null|losartan|Drug|false|false||losartannull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Daily|Time|false|false||dailynull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|clopidogrel|Drug|false|false||Clopidogrel
null|clopidogrel|Drug|false|false||Clopidogrelnull|Daily|Time|false|false||DAILYnull|fluticasone propionate|Drug|false|false||Fluticasone Propionate
null|fluticasone propionate|Drug|false|false||Fluticasone Propionatenull|fluticasone|Drug|false|false||Fluticasone
null|fluticasone|Drug|false|false||Fluticasonenull|propionate|Drug|false|false||Propionate
null|Propionates|Drug|false|false||Propionatenull|Puff Dosing Unit|LabModifier|false|false||PUFF
null|Picofarad|LabModifier|false|false||PUFFnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|True primary (qualifier value)|Time|false|false||Primarynull|Primary|Modifier|false|false||Primarynull|Elevation procedure|Procedure|false|false||elevationnull|Elevation|Modifier|false|false||elevationnull|Coronary Artery Disease|Disorder|false|false||coronary artery disease
null|Coronary Arteriosclerosis|Disorder|false|false||coronary artery diseasenull|Coronary artery|Anatomy|false|false||coronary arterynull|Heart|Anatomy|false|false||coronarynull|Coronary|Modifier|false|false||coronarynull|Arteriopathic disease|Disorder|false|false||artery diseasenull|Arterial system|Anatomy|false|false||artery
null|Arteries|Anatomy|false|false||arterynull|Disease|Disorder|false|false||diseasenull|Neoplasm Metastasis|Disorder|false|false||Secondarynull|metastatic qualifier|Finding|false|false||Secondarynull|Secondary to|Modifier|false|false||Secondarynull|second (number)|LabModifier|false|false||Secondarynull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||diabetes mellitus type 2null|Diabetes Mellitus|Disorder|false|false||diabetes mellitusnull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||diabetes
null|Diabetes|Disorder|false|false||diabetes
null|Diabetes Mellitus|Disorder|false|false||diabetesnull|Type 2|Finding|false|false||type 2null|Type - ParameterizedDataType|Finding|false|false||type
null|SGCG gene|Finding|false|false||typenull|null|Modifier|false|false||typenull|Hypertensive disease|Disorder|false|false||hypertensionnull|Hyperlipidemia|Disorder|false|false||hyperlipidemia
null|Hyperlipoproteinemias|Disorder|false|false||hyperlipidemianull|Serum lipids high (finding)|Finding|false|false||hyperlipidemianull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Disease|Disorder|false|false||Conditionnull|Logical Condition|Finding|false|false||Conditionnull|null|Attribute|false|false||Conditionnull|Condition|Modifier|false|false||Conditionnull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Coordination of Benefits - Independent|Finding|false|false||Independent
null|Religious Affiliation - Independent|Finding|false|false||Independent
null|Independence|Finding|false|false||Independent
null|Independently able|Finding|false|false||Independentnull|Discharge instructions|Finding|false|false||Discharge Instructionsnull|hospital discharge instructions (treatment)|Procedure|false|false||Discharge Instructionsnull|null|Attribute|false|false||Discharge Instructionsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructionsnull|Production Class Code - Pleasure|Finding|false|false||pleasure
null|pleasurable emotion|Finding|false|false||pleasurenull|Pleasure - Animals raised for recreation|Entity|false|false||pleasurenull|care of - AddressPartType|Finding|false|false||care ofnull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Recent|Time|false|false||recentnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Chest Pain|Finding|false|false||chest painnull|null|Attribute|false|false||chest painnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|Myocardial Infarction|Disorder|false|false||heart attacknull|Malignant neoplasm of heart|Disorder|false|false||heart
null|benign neoplasm of heart|Disorder|false|false||heartnull|HEART PROBLEM|Finding|false|false||heartnull|Chest>Heart|Anatomy|false|false||heart
null|Heart|Anatomy|false|false||heartnull|Attack (finding)|Finding|false|false||attack
null|Attack behavior|Finding|false|false||attacknull|Attack device|Device|false|false||attacknull|Cardiac catheterisation as the cause of abnormal reaction of the patient, or of later complication, without mention of misadventure at the time of the procedure|Disorder|false|false||cardiac catheterizationnull|Diagnostic Service Section ID - Cardiac Catheterization|Finding|false|false||cardiac catheterizationnull|Consent Type - Cardiac Catheterization|Procedure|false|false||cardiac catheterization
null|Cardiac Catheterization Procedures|Procedure|false|false||cardiac catheterizationnull|Cardiac attachment|Finding|false|false||cardiacnull|Heart|Anatomy|false|false||cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||cardiacnull|Catheterization|Procedure|false|false||catheterizationnull|Graft material|Drug|false|false||graftsnull|Transplanted tissue|Anatomy|false|false||graftsnull|grafting qualifier|Modifier|false|false||graftsnull|Recent|Time|true|false||recentnull|Cardiac attachment|Finding|true|false||cardiacnull|Heart|Anatomy|true|false||cardiacnull|Cardiac - anatomy qualifier|Modifier|true|false||cardiacnull|Bypass surgery|Procedure|true|false||bypass surgerynull|Creation of shunt|Procedure|true|false||bypassnull|Level of Care - Surgery|Finding|true|false||surgery
null|Surgical procedure finding|Finding|true|false||surgery
null|Surgical aspects|Finding|true|false||surgerynull|Operative Surgical Procedures|Procedure|true|false||surgerynull|General surgery specialty|Title|true|false||surgery
null|Surgery specialty|Title|true|false||surgerynull|Diagnosis Type - Working|Finding|true|false||workingnull|Work|Event|true|false||workingnull|Working animal|Entity|true|false||workingnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|Start brand of breakfast cereal|Drug|false|false||STARTnull|start - HtmlLinkType|Finding|false|false||STARTnull|Collagen Tile Brachytherapy|Procedure|false|false||STARTnull|Beginning|Time|false|false||STARTnull|losartan|Drug|false|false||losartan
null|losartan|Drug|false|false||losartannull|Start brand of breakfast cereal|Drug|false|false||STARTnull|start - HtmlLinkType|Finding|false|false||STARTnull|Collagen Tile Brachytherapy|Procedure|false|false||STARTnull|Beginning|Time|false|false||STARTnull|isosorbide mononitrate|Drug|false|false||isosorbide mononitrate
null|isosorbide mononitrate|Drug|false|false||isosorbide mononitratenull|isosorbide|Drug|false|false||isosorbide
null|isosorbide|Drug|false|false||isosorbidenull|Increase|Finding|false|false||INCREASEnull|atorvastatin|Drug|false|false||atorvastatin
null|atorvastatin|Drug|false|false||atorvastatinnull|Increase|Finding|false|false||INCREASEnull|metoprolol|Drug|false|false||metoprolol
null|metoprolol|Drug|false|false||metoprololnull|Reduced|Finding|false|false||DECREASEnull|Decrease|LabModifier|false|false||DECREASEnull|aspirin|Drug|false|false||aspirin
null|aspirin|Drug|false|false||aspirinnull|Reduced|Finding|false|false||DECREASEnull|Decrease|LabModifier|false|false||DECREASEnull|pantoprazole|Drug|false|false||pantoprazole
null|pantoprazole|Drug|false|false||pantoprazolenull|Stop brand of fluoride|Drug|false|false||STOP
null|Stop brand of fluoride|Drug|false|false||STOPnull|MAP6 gene|Finding|false|false||STOPnull|Stop (Instruction Imperative)|Event|false|false||STOPnull|Stop (qualifier value)|Time|false|false||STOPnull|ibuprofen|Drug|false|false||ibuprofen
null|ibuprofen|Drug|false|false||ibuprofennull|Too much|Finding|false|false||too muchnull|Much|Finding|false|false||muchnull|Tylenol|Drug|false|false||tylenol
null|Tylenol|Drug|false|false||tylenolnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Further|Modifier|false|false||furthernull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Collection Object - UML Entity|Finding|false|false||collection
null|Item Collection|Finding|false|false||collection
null|Collections (publication)|Finding|false|false||collection
null|Collection (action)|Finding|false|false||collectionnull|Left lung|Anatomy|false|false||left lungnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Lung diseases|Disorder|false|false||lungnull|Lung Problem|Finding|false|false||lungnull|Chest>Lung|Anatomy|false|false||lung
null|Lung|Anatomy|false|false||lungnull|Observation Interpretation - better|Finding|false|false||betternull|Better|Modifier|false|false||betternull|Disease Management|Procedure|false|false||managementnull|Management Occupations|Subject|false|false||managementnull|Management procedure|Event|false|false||management
null|Administration occupational activities|Event|false|false||managementnull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||diabetes
null|Diabetes|Disorder|false|false||diabetes
null|Diabetes Mellitus|Disorder|false|false||diabetesnull|Help document|Finding|false|false||helpnull|Assisted (qualifier value)|Modifier|false|false||helpnull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions