CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Pharmaceutical Preparations|Drug|false|false||MEDICINEnull|Medicine|Title|false|false||MEDICINEnull|Known|Modifier|false|false||Knownnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|Adverse reaction to drug|Finding|true|false||Adverse Drug Reactionsnull|Adverse reaction to drug|Finding|true|false||Drug Reactionsnull|Pharmaceutical Preparations|Drug|false|false||Drug
null|Pharmacologic Substance|Drug|false|false||Drugnull|Drug problem|Finding|false|false||Drugnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Chest Pain|Finding|false|false||Chest Painnull|null|Attribute|false|false||Chest Painnull|Chest problem|Finding|false|false||Chestnull|Chest|Anatomy|false|false||Chest
null|Anterior thoracic region|Anatomy|false|false||Chestnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Females|Subject|false|false||female
null|Woman|Subject|false|false||femalenull|Female, Self-Report|Modifier|false|false||female
null|Female Phenotype|Modifier|false|false||femalenull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Hypertensive disease|Disorder|false|false||hypertensionnull|Asthma|Disorder|false|false||asthmanull|Recent|Time|false|false||recentnull|Diagnosis Classification - Diagnosis|Finding|false|false||diagnosis
null|diagnosis aspects|Finding|false|false||diagnosisnull|Diagnosis|Procedure|false|false||diagnosisnull|null|Attribute|false|false||diagnosisnull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Stress bismuth subsalicylate|Drug|false|false||stress
null|Stress bismuth subsalicylate|Drug|false|false||stressnull|Stress|Finding|false|false||stressnull|W stress|Attribute|false|false||stressnull|ECHO protocol|Procedure|false|false||echo
null|Extension for Community Healthcare Outcomes|Procedure|false|false||echonull|Echo <Calopterygidae>|Entity|false|false||echonull|Thought|Finding|false|false||thought
null|null|Finding|false|false||thoughtnull|Single vessel disease|Disorder|false|false||single vessel diseasenull|Marital Status - Single|Finding|false|false||single
null|Unmarried|Finding|false|false||singlenull|Singular|LabModifier|false|false||singlenull|Vessel Positions|Anatomy|false|false||vessel
null|Blood Vessel|Anatomy|false|false||vesselnull|Vessel (unit of presentation)|LabModifier|false|false||vesselnull|Disease|Disorder|false|false||diseasenull|Intermittent|Time|false|false||intermittentnull|Chest Pain|Finding|false|false||chest painnull|null|Attribute|false|false||chest painnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Recent|Time|false|false||recentnull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|History of recent hospitalization|Finding|false|false||recent hospitalizationnull|Recent|Time|false|false||recentnull|Hospitalization|Procedure|false|false||hospitalizationnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Cardiac enzymes|Drug|false|false||cardiac enzymes
null|Cardiac enzymes|Drug|false|false||cardiac enzymesnull|Cardiac enzymes/isoenzymes measurement|Procedure|false|false||cardiac enzymesnull|null|Attribute|false|false||cardiac enzymesnull|Cardiac attachment|Finding|false|false||cardiacnull|Heart|Anatomy|false|false||cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||cardiacnull|Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM|Drug|false|false||enzymes
null|Enzymes, peripheral vasodilators|Drug|false|false||enzymes
null|Enzymes, peripheral vasodilators|Drug|false|false||enzymes
null|Enzymes, peripheral vasodilators|Drug|false|false||enzymes
null|Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM|Drug|false|false||enzymes
null|Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM|Drug|false|false||enzymes
null|Enzymes, antithrombotic|Drug|false|false||enzymes
null|Enzymes, antithrombotic|Drug|false|false||enzymes
null|Enzymes, antithrombotic|Drug|false|false||enzymes
null|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS|Drug|false|false||enzymes
null|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS|Drug|false|false||enzymes
null|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS|Drug|false|false||enzymes
null|Enzymes, hematological|Drug|false|false||enzymes
null|Enzymes, hematological|Drug|false|false||enzymes
null|Enzymes, hematological|Drug|false|false||enzymes
null|Enzymes|Drug|false|false||enzymes
null|Enzymes|Drug|false|false||enzymes
null|Enzymes for ALIMENTARY TRACT AND METABOLISM|Drug|false|false||enzymes
null|Enzymes for ALIMENTARY TRACT AND METABOLISM|Drug|false|false||enzymes
null|Enzymes for ALIMENTARY TRACT AND METABOLISM|Drug|false|false||enzymesnull|enzymology|Finding|false|false||enzymesnull|Echocardiography, Stress|Procedure|false|false||stress echonull|Stress bismuth subsalicylate|Drug|false|false||stress
null|Stress bismuth subsalicylate|Drug|false|false||stressnull|Stress|Finding|false|false||stressnull|W stress|Attribute|false|false||stressnull|ECHO protocol|Procedure|false|false||echo
null|Extension for Community Healthcare Outcomes|Procedure|false|false||echonull|Echo <Calopterygidae>|Entity|false|false||echonull|Induce (action)|Finding|false|false||induciblenull|Ischemia|Finding|false|false||ischemianull|Ischemia Procedure|Procedure|false|false||ischemianull|Achieved|Finding|false|false||achievednull|Workload|LabModifier|false|false||workloadnull|Thought|Finding|false|false||thought
null|null|Finding|false|false||thoughtnull|Single vessel disease|Disorder|false|false||single vessel diseasenull|Marital Status - Single|Finding|false|false||single
null|Unmarried|Finding|false|false||singlenull|Singular|LabModifier|false|false||singlenull|Vessel Positions|Anatomy|false|false||vessel
null|Blood Vessel|Anatomy|false|false||vesselnull|Vessel (unit of presentation)|LabModifier|false|false||vesselnull|Disease|Disorder|false|false||diseasenull|ECHO protocol|Procedure|false|false||echo
null|Extension for Community Healthcare Outcomes|Procedure|false|false||echonull|Echo <Calopterygidae>|Entity|false|false||echonull|Report (document)|Finding|false|false||reportnull|Reporting|Procedure|false|false||reportnull|null|Attribute|false|false||reportnull|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Infantile Neuroaxonal Dystrophy|Disorder|false|false||plannull|Treatment Plan|Finding|false|false||plan
null|Planned|Finding|false|false||plan
null|null|Finding|false|false||plannull|Medical referral type|Finding|false|false||medical
null|Medical|Finding|false|false||medical
null|Medical school type|Finding|false|false||medicalnull|Medical service|Procedure|false|false||medicalnull|Disease Management|Procedure|false|false||managementnull|Management Occupations|Subject|false|false||managementnull|Management procedure|Event|false|false||management
null|Administration occupational activities|Event|false|false||managementnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Lung diseases|Disorder|false|false||pulmonary diseasenull|History of - respiratory disease|Finding|false|false||pulmonary diseasenull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Disease|Disorder|false|false||diseasenull|Adrenergic beta-Antagonists|Drug|false|false||beta blockernull|Beta adrenergic receptor antagonist (disposition)|Modifier|false|false||beta blockernull|Greek letter beta|Finding|false|false||betanull|Beta <eudicots>|Entity|false|false||betanull|Beta Distribution|LabModifier|false|false||betanull|diltiazem|Drug|false|false||diltiazem
null|diltiazem|Drug|false|false||diltiazemnull|Daily|Time|false|false||dailynull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Intermittent|Time|false|false||intermittentnull|Episode of|Time|false|false||episodesnull|Multinational Association of Supportive Care in Cancer Antiemesis Tool|Finding|false|false||MAT
null|MAT1A wt Allele|Finding|false|false||MAT
null|[acyl-carrier-protein] S-malonyltransferase activity|Finding|false|false||MAT
null|Multifocal atrial tachycardia|Finding|false|false||MAT
null|ACAT1 wt Allele|Finding|false|false||MAT
null|ACAT1 gene|Finding|false|false||MAT
null|MAT1A gene|Finding|false|false||MATnull|Mats|Device|false|false||MATnull|MAT Format|Modifier|false|false||MATnull|Authorization Mode - Phone|Finding|false|false||phone
null|Visit User Code - Phone|Finding|false|false||phone
null|Telephone Number|Finding|false|false||phone
null|MDFAttributeType - Phone|Finding|false|false||phonenull|Telephone|Device|false|false||phonenull|Person location type - Phone|Modifier|false|false||phonenull|Transaction counts and value totals - year|Finding|false|false||year
null|Precision - year|Finding|false|false||yearnull|year|Time|false|false||yearnull|Old|Time|false|false||oldnull|Aunt|Subject|false|false||auntnull|Very hard|Finding|false|false||very hardnull|Very|Modifier|false|false||verynull|Hardness|Modifier|false|false||hardnull|outcomes otolaryngology hearing|Finding|false|false||hearing
null|Hearing finding|Finding|false|false||hearing
null|Hearing|Finding|false|false||hearingnull|Aunt|Subject|false|false||auntnull|Authorization Mode - Phone|Finding|false|false||phone
null|Visit User Code - Phone|Finding|false|false||phone
null|Telephone Number|Finding|false|false||phone
null|MDFAttributeType - Phone|Finding|false|false||phonenull|Telephone|Device|false|false||phonenull|Person location type - Phone|Modifier|false|false||phonenull|Chest Pain|Finding|false|false||chest painnull|null|Attribute|false|false||chest painnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Dull pain|Finding|false|false||dull painnull|Dull pain|Finding|false|false||dullnull|Dull sensation quality|Modifier|false|false||dull
null|Dull|Modifier|false|false||dullnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Examination of shoulder(s)|Procedure|false|false||shoulder
null|Procedures on Shoulder|Procedure|false|false||shouldernull|Upper extremity>Shoulder|Anatomy|false|false||shoulder
null|Shoulder|Anatomy|false|false||shouldernull|Left breast|Anatomy|false|false||left breastnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false||breastnull|Breast problem|Finding|false|false||breastnull|Procedures on breast|Procedure|false|false||breastnull|Breast|Anatomy|false|false||breastnull|Worst|Modifier|false|false||worstnull|At home|Finding|false|false||at homenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|minor (disease)|Disorder|false|false||minornull|NR4A3 wt Allele|Finding|false|false||minor
null|NR4A3 gene|Finding|false|false||minornull|Minor (person)|Subject|false|false||minornull|Minor (value)|Modifier|false|false||minornull|Improvement|Finding|false|false||improvementnull|Associated with|Modifier|false|false||associatednull|Dyspnea|Finding|false|false||SOBnull|Nausea and vomiting|Finding|false|false||nausea/vomitingnull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|Vomiting|Finding|false|false||vomitingnull|sleeping upright or using specific number of extra pillows (orthopnea)|Finding|true|false||orthopnea
null|Orthopnea|Finding|true|false||orthopneanull|Paroxysmal nocturnal dyspnea|Disorder|true|false||PNDnull|NPPA wt Allele|Finding|true|false||PND
null|NPPA gene|Finding|true|false||PNDnull|Edema|Finding|true|false||edemanull|null|Attribute|true|false||edemanull|Palpitations|Finding|false|false||palpitationsnull|Initial (abbreviation)|Finding|false|false||initialnull|Initially|Time|false|false||initialnull|Firstly|Modifier|false|false||initialnull|Electrocardiogram image|Finding|false|false||EKG
null|Electrocardiogram|Finding|false|false||EKGnull|Electrocardiography|Procedure|false|false||EKGnull|Left Bundle-Branch Block|Disorder|false|false||LBBBnull|null|Lab|false|false||LBBBnull|null|Finding|false|false||unchangednull|About The Same|Modifier|false|false||unchangednull|null|Time|false|false||priornull|Plain chest X-ray|Procedure|false|false||CXRnull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Process Pharmacologic Substance|Drug|false|false||processnull|Process (qualifier value)|Finding|false|false||processnull|bony process|Anatomy|false|false||processnull|Process|Phenomenon|false|false||processnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|aspirin|Drug|false|false||aspirin
null|aspirin|Drug|false|false||aspirinnull|aspirin|Drug|false|false||aspirin
null|aspirin|Drug|false|false||aspirinnull|At home|Finding|false|false||at homenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Episode of|Time|false|false||episodesnull|Chest Pain|Finding|false|false||chest painnull|null|Attribute|false|false||chest painnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Further|Modifier|false|false||furthernull|Intervention regimes|Procedure|false|false||intervention
null|Nursing interventions|Procedure|false|false||intervention
null|Interventional procedure|Procedure|false|false||interventionnull|Transfer - product ownership|Finding|false|false||transfer
null|Transfer Technique|Finding|false|false||transfer
null|ActClass - transfer|Finding|false|false||transfer
null|null|Finding|false|false||transfernull|Transfer (immobility management)|Procedure|false|false||transfernull|arrival - ActRelationshipType|Finding|false|false||arrivalnull|null|Event|false|false||arrivalnull|Floor (anatomic)|Anatomy|false|false||floornull|floor (object)|Device|false|false||floornull|Floor - story of building|Entity|false|false||floornull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Initial (abbreviation)|Finding|false|false||initialnull|Initially|Time|false|false||initialnull|Firstly|Modifier|false|false||initialnull|Current (present time)|Time|false|false||currentlynull|A little bit|Finding|false|false||a little bitnull|A little bit|Finding|false|false||a little
null|Only a Little|Finding|false|false||a littlenull|Little's Disease|Disorder|false|false||littlenull|Only a Little|Finding|false|false||littlenull|Smallest|LabModifier|false|false||little
null|Small|LabModifier|false|false||littlenull|2-(4-ethoxybenzyl)-1-diethylaminoethyl-5-isothiocyanatobenzimidazole|Drug|false|false||bit
null|2-(4-ethoxybenzyl)-1-diethylaminoethyl-5-isothiocyanatobenzimidazole|Drug|false|false||bit
null|PTPNS1 protein, human|Drug|false|false||bitnull|Breast-Impact of Treatment Scale|Finding|false|false||bit
null|PTPNS1 protein, human|Finding|false|false||bit
null|SIRPA gene|Finding|false|false||bit
null|SIRPA wt Allele|Finding|false|false||bitnull|bit - unit of measure|LabModifier|false|false||bitnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Complaint (finding)|Finding|false|false||complaintsnull|Hypertensive disease|Disorder|false|false||HTNnull|Asthma|Disorder|false|false||Asthmanull|Diverticulitis|Disorder|false|false||Diverticulitisnull|Several|LabModifier|false|false||severalnull|year|Time|false|false||yearsnull|FBXW7 wt Allele|Finding|false|false||ago
null|FBXW7 gene|Finding|false|false||agonull|Right hip region structure|Anatomy|false|false||R hipnull|Prosthetic arthroplasty of hip (procedure)|Procedure|false|false||hip replacementnull|heme iron polypeptide|Drug|false|false||hip
null|ST13 protein, human|Drug|false|false||hip
null|ST13 protein, human|Drug|false|false||hip
null|RPL29 protein, human|Drug|false|false||hip
null|RPL29 protein, human|Drug|false|false||hip
null|HHIP protein, human|Drug|false|false||hip
null|HHIP protein, human|Drug|false|false||hip
null|heme iron polypeptide|Drug|false|false||hipnull|RPL29 wt Allele|Finding|false|false||hip
null|REG3A gene|Finding|false|false||hip
null|RPL29 gene|Finding|false|false||hip
null|ST13 wt Allele|Finding|false|false||hip
null|ST13 gene|Finding|false|false||hip
null|HHIP gene|Finding|false|false||hip
null|HHIP wt Allele|Finding|false|false||hip
null|REG3A wt Allele|Finding|false|false||hipnull|Procedure on hip|Procedure|false|false||hipnull|Lower extremity>Hip|Anatomy|false|false||hip
null|Hip structure|Anatomy|false|false||hip
null|Structure of habenulopeduncular tract|Anatomy|false|false||hip
null|Bone structure of ischium|Anatomy|false|false||hipnull|Replacement|Finding|false|false||replacementnull|Replacement - supply|Procedure|false|false||replacement
null|Surgical Replantation|Procedure|false|false||replacementnull|exercise induced|Finding|false|false||Exertionalnull|Atypical chest pain|Finding|false|false||Atypical Chest Painnull|atypia morphology|Finding|false|false||Atypicalnull|Atypical|Modifier|false|false||Atypicalnull|Chest Pain|Finding|false|false||Chest Painnull|null|Attribute|false|false||Chest Painnull|Chest problem|Finding|false|false||Chestnull|Chest|Anatomy|false|false||Chest
null|Anterior thoracic region|Anatomy|false|false||Chestnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Relationship - Mother|Finding|false|false||Mothernull|Mother (person)|Subject|false|false||Mothernull|Hypertensive disease|Disorder|false|false||HTNnull|Indirect exposure mechanism - Father|Finding|false|false||Father
null|Relationship - Father|Finding|false|false||Father
null|Father - courtesy title|Finding|false|false||Fathernull|Father (person)|Subject|false|false||Fathernull|Brother - courtesy title|Finding|false|false||Brother
null|Relationship - Brother|Finding|false|false||Brothernull|Brothers|Subject|false|false||Brothernull|Brother - courtesy title|Finding|false|false||Brother
null|Relationship - Brother|Finding|false|false||Brothernull|Brothers|Subject|false|false||Brothernull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|On admission|Time|false|false||On Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||GENERALnull|General medical service|Procedure|false|false||GENERALnull|Generalized|Modifier|false|false||GENERALnull|Females|Subject|false|false||female
null|Woman|Subject|false|false||femalenull|Female, Self-Report|Modifier|false|false||female
null|Female Phenotype|Modifier|false|false||femalenull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|Oriented to place|Finding|false|false||Orientednull|Orientation, Spatial|Modifier|false|false||Orientednull|Mood (psychological function)|Finding|false|false||Mood
null|mood (physical finding)|Finding|false|false||Mood
null|Mood (attribute)|Finding|false|false||Moodnull|null|Attribute|false|false||Moodnull|Affect (mental function)|Finding|false|false||affectnull|assessment of affect|Procedure|false|false||affectnull|Appropriate|Modifier|false|false||appropriatenull|HEENT|Anatomy|false|false||HEENTnull|Scleral Diseases|Disorder|false|false||Scleranull|examination of sclera|Procedure|false|false||Scleranull|Sclera|Anatomy|false|false||Scleranull|Anicteric|Finding|false|false||anictericnull|Malignant neoplasm of conjunctiva|Disorder|false|false||Conjunctiva
null|Benign neoplasm of conjunctiva|Disorder|false|false||Conjunctiva
null|Conjunctival Diseases|Disorder|false|false||Conjunctivanull|Specimen Type - Conjunctiva|Finding|false|false||Conjunctiva
null|null|Finding|false|false||Conjunctivanull|examination of conjunctiva|Procedure|false|false||Conjunctiva
null|Procedure on conjunctiva|Procedure|false|false||Conjunctivanull|Structure of palpebral conjunctiva|Anatomy|false|false||Conjunctiva
null|conjunctiva|Anatomy|false|false||Conjunctivanull|Pink color|Modifier|false|false||pinknull|Pallor of skin|Finding|true|false||pallornull|Cyanosis|Finding|false|false||cyanosisnull|Oral mucous membrane structure|Anatomy|false|false||oral mucosanull|Oral Dosage Form|Drug|false|false||oralnull|Oral Route of Administration|Finding|false|false||oral
null|Oral (intended site)|Finding|false|false||oralnull|Oral cavity|Anatomy|false|false||oralnull|Oral|Modifier|false|false||oralnull|null|Finding|false|false||mucosanull|Mucous Membrane|Anatomy|false|false||mucosanull|Passive joint movement of neck (finding)|Finding|false|false||NECK
null|Neck problem|Finding|false|false||NECKnull|dendritic spine neck|Anatomy|false|false||NECK
null|Neck|Anatomy|false|false||NECKnull|Supple|Finding|false|false||Supplenull|Cardiac attachment|Finding|false|false||CARDIACnull|Heart|Anatomy|false|false||CARDIACnull|Cardiac - anatomy qualifier|Modifier|false|false||CARDIACnull|Cardiac thrill (finding)|Finding|true|false||thrillsnull|hoist [device]|Device|true|false||liftsnull|Lung|Anatomy|false|false||LUNGSnull|Deformity of chest wall|Disorder|true|false||chest wall deformitiesnull|Chest wall structure|Anatomy|false|false||chest wall
null|Chest>Chest wall|Anatomy|false|false||chest wallnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Walls of a building|Device|false|false||wallnull|Congenital Abnormality|Disorder|true|false||deformitiesnull|deformities qualifier|Modifier|false|false||deformitiesnull|Congenital scoliosis|Disorder|true|false||scoliosis
null|null|Disorder|true|false||scoliosis
null|Acquired scoliosis|Disorder|true|false||scoliosisnull|Kyphosis deformity of spine|Disorder|true|false||kyphosis
null|Acquired kyphosis|Disorder|true|false||kyphosis
null|Congenital kyphosis|Disorder|true|false||kyphosisnull|kyphosis|Finding|true|false||kyphosisnull|Respiratory, thoracic and mediastinal disorders|Disorder|false|false||Respnull|Respiratory rate|Attribute|false|false||Respnull|Unlabored|Finding|false|false||unlaborednull|Use of accessory muscles|Finding|true|false||accessory muscle usenull|Accessory skeletal muscle|Disorder|true|false||accessory musclenull|Accessory|Device|true|false||accessorynull|Muscle (organ)|Anatomy|false|false||muscle
null|Muscle Tissue|Anatomy|false|false||musclenull|Use - dosing instruction imperative|Finding|true|false||use
null|utilization qualifier|Finding|true|false||use
null|Usage|Finding|true|false||usenull|Decreased breath sounds|Finding|false|false||decreased breath soundsnull|null|Attribute|false|false||breath sounds
null|Respiratory Sounds|Attribute|false|false||breath soundsnull|Breath|Finding|false|false||breathnull|null|Device|false|false||soundsnull|null|Phenomenon|false|false||soundsnull|Cancer/Testis Antigen|Drug|false|false||CTAnull|PCYT1A wt Allele|Finding|false|false||CTA
null|CERNA3 gene|Finding|false|false||CTAnull|Cardiac Computerized Tomographic Angiography|Procedure|false|false||CTAnull|Basilar Rales|Finding|true|false||crackles
null|Rales|Finding|true|false||cracklesnull|Wheezing|Finding|true|false||wheezesnull|Rhonchi|Finding|true|false||rhonchinull|Malignant neoplasm of abdomen|Disorder|false|false||ABDOMENnull|Abdomen problem|Finding|false|false||ABDOMENnull|Abdomen|Anatomy|false|false||ABDOMEN
null|Abdominal Cavity|Anatomy|false|false||ABDOMENnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||Softnull|Soft|Modifier|false|false||Softnull|Emotional tenderness|Finding|true|false||tenderness
null|Sore to touch|Finding|true|false||tendernessnull|All extremities|Anatomy|false|false||EXTREMITIES
null|Limb structure|Anatomy|false|false||EXTREMITIESnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false||SKIN
null|Skin and subcutaneous tissue disorders|Disorder|false|false||SKINnull|Skin Specimen Source Code|Finding|false|false||SKIN
null|Skin Specimen|Finding|false|false||SKINnull|Skin, Human|Anatomy|false|false||SKIN
null|Skin|Anatomy|false|false||SKINnull|Stasis dermatitis|Disorder|true|false||stasis dermatitisnull|Stasis|Finding|false|false||stasisnull|Dermatitis|Disorder|true|false||dermatitisnull|Ulcer|Finding|true|false||ulcersnull|Scar Tissue|Finding|true|false||scars
null|Cicatrix|Finding|true|false||scarsnull|Xanthoma|Disorder|true|false||xanthomasnull|null|Drug|false|false||PULSESnull|Physiologic pulse|Finding|false|false||PULSESnull|Pulse taking|Procedure|false|false||PULSESnull|Table Cell Horizontal Align - right|Finding|false|false||Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|Table Cell Horizontal Align - left|Finding|false|false||Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Primed lymphocyte test|Procedure|false|false||PLTnull|Count Dosing Unit|LabModifier|false|false||COUNT
null|Count|LabModifier|false|false||COUNTnull|Monos|Drug|false|false||MONOS
null|Mono-S|Drug|false|false||MONOS
null|Monos|Drug|false|false||MONOSnull|SARCOIDOSIS, EARLY-ONSET|Disorder|false|false||EOS
null|Familial eosinophilia|Disorder|false|false||EOSnull|PRSS33 gene|Finding|false|false||EOS
null|IKZF4 gene|Finding|false|false||EOSnull|Eos <Loriini>|Entity|false|false||EOSnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||HGB
null|Hemoglobin|Drug|false|false||HGBnull|CYGB gene|Finding|false|false||HGBnull|Hemoglobin concentration|Lab|false|false||HGBnull|Hemopoietic stem cell transplant|Procedure|false|false||HCT
null|Hematocrit Measurement|Procedure|false|false||HCTnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSEnull|Glucose measurement|Procedure|false|false||GLUCOSEnull|Glucose^1.5H post dose glucagon|Lab|false|false||GLUCOSEnull|urea|Drug|false|false||UREA
null|urea|Drug|false|false||UREA
null|urea|Drug|false|false||UREAnull|Urea measurement|Procedure|false|false||UREAnull|Sodium supplements|Drug|false|false||SODIUM
null|sodium|Drug|false|false||SODIUM
null|sodium|Drug|false|false||SODIUM
null|Sodium Drug Class|Drug|false|false||SODIUMnull|Sodium metabolic function|Finding|false|false||SODIUMnull|Sodium measurement|Procedure|false|false||SODIUMnull|Potassium Drug Class|Drug|false|false||POTASSIUM
null|Dietary Potassium|Drug|false|false||POTASSIUM
null|potassium|Drug|false|false||POTASSIUM
null|potassium|Drug|false|false||POTASSIUM
null|potassium|Drug|false|false||POTASSIUM
null|Potassium supplement|Drug|false|false||POTASSIUM
null|Potassium supplement|Drug|false|false||POTASSIUMnull|Potassium metabolic function|Finding|false|false||POTASSIUMnull|Potassium measurement|Procedure|false|false||POTASSIUMnull|chloride ion|Drug|false|false||CHLORIDE
null|Chlorides|Drug|false|false||CHLORIDEnull|Chloride metabolic function|Finding|false|false||CHLORIDEnull|Chloride measurement|Procedure|false|false||CHLORIDEnull|Total|Modifier|false|false||TOTALnull|carbon dioxide|Drug|false|false||CO2
null|carbon dioxide|Drug|false|false||CO2null|MT-CO2 gene|Finding|false|false||CO2
null|null|Finding|false|false||CO2
null|C2 wt Allele|Finding|false|false||CO2null|blood anion gap (lab test)|Procedure|false|false||ANION GAP
null|Anion gap measurement|Procedure|false|false||ANION GAPnull|Anion Gap|Attribute|false|false||ANION GAPnull|Anion gap result|Lab|false|false||ANION GAPnull|Anions|Drug|false|false||ANIONnull|Ras GTPase-Activating Protein 1, Human|Drug|false|false||GAP
null|Ras GTPase-Activating Protein 1, Human|Drug|false|false||GAP
null|GTPase-Activating Proteins|Drug|false|false||GAP
null|GTPase-Activating Proteins|Drug|false|false||GAPnull|RASA1 wt Allele|Finding|false|false||GAP
null|RASA1 gene|Finding|false|false||GAPnull|Gap (space)|Modifier|false|false||GAPnull|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSEnull|Glucose measurement|Procedure|false|false||GLUCOSEnull|Glucose^1.5H post dose glucagon|Lab|false|false||GLUCOSEnull|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MB
null|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MBnull|creatine kinase activity|Finding|false|false||CK-MBnull|Serum creatine phosphokinase MB isoenzyme measurement|Procedure|false|false||CK-MB
null|Creatine kinase MB measurement|Procedure|false|false||CK-MBnull|MB 3|Drug|false|false||MB-3null|Creatine Kinase|Drug|false|false||CPK
null|Creatine Kinase|Drug|false|false||CPKnull|PIK3C2A gene|Finding|false|false||CPKnull|Creatine kinase measurement|Procedure|false|false||CPKnull|Plain chest X-ray|Procedure|false|false||CXRnull|Pulmonary Emphysema|Disorder|false|false||Emphysemanull|Pathological accumulation of air in tissues|Finding|false|false||Emphysemanull|Pneumonia|Disorder|true|false||pneumonianull|Congestive heart failure|Disorder|true|false||CHFnull|Choroidal fissure|Anatomy|false|false||CHFnull|Knowledge acquisition using a method of assessment|Finding|false|false||ASSESSMENTnull|assessment of cognitive functions|Procedure|false|false||ASSESSMENT
null|Physical Examination|Procedure|false|false||ASSESSMENT
null|Nutrition Assessment|Procedure|false|false||ASSESSMENT
null|null|Procedure|false|false||ASSESSMENT
null|null|Procedure|false|false||ASSESSMENT
null|null|Procedure|false|false||ASSESSMENT
null|null|Procedure|false|false||ASSESSMENT
null|Personal care assessment|Procedure|false|false||ASSESSMENT
null|null|Procedure|false|false||ASSESSMENT
null|null|Procedure|false|false||ASSESSMENT
null|null|Procedure|false|false||ASSESSMENT
null|Evaluation procedure|Procedure|false|false||ASSESSMENT
null|Evaluation|Procedure|false|false||ASSESSMENT
null|null|Procedure|false|false||ASSESSMENT
null|null|Procedure|false|false||ASSESSMENT
null|null|Procedure|false|false||ASSESSMENT
null|null|Procedure|false|false||ASSESSMENT
null|null|Procedure|false|false||ASSESSMENTnull|Assessed|Event|false|false||ASSESSMENTnull|Infantile Neuroaxonal Dystrophy|Disorder|false|false||PLANnull|Treatment Plan|Finding|false|false||PLAN
null|Planned|Finding|false|false||PLAN
null|null|Finding|false|false||PLANnull|Transaction counts and value totals - year|Finding|false|false||year
null|Precision - year|Finding|false|false||yearnull|year|Time|false|false||yearnull|Old|Time|false|false||oldnull|Females|Subject|false|false||female
null|Woman|Subject|false|false||femalenull|Female, Self-Report|Modifier|false|false||female
null|Female Phenotype|Modifier|false|false||femalenull|Recent|Time|false|false||recentnull|Diagnosis Classification - Diagnosis|Finding|false|false||diagnosis
null|diagnosis aspects|Finding|false|false||diagnosisnull|Diagnosis|Procedure|false|false||diagnosisnull|null|Attribute|false|false||diagnosisnull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Hypertensive disease|Disorder|false|false||HTNnull|Asthma|Disorder|false|false||asthmanull|Intermittent|Time|false|false||intermittentnull|Episode of|Time|false|false||episodesnull|Chest Pain|Finding|false|false||chest painnull|null|Attribute|false|false||chest painnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Recent|Time|false|false||recentnull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Intermittent|Time|false|false||intermittentnull|Episode of|Time|false|false||episodesnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Burning sensation|Finding|false|false||burningnull|Burning sensation quality|Modifier|false|false||burningnull|Usual|Modifier|false|false||typicalnull|Angina Pectoris|Finding|true|false||angina
null|null|Finding|true|false||anginanull|null|Attribute|true|false||anginanull|Intervention regimes|Procedure|true|false||intervention
null|Nursing interventions|Procedure|true|false||intervention
null|Interventional procedure|Procedure|true|false||interventionnull|Relationship by association|Finding|false|false||association
null|Mental association|Finding|false|false||association
null|NCI Thesaurus Association|Finding|false|false||association
null|Association Class|Finding|false|false||associationnull|Chemical Association|Phenomenon|false|false||associationnull|Relationships|Modifier|false|false||associationnull|Exercise|Finding|false|false||exercisenull|Exercise Pain Management|Procedure|false|false||exercisenull|findings aspects|Finding|false|false||findingsnull|null|Attribute|false|false||findingsnull|Recent|Time|false|false||recentnull|Echocardiography, Stress|Procedure|false|false||stress echonull|Stress bismuth subsalicylate|Drug|false|false||stress
null|Stress bismuth subsalicylate|Drug|false|false||stressnull|Stress|Finding|false|false||stressnull|W stress|Attribute|false|false||stressnull|ECHO protocol|Procedure|false|false||echo
null|Extension for Community Healthcare Outcomes|Procedure|false|false||echonull|Echo <Calopterygidae>|Entity|false|false||echonull|Induce (action)|Finding|false|false||induciblenull|Ischemia|Finding|false|false||ischemianull|Ischemia Procedure|Procedure|false|false||ischemianull|Electrical Current|Phenomenon|false|false||currentnull|Current (present time)|Time|false|false||currentnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Underlying|Finding|false|false||underlyingnull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Troponin|Drug|false|false||troponins
null|Troponin|Drug|false|false||troponinsnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Hospital Stay|Time|false|false||hospital staynull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Imdur|Drug|false|false||Imdur
null|Imdur|Drug|false|false||Imdurnull|In addition to|Finding|false|false||in addition tonull|In addition to|Finding|false|false||addition
null|Add - instruction imperative|Finding|false|false||additionnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Last|Modifier|false|false||lastnull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Observation Interpretation - better|Finding|false|false||betternull|Better|Modifier|false|false||betternull|Medical referral type|Finding|false|false||medical
null|Medical|Finding|false|false||medical
null|Medical school type|Finding|false|false||medicalnull|Medical service|Procedure|false|false||medicalnull|Disease Management|Procedure|false|false||managementnull|Management Occupations|Subject|false|false||managementnull|Management procedure|Event|false|false||management
null|Administration occupational activities|Event|false|false||managementnull|null|Time|false|false||prior tonull|null|Time|false|false||priornull|SERPINA5 protein, human|Drug|false|false||PCI
null|SERPINA5 protein, human|Drug|false|false||PCInull|Peritoneal Cancer Index|Finding|false|false||PCI
null|SERPINA5 wt Allele|Finding|false|false||PCI
null|SERPINA5 gene|Finding|false|false||PCInull|Percutaneous Coronary Intervention|Procedure|false|false||PCI
null|photochemical internalization|Procedure|false|false||PCI
null|Prophylactic Cranial Irradiation|Procedure|false|false||PCInull|Picocurie|LabModifier|false|false||PCInull|Future|Time|false|false||futurenull|Administration (procedure)|Procedure|false|false||administrationnull|Administration occupational activities|Event|false|false||administrationnull|Imdur|Drug|false|false||IMDUR
null|Imdur|Drug|false|false||IMDURnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Several|LabModifier|false|false||severalnull|Prior functioning.stairs|Finding|false|false||stairsnull|Dyspnea|Finding|false|false||short of breathnull|Shortened|Modifier|false|false||shortnull|Short Value|LabModifier|false|false||short
null|Short|LabModifier|false|false||shortnull|Breath|Finding|false|false||breathnull|Cardiac attachment|Finding|false|false||cardiacnull|Heart|Anatomy|false|false||cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||cardiacnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|FACT Complex|Drug|false|false||fact
null|FACT Complex|Drug|false|false||factnull|SSRP1 wt Allele|Finding|false|false||fact
null|SUPT16H gene|Finding|false|false||factnull|Foundation for the Accreditation of Cellular Therapy|Subject|false|false||factnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Rhythm|Finding|false|false||RHYTHM
null|rhythmic process (biological)|Finding|false|false||RHYTHMnull|Left Bundle-Branch Block|Disorder|false|false||LBBBnull|null|Lab|false|false||LBBBnull|Electrocardiogram image|Finding|false|false||EKG
null|Electrocardiogram|Finding|false|false||EKGnull|Electrocardiography|Procedure|false|false||EKGnull|Regular|Modifier|false|false||regularnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|New diagnosis (finding)|Finding|false|false||new diagnosisnull|New Diagnosis Procedure|Procedure|false|false||new diagnosisnull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|Diagnosis Classification - Diagnosis|Finding|false|false||diagnosis
null|diagnosis aspects|Finding|false|false||diagnosisnull|Diagnosis|Procedure|false|false||diagnosisnull|null|Attribute|false|false||diagnosisnull|Multinational Association of Supportive Care in Cancer Antiemesis Tool|Finding|false|false||MAT
null|MAT1A wt Allele|Finding|false|false||MAT
null|[acyl-carrier-protein] S-malonyltransferase activity|Finding|false|false||MAT
null|Multifocal atrial tachycardia|Finding|false|false||MAT
null|ACAT1 wt Allele|Finding|false|false||MAT
null|ACAT1 gene|Finding|false|false||MAT
null|MAT1A gene|Finding|false|false||MATnull|Mats|Device|false|false||MATnull|MAT Format|Modifier|false|false||MATnull|Last|Modifier|false|false||lastnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|diltiazem|Drug|false|false||Diltiazem
null|diltiazem|Drug|false|false||Diltiazemnull|Several|LabModifier|false|false||severalnull|Episode of|Time|false|false||episodesnull|Multinational Association of Supportive Care in Cancer Antiemesis Tool|Finding|false|false||MAT
null|MAT1A wt Allele|Finding|false|false||MAT
null|[acyl-carrier-protein] S-malonyltransferase activity|Finding|false|false||MAT
null|Multifocal atrial tachycardia|Finding|false|false||MAT
null|ACAT1 wt Allele|Finding|false|false||MAT
null|ACAT1 gene|Finding|false|false||MAT
null|MAT1A gene|Finding|false|false||MATnull|Mats|Device|false|false||MATnull|MAT Format|Modifier|false|false||MATnull|Telephone Number|Finding|false|false||tele
null|TCAP gene|Finding|false|false||telenull|Asymptomatic diagnosis of|Finding|false|false||asymptomatic
null|Asymptomatic (finding)|Finding|false|false||asymptomaticnull|Frequently|Time|false|false||frequentnull|Fenamole|Drug|false|false||PAT
null|Fenamole|Drug|false|false||PATnull|Paroxysmal atrial tachycardia|Disorder|false|false||PATnull|glutamate-prephenate aminotransferase activity|Finding|false|false||PAT
null|aspartate-prephenate aminotransferase activity|Finding|false|false||PAT
null|protein acetyltransferase activity|Finding|false|false||PATnull|Thermoacoustic Computed Tomography|Procedure|false|false||PATnull|Heart|Anatomy|false|false||Heartsnull|Monitor brand of insecticide|Drug|false|false||monitor
null|Monitor brand of insecticide|Drug|false|false||monitornull|Monitor Device|Device|false|false||monitor
null|Monitoring Device|Device|false|false||monitornull|Monitor, occupation|Subject|false|false||monitornull|On discharge|Time|false|false||on dischargenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Tachyarrhythmia|Finding|false|false||tachyarrhythmianull|Immunization Registry Status - Inactive|Finding|false|false||Inactive
null|Physical Inactivity|Finding|false|false||Inactive
null|Inactive Healthcare Coverage|Finding|false|false||Inactive
null|Certificate Status - Inactive|Finding|false|false||Inactive
null|Inactive - answer to question|Finding|false|false||Inactive
null|Edit Status - Inactive|Finding|false|false||Inactivenull|Inactive Entity|Modifier|false|false||Inactive
null|Sedentary|Modifier|false|false||Inactivenull|Hypertensive disease|Disorder|false|false||Hypertensionnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|hydrochlorothiazide|Drug|false|false||HCTZ
null|hydrochlorothiazide|Drug|false|false||HCTZnull|diltiazem|Drug|false|false||diltiazem
null|diltiazem|Drug|false|false||diltiazemnull|Asthma|Disorder|false|false||Asthmanull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Gastroesophageal reflux disease|Disorder|false|false||GERDnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|omeprazole|Drug|false|false||omeprazole
null|omeprazole|Drug|false|false||omeprazolenull|Full|Modifier|false|false||fullnull|MDF Attribute Type - Code|Finding|false|false||code
null|A Codes|Finding|false|false||code
null|Code|Finding|false|false||codenull|Coding|Event|false|false||codenull|Marketing basis - Transitional|Finding|false|false||Transitionalnull|Transitional cell morphology|Modifier|false|false||Transitionalnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Imdur|Drug|false|false||Imdur
null|Imdur|Drug|false|false||Imdurnull|Daily|Time|false|false||dailynull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Coronary Artery Disease|Disorder|false|false||coronary artery disease
null|Coronary Arteriosclerosis|Disorder|false|false||coronary artery diseasenull|Coronary artery|Anatomy|false|false||coronary arterynull|Heart|Anatomy|false|false||coronarynull|Coronary|Modifier|false|false||coronarynull|Arteriopathic disease|Disorder|false|false||artery diseasenull|Arterial system|Anatomy|false|false||artery
null|Arteries|Anatomy|false|false||arterynull|Disease|Disorder|false|false||diseasenull|Candidate|Finding|false|false||candidatenull|SERPINA5 protein, human|Drug|false|false||PCI
null|SERPINA5 protein, human|Drug|false|false||PCInull|Peritoneal Cancer Index|Finding|false|false||PCI
null|SERPINA5 wt Allele|Finding|false|false||PCI
null|SERPINA5 gene|Finding|false|false||PCInull|Percutaneous Coronary Intervention|Procedure|false|false||PCI
null|photochemical internalization|Procedure|false|false||PCI
null|Prophylactic Cranial Irradiation|Procedure|false|false||PCInull|Picocurie|LabModifier|false|false||PCInull|Future|Time|false|false||futurenull|Chest Pain|Finding|false|false||chest painnull|null|Attribute|false|false||chest painnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Return to (contextual qualifier) (qualifier value)|Modifier|false|false||returnnull|Event|Event|false|false||eventnull|Monitor brand of insecticide|Drug|false|false||monitor
null|Monitor brand of insecticide|Drug|false|false||monitornull|Monitor Device|Device|false|false||monitor
null|Monitoring Device|Device|false|false||monitornull|Monitor, occupation|Subject|false|false||monitornull|Processing type - Evaluation|Finding|false|false||evaluationnull|Evaluation procedure|Procedure|false|false||evaluation
null|Evaluation|Procedure|false|false||evaluationnull|Cardiac Arrhythmia|Disorder|false|false||arrhythmiasnull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|Acetaminophen [EPC]|Drug|false|false||acetaminophen
null|acetaminophen|Drug|false|false||acetaminophen
null|acetaminophen|Drug|false|false||acetaminophennull|Acetaminophen measurement|Procedure|false|false||acetaminophennull|Every four hours|Time|false|false||Q4Hnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|albuterol sulfate|Drug|false|false||albuterol sulfate
null|albuterol sulfate|Drug|false|false||albuterol sulfatenull|albuterol|Drug|false|false||albuterol
null|albuterol|Drug|false|false||albuterolnull|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||sulfate
null|Sulfates, Inorganic|Drug|false|false||sulfate
null|sulfate ion|Drug|false|false||sulfate
null|sulfate ion|Drug|false|false||sulfate
null|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||sulfatenull|microgram|LabModifier|false|false||mcgnull|Puff Dosing Unit|LabModifier|false|false||Puff
null|Picofarad|LabModifier|false|false||Puffnull|Inhalation Route of Administration|Finding|false|false||Inhalation
null|Inspiration (function)|Finding|false|false||Inhalationnull|Inhalation Dosing Unit|LabModifier|false|false||Inhalationnull|Every six hours|Time|false|false||Q6Hnull|Hour|Time|false|false||hoursnull|Dyspnea|Finding|false|false||SOBnull|Wheezing|Finding|false|false||wheezenull|fluticasone / salmeterol|Drug|false|false||fluticasone-salmeterolnull|fluticasone|Drug|false|false||fluticasone
null|fluticasone|Drug|false|false||fluticasonenull|salmeterol|Drug|false|false||salmeterol
null|salmeterol|Drug|false|false||salmeterolnull|microgram|LabModifier|false|false||mcgnull|Inhalation Route of Administration|Finding|false|false||Inhalation
null|Inspiration (function)|Finding|false|false||Inhalationnull|Inhalation Dosing Unit|LabModifier|false|false||Inhalationnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|fluticasone|Drug|false|false||fluticasone
null|fluticasone|Drug|false|false||fluticasonenull|microgram|LabModifier|false|false||mcgnull|Nasal brand of oxymetazoline|Drug|false|false||Nasal
null|Nasal brand of oxymetazoline|Drug|false|false||Nasal
null|Nasal dosage form|Drug|false|false||Nasalnull|Nasal Route of Administration|Finding|false|false||Nasal
null|Nasal (intended site)|Finding|false|false||Nasalnull|null|Anatomy|false|false||Nasalnull|Once A Day|Drug|false|false||once a daynull|Once daily|Time|false|false||once a daynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|hydrochlorothiazide|Drug|false|false||hydrochlorothiazide
null|hydrochlorothiazide|Drug|false|false||hydrochlorothiazidenull|Once A Day|Drug|false|false||once a daynull|Once daily|Time|false|false||once a daynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|omeprazole|Drug|false|false||omeprazole
null|omeprazole|Drug|false|false||omeprazolenull|Daily|Time|false|false||DAILYnull|simvastatin|Drug|false|false||simvastatin
null|simvastatin|Drug|false|false||simvastatinnull|Once A Day|Drug|false|false||once a daynull|Once daily|Time|false|false||once a daynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|tiotropium bromide|Drug|false|false||tiotropium bromide
null|tiotropium bromide|Drug|false|false||tiotropium bromidenull|tiotropium|Drug|false|false||tiotropium
null|tiotropium|Drug|false|false||tiotropiumnull|Bromides|Drug|false|false||bromidenull|Bromides measurement|Procedure|false|false||bromidenull|microgram|LabModifier|false|false||mcgnull|Daily|Time|false|false||DAILYnull|aspirin|Drug|false|false||aspirin
null|aspirin|Drug|false|false||aspirinnull|Once A Day|Drug|false|false||once a daynull|Once daily|Time|false|false||once a daynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Multivitamin preparation|Drug|false|false||multivitamin
null|Multivitamin preparation|Drug|false|false||multivitamin
null|Multivitamin preparation|Drug|false|false||multivitaminnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Daily|Time|false|false||DAILYnull|diltiazem hydrochloride|Drug|false|false||diltiazem HCl
null|diltiazem hydrochloride|Drug|false|false||diltiazem HClnull|diltiazem|Drug|false|false||diltiazem
null|diltiazem|Drug|false|false||diltiazemnull|Flinders medical centre-7 marker|Drug|false|false||HCl
null|hydrochloride|Drug|false|false||HCl
null|hydrochloride|Drug|false|false||HClnull|Hairy Cell Leukemia|Disorder|false|false||HClnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Daily|Time|false|false||dailynull|Singulair|Drug|false|false||singulair
null|Singulair|Drug|false|false||singulairnull|Once a day, at bedtime|Time|false|false||QHSnull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|Acetaminophen [EPC]|Drug|false|false||acetaminophen
null|acetaminophen|Drug|false|false||acetaminophen
null|acetaminophen|Drug|false|false||acetaminophennull|Acetaminophen measurement|Procedure|false|false||acetaminophennull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Hour|Time|false|false||hoursnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|albuterol sulfate|Drug|false|false||albuterol sulfate
null|albuterol sulfate|Drug|false|false||albuterol sulfatenull|albuterol|Drug|false|false||albuterol
null|albuterol|Drug|false|false||albuterolnull|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||sulfate
null|Sulfates, Inorganic|Drug|false|false||sulfate
null|sulfate ion|Drug|false|false||sulfate
null|sulfate ion|Drug|false|false||sulfate
null|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||sulfatenull|mcg/actuation|LabModifier|false|false||mcg/Actuationnull|microgram|LabModifier|false|false||mcgnull|Actuation (unit of presentation)|LabModifier|false|false||Actuationnull|Facial Hemiatrophy|Disorder|false|false||HFAnull|High frequency audiometry|Procedure|false|false||HFAnull|Inhalers, Aerosol|Device|false|false||Aerosol Inhalernull|Aerosol Dose Form|Drug|false|false||Aerosolnull|Aerosols|Device|false|false||Aerosolnull|Inhaler (unit of presentation)|Finding|false|false||Inhalernull|Inhaler|Device|false|false||Inhalernull|Inhaler Dosing Unit|LabModifier|false|false||Inhalernull|Puff Dosing Unit|LabModifier|false|false||Puff
null|Picofarad|LabModifier|false|false||Puffnull|Inhalation Route of Administration|Finding|false|false||Inhalation
null|Inspiration (function)|Finding|false|false||Inhalationnull|Inhalation Dosing Unit|LabModifier|false|false||Inhalationnull|Every six hours|Time|false|false||Q6Hnull|6 Hours|Time|false|false||6 hoursnull|Hour|Time|false|false||hoursnull|Dyspnea|Finding|false|false||sobnull|Wheezing|Finding|false|false||wheezingnull|fluticasone / salmeterol|Drug|false|false||fluticasone-salmeterolnull|fluticasone|Drug|false|false||fluticasone
null|fluticasone|Drug|false|false||fluticasonenull|salmeterol|Drug|false|false||salmeterol
null|salmeterol|Drug|false|false||salmeterolnull|microgram|LabModifier|false|false||mcgnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Disk Drug Form|Drug|false|false||Disknull|Disc - Body Part|Anatomy|false|false||Disknull|Disk Device|Device|false|false||Disk
null|Disk - package|Device|false|false||Disknull|Disk Shape|Modifier|false|false||Disknull|Disk Dosing Unit|LabModifier|false|false||Disknull|Participation Type - device|Finding|false|false||Devicenull|Medical Devices|Device|false|false||Device
null|Devices|Device|false|false||Devicenull|Kind of quantity - Device|LabModifier|false|false||Devicenull|Receptors, Antigen, B-Cell|Drug|false|false||Sig
null|Receptors, Antigen, B-Cell|Drug|false|false||Signull|Receptors, Antigen, B-Cell|Finding|false|false||Signull|Short insular gyrus|Anatomy|false|false||Signull|Surveillance Implementation Group|Entity|false|false||Sig
null|Staphylococcus intermedius group|Entity|false|false||Signull|Disk Drug Form|Drug|false|false||Disknull|Disc - Body Part|Anatomy|false|false||Disknull|Disk Device|Device|false|false||Disk
null|Disk - package|Device|false|false||Disknull|Disk Shape|Modifier|false|false||Disknull|Disk Dosing Unit|LabModifier|false|false||Disknull|Participation Type - device|Finding|false|false||Devicenull|Medical Devices|Device|false|false||Device
null|Devices|Device|false|false||Devicenull|Kind of quantity - Device|LabModifier|false|false||Devicenull|Inhalation Route of Administration|Finding|false|false||Inhalation
null|Inspiration (function)|Finding|false|false||Inhalationnull|Inhalation Dosing Unit|LabModifier|false|false||Inhalationnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|2 times|Finding|false|false||2 timesnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|fluticasone|Drug|false|false||fluticasone
null|fluticasone|Drug|false|false||fluticasonenull|mcg/actuation|LabModifier|false|false||mcg/Actuationnull|microgram|LabModifier|false|false||mcgnull|Actuation (unit of presentation)|LabModifier|false|false||Actuationnull|SPRAY, SUSPENSION|Drug|false|false||Spray, Suspensionnull|Spray Dosage Form|Drug|false|false||Spraynull|Spray (administration method)|Finding|false|false||Spraynull|Spray (action)|Event|false|false||Spraynull|Spray Dosing Unit|LabModifier|false|false||Spraynull|Suspension substance|Drug|false|false||Suspension
null|Suspensions|Drug|false|false||Suspensionnull|Suspension (action)|Finding|false|false||Suspensionnull|Spray Dosage Form|Drug|false|false||Spraynull|Spray (administration method)|Finding|false|false||Spraynull|Spray (action)|Event|false|false||Spraynull|Spray Dosing Unit|LabModifier|false|false||Spraynull|Nasal brand of oxymetazoline|Drug|false|false||Nasal
null|Nasal brand of oxymetazoline|Drug|false|false||Nasal
null|Nasal dosage form|Drug|false|false||Nasalnull|Nasal Route of Administration|Finding|false|false||Nasal
null|Nasal (intended site)|Finding|false|false||Nasalnull|null|Anatomy|false|false||Nasalnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|hydrochlorothiazide|Drug|false|false||hydrochlorothiazide
null|hydrochlorothiazide|Drug|false|false||hydrochlorothiazidenull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Once A Day|Drug|false|false||once a daynull|Once daily|Time|false|false||once a daynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|omeprazole|Drug|false|false||omeprazole
null|omeprazole|Drug|false|false||omeprazolenull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Delayed Release Dosage Form|Drug|false|false||Delayed Releasenull|Views delayed|Attribute|false|false||Delayednull|Deferred|Time|false|false||Delayednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Delayed Release Dosage Form|Drug|false|false||Delayed Releasenull|Views delayed|Attribute|false|false||Delayednull|Deferred|Time|false|false||Delayednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|simvastatin|Drug|false|false||simvastatin
null|simvastatin|Drug|false|false||simvastatinnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Once A Day|Drug|false|false||once a daynull|Once daily|Time|false|false||once a daynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|tiotropium bromide|Drug|false|false||tiotropium bromide
null|tiotropium bromide|Drug|false|false||tiotropium bromidenull|tiotropium|Drug|false|false||tiotropium
null|tiotropium|Drug|false|false||tiotropiumnull|Bromides|Drug|false|false||bromidenull|Bromides measurement|Procedure|false|false||bromidenull|microgram|LabModifier|false|false||mcgnull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Inhalation Devices|Device|false|false||Inhalation Devicenull|Inhalation Route of Administration|Finding|false|false||Inhalation
null|Inspiration (function)|Finding|false|false||Inhalationnull|Inhalation Dosing Unit|LabModifier|false|false||Inhalationnull|Participation Type - device|Finding|false|false||Devicenull|Medical Devices|Device|false|false||Device
null|Devices|Device|false|false||Devicenull|Kind of quantity - Device|LabModifier|false|false||Devicenull|capsule (pharmacologic)|Drug|false|false||Capnull|CATARACT, ANTERIOR POLAR|Disorder|false|false||Capnull|BRD4 wt Allele|Finding|false|false||Cap
null|HACD1 gene|Finding|false|false||Cap
null|SERPINB6 gene|Finding|false|false||Cap
null|BRD4 gene|Finding|false|false||Cap
null|CAP1 gene|Finding|false|false||Cap
null|SORBS1 gene|Finding|false|false||Cap
null|LNPEP gene|Finding|false|false||Capnull|CAP Regimen|Procedure|false|false||Cap
null|cisplatin/cyclophosphamide/doxorubicin protocol|Procedure|false|false||Cap
null|cyclophosphamide/doxorubicin/prednisone protocol|Procedure|false|false||Capnull|Cap (physical object)|Device|false|false||Cap
null|Syringe Caps|Device|false|false||Cap
null|Cap device|Device|false|false||Capnull|College of American Pathologists|Subject|false|false||Capnull|Controlled Attenuation Parameter|Modifier|false|false||Capnull|Capsule Dosing Unit|LabModifier|false|false||Capnull|Inhalation Route of Administration|Finding|false|false||Inhalation
null|Inspiration (function)|Finding|false|false||Inhalationnull|Inhalation Dosing Unit|LabModifier|false|false||Inhalationnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|aspirin|Drug|false|false||aspirin
null|aspirin|Drug|false|false||aspirinnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Once A Day|Drug|false|false||once a daynull|Once daily|Time|false|false||once a daynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Multivitamin tablet|Drug|false|false||multivitamin     Tabletnull|Multivitamin preparation|Drug|false|false||multivitamin
null|Multivitamin preparation|Drug|false|false||multivitamin
null|Multivitamin preparation|Drug|false|false||multivitaminnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|montelukast|Drug|false|false||montelukast
null|montelukast|Drug|false|false||montelukastnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Once a day, at bedtime|Time|false|false||QHSnull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Once a day, at bedtime|Time|false|false||at bedtimenull|Once a day, at bedtime|Time|false|false||bedtime
null|Bedtime (qualifier value)|Time|false|false||bedtimenull|isosorbide mononitrate|Drug|false|false||isosorbide mononitrate
null|isosorbide mononitrate|Drug|false|false||isosorbide mononitratenull|isosorbide|Drug|false|false||isosorbide
null|isosorbide|Drug|false|false||isosorbidenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Once A Day|Drug|false|false||once a daynull|Once daily|Time|false|false||once a daynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|refill|Finding|false|false||Refillsnull|diltiazem hydrochloride|Drug|false|false||diltiazem HCl
null|diltiazem hydrochloride|Drug|false|false||diltiazem HClnull|diltiazem|Drug|false|false||diltiazem
null|diltiazem|Drug|false|false||diltiazemnull|Flinders medical centre-7 marker|Drug|false|false||HCl
null|hydrochloride|Drug|false|false||HCl
null|hydrochloride|Drug|false|false||HClnull|Hairy Cell Leukemia|Disorder|false|false||HClnull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Once A Day|Drug|false|false||once a daynull|Once daily|Time|false|false||once a daynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|refill|Finding|false|false||Refillsnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|True primary (qualifier value)|Time|false|false||PRIMARYnull|Primary|Modifier|false|false||PRIMARYnull|Atypical chest pain|Finding|false|false||atypical chest painnull|atypia morphology|Finding|false|false||atypicalnull|Atypical|Modifier|false|false||atypicalnull|Chest Pain|Finding|false|false||chest painnull|null|Attribute|false|false||chest painnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Neoplasm Metastasis|Disorder|false|false||Secondarynull|metastatic qualifier|Finding|false|false||Secondarynull|Secondary to|Modifier|false|false||Secondarynull|second (number)|LabModifier|false|false||Secondarynull|Hypertensive disease|Disorder|false|false||Hypertensionnull|Asthma|Disorder|false|false||Asthmanull|Diverticulitis|Disorder|false|false||Diverticulitisnull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Coordination of Benefits - Independent|Finding|false|false||Independent
null|Religious Affiliation - Independent|Finding|false|false||Independent
null|Independence|Finding|false|false||Independent
null|Independently able|Finding|false|false||Independentnull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Atypical chest pain|Finding|false|false||atypical chest painnull|atypia morphology|Finding|false|false||atypicalnull|Atypical|Modifier|false|false||atypicalnull|Chest Pain|Finding|false|false||chest painnull|null|Attribute|false|false||chest painnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Telemetry|Procedure|false|false||telemetrynull|Electrocardiogram image|Finding|false|false||EKG
null|Electrocardiogram|Finding|false|false||EKGnull|Electrocardiography|Procedure|false|false||EKGnull|null|Finding|false|false||unchangednull|About The Same|Modifier|false|false||unchangednull|Cardiac enzymes|Drug|false|false||cardiac enzymes
null|Cardiac enzymes|Drug|false|false||cardiac enzymesnull|Cardiac enzymes/isoenzymes measurement|Procedure|false|false||cardiac enzymesnull|null|Attribute|false|false||cardiac enzymesnull|Cardiac attachment|Finding|false|false||cardiacnull|Heart|Anatomy|false|false||cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||cardiacnull|Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM|Drug|false|false||enzymes
null|Enzymes, peripheral vasodilators|Drug|false|false||enzymes
null|Enzymes, peripheral vasodilators|Drug|false|false||enzymes
null|Enzymes, peripheral vasodilators|Drug|false|false||enzymes
null|Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM|Drug|false|false||enzymes
null|Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM|Drug|false|false||enzymes
null|Enzymes, antithrombotic|Drug|false|false||enzymes
null|Enzymes, antithrombotic|Drug|false|false||enzymes
null|Enzymes, antithrombotic|Drug|false|false||enzymes
null|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS|Drug|false|false||enzymes
null|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS|Drug|false|false||enzymes
null|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS|Drug|false|false||enzymes
null|Enzymes, hematological|Drug|false|false||enzymes
null|Enzymes, hematological|Drug|false|false||enzymes
null|Enzymes, hematological|Drug|false|false||enzymes
null|Enzymes|Drug|false|false||enzymes
null|Enzymes|Drug|false|false||enzymes
null|Enzymes for ALIMENTARY TRACT AND METABOLISM|Drug|false|false||enzymes
null|Enzymes for ALIMENTARY TRACT AND METABOLISM|Drug|false|false||enzymes
null|Enzymes for ALIMENTARY TRACT AND METABOLISM|Drug|false|false||enzymesnull|enzymology|Finding|false|false||enzymesnull|Evidence of (contextual qualifier)|Finding|true|false||evidence fornull|Evidence|Finding|true|false||evidencenull|Malignant neoplasm of heart|Disorder|true|false||heart
null|benign neoplasm of heart|Disorder|true|false||heartnull|HEART PROBLEM|Finding|true|false||heartnull|Chest>Heart|Anatomy|false|false||heart
null|Heart|Anatomy|false|false||heartnull|Tissue damage|Disorder|true|false||damagenull|Damage|Finding|true|false||damage
null|MAGEE1 gene|Finding|true|false||damagenull|Myocardial Infarction|Disorder|false|false||heart attacknull|Malignant neoplasm of heart|Disorder|false|false||heart
null|benign neoplasm of heart|Disorder|false|false||heartnull|HEART PROBLEM|Finding|false|false||heartnull|Chest>Heart|Anatomy|false|false||heart
null|Heart|Anatomy|false|false||heartnull|Attack (finding)|Finding|false|false||attack
null|Attack behavior|Finding|false|false||attacknull|Attack device|Device|false|false||attacknull|Long Variable|Modifier|false|false||long
null|Long|Modifier|false|false||longnull|nitrate ion|Drug|false|false||nitrate
null|nitrate ion|Drug|false|false||nitrate
null|Nitrate|Drug|false|false||nitrate
null|Nitrates|Drug|false|false||nitratenull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Chest Pain|Finding|false|false||chest painnull|null|Attribute|false|false||chest painnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Pain|Finding|false|false||pain symptomsnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|diltiazem|Drug|false|false||diltiazem
null|diltiazem|Drug|false|false||diltiazemnull|Observation Interpretation - better|Finding|false|false||betternull|Better|Modifier|false|false||betternull|Blood pressure finding|Finding|false|false||blood pressure
null|Systemic arterial pressure|Finding|false|false||blood pressure
null|Blood Pressure|Finding|false|false||blood pressurenull|Blood pressure determination|Procedure|false|false||blood pressurenull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|Malignant neoplasm of heart|Disorder|false|false||heart
null|benign neoplasm of heart|Disorder|false|false||heartnull|HEART PROBLEM|Finding|false|false||heartnull|Chest>Heart|Anatomy|false|false||heart
null|Heart|Anatomy|false|false||heartnull|rate control|Finding|false|false||rate controlnull|Amount type - Rate|Finding|false|false||ratenull|Rating (action)|Event|false|false||ratenull|Rate|LabModifier|false|false||ratenull|Control brand of phenylpropanolamine|Drug|false|false||control
null|CONTROL veterinary product|Drug|false|false||control
null|control substance|Drug|false|false||control
null|Control brand of phenylpropanolamine|Drug|false|false||controlnull|Control - Relationship modifier|Finding|false|false||control
null|Control function|Finding|false|false||control
null|Scientific Control|Finding|false|false||controlnull|Control Groups|Subject|false|false||controlnull|True Control Status|Modifier|false|false||control
null|control aspects|Modifier|false|false||controlnull|48 hours|Time|false|false||48 hournull|Hour|Time|false|false||hournull|Holter Electrocardiography|Procedure|false|false||holter monitornull|Holter Monitors|Device|false|false||holter monitornull|Monitor brand of insecticide|Drug|false|false||monitor
null|Monitor brand of insecticide|Drug|false|false||monitornull|Monitor Device|Device|false|false||monitor
null|Monitoring Device|Device|false|false||monitornull|Monitor, occupation|Subject|false|false||monitornull|Observation Interpretation - better|Finding|false|false||betternull|Better|Modifier|false|false||betternull|Idea|Entity|false|false||ideanull|Cardiac rhythm type|Finding|false|false||heart rhythmnull|Malignant neoplasm of heart|Disorder|false|false||heart
null|benign neoplasm of heart|Disorder|false|false||heartnull|HEART PROBLEM|Finding|false|false||heartnull|Chest>Heart|Anatomy|false|false||heart
null|Heart|Anatomy|false|false||heartnull|Rhythm|Finding|false|false||rhythm
null|rhythmic process (biological)|Finding|false|false||rhythmnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Cardiovascular system|Anatomy|false|false||cardiologynull|cardiology (field)|Title|false|false||cardiologynull|Cardiology service|Entity|false|false||cardiologynull|Appointments|Event|false|false||appointmentnull|Pharmaceutical Preparations|Drug|false|false||MEDICATIONnull|medication - HL7 publishing domain|Finding|false|false||MEDICATION
null|Medications|Finding|false|false||MEDICATIONnull|Changing|Finding|false|false||CHANGESnull|Changed status|LabModifier|false|false||CHANGESnull|Start brand of breakfast cereal|Drug|false|false||STARTnull|start - HtmlLinkType|Finding|false|false||STARTnull|Collagen Tile Brachytherapy|Procedure|false|false||STARTnull|Beginning|Time|false|false||STARTnull|Daily|Time|false|false||dailynull|Increase|Finding|false|false||INCREASEnull|diltiazem|Drug|false|false||diltiazem
null|diltiazem|Drug|false|false||diltiazemnull|Daily|Time|false|false||dailynull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Medical referral type|Finding|false|false||medical
null|Medical|Finding|false|false||medical
null|Medical school type|Finding|false|false||medicalnull|Medical service|Procedure|false|false||medicalnull|Attention - G-code|Finding|false|false||attention
null|Attention|Finding|false|false||attentionnull|Chest Pain|Finding|false|false||chest painnull|null|Attribute|false|false||chest painnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Dyspnea|Finding|false|false||shortness of breathnull|null|Attribute|false|false||shortness of breathnull|Breath|Finding|false|false||breathnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions