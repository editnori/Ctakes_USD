 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
_|27,28
_|28,29
_|29,30
No|31,33
:|33,34
_|37,38
_|38,39
_|39,40
<EOL>|40,41
<EOL>|42,43
Admission|43,52
Date|53,57
:|57,58
_|60,61
_|61,62
_|62,63
Discharge|77,86
Date|87,91
:|91,92
_|95,96
_|96,97
_|97,98
<EOL>|98,99
<EOL>|100,101
Date|101,105
of|106,108
Birth|109,114
:|114,115
_|117,118
_|118,119
_|119,120
Sex|133,136
:|136,137
F|140,141
<EOL>|141,142
<EOL>|143,144
Service|144,151
:|151,152
MEDICINE|153,161
<EOL>|161,162
<EOL>|163,164
Allergies|164,173
:|173,174
<EOL>|175,176
No|176,178
Known|179,184
Allergies|185,194
/|195,196
Adverse|197,204
Drug|205,209
Reactions|210,219
<EOL>|219,220
<EOL>|221,222
Attending|222,231
:|231,232
_|233,234
_|234,235
_|235,236
.|236,237
<EOL>|237,238
<EOL>|239,240
Chief|240,245
Complaint|246,255
:|255,256
<EOL>|256,257
Diarrhea|257,265
-|266,267
Transfer|268,276
to|277,279
MICU|280,284
for|285,288
Hypoxia|289,296
<EOL>|296,297
<EOL>|298,299
Major|299,304
Surgical|305,313
or|314,316
Invasive|317,325
Procedure|326,335
:|335,336
<EOL>|336,337
_|337,338
_|338,339
_|339,340
line|341,345
placement|346,355
<EOL>|355,356
Right|356,361
pigtail|362,369
pleural|370,377
catheter|378,386
placement|387,396
<EOL>|396,397
<EOL>|398,399
History|399,406
of|407,409
Present|410,417
Illness|418,425
:|425,426
<EOL>|426,427
Pt|427,429
is|430,432
an|433,435
_|436,437
_|437,438
_|438,439
year|440,444
-|444,445
old|445,448
female|449,455
with|456,460
h|461,462
/|462,463
o|463,464
Sjogren|465,472
's|472,474
syndrome|475,483
,|483,484
IBS|485,488
,|488,489
<EOL>|490,491
who|491,494
presents|495,503
with|504,508
diarrhea|509,517
and|518,521
fever|522,527
.|527,528
Patietn|529,536
starting|537,545
having|546,552
<EOL>|553,554
non-bloody|554,564
,|564,565
watery|566,572
diarreha|573,581
approximately|582,595
three|596,601
weeks|602,607
ago|608,611
.|611,612
This|613,617
<EOL>|618,619
has|619,622
been|623,627
persistent|628,638
since|639,644
that|645,649
time|650,654
.|654,655
For|656,659
the|660,663
past|664,668
several|669,676
days|677,681
,|681,682
<EOL>|683,684
she|684,687
has|688,691
been|692,696
experiencing|697,709
crampy|710,716
b|717,718
/|718,719
l|719,720
lower|721,726
quadrant|727,735
abdominal|736,745
<EOL>|746,747
pain|747,751
and|752,755
distension|756,766
.|766,767
Today|768,773
she|774,777
developed|778,787
subjective|788,798
fever|799,804
and|805,808
<EOL>|809,810
rigors|810,816
at|817,819
home|820,824
.|824,825
Denies|826,832
nausea|833,839
,|839,840
vomiting|841,849
,|849,850
dysuria|851,858
.|858,859
Decreased|860,869
<EOL>|870,871
appetite|871,879
over|880,884
same|885,889
time|890,894
course|895,901
.|901,902
<EOL>|902,903
In|903,905
the|906,909
ED|910,912
,|912,913
initial|914,921
vs|922,924
were|925,929
:|929,930
98.5|931,935
125|936,939
111|940,943
/|943,944
63|944,946
22|947,949
100|950,953
%|953,954
.|954,955
Patient|956,963
<EOL>|964,965
AAOx3|965,970
.|970,971
Subsequently|972,984
febrile|985,992
to|993,995
101.0|996,1001
.|1001,1002
Exam|1003,1007
remarkable|1008,1018
for|1019,1022
mild|1023,1027
<EOL>|1028,1029
discomfort|1029,1039
to|1040,1042
palpation|1043,1052
in|1053,1055
RLQ|1056,1059
/|1059,1060
LLQ|1060,1063
.|1063,1064
Labs|1065,1069
notable|1070,1077
for|1078,1081
WBC|1082,1085
20.2|1086,1090
<EOL>|1091,1092
with|1092,1096
93.6|1097,1101
%|1101,1102
PMNs|1103,1107
(|1108,1109
no|1109,1111
bands|1112,1117
)|1117,1118
,|1118,1119
Na|1120,1122
127|1123,1126
,|1126,1127
lactate|1128,1135
2.2|1136,1139
,|1139,1140
normal|1141,1147
LFTs|1148,1152
.|1152,1153
UA|1154,1156
<EOL>|1157,1158
showed|1158,1164
5|1165,1166
hyaline|1167,1174
casts|1175,1180
,|1180,1181
no|1182,1184
mucus|1185,1190
/|1190,1191
WBC|1191,1194
/|1194,1195
RBC|1195,1198
etc|1199,1202
.|1202,1203
BCx|1204,1207
and|1208,1211
UCx|1212,1215
drawn|1216,1221
.|1221,1222
<EOL>|1223,1224
CT|1224,1226
_|1227,1228
_|1228,1229
_|1229,1230
with|1231,1235
contrast|1236,1244
showed|1245,1251
pancolitis|1252,1262
without|1263,1270
<EOL>|1271,1272
perforation|1272,1283
or|1284,1286
obstruction|1287,1298
,|1298,1299
intrahepatic|1300,1312
biliary|1313,1320
duct|1321,1325
dilatation|1326,1336
<EOL>|1337,1338
and|1338,1341
prominent|1342,1351
CBD|1352,1355
,|1355,1356
right|1357,1362
lung|1363,1367
base|1368,1372
consolidation|1373,1386
.|1386,1387
CXR|1388,1391
showed|1392,1398
<EOL>|1399,1400
bibasilar|1400,1409
opacities|1410,1419
+|1420,1421
/|1421,1422
-|1422,1423
pulm|1424,1428
edema|1429,1434
and|1435,1438
multiple|1439,1447
dilated|1448,1455
small|1456,1461
<EOL>|1462,1463
bowel|1463,1468
loops|1469,1474
.|1474,1475
Patient|1476,1483
given|1484,1489
2L|1490,1492
NS|1493,1495
,|1495,1496
2L|1497,1499
LR|1500,1502
,|1502,1503
IV|1504,1506
Cipro|1507,1512
,|1512,1513
IV|1514,1516
Flagyl|1517,1523
and|1524,1527
<EOL>|1528,1529
Tylenol|1529,1536
.|1536,1537
Patient|1538,1545
was|1546,1549
initially|1550,1559
admitted|1560,1568
to|1569,1571
medicine|1572,1580
floor|1581,1586
,|1586,1587
but|1588,1591
<EOL>|1592,1593
developed|1593,1602
hypoxia|1603,1610
while|1611,1616
in|1617,1619
ED|1620,1622
and|1623,1626
had|1627,1630
new|1631,1634
5L|1635,1637
O2|1638,1640
requirement|1641,1652
.|1652,1653
She|1654,1657
<EOL>|1658,1659
had|1659,1662
a|1663,1664
repeat|1665,1671
CXR|1672,1675
showing|1676,1683
possible|1684,1692
pneumonia|1693,1702
vs|1703,1705
.|1705,1706
pulmonary|1707,1716
edema|1717,1722
.|1722,1723
<EOL>|1724,1725
She|1725,1728
received|1729,1737
ceftriaxone|1738,1749
for|1750,1753
possible|1754,1762
pneumonia|1763,1772
and|1773,1776
was|1777,1780
<EOL>|1781,1782
transferred|1782,1793
to|1794,1796
MICU|1797,1801
.|1801,1802
<EOL>|1802,1803
.|1803,1804
<EOL>|1804,1805
On|1805,1807
arrival|1808,1815
to|1816,1818
the|1819,1822
MICU|1823,1827
,|1827,1828
patient|1829,1836
appears|1837,1844
uncomfortable|1845,1858
and|1859,1862
is|1863,1865
<EOL>|1866,1867
rigoring|1867,1875
.|1875,1876
She|1877,1880
reports|1881,1888
crampy|1889,1895
abdominal|1896,1905
pain|1906,1910
in|1911,1913
her|1914,1917
lower|1918,1923
<EOL>|1924,1925
abdomen|1925,1932
,|1932,1933
fevers|1934,1940
,|1940,1941
and|1942,1945
rigors|1946,1952
.|1952,1953
She|1954,1957
continues|1958,1967
to|1968,1970
have|1971,1975
diarrhea|1976,1984
,|1984,1985
but|1986,1989
<EOL>|1990,1991
no|1991,1993
nausea|1994,2000
or|2001,2003
vomiting|2004,2012
.|2012,2013
Mild|2014,2018
cough|2019,2024
productive|2025,2035
of|2036,2038
white|2039,2044
sputum|2045,2051
.|2051,2052
Of|2053,2055
<EOL>|2056,2057
note|2057,2061
,|2061,2062
patient|2063,2070
last|2071,2075
received|2076,2084
antibiotics|2085,2096
in|2097,2099
_|2100,2101
_|2101,2102
_|2102,2103
<EOL>|2104,2105
(|2105,2106
azithromycin|2106,2118
for|2119,2122
CAP|2123,2126
)|2126,2127
.|2127,2128
<EOL>|2128,2129
.|2129,2130
<EOL>|2130,2131
Review|2131,2137
of|2138,2140
systems|2141,2148
:|2148,2149
<EOL>|2149,2150
(|2150,2151
+|2151,2152
)|2152,2153
Per|2154,2157
HPI|2158,2161
<EOL>|2161,2162
(|2162,2163
-|2163,2164
)|2164,2165
Denies|2166,2172
night|2173,2178
sweats|2179,2185
.|2185,2186
Denies|2187,2193
headache|2194,2202
,|2202,2203
sinus|2204,2209
tenderness|2210,2220
,|2220,2221
<EOL>|2222,2223
rhinorrhea|2223,2233
or|2234,2236
congestion|2237,2247
.|2247,2248
Denies|2249,2255
shortness|2256,2265
of|2266,2268
breath|2269,2275
,|2275,2276
or|2277,2279
<EOL>|2280,2281
wheezing|2281,2289
.|2289,2290
Denies|2291,2297
chest|2298,2303
pain|2304,2308
,|2308,2309
chest|2310,2315
pressure|2316,2324
,|2324,2325
palpitations|2326,2338
,|2338,2339
or|2340,2342
<EOL>|2343,2344
weakness|2344,2352
.|2352,2353
Denies|2354,2360
nausea|2361,2367
,|2367,2368
vomiting|2369,2377
.|2377,2378
Denies|2379,2385
dysuria|2386,2393
,|2393,2394
frequency|2395,2404
,|2404,2405
or|2406,2408
<EOL>|2409,2410
urgency|2410,2417
.|2417,2418
Denies|2419,2425
arthralgias|2426,2437
or|2438,2440
myalgias|2441,2449
.|2449,2450
Denies|2451,2457
rashes|2458,2464
or|2465,2467
skin|2468,2472
<EOL>|2473,2474
changes|2474,2481
<EOL>|2481,2482
<EOL>|2483,2484
Past|2484,2488
Medical|2489,2496
History|2497,2504
:|2504,2505
<EOL>|2505,2506
Anemia|2506,2512
<EOL>|2512,2513
Borderline|2513,2523
cholesterol|2524,2535
<EOL>|2535,2536
C.|2536,2538
Diff|2539,2543
<EOL>|2543,2544
Heart|2544,2549
Murmur|2550,2556
<EOL>|2556,2557
Hypertension|2557,2569
<EOL>|2569,2570
Hypothyroidism|2570,2584
<EOL>|2584,2585
Mitral|2585,2591
Regurgitation|2592,2605
<EOL>|2605,2606
Osteoporosis|2606,2618
<EOL>|2618,2619
Pneumonia|2619,2628
<EOL>|2628,2629
Sinusitis|2629,2638
<EOL>|2638,2639
_|2639,2640
_|2640,2641
_|2641,2642
<EOL>|2643,2644
<EOL>|2645,2646
Social|2646,2652
History|2653,2660
:|2660,2661
<EOL>|2661,2662
_|2662,2663
_|2663,2664
_|2664,2665
<EOL>|2665,2666
Family|2666,2672
History|2673,2680
:|2680,2681
<EOL>|2681,2682
Long|2682,2686
history|2687,2694
of|2695,2697
hypertension|2698,2710
in|2711,2713
her|2714,2717
family|2718,2724
.|2724,2725
She|2727,2730
does|2731,2735
report|2736,2742
<EOL>|2743,2744
that|2744,2748
her|2749,2752
father|2753,2759
's|2759,2761
family|2762,2768
has|2769,2772
a|2773,2774
history|2775,2782
of|2783,2785
multiple|2786,2794
cancers|2795,2802
.|2802,2803
She|2805,2808
<EOL>|2809,2810
has|2810,2813
a|2814,2815
grandfather|2816,2827
with|2828,2832
a|2833,2834
history|2835,2842
of|2843,2845
stomach|2846,2853
cancer|2854,2860
and|2861,2864
an|2865,2867
uncle|2868,2873
<EOL>|2874,2875
with|2875,2879
a|2880,2881
history|2882,2889
of|2890,2892
throat|2893,2899
cancer|2900,2906
.|2906,2907
She|2909,2912
denies|2913,2919
any|2920,2923
history|2924,2931
of|2932,2934
<EOL>|2935,2936
colon|2936,2941
cancers|2942,2949
.|2949,2950
Father|2951,2957
had|2958,2961
stroke|2962,2968
.|2968,2969
No|2970,2972
family|2973,2979
h|2980,2981
/|2981,2982
o|2982,2983
MI|2984,2986
.|2986,2987
Mother|2988,2994
had|2995,2998
a|2999,3000
<EOL>|3001,3002
heart|3002,3007
valve|3008,3013
replaced|3014,3022
(|3023,3024
pt|3024,3026
not|3027,3030
sure|3031,3035
which|3036,3041
one|3042,3045
)|3045,3046
.|3046,3047
<EOL>|3047,3048
<EOL>|3048,3049
<EOL>|3050,3051
Physical|3051,3059
Exam|3060,3064
:|3064,3065
<EOL>|3065,3066
Admission|3066,3075
Exam|3076,3080
:|3080,3081
<EOL>|3081,3082
General|3082,3089
:|3089,3090
Alert|3091,3096
,|3096,3097
oriented|3098,3106
,|3106,3107
rigoring|3108,3116
,|3116,3117
appears|3118,3125
uncomfortable|3126,3139
<EOL>|3139,3140
HEENT|3140,3145
:|3145,3146
Sclera|3147,3153
anicteric|3154,3163
,|3163,3164
dry|3165,3168
mucus|3169,3174
membranes|3175,3184
,|3184,3185
EOMI|3186,3190
,|3190,3191
PERRL|3192,3197
<EOL>|3197,3198
Neck|3198,3202
:|3202,3203
supple|3204,3210
,|3210,3211
JVP|3212,3215
not|3216,3219
elevated|3220,3228
,|3228,3229
no|3230,3232
LAD|3233,3236
<EOL>|3236,3237
CV|3237,3239
:|3239,3240
Tachy|3241,3246
,|3246,3247
S1|3248,3250
,|3250,3251
S2|3252,3254
,|3254,3255
II|3256,3258
/|3258,3259
VI|3259,3261
holosystolic|3262,3274
murmur|3275,3281
at|3282,3284
apex|3285,3289
<EOL>|3289,3290
Lungs|3290,3295
:|3295,3296
Diffuse|3297,3304
rhonchi|3305,3312
,|3312,3313
no|3314,3316
wheezes|3317,3324
<EOL>|3324,3325
Abdomen|3325,3332
:|3332,3333
+|3334,3335
BP|3335,3337
,|3337,3338
Firm|3339,3343
,|3343,3344
distended|3345,3354
,|3354,3355
tender|3356,3362
to|3363,3365
palpation|3366,3375
in|3376,3378
right|3379,3384
and|3385,3388
<EOL>|3389,3390
left|3390,3394
lower|3395,3400
quadrant|3401,3409
,|3409,3410
no|3411,3413
rebound|3414,3421
/|3421,3422
guarding|3422,3430
<EOL>|3430,3431
GU|3431,3433
:|3433,3434
foley|3435,3440
in|3441,3443
place|3444,3449
<EOL>|3449,3450
Ext|3450,3453
:|3453,3454
warm|3455,3459
,|3459,3460
well|3461,3465
perfused|3466,3474
,|3474,3475
2|3476,3477
+|3477,3478
pulses|3479,3485
,|3485,3486
no|3487,3489
clubbing|3490,3498
,|3498,3499
cyanosis|3500,3508
or|3509,3511
<EOL>|3512,3513
edema|3513,3518
<EOL>|3518,3519
Neuro|3519,3524
:|3524,3525
CNII|3526,3530
-|3530,3531
XII|3531,3534
intact|3535,3541
,|3541,3542
moving|3543,3549
all|3550,3553
extremities|3554,3565
<EOL>|3566,3567
<EOL>|3567,3568
Discharge|3568,3577
exam|3578,3582
-|3583,3584
unchanged|3585,3594
from|3595,3599
above|3600,3605
,|3605,3606
except|3607,3613
as|3614,3616
below|3617,3622
:|3622,3623
<EOL>|3623,3624
General|3624,3631
:|3631,3632
tired|3633,3638
but|3639,3642
arousable|3643,3652
to|3653,3655
voice|3656,3661
,|3661,3662
appropriate|3663,3674
<EOL>|3674,3675
CV|3675,3677
:|3677,3678
RRR|3679,3682
,|3682,3683
_|3684,3685
_|3685,3686
_|3686,3687
systolic|3688,3696
murmur|3697,3703
at|3704,3706
the|3707,3710
apex|3711,3715
<EOL>|3715,3716
Lungs|3716,3721
:|3721,3722
Slightly|3723,3731
decreased|3732,3741
breath|3742,3748
sounds|3749,3755
at|3756,3758
the|3759,3762
lung|3763,3767
bases|3768,3773
,|3773,3774
right|3775,3780
<EOL>|3781,3782
pigtail|3782,3789
catheter|3790,3798
in|3799,3801
place|3802,3807
<EOL>|3807,3808
Abd|3808,3811
:|3811,3812
Hypoactive|3813,3823
BS|3824,3826
,|3826,3827
soft|3828,3832
,|3832,3833
non-tender|3834,3844
,|3844,3845
mildly|3846,3852
distended|3853,3862
<EOL>|3862,3863
Extr|3863,3867
:|3867,3868
2|3869,3870
+|3870,3871
edema|3872,3877
to|3878,3880
the|3881,3884
thigh|3885,3890
bilaterally|3891,3902
<EOL>|3902,3903
<EOL>|3904,3905
Pertinent|3905,3914
Results|3915,3922
:|3922,3923
<EOL>|3923,3924
Admission|3924,3933
Labs|3934,3938
:|3938,3939
<EOL>|3939,3940
_|3940,3941
_|3941,3942
_|3942,3943
10|3944,3946
:|3946,3947
20AM|3947,3951
BLOOD|3952,3957
WBC|3958,3961
-|3961,3962
20|3962,3964
.|3964,3965
2|3965,3966
*|3966,3967
#|3967,3968
RBC|3969,3972
-|3972,3973
3|3973,3974
.|3974,3975
76|3975,3977
*|3977,3978
Hgb|3979,3982
-|3982,3983
11|3983,3985
.|3985,3986
6|3986,3987
*|3987,3988
Hct|3989,3992
-|3992,3993
36.1|3993,3997
<EOL>|3998,3999
MCV|3999,4002
-|4002,4003
96|4003,4005
MCH|4006,4009
-|4009,4010
30.9|4010,4014
MCHC|4015,4019
-|4019,4020
32.3|4020,4024
RDW|4025,4028
-|4028,4029
12.8|4029,4033
Plt|4034,4037
_|4038,4039
_|4039,4040
_|4040,4041
<EOL>|4041,4042
_|4042,4043
_|4043,4044
_|4044,4045
10|4046,4048
:|4048,4049
20AM|4049,4053
BLOOD|4054,4059
Neuts|4060,4065
-|4065,4066
93|4066,4068
.|4068,4069
6|4069,4070
*|4070,4071
Lymphs|4072,4078
-|4078,4079
3|4079,4080
.|4080,4081
6|4081,4082
*|4082,4083
Monos|4084,4089
-|4089,4090
2.4|4090,4093
Eos|4094,4097
-|4097,4098
0.1|4098,4101
<EOL>|4102,4103
Baso|4103,4107
-|4107,4108
0.2|4108,4111
<EOL>|4111,4112
_|4112,4113
_|4113,4114
_|4114,4115
07|4116,4118
:|4118,4119
24PM|4119,4123
BLOOD|4124,4129
_|4130,4131
_|4131,4132
_|4132,4133
PTT|4134,4137
-|4137,4138
26.9|4138,4142
_|4143,4144
_|4144,4145
_|4145,4146
<EOL>|4146,4147
_|4147,4148
_|4148,4149
_|4149,4150
10|4151,4153
:|4153,4154
20AM|4154,4158
BLOOD|4159,4164
Glucose|4165,4172
-|4172,4173
121|4173,4176
*|4176,4177
UreaN|4178,4183
-|4183,4184
15|4184,4186
Creat|4187,4192
-|4192,4193
1.1|4193,4196
Na|4197,4199
-|4199,4200
127|4200,4203
*|4203,4204
<EOL>|4205,4206
K|4206,4207
-|4207,4208
4.3|4208,4211
Cl|4212,4214
-|4214,4215
89|4215,4217
*|4217,4218
HCO3|4219,4223
-|4223,4224
25|4224,4226
AnGap|4227,4232
-|4232,4233
17|4233,4235
<EOL>|4235,4236
_|4236,4237
_|4237,4238
_|4238,4239
10|4240,4242
:|4242,4243
20AM|4243,4247
BLOOD|4248,4253
ALT|4254,4257
-|4257,4258
26|4258,4260
AST|4261,4264
-|4264,4265
30|4265,4267
AlkPhos|4268,4275
-|4275,4276
78|4276,4278
TotBili|4279,4286
-|4286,4287
0.5|4287,4290
<EOL>|4290,4291
_|4291,4292
_|4292,4293
_|4293,4294
10|4295,4297
:|4297,4298
20AM|4298,4302
BLOOD|4303,4308
Lipase|4309,4315
-|4315,4316
21|4316,4318
<EOL>|4318,4319
_|4319,4320
_|4320,4321
_|4321,4322
07|4323,4325
:|4325,4326
24PM|4326,4330
BLOOD|4331,4336
Calcium|4337,4344
-|4344,4345
7|4345,4346
.|4346,4347
4|4347,4348
*|4348,4349
Phos|4350,4354
-|4354,4355
2|4355,4356
.|4356,4357
2|4357,4358
*|4358,4359
Mg|4360,4362
-|4362,4363
1.4|4363,4366
*|4366,4367
<EOL>|4367,4368
_|4368,4369
_|4369,4370
_|4370,4371
10|4372,4374
:|4374,4375
20AM|4375,4379
BLOOD|4380,4385
Albumin|4386,4393
-|4393,4394
4.1|4394,4397
<EOL>|4397,4398
_|4398,4399
_|4399,4400
_|4400,4401
10|4402,4404
:|4404,4405
29AM|4405,4409
BLOOD|4410,4415
Lactate|4416,4423
-|4423,4424
2|4424,4425
.|4425,4426
2|4426,4427
*|4427,4428
<EOL>|4428,4429
<EOL>|4429,4430
Discharge|4430,4439
Labs|4440,4444
:|4444,4445
<EOL>|4445,4446
_|4446,4447
_|4447,4448
_|4448,4449
07|4450,4452
:|4452,4453
30AM|4453,4457
BLOOD|4458,4463
WBC|4464,4467
-|4467,4468
7.1|4468,4471
RBC|4472,4475
-|4475,4476
3|4476,4477
.|4477,4478
11|4478,4480
*|4480,4481
Hgb|4482,4485
-|4485,4486
9|4486,4487
.|4487,4488
3|4488,4489
*|4489,4490
Hct|4491,4494
-|4494,4495
30|4495,4497
.|4497,4498
3|4498,4499
*|4499,4500
<EOL>|4501,4502
MCV|4502,4505
-|4505,4506
97|4506,4508
MCH|4509,4512
-|4512,4513
29.9|4513,4517
MCHC|4518,4522
-|4522,4523
30|4523,4525
.|4525,4526
7|4526,4527
*|4527,4528
RDW|4529,4532
-|4532,4533
14.0|4533,4537
Plt|4538,4541
_|4542,4543
_|4543,4544
_|4544,4545
<EOL>|4545,4546
_|4546,4547
_|4547,4548
_|4548,4549
07|4550,4552
:|4552,4553
30AM|4553,4557
BLOOD|4558,4563
Glucose|4564,4571
-|4571,4572
122|4572,4575
*|4575,4576
UreaN|4577,4582
-|4582,4583
20|4583,4585
Creat|4586,4591
-|4591,4592
0|4592,4593
.|4593,4594
3|4594,4595
*|4595,4596
Na|4597,4599
-|4599,4600
133|4600,4603
<EOL>|4604,4605
K|4605,4606
-|4606,4607
4.0|4607,4610
Cl|4611,4613
-|4613,4614
92|4614,4616
*|4616,4617
HCO3|4618,4622
-|4622,4623
39|4623,4625
*|4625,4626
AnGap|4627,4632
-|4632,4633
6|4633,4634
*|4634,4635
<EOL>|4635,4636
<EOL>|4636,4637
Micro|4637,4642
:|4642,4643
<EOL>|4643,4644
Stool|4644,4649
Culture|4650,4657
(|4658,4659
_|4659,4660
_|4660,4661
_|4661,4662
)|4662,4663
:|4663,4664
<EOL>|4664,4665
C.|4668,4670
difficile|4671,4680
DNA|4681,4684
amplification|4685,4698
assay|4699,4704
(|4705,4706
Final|4706,4711
_|4712,4713
_|4713,4714
_|4714,4715
:|4715,4716
<EOL>|4717,4718
Reported|4724,4732
to|4733,4735
and|4736,4739
read|4740,4744
back|4745,4749
by|4750,4752
_|4753,4754
_|4754,4755
_|4755,4756
-|4757,4758
-|4758,4759
CC7D|4759,4763
-|4763,4764
-|4764,4765
@|4766,4767
09|4768,4770
:|4770,4771
40|4771,4773
<EOL>|4774,4775
_|4775,4776
_|4776,4777
_|4777,4778
.|4778,4779
<EOL>|4780,4781
CLOSTRIDIUM|4787,4798
DIFFICILE|4799,4808
.|4808,4809
<EOL>|4810,4811
Positive|4820,4828
for|4829,4832
toxigenic|4833,4842
C.|4843,4845
difficile|4846,4855
by|4856,4858
the|4859,4862
Illumigene|4863,4873
<EOL>|4874,4875
DNA|4875,4878
<EOL>|4878,4879
amplification|4888,4901
.|4901,4902
(|4914,4915
Reference|4915,4924
Range|4925,4930
-|4930,4931
Negative|4931,4939
)|4939,4940
.|4940,4941
<EOL>|4942,4943
<EOL>|4943,4944
FECAL|4947,4952
CULTURE|4953,4960
(|4961,4962
Final|4962,4967
_|4968,4969
_|4969,4970
_|4970,4971
:|4971,4972
NO|4976,4978
SALMONELLA|4979,4989
OR|4990,4992
SHIGELLA|4993,5001
<EOL>|5002,5003
FOUND|5003,5008
.|5008,5009
<EOL>|5010,5011
<EOL>|5011,5012
CAMPYLOBACTER|5015,5028
CULTURE|5029,5036
(|5037,5038
Final|5038,5043
_|5044,5045
_|5045,5046
_|5046,5047
:|5047,5048
NO|5052,5054
CAMPYLOBACTER|5055,5068
<EOL>|5069,5070
FOUND|5070,5075
.|5075,5076
<EOL>|5076,5077
<EOL>|5077,5078
_|5078,5079
_|5079,5080
_|5080,5081
12|5082,5084
:|5084,5085
50|5085,5087
pm|5088,5090
Mini-BAL|5091,5099
<EOL>|5099,5100
<EOL>|5100,5101
*|5129,5130
*|5130,5131
FINAL|5131,5136
REPORT|5137,5143
_|5144,5145
_|5145,5146
_|5146,5147
<EOL>|5147,5148
<EOL>|5148,5149
GRAM|5152,5156
STAIN|5157,5162
(|5163,5164
Final|5164,5169
_|5170,5171
_|5171,5172
_|5172,5173
:|5173,5174
<EOL>|5175,5176
4|5182,5183
+|5183,5184
(|5187,5188
>|5188,5189
10|5189,5191
per|5192,5195
1000X|5196,5201
FIELD|5202,5207
)|5207,5208
:|5208,5209
POLYMORPHONUCLEAR|5212,5229
<EOL>|5230,5231
LEUKOCYTES|5231,5241
.|5241,5242
<EOL>|5243,5244
NO|5250,5252
MICROORGANISMS|5253,5267
SEEN|5268,5272
.|5272,5273
<EOL>|5274,5275
<EOL>|5275,5276
RESPIRATORY|5279,5290
CULTURE|5291,5298
(|5299,5300
Final|5300,5305
_|5306,5307
_|5307,5308
_|5308,5309
:|5309,5310
NO|5314,5316
GROWTH|5317,5323
,|5323,5324
<|5325,5326
1000|5326,5330
<EOL>|5331,5332
CFU|5332,5335
/|5335,5336
ml|5336,5338
.|5338,5339
<EOL>|5340,5341
<EOL>|5341,5342
_|5342,5343
_|5343,5344
_|5344,5345
10|5346,5348
:|5348,5349
42|5349,5351
am|5352,5354
PLEURAL|5355,5362
FLUID|5363,5368
PLEURAL|5374,5381
FLUID|5382,5387
.|5387,5388
<EOL>|5389,5390
<EOL>|5390,5391
GRAM|5394,5398
STAIN|5399,5404
(|5405,5406
Final|5406,5411
_|5412,5413
_|5413,5414
_|5414,5415
:|5415,5416
<EOL>|5417,5418
2|5424,5425
+|5425,5426
_|5429,5430
_|5430,5431
_|5431,5432
per|5433,5436
1000X|5437,5442
FIELD|5443,5448
)|5448,5449
:|5449,5450
POLYMORPHONUCLEAR|5453,5470
<EOL>|5471,5472
LEUKOCYTES|5472,5482
.|5482,5483
<EOL>|5484,5485
NO|5491,5493
MICROORGANISMS|5494,5508
SEEN|5509,5513
.|5513,5514
<EOL>|5515,5516
This|5522,5526
is|5527,5529
a|5530,5531
concentrated|5532,5544
smear|5545,5550
made|5551,5555
by|5556,5558
cytospin|5559,5567
method|5568,5574
,|5574,5575
<EOL>|5576,5577
please|5577,5583
refer|5584,5589
to|5590,5592
<EOL>|5592,5593
hematology|5599,5609
for|5610,5613
a|5614,5615
quantitative|5616,5628
white|5629,5634
blood|5635,5640
cell|5641,5645
count|5646,5651
.|5651,5652
.|5652,5653
<EOL>|5654,5655
<EOL>|5655,5656
FLUID|5659,5664
CULTURE|5665,5672
(|5673,5674
Final|5674,5679
_|5680,5681
_|5681,5682
_|5682,5683
:|5683,5684
NO|5688,5690
GROWTH|5691,5697
.|5697,5698
<EOL>|5699,5700
<EOL>|5700,5701
ANAEROBIC|5704,5713
CULTURE|5714,5721
(|5722,5723
Preliminary|5723,5734
)|5734,5735
:|5735,5736
NO|5740,5742
GROWTH|5743,5749
.|5749,5750
<EOL>|5751,5752
<EOL>|5752,5753
Legionella|5753,5763
Urinary|5764,5771
Antigen|5772,5779
(|5780,5781
_|5781,5782
_|5782,5783
_|5783,5784
)|5784,5785
:|5785,5786
NEG|5787,5790
FOR|5791,5794
LEGIONELLA|5795,5805
<EOL>|5806,5807
SEROGROUP|5807,5816
1|5817,5818
AG|5819,5821
<EOL>|5824,5825
<EOL>|5825,5826
Urine|5826,5831
Culture|5832,5839
:|5839,5840
negative|5841,5849
or|5850,5852
yeast|5853,5858
in|5859,5861
multiple|5862,5870
cultures|5871,5879
<EOL>|5879,5880
<EOL>|5880,5881
Blood|5881,5886
Cultures|5887,5895
:|5895,5896
NGTD|5897,5901
or|5902,5904
negative|5905,5913
in|5914,5916
multiple|5917,5925
cultures|5926,5934
<EOL>|5934,5935
<EOL>|5935,5936
Imaging|5936,5943
:|5943,5944
<EOL>|5944,5945
CT|5945,5947
Abd|5948,5951
/|5951,5952
Plevis|5952,5958
with|5959,5963
Contrast|5964,5972
(|5973,5974
_|5974,5975
_|5975,5976
_|5976,5977
)|5977,5978
:|5978,5979
<EOL>|5979,5980
IMPRESSION|5980,5990
:|5990,5991
<EOL>|5991,5992
1.|5992,5994
Diffuse|5996,6003
colonic|6004,6011
mucosal|6012,6019
hyperenhancement|6020,6036
and|6037,6040
bowel|6041,6046
wall|6047,6051
<EOL>|6052,6053
thickening|6053,6063
is|6064,6066
<EOL>|6066,6067
consistent|6067,6077
with|6078,6082
pancolitis|6083,6093
.|6093,6094
<EOL>|6094,6095
2.|6095,6097
Ground|6099,6105
-|6105,6106
glass|6106,6111
opacities|6112,6121
within|6122,6128
the|6129,6132
right|6133,6138
middle|6139,6145
and|6146,6149
right|6150,6155
<EOL>|6156,6157
lower|6157,6162
lobes|6163,6168
<EOL>|6168,6169
compatible|6169,6179
with|6180,6184
acute|6185,6190
infection|6191,6200
and|6201,6204
/|6204,6205
or|6205,6207
aspiration|6208,6218
.|6218,6219
Possible|6221,6229
<EOL>|6230,6231
mild|6231,6235
pulmonary|6236,6245
<EOL>|6245,6246
edema|6246,6251
.|6251,6252
<EOL>|6252,6253
3.|6253,6255
Intrahepatic|6257,6269
biliary|6270,6277
ductal|6278,6284
dilatation|6285,6295
and|6296,6299
prominence|6300,6310
of|6311,6313
the|6314,6317
<EOL>|6318,6319
common|6319,6325
bile|6326,6330
and|6331,6334
pancreatic|6335,6345
ducts|6346,6351
could|6352,6357
be|6358,6360
better|6361,6367
characterized|6368,6381
<EOL>|6382,6383
with|6383,6387
non-emergent|6388,6400
MRCP|6401,6405
.|6405,6406
<EOL>|6406,6407
<EOL>|6407,6408
CXR|6408,6411
(|6412,6413
_|6413,6414
_|6414,6415
_|6415,6416
)|6416,6417
:|6417,6418
<EOL>|6418,6419
IMPRESSION|6419,6429
:|6429,6430
<EOL>|6430,6431
1.|6431,6433
Bibasilar|6435,6444
opacities|6445,6454
would|6455,6460
be|6461,6463
consistent|6464,6474
with|6475,6479
pneumonia|6480,6489
<EOL>|6490,6491
and|6491,6494
/|6494,6495
or|6495,6497
aspiration|6498,6508
in|6509,6511
the|6512,6515
right|6516,6521
clinical|6522,6530
setting|6531,6538
.|6538,6539
Likely|6541,6547
some|6548,6552
<EOL>|6553,6554
component|6554,6563
of|6564,6566
pulmonary|6567,6576
edema|6577,6582
given|6583,6588
the|6589,6592
interstitial|6593,6605
thickening|6606,6616
.|6616,6617
<EOL>|6617,6618
2.|6618,6620
Multiple|6622,6630
dilated|6631,6638
loops|6639,6644
of|6645,6647
small|6648,6653
bowel|6654,6659
may|6660,6663
represent|6664,6673
ileus|6674,6679
or|6680,6682
<EOL>|6683,6684
obstruction|6684,6695
.|6695,6696
Dedicated|6697,6706
abdominal|6707,6716
radiograph|6717,6727
may|6728,6731
be|6732,6734
performed|6735,6744
for|6745,6748
<EOL>|6749,6750
better|6750,6756
characterization|6757,6773
.|6773,6774
<EOL>|6774,6775
<EOL>|6775,6776
ECHO|6776,6780
(|6781,6782
_|6782,6783
_|6783,6784
_|6784,6785
)|6785,6786
:|6786,6787
<EOL>|6787,6788
Left|6788,6792
ventricular|6793,6804
wall|6805,6809
thicknesses|6810,6821
are|6822,6825
normal|6826,6832
.|6832,6833
Left|6834,6838
ventricular|6839,6850
<EOL>|6851,6852
systolic|6852,6860
function|6861,6869
is|6870,6872
hyperdynamic|6873,6885
(|6886,6887
EF|6887,6889
>|6889,6890
75|6890,6892
%|6892,6893
)|6893,6894
.|6894,6895
There|6896,6901
is|6902,6904
a|6905,6906
mild|6907,6911
<EOL>|6912,6913
resting|6913,6920
left|6921,6925
ventricular|6926,6937
outflow|6938,6945
tract|6946,6951
obstruction|6952,6963
.|6963,6964
Right|6965,6970
<EOL>|6971,6972
ventricular|6972,6983
chamber|6984,6991
size|6992,6996
and|6997,7000
free|7001,7005
wall|7006,7010
motion|7011,7017
are|7018,7021
normal|7022,7028
.|7028,7029
The|7030,7033
<EOL>|7034,7035
aortic|7035,7041
valve|7042,7047
leaflets|7048,7056
(|7057,7058
3|7058,7059
)|7059,7060
are|7061,7064
mildly|7065,7071
thickened|7072,7081
.|7081,7082
The|7083,7086
mitral|7087,7093
valve|7094,7099
<EOL>|7100,7101
leaflets|7101,7109
are|7110,7113
mildly|7114,7120
thickened|7121,7130
.|7130,7131
There|7132,7137
is|7138,7140
severe|7141,7147
mitral|7148,7154
annular|7155,7162
<EOL>|7163,7164
calcification|7164,7177
.|7177,7178
There|7179,7184
is|7185,7187
moderate|7188,7196
functional|7197,7207
mitral|7208,7214
stenosis|7215,7223
<EOL>|7224,7225
(|7225,7226
mean|7226,7230
gradient|7231,7239
XXmmHg|7240,7246
)|7246,7247
due|7248,7251
to|7252,7254
mitral|7255,7261
annular|7262,7269
calcification|7270,7283
.|7283,7284
Mild|7285,7289
<EOL>|7290,7291
to|7291,7293
moderate|7294,7302
(|7303,7304
_|7304,7305
_|7305,7306
_|7306,7307
)|7307,7308
mitral|7309,7315
regurgitation|7316,7329
is|7330,7332
seen|7333,7337
.|7337,7338
[|7339,7340
Due|7340,7343
to|7344,7346
<EOL>|7347,7348
acoustic|7348,7356
shadowing|7357,7366
,|7366,7367
the|7368,7371
severity|7372,7380
of|7381,7383
mitral|7384,7390
regurgitation|7391,7404
may|7405,7408
be|7409,7411
<EOL>|7412,7413
significantly|7413,7426
UNDERestimated|7427,7441
.|7441,7442
]|7442,7443
The|7444,7447
left|7448,7452
ventricular|7453,7464
inflow|7465,7471
<EOL>|7472,7473
pattern|7473,7480
suggests|7481,7489
impaired|7490,7498
relaxation|7499,7509
.|7509,7510
The|7511,7514
tricuspid|7515,7524
valve|7525,7530
<EOL>|7531,7532
leaflets|7532,7540
are|7541,7544
mildly|7545,7551
thickened|7552,7561
.|7561,7562
Moderate|7563,7571
[|7572,7573
2|7573,7574
+|7574,7575
]|7575,7576
tricuspid|7577,7586
<EOL>|7587,7588
regurgitation|7588,7601
is|7602,7604
seen|7605,7609
.|7609,7610
There|7611,7616
is|7617,7619
mild|7620,7624
pulmonary|7625,7634
artery|7635,7641
systolic|7642,7650
<EOL>|7651,7652
hypertension|7652,7664
.|7664,7665
There|7666,7671
is|7672,7674
no|7675,7677
pericardial|7678,7689
effusion|7690,7698
.|7698,7699
<EOL>|7699,7700
<EOL>|7700,7701
Compared|7701,7709
with|7710,7714
the|7715,7718
prior|7719,7724
study|7725,7730
(|7731,7732
images|7732,7738
reviewed|7739,7747
)|7747,7748
of|7749,7751
_|7752,7753
_|7753,7754
_|7754,7755
,|7755,7756
<EOL>|7757,7758
mitral|7758,7764
regurgitation|7765,7778
is|7779,7781
now|7782,7785
less|7786,7790
prominent|7791,7800
.|7800,7801
The|7802,7805
mitral|7806,7812
inflow|7813,7819
<EOL>|7820,7821
gradient|7821,7829
is|7830,7832
similar|7833,7840
(|7841,7842
although|7842,7850
not|7851,7854
reported|7855,7863
in|7864,7866
the|7867,7870
previous|7871,7879
<EOL>|7880,7881
report|7881,7887
)|7887,7888
.|7888,7889
<EOL>|7890,7891
<EOL>|7891,7892
AXR|7892,7895
(|7896,7897
_|7897,7898
_|7898,7899
_|7899,7900
)|7900,7901
:|7901,7902
<EOL>|7902,7903
There|7903,7908
is|7909,7911
no|7912,7914
subdiaphragmatic|7915,7931
free|7932,7936
air|7937,7940
.|7940,7941
There|7943,7948
are|7949,7952
multiple|7953,7961
<EOL>|7962,7963
distended|7963,7972
loops|7973,7978
of|7979,7981
bowel|7982,7987
,|7987,7988
most|7989,7993
likely|7994,8000
representing|8001,8013
both|8014,8018
colon|8019,8024
<EOL>|8025,8026
and|8026,8029
small|8030,8035
bowel|8036,8041
.|8041,8042
Findings|8044,8052
are|8053,8056
most|8057,8061
consistent|8062,8072
with|8073,8077
an|8078,8080
ileus|8081,8086
.|8086,8087
<EOL>|8089,8090
Air|8090,8093
-|8093,8094
fluid|8094,8099
levels|8100,8106
are|8107,8110
seen|8111,8115
on|8116,8118
the|8119,8122
left|8123,8127
lateral|8128,8135
decubitus|8136,8145
view|8146,8150
.|8150,8151
<EOL>|8151,8152
IMPRESSION|8152,8162
:|8162,8163
Dilated|8165,8172
colon|8173,8178
and|8179,8182
small|8183,8188
bowel|8189,8194
consistent|8195,8205
with|8206,8210
<EOL>|8211,8212
ileus|8212,8217
.|8217,8218
<EOL>|8218,8219
<EOL>|8219,8220
Head|8220,8224
CT|8225,8227
(|8228,8229
_|8229,8230
_|8230,8231
_|8231,8232
)|8232,8233
:|8233,8234
IMPRESSION|8235,8245
:|8245,8246
No|8248,8250
acute|8251,8256
intracranial|8257,8269
process|8270,8277
.|8277,8278
<EOL>|8278,8279
<EOL>|8279,8280
ECHO|8280,8284
(|8285,8286
_|8286,8287
_|8287,8288
_|8288,8289
)|8289,8290
:|8290,8291
<EOL>|8291,8292
The|8292,8295
left|8296,8300
atrium|8301,8307
is|8308,8310
normal|8311,8317
in|8318,8320
size|8321,8325
.|8325,8326
There|8327,8332
is|8333,8335
mild|8336,8340
symmetric|8341,8350
left|8351,8355
<EOL>|8356,8357
ventricular|8357,8368
hypertrophy|8369,8380
.|8380,8381
The|8382,8385
left|8386,8390
ventricular|8391,8402
cavity|8403,8409
is|8410,8412
<EOL>|8413,8414
unusually|8414,8423
small|8424,8429
.|8429,8430
Left|8431,8435
ventricular|8436,8447
systolic|8448,8456
function|8457,8465
is|8466,8468
<EOL>|8469,8470
hyperdynamic|8470,8482
(|8483,8484
EF|8484,8486
80|8487,8489
%|8489,8490
)|8490,8491
.|8491,8492
Right|8493,8498
ventricular|8499,8510
chamber|8511,8518
size|8519,8523
and|8524,8527
free|8528,8532
<EOL>|8533,8534
wall|8534,8538
motion|8539,8545
are|8546,8549
normal|8550,8556
.|8556,8557
There|8558,8563
is|8564,8566
mild|8567,8571
aortic|8572,8578
valve|8579,8584
stenosis|8585,8593
<EOL>|8594,8595
(|8595,8596
valve|8596,8601
area|8602,8606
1.6|8607,8610
cm2|8611,8614
)|8614,8615
.|8615,8616
Due|8617,8620
to|8621,8623
the|8624,8627
technically|8628,8639
suboptimal|8640,8650
nature|8651,8657
<EOL>|8658,8659
of|8659,8661
this|8662,8666
study|8667,8672
,|8672,8673
LVOT|8674,8678
obstruction|8679,8690
can|8691,8694
not|8694,8697
be|8698,8700
excluded|8701,8709
with|8710,8714
<EOL>|8715,8716
certainty|8716,8725
.|8725,8726
The|8727,8730
mitral|8731,8737
valve|8738,8743
leaflets|8744,8752
are|8753,8756
mildly|8757,8763
thickened|8764,8773
.|8773,8774
There|8775,8780
<EOL>|8781,8782
is|8782,8784
severe|8785,8791
mitral|8792,8798
annular|8799,8806
calcification|8807,8820
(|8821,8822
can|8822,8825
not|8825,8828
exclude|8829,8836
posterior|8837,8846
<EOL>|8847,8848
leaflet|8848,8855
MVP|8856,8859
)|8859,8860
.|8860,8861
Moderate|8862,8870
(|8871,8872
2|8872,8873
+|8873,8874
)|8874,8875
mitral|8876,8882
regurgitation|8883,8896
is|8897,8899
seen|8900,8904
.|8904,8905
[|8906,8907
Due|8907,8910
<EOL>|8911,8912
to|8912,8914
acoustic|8915,8923
shadowing|8924,8933
,|8933,8934
the|8935,8938
severity|8939,8947
of|8948,8950
mitral|8951,8957
regurgitation|8958,8971
may|8972,8975
<EOL>|8976,8977
be|8977,8979
significantly|8980,8993
UNDERestimated|8994,9008
.|9008,9009
]|9009,9010
There|9011,9016
is|9017,9019
no|9020,9022
pericardial|9023,9034
<EOL>|9035,9036
effusion|9036,9044
.|9044,9045
<EOL>|9046,9047
<EOL>|9047,9048
Repeat|9048,9054
CT|9055,9057
Abd|9058,9061
/|9061,9062
Pelvis|9062,9068
(|9069,9070
_|9070,9071
_|9071,9072
_|9072,9073
)|9073,9074
:|9074,9075
<EOL>|9075,9076
IMPRESSION|9076,9086
:|9086,9087
Interval|9089,9097
increase|9098,9106
in|9107,9109
bilateral|9110,9119
pleural|9120,9127
effusions|9128,9137
,|9137,9138
<EOL>|9139,9140
and|9140,9143
in|9144,9146
<EOL>|9147,9148
abdominal|9148,9157
ascites|9158,9165
.|9165,9166
The|9168,9171
colon|9172,9177
remains|9178,9185
dilated|9186,9193
and|9194,9197
ahaustral|9198,9207
,|9207,9208
in|9209,9211
<EOL>|9212,9213
keeping|9213,9220
with|9221,9225
C.|9226,9228
difficile|9229,9238
colitis|9239,9246
.|9246,9247
<EOL>|9248,9249
<EOL>|9249,9250
CXR|9250,9253
(|9254,9255
_|9255,9256
_|9256,9257
_|9257,9258
)|9258,9259
:|9259,9260
<EOL>|9260,9261
There|9261,9266
is|9267,9269
a|9270,9271
Dobbhoff|9272,9280
tube|9281,9285
whose|9286,9291
distal|9292,9298
tip|9299,9302
is|9303,9305
in|9306,9308
the|9309,9312
body|9313,9317
of|9318,9320
the|9321,9324
<EOL>|9325,9326
stomach|9326,9333
.|9333,9334
<EOL>|9336,9337
There|9337,9342
are|9343,9346
bilateral|9347,9356
pleural|9357,9364
effusions|9365,9374
.|9374,9375
There|9377,9382
is|9383,9385
a|9386,9387
right|9388,9393
-|9393,9394
sided|9394,9399
<EOL>|9400,9401
pleural|9401,9408
-|9408,9409
based|9409,9414
catheter|9415,9423
.|9423,9424
There|9426,9431
is|9432,9434
no|9435,9437
pneumothoraces|9438,9452
or|9453,9455
signs|9456,9461
for|9462,9465
<EOL>|9466,9467
overt|9467,9472
pulmonary|9473,9482
edema|9483,9488
.|9488,9489
Overall|9491,9498
,|9498,9499
these|9500,9505
findings|9506,9514
are|9515,9518
stable|9519,9525
since|9526,9531
<EOL>|9532,9533
prior|9533,9538
study|9539,9544
from|9545,9549
_|9550,9551
_|9551,9552
_|9552,9553
.|9553,9554
<EOL>|9555,9556
<EOL>|9556,9557
<EOL>|9558,9559
Brief|9559,9564
Hospital|9565,9573
Course|9574,9580
:|9580,9581
<EOL>|9581,9582
Pt|9582,9584
is|9585,9587
an|9588,9590
_|9591,9592
_|9592,9593
_|9593,9594
year|9595,9599
-|9599,9600
old|9600,9603
woman|9604,9609
with|9610,9614
history|9615,9622
of|9623,9625
Sjogren|9626,9633
's|9633,9635
syndrome|9636,9644
<EOL>|9645,9646
and|9646,9649
IBS|9650,9653
presenting|9654,9664
with|9665,9669
fevers|9670,9676
,|9676,9677
diarrhea|9678,9686
,|9686,9687
tachycardia|9688,9699
,|9699,9700
<EOL>|9701,9702
hypotension|9702,9713
,|9713,9714
leukocytosis|9715,9727
,|9727,9728
hypoxia|9729,9736
,|9736,9737
found|9738,9743
to|9744,9746
have|9747,9751
pancolitis|9752,9762
and|9763,9766
<EOL>|9767,9768
pneumonia|9768,9777
.|9777,9778
<EOL>|9778,9779
<EOL>|9779,9780
#|9780,9781
Septic|9782,9788
Shock|9789,9794
due|9795,9798
to|9799,9801
Cdiff|9802,9807
Colitis|9808,9815
:|9815,9816
On|9817,9819
admission|9820,9829
meet|9830,9834
criteria|9835,9843
<EOL>|9844,9845
for|9845,9848
sepsis|9849,9855
given|9856,9861
fever|9862,9867
,|9867,9868
tachycardia|9869,9880
,|9880,9881
leukocytosis|9882,9894
and|9895,9898
likely|9899,9905
<EOL>|9906,9907
source|9907,9913
being|9914,9919
colitis|9920,9927
.|9927,9928
BP|9929,9931
remained|9932,9940
low|9941,9944
and|9945,9948
patient|9949,9956
remained|9957,9965
<EOL>|9966,9967
mildly|9967,9973
tachycardic|9974,9985
for|9986,9989
next|9990,9994
_|9995,9996
_|9996,9997
_|9997,9998
requiring|9999,10008
aggressive|10009,10019
IVF|10020,10023
<EOL>|10024,10025
(|10025,10026
roughly|10026,10033
20L|10034,10037
in|10038,10040
first|10041,10046
72hrs|10047,10052
)|10052,10053
.|10053,10054
Initially|10055,10064
started|10065,10072
on|10073,10075
IV|10076,10078
flagyl|10079,10085
/|10085,10086
PO|10086,10088
<EOL>|10089,10090
vanco|10090,10095
emperically|10096,10107
for|10108,10111
possible|10112,10120
Cdiff|10121,10126
as|10127,10129
well|10130,10134
as|10135,10137
levofloxacin|10138,10150
<EOL>|10151,10152
over|10152,10156
concern|10157,10164
for|10165,10168
PNA|10169,10172
.|10172,10173
Bcx|10174,10177
,|10177,10178
Ucx|10179,10182
unrevealing|10183,10194
.|10194,10195
Stool|10196,10201
for|10202,10205
Cdiff|10206,10211
<EOL>|10212,10213
ultimately|10213,10223
positive|10224,10232
and|10233,10236
levofloxacin|10237,10249
changed|10250,10257
to|10258,10260
CTX|10261,10264
/|10264,10265
Azithro|10265,10272
.|10272,10273
PCP|10274,10277
<EOL>|10278,10279
(|10279,10280
Dr|10280,10282
.|10282,10283
_|10284,10285
_|10285,10286
_|10286,10287
visited|10288,10295
and|10296,10299
said|10300,10304
that|10305,10309
pt|10310,10312
always|10313,10319
has|10320,10323
CXR|10324,10327
infiltrate|10328,10338
<EOL>|10339,10340
so|10340,10342
abx|10343,10346
for|10347,10350
CTX|10351,10354
/|10354,10355
Azithro|10355,10362
for|10363,10366
pneumonia|10367,10376
stopped|10377,10384
after|10385,10390
pt|10391,10393
had|10394,10397
<EOL>|10398,10399
received|10399,10407
total|10408,10413
of|10414,10416
3|10417,10418
days|10419,10423
PNA|10424,10427
treatment|10428,10437
.|10437,10438
Lactate|10439,10446
and|10447,10450
WBC|10451,10454
count|10455,10460
<EOL>|10461,10462
trended|10462,10469
up|10470,10472
in|10473,10475
first|10476,10481
48hrs|10482,10487
and|10488,10491
patient|10492,10499
developed|10500,10509
ileus|10510,10515
on|10516,10518
<EOL>|10519,10520
abdominal|10520,10529
imaging|10530,10537
with|10538,10542
worsening|10543,10552
distension|10553,10563
.|10563,10564
GI|10565,10567
and|10568,10571
Gen|10572,10575
Surg|10576,10580
<EOL>|10581,10582
followed|10582,10590
and|10591,10594
pt|10595,10597
kept|10598,10602
NPO|10603,10606
initially|10607,10616
,|10616,10617
but|10618,10621
ultimately|10622,10632
illness|10633,10640
<EOL>|10641,10642
turned|10642,10648
around|10649,10655
with|10656,10660
just|10661,10665
Abx|10666,10669
and|10670,10673
IVF|10674,10677
.|10677,10678
By|10679,10681
time|10682,10686
of|10687,10689
ICU|10690,10693
call|10694,10698
-|10698,10699
out|10699,10702
,|10702,10703
BP|10704,10706
<EOL>|10707,10708
had|10708,10711
stabilized|10712,10722
without|10723,10730
requiring|10731,10740
fluids|10741,10747
and|10748,10751
abdominal|10752,10761
exam|10762,10766
was|10767,10770
<EOL>|10771,10772
improving|10772,10781
with|10782,10786
downtrending|10787,10799
WBC|10800,10803
.|10803,10804
Came|10805,10809
back|10810,10814
to|10815,10817
ICU|10818,10821
on|10822,10824
_|10825,10826
_|10826,10827
_|10827,10828
due|10829,10832
to|10833,10835
<EOL>|10836,10837
respiratory|10837,10848
distress|10849,10857
and|10858,10861
hypoxia|10862,10869
.|10869,10870
Also|10871,10875
had|10876,10879
to|10880,10882
be|10883,10885
started|10886,10893
back|10894,10898
on|10899,10901
<EOL>|10902,10903
pressors|10903,10911
,|10911,10912
initially|10913,10922
phenylephrine|10923,10936
but|10937,10940
then|10941,10945
this|10946,10950
was|10951,10954
stopped|10955,10962
as|10963,10965
<EOL>|10966,10967
extremities|10967,10978
were|10979,10983
cold|10984,10988
and|10989,10992
mottled|10993,11000
.|11000,11001
Pressors|11002,11010
changed|11011,11018
to|11019,11021
<EOL>|11022,11023
Norepinephrine|11023,11037
and|11038,11041
mottling|11042,11050
of|11051,11053
ext|11054,11057
quickly|11058,11065
resolved|11066,11074
.|11074,11075
SVO2|11076,11080
and|11081,11084
<EOL>|11085,11086
ECHO|11086,11090
not|11091,11094
consistent|11095,11105
with|11106,11110
cardiogenic|11111,11122
shock|11123,11128
and|11129,11132
EKG|11133,11136
/|11136,11137
Trops|11137,11142
were|11143,11147
<EOL>|11148,11149
negative|11149,11157
.|11157,11158
ID|11159,11161
saw|11162,11165
in|11166,11168
consult|11169,11176
and|11177,11180
recommended|11181,11192
starting|11193,11201
Tigecycline|11202,11213
<EOL>|11214,11215
to|11215,11217
help|11218,11222
cover|11223,11228
Cdiff|11229,11234
which|11235,11240
she|11241,11244
completed|11245,11254
an|11255,11257
8|11258,11259
day|11260,11263
course|11264,11270
of|11271,11273
.|11273,11274
<EOL>|11275,11276
Abdominal|11276,11285
exam|11286,11290
improved|11291,11299
and|11300,11303
ileus|11304,11309
resolved|11310,11318
.|11318,11319
Doboff|11320,11326
was|11327,11330
placed|11331,11337
on|11338,11340
<EOL>|11341,11342
_|11342,11343
_|11343,11344
_|11344,11345
and|11346,11349
tube|11350,11354
feeds|11355,11360
were|11361,11365
started|11366,11373
due|11374,11377
poor|11378,11382
ability|11383,11390
to|11391,11393
keep|11394,11398
with|11399,11403
<EOL>|11404,11405
with|11405,11409
nutritional|11410,11421
requirements|11422,11434
.|11434,11435
Metronidazole|11436,11449
d|11450,11451
/|11451,11452
c|11452,11453
'd|11453,11455
on|11456,11458
_|11459,11460
_|11460,11461
_|11461,11462
.|11462,11463
Plan|11464,11468
<EOL>|11469,11470
to|11470,11472
continue|11473,11481
Vancomycin|11482,11492
500mg|11493,11498
PO|11499,11501
Q6|11502,11504
for|11505,11508
a|11509,11510
total|11511,11516
of|11517,11519
2|11520,11521
weeks|11522,11527
after|11528,11533
<EOL>|11534,11535
all|11535,11538
other|11539,11544
antibiotics|11545,11556
were|11557,11561
stopped|11562,11569
(|11570,11571
last|11571,11575
day|11576,11579
_|11580,11581
_|11581,11582
_|11582,11583
.|11583,11584
<EOL>|11584,11585
<EOL>|11585,11586
#|11586,11587
Hypoxia|11588,11595
:|11595,11596
No|11597,11599
breathing|11600,11609
issues|11610,11616
at|11617,11619
baseline|11620,11628
but|11629,11632
developed|11633,11642
hypoxia|11643,11650
<EOL>|11651,11652
requiring|11652,11661
5L|11662,11664
NC|11665,11667
while|11668,11673
in|11674,11676
ED|11677,11679
so|11680,11682
was|11683,11686
admitted|11687,11695
to|11696,11698
the|11699,11702
ICU|11703,11706
.|11706,11707
Initial|11708,11715
<EOL>|11716,11717
concern|11717,11724
for|11725,11728
RLL|11729,11732
PNA|11733,11736
on|11737,11739
CXR|11740,11743
and|11744,11747
received|11748,11756
3|11757,11758
days|11759,11763
of|11764,11766
Abx|11767,11770
as|11771,11773
noted|11774,11779
<EOL>|11780,11781
above|11781,11786
until|11787,11792
PCP|11793,11796
informed|11797,11805
MICU|11806,11810
team|11811,11815
that|11816,11820
infiltrate|11821,11831
had|11832,11835
been|11836,11840
<EOL>|11841,11842
present|11842,11849
for|11850,11853
some|11854,11858
time|11859,11863
.|11863,11864
Thought|11865,11872
that|11873,11877
hypoxia|11878,11885
developed|11886,11895
in|11896,11898
setting|11899,11906
<EOL>|11907,11908
of|11908,11910
aggressive|11911,11921
fluids|11922,11928
in|11929,11931
patient|11932,11939
with|11940,11944
significant|11945,11956
mitral|11957,11963
regurg|11964,11970
<EOL>|11971,11972
(|11972,11973
got|11973,11976
4L|11977,11979
in|11980,11982
ED|11983,11985
and|11986,11989
then|11990,11994
aggressive|11995,12005
IVF|12006,12009
in|12010,12012
first|12013,12018
72hrs|12019,12024
)|12024,12025
and|12026,12029
the|12030,12033
<EOL>|12034,12035
development|12035,12046
of|12047,12049
pleural|12050,12057
effusions|12058,12067
.|12067,12068
Had|12069,12072
started|12073,12080
diuresis|12081,12089
by|12090,12092
MICU|12093,12097
<EOL>|12098,12099
callout|12099,12106
on|12107,12109
_|12110,12111
_|12111,12112
_|12112,12113
but|12114,12117
then|12118,12122
after|12123,12128
couple|12129,12135
days|12136,12140
on|12141,12143
floor|12144,12149
,|12149,12150
triggered|12151,12160
<EOL>|12161,12162
for|12162,12165
hypoxia|12166,12173
and|12174,12177
increased|12178,12187
work|12188,12192
of|12193,12195
breathing|12196,12205
on|12206,12208
_|12209,12210
_|12210,12211
_|12211,12212
.|12212,12213
Found|12214,12219
to|12220,12222
<EOL>|12223,12224
have|12224,12228
significant|12229,12240
worsening|12241,12250
of|12251,12253
R|12254,12255
pleural|12256,12263
effusion|12264,12272
and|12273,12276
development|12277,12288
<EOL>|12289,12290
of|12290,12292
L|12293,12294
pleural|12295,12302
effusion|12303,12311
.|12311,12312
Required|12313,12321
intubation|12322,12332
for|12333,12336
respiratory|12337,12348
state|12349,12354
<EOL>|12355,12356
on|12356,12358
_|12359,12360
_|12360,12361
_|12361,12362
.|12362,12363
Cardiac|12364,12371
w|12372,12373
/|12373,12374
u|12374,12375
showed|12376,12382
no|12383,12385
cardiogenic|12386,12397
component|12398,12407
and|12408,12411
when|12412,12416
<EOL>|12417,12418
spiked|12418,12424
fever|12425,12430
on|12431,12433
_|12434,12435
_|12435,12436
_|12436,12437
started|12438,12445
on|12446,12448
empiric|12449,12456
HCAP|12457,12461
coverage|12462,12470
after|12471,12476
<EOL>|12477,12478
mini-BAL|12478,12486
was|12487,12490
performed|12491,12500
.|12500,12501
Interventional|12502,12516
pulmonary|12517,12526
(|12527,12528
IP|12528,12530
)|12530,12531
consulted|12532,12541
<EOL>|12542,12543
on|12543,12545
_|12546,12547
_|12547,12548
_|12548,12549
and|12550,12553
performed|12554,12563
right|12564,12569
sided|12570,12575
thoracentesis|12576,12589
with|12590,12594
pigtail|12595,12602
<EOL>|12603,12604
placement|12604,12613
.|12613,12614
ID|12615,12617
saw|12618,12621
on|12622,12624
_|12625,12626
_|12626,12627
_|12627,12628
and|12629,12632
recommended|12633,12644
stopping|12645,12653
<EOL>|12654,12655
Vanco|12655,12660
/|12660,12661
cefepime|12661,12669
as|12670,12672
unclear|12673,12680
if|12681,12683
actual|12684,12690
pneumonia|12691,12700
and|12701,12704
starting|12705,12713
<EOL>|12714,12715
Tigecycline|12715,12726
as|12727,12729
would|12730,12735
cover|12736,12741
many|12742,12746
HCAP|12747,12751
organisms|12752,12761
and|12762,12765
also|12766,12770
treat|12771,12776
<EOL>|12777,12778
Cdiff|12778,12783
.|12783,12784
Mini-BAL|12785,12793
and|12794,12797
pleural|12798,12805
fluid|12806,12811
with|12812,12816
negative|12817,12825
cultures|12826,12834
.|12834,12835
<EOL>|12836,12837
Started|12837,12844
diuresis|12845,12853
again|12854,12859
on|12860,12862
_|12863,12864
_|12864,12865
_|12865,12866
as|12867,12869
she|12870,12873
was|12874,12877
weaned|12878,12884
off|12885,12888
pressors|12889,12897
<EOL>|12898,12899
and|12899,12902
extubated|12903,12912
.|12912,12913
She|12914,12917
was|12918,12921
weaned|12922,12928
off|12929,12932
all|12933,12936
oxygen|12937,12943
at|12944,12946
the|12947,12950
time|12951,12955
of|12956,12958
<EOL>|12959,12960
discharge|12960,12969
and|12970,12973
right|12974,12979
pigtail|12980,12987
still|12988,12993
draining|12994,13002
400|13003,13006
-|13006,13007
700cc|13007,13012
per|13013,13016
day|13017,13020
,|13020,13021
<EOL>|13022,13023
will|13023,13027
follow|13028,13034
-|13034,13035
up|13035,13037
with|13038,13042
IP|13043,13045
after|13046,13051
discharge|13052,13061
.|13061,13062
She|13064,13067
will|13068,13072
require|13073,13080
<EOL>|13081,13082
ongoing|13082,13089
diuresis|13090,13098
given|13099,13104
her|13105,13108
significant|13109,13120
volume|13121,13127
overload|13128,13136
,|13136,13137
she|13138,13141
<EOL>|13142,13143
responds|13143,13151
well|13152,13156
to|13157,13159
_|13160,13161
_|13161,13162
_|13162,13163
IV|13164,13166
Lasix|13167,13172
and|13173,13176
had|13177,13180
been|13181,13185
_|13186,13187
_|13187,13188
_|13188,13189
negative|13190,13198
<EOL>|13199,13200
in|13200,13202
the|13203,13206
days|13207,13211
leading|13212,13219
up|13220,13222
to|13223,13225
discharge|13226,13235
.|13235,13236
<EOL>|13236,13237
<EOL>|13237,13238
#|13238,13239
Altered|13240,13247
Mental|13248,13254
Status|13255,13261
:|13261,13262
<EOL>|13263,13264
In|13264,13266
setting|13267,13274
of|13275,13277
trigger|13278,13285
for|13286,13289
hypoxia|13290,13297
and|13298,13301
MICU|13302,13306
transfer|13307,13315
on|13316,13318
_|13319,13320
_|13320,13321
_|13321,13322
,|13322,13323
<EOL>|13324,13325
there|13325,13330
was|13331,13334
concern|13335,13342
that|13343,13347
she|13348,13351
was|13352,13355
less|13356,13360
responsive|13361,13371
with|13372,13376
concern|13377,13384
for|13385,13388
<EOL>|13389,13390
focal|13390,13395
defecits|13396,13404
.|13404,13405
Stat|13406,13410
head|13411,13415
CT|13416,13418
without|13419,13426
evidence|13427,13435
of|13436,13438
stroke|13439,13445
or|13446,13448
<EOL>|13449,13450
bleed|13450,13455
.|13455,13456
Neuro|13457,13462
was|13463,13466
consulted|13467,13476
and|13477,13480
said|13481,13485
nothing|13486,13493
to|13494,13496
do|13497,13499
and|13500,13503
deficits|13504,13512
<EOL>|13513,13514
resolved|13514,13522
over|13523,13527
next|13528,13532
_|13533,13534
_|13534,13535
_|13535,13536
.|13536,13537
EEG|13538,13541
initially|13542,13551
ordered|13552,13559
but|13560,13563
then|13564,13568
<EOL>|13569,13570
canceled|13570,13578
after|13579,13584
discussion|13585,13595
with|13596,13600
neuro|13601,13606
.|13606,13607
Rest|13608,13612
of|13613,13615
ICU|13616,13619
stay|13620,13624
had|13625,13628
<EOL>|13629,13630
intermittent|13630,13642
delerium|13643,13651
in|13652,13654
the|13655,13658
evenings|13659,13667
requiring|13668,13677
some|13678,13682
doses|13683,13688
of|13689,13691
<EOL>|13692,13693
Olanzapine|13693,13703
.|13703,13704
Delerium|13705,13713
had|13714,13717
improved|13718,13726
by|13727,13729
time|13730,13734
of|13735,13737
ICU|13738,13741
callout|13742,13749
but|13750,13753
<EOL>|13754,13755
still|13755,13760
with|13761,13765
some|13766,13770
sundowning|13771,13781
.|13781,13782
<EOL>|13782,13783
<EOL>|13783,13784
#|13784,13785
Hyponatremia|13786,13798
:|13798,13799
Patient|13800,13807
with|13808,13812
Na|13813,13815
of|13816,13818
127|13819,13822
in|13823,13825
ED|13826,13828
.|13828,13829
Likely|13830,13836
hypovolemic|13837,13848
<EOL>|13849,13850
hyponatremia|13850,13862
in|13863,13865
setting|13866,13873
of|13874,13876
diarrhea|13877,13885
/|13885,13886
poor|13886,13890
PO|13891,13893
intake|13894,13900
.|13900,13901
Could|13902,13907
also|13908,13912
<EOL>|13913,13914
be|13914,13916
SIADH|13917,13922
given|13923,13928
pneumonia|13929,13938
,|13938,13939
pain|13940,13944
.|13944,13945
Upon|13946,13950
review|13951,13957
of|13958,13960
old|13961,13964
labs|13965,13969
,|13969,13970
patient|13971,13978
<EOL>|13979,13980
often|13980,13985
hyponatremic|13986,13998
as|13999,14001
outpatient|14002,14012
as|14013,14015
well|14016,14020
.|14020,14021
Urine|14022,14027
lytes|14028,14033
confusing|14034,14043
<EOL>|14044,14045
in|14045,14047
setting|14048,14055
of|14056,14058
shock|14059,14064
as|14065,14067
urine|14068,14073
Na|14074,14076
elevated|14077,14085
in|14086,14088
_|14089,14090
_|14090,14091
_|14091,14092
so|14093,14095
some|14096,14100
question|14101,14109
<EOL>|14110,14111
of|14111,14113
sodium|14114,14120
wasting|14121,14128
renal|14129,14134
injury|14135,14141
.|14141,14142
Hyponatremia|14143,14155
started|14156,14163
to|14164,14166
resolve|14167,14174
<EOL>|14175,14176
as|14176,14178
overall|14179,14186
condition|14187,14196
improved|14197,14205
and|14206,14209
did|14210,14213
not|14214,14217
re-develop|14218,14228
even|14229,14233
in|14234,14236
<EOL>|14237,14238
setting|14238,14245
of|14246,14248
_|14249,14250
_|14250,14251
_|14251,14252
ICU|14253,14256
readmission|14257,14268
for|14269,14272
hypoxia|14273,14280
.|14280,14281
<EOL>|14281,14282
<EOL>|14282,14283
#|14283,14284
_|14285,14286
_|14286,14287
_|14287,14288
:|14288,14289
Patient|14290,14297
with|14298,14302
creatinine|14303,14313
of|14314,14316
1.1|14317,14320
at|14321,14323
admission|14324,14333
up|14334,14336
from|14337,14341
<EOL>|14342,14343
recent|14343,14349
baseline|14350,14358
of|14359,14361
0.7|14362,14365
-|14366,14367
0.8|14368,14371
.|14371,14372
Likely|14373,14379
pre-renal|14380,14389
etiology|14390,14398
in|14399,14401
<EOL>|14402,14403
setting|14403,14410
of|14411,14413
infection|14414,14423
,|14423,14424
diarrhea|14425,14433
,|14433,14434
poor|14435,14439
PO|14440,14442
intake|14443,14449
.|14449,14450
Trended|14451,14458
up|14459,14461
<EOL>|14462,14463
slightly|14463,14471
to|14472,14474
1.3|14475,14478
after|14479,14484
a|14485,14486
few|14487,14490
days|14491,14495
likely|14496,14502
with|14503,14507
mild|14508,14512
ATN|14513,14516
in|14517,14519
setting|14520,14527
<EOL>|14528,14529
of|14529,14531
persistent|14532,14542
boarderline|14543,14554
hypotension|14555,14566
.|14566,14567
Lisinopril|14568,14578
was|14579,14582
held|14583,14587
while|14588,14593
<EOL>|14594,14595
in|14595,14597
ICU|14598,14601
for|14602,14605
this|14606,14610
and|14611,14614
hypotension|14615,14626
.|14626,14627
Cr|14628,14630
trended|14631,14638
back|14639,14643
down|14644,14648
to|14649,14651
roughly|14652,14659
<EOL>|14660,14661
0.5|14661,14664
and|14665,14668
stayed|14669,14675
there|14676,14681
for|14682,14685
rest|14686,14690
of|14691,14693
hospitalization|14694,14709
even|14710,14714
in|14715,14717
setting|14718,14725
<EOL>|14726,14727
of|14727,14729
second|14730,14736
ICU|14737,14740
readmission|14741,14752
.|14752,14753
<EOL>|14753,14754
<EOL>|14754,14755
-|14755,14756
-|14756,14757
Inactive|14757,14765
issues|14766,14772
-|14772,14773
-|14773,14774
<EOL>|14774,14775
<EOL>|14775,14776
#|14776,14777
Hypothyroidism|14778,14792
:|14792,14793
Continued|14794,14803
levothyroxine|14804,14817
50|14818,14820
mcg|14821,14824
daily|14825,14830
<EOL>|14830,14831
<EOL>|14831,14832
#|14832,14833
Hypertension|14834,14846
:|14846,14847
Due|14848,14851
to|14852,14854
hypotension|14855,14866
with|14867,14871
sepsis|14872,14878
,|14878,14879
lisinopril|14880,14890
was|14891,14894
<EOL>|14895,14896
held|14896,14900
.|14900,14901
BP|14903,14905
remained|14906,14914
well|14915,14919
controlled|14920,14930
and|14931,14934
this|14935,14939
will|14940,14944
continue|14945,14953
to|14954,14956
be|14957,14959
<EOL>|14960,14961
held|14961,14965
at|14966,14968
discharge|14969,14978
.|14978,14979
<EOL>|14979,14980
<EOL>|14980,14981
#|14981,14982
GERD|14983,14987
:|14987,14988
Omeprazole|14989,14999
stopped|15000,15007
when|15008,15012
Cdiff|15013,15018
came|15019,15023
back|15024,15028
positive|15029,15037
.|15037,15038
For|15039,15042
<EOL>|15043,15044
time|15044,15048
was|15049,15052
put|15053,15056
on|15057,15059
H2|15060,15062
blocker|15063,15070
for|15071,15074
GI|15075,15077
prophylaxis|15078,15089
but|15090,15093
this|15094,15098
stopped|15099,15106
<EOL>|15107,15108
again|15108,15113
when|15114,15118
delerious|15119,15128
and|15129,15132
started|15133,15140
feeeding|15141,15149
.|15149,15150
<EOL>|15150,15151
<EOL>|15151,15152
#|15152,15153
Code|15154,15158
:|15158,15159
Full|15160,15164
(|15165,15166
confirmed|15166,15175
with|15176,15180
patient|15181,15188
,|15188,15189
son|15190,15193
-|15193,15194
in|15194,15196
-|15196,15197
law|15197,15200
)|15200,15201
<EOL>|15201,15202
<EOL>|15202,15203
#|15203,15204
Transitional|15205,15217
issues|15218,15224
<EOL>|15224,15225
-|15225,15226
Right|15226,15231
pigtail|15232,15239
pleural|15240,15247
catheter|15248,15256
in|15257,15259
place|15260,15265
at|15266,15268
discharge|15269,15278
,|15278,15279
she|15280,15283
will|15284,15288
<EOL>|15289,15290
follow|15290,15296
-|15296,15297
up|15297,15299
with|15300,15304
interventional|15305,15319
pulmonary|15320,15329
after|15330,15335
discharge|15336,15345
.|15345,15346
Tube|15347,15351
<EOL>|15352,15353
can|15353,15356
be|15357,15359
removed|15360,15367
when|15368,15372
output|15373,15379
is|15380,15382
<|15383,15384
200cc|15384,15389
per|15390,15393
day|15394,15397
.|15397,15398
<EOL>|15398,15399
-|15399,15400
Will|15400,15404
need|15405,15409
ongoing|15410,15417
diuresis|15418,15426
given|15427,15432
large|15433,15438
volume|15439,15445
of|15446,15448
fluids|15449,15455
she|15456,15459
<EOL>|15460,15461
received|15461,15469
in|15470,15472
the|15473,15476
ICU|15477,15480
this|15481,15485
admission|15486,15495
,|15495,15496
she|15497,15500
responds|15501,15509
well|15510,15514
to|15515,15517
Lasix|15518,15523
<EOL>|15524,15525
10mg|15525,15529
IV|15530,15532
.|15532,15533
Goal|15534,15538
_|15539,15540
_|15540,15541
_|15541,15542
negative|15543,15551
as|15552,15554
BP|15555,15557
tolerates|15558,15567
.|15567,15568
<EOL>|15568,15569
-|15569,15570
Will|15570,15574
continue|15575,15583
on|15584,15586
high|15587,15591
dose|15592,15596
PO|15597,15599
vancomycin|15600,15610
through|15611,15618
_|15619,15620
_|15620,15621
_|15621,15622
(|15623,15624
_|15624,15625
_|15625,15626
_|15626,15627
fter|15627,15631
other|15632,15637
abx|15638,15641
stopped|15642,15649
)|15649,15650
<EOL>|15650,15651
-|15651,15652
She|15652,15655
should|15656,15662
continue|15663,15671
tube|15672,15676
feeds|15677,15682
until|15683,15688
taking|15689,15695
adequate|15696,15704
PO|15705,15707
,|15707,15708
would|15709,15714
<EOL>|15715,15716
benefit|15716,15723
from|15724,15728
ongoing|15729,15736
nutrition|15737,15746
evaluation|15747,15757
<EOL>|15757,15758
<EOL>|15759,15760
Medications|15760,15771
on|15772,15774
Admission|15775,15784
:|15784,15785
<EOL>|15785,15786
fluticasone|15786,15797
50|15798,15800
mcg|15801,15804
1|15805,15806
-|15807,15808
2|15809,15810
nasal|15811,15816
sprays|15817,15823
BID|15824,15827
PRN|15828,15831
allergies|15832,15841
<EOL>|15841,15842
levothyroxine|15842,15855
50|15856,15858
mcg|15859,15862
daily|15863,15868
<EOL>|15868,15869
lisinopril|15869,15879
10|15880,15882
mg|15883,15885
daily|15886,15891
<EOL>|15891,15892
tiotropum|15892,15901
bromide|15902,15909
18|15910,15912
mcg|15913,15916
daily|15917,15922
<EOL>|15922,15923
Calcium|15923,15930
<EOL>|15930,15931
multivitamin|15931,15943
<EOL>|15943,15944
omeprazole|15944,15954
20|15955,15957
mg|15958,15960
daily|15961,15966
<EOL>|15966,15967
acetaminophen|15967,15980
PRN|15981,15984
pain|15985,15989
<EOL>|15990,15991
<EOL>|15992,15993
Discharge|15993,16002
Medications|16003,16014
:|16014,16015
<EOL>|16015,16016
1.|16016,16018
fluticasone|16019,16030
50|16031,16033
mcg|16034,16037
/|16037,16038
actuation|16038,16047
Spray|16048,16053
,|16053,16054
Suspension|16055,16065
Sig|16066,16069
:|16069,16070
_|16071,16072
_|16072,16073
_|16073,16074
puffs|16075,16080
<EOL>|16081,16082
Nasal|16082,16087
twice|16088,16093
a|16094,16095
day|16096,16099
as|16100,16102
needed|16103,16109
for|16110,16113
allergies|16114,16123
.|16123,16124
<EOL>|16126,16127
2.|16127,16129
levothyroxine|16130,16143
50|16144,16146
mcg|16147,16150
Tablet|16151,16157
Sig|16158,16161
:|16161,16162
One|16163,16166
(|16167,16168
1|16168,16169
)|16169,16170
Tablet|16171,16177
PO|16178,16180
DAILY|16181,16186
<EOL>|16187,16188
(|16188,16189
Daily|16189,16194
)|16194,16195
.|16195,16196
<EOL>|16198,16199
3.|16199,16201
acetaminophen|16202,16215
325|16216,16219
mg|16220,16222
Tablet|16223,16229
Sig|16230,16233
:|16233,16234
_|16235,16236
_|16236,16237
_|16237,16238
Tablets|16239,16246
PO|16247,16249
every|16250,16255
four|16256,16260
<EOL>|16261,16262
(|16262,16263
4|16263,16264
)|16264,16265
hours|16266,16271
as|16272,16274
needed|16275,16281
for|16282,16285
pain|16286,16290
.|16290,16291
<EOL>|16293,16294
4.|16294,16296
polyvinyl|16297,16306
alcohol|16307,16314
1.4|16315,16318
%|16319,16320
Drops|16321,16326
Sig|16327,16330
:|16330,16331
One|16332,16335
(|16336,16337
1|16337,16338
)|16338,16339
drop|16340,16344
Ophthalmic|16345,16355
<EOL>|16356,16357
every|16357,16362
four|16363,16367
(|16368,16369
4|16369,16370
)|16370,16371
hours|16372,16377
as|16378,16380
needed|16381,16387
for|16388,16391
dry|16392,16395
eyes|16396,16400
.|16400,16401
<EOL>|16403,16404
5.|16404,16406
heparin|16407,16414
,|16414,16415
porcine|16416,16423
(|16424,16425
PF|16425,16427
)|16427,16428
10|16429,16431
unit|16432,16436
/|16436,16437
mL|16437,16439
Syringe|16440,16447
Sig|16448,16451
:|16451,16452
Two|16453,16456
(|16457,16458
2|16458,16459
)|16459,16460
ML|16461,16463
<EOL>|16464,16465
Intravenous|16465,16476
PRN|16477,16480
(|16481,16482
as|16482,16484
needed|16485,16491
)|16491,16492
as|16493,16495
needed|16496,16502
for|16503,16506
line|16507,16511
flush|16512,16517
.|16517,16518
<EOL>|16520,16521
6.|16521,16523
heparin|16524,16531
(|16532,16533
porcine|16533,16540
)|16540,16541
5,000|16542,16547
unit|16548,16552
/|16552,16553
mL|16553,16555
Solution|16556,16564
Sig|16565,16568
:|16568,16569
5000|16570,16574
(|16575,16576
5000|16576,16580
)|16580,16581
<EOL>|16582,16583
units|16583,16588
Injection|16589,16598
twice|16599,16604
a|16605,16606
day|16607,16610
.|16610,16611
<EOL>|16613,16614
7.|16614,16616
insulin|16617,16624
lispro|16625,16631
100|16632,16635
unit|16636,16640
/|16640,16641
mL|16641,16643
Solution|16644,16652
Sig|16653,16656
:|16656,16657
sliding|16658,16665
scale|16666,16671
units|16672,16677
<EOL>|16678,16679
Subcutaneous|16679,16691
three|16692,16697
times|16698,16703
a|16704,16705
day|16706,16709
:|16709,16710
Sliding|16711,16718
scale|16719,16724
:|16724,16725
<EOL>|16726,16727
150|16727,16730
-|16730,16731
200|16731,16734
-|16735,16736
2|16737,16738
units|16739,16744
;|16744,16745
<EOL>|16745,16746
201|16746,16749
-|16749,16750
250|16750,16753
-|16754,16755
4|16756,16757
units|16758,16763
;|16763,16764
<EOL>|16764,16765
251|16765,16768
-|16768,16769
300|16769,16772
-|16773,16774
6|16775,16776
units|16777,16782
;|16782,16783
<EOL>|16783,16784
301|16784,16787
-|16787,16788
350|16788,16791
-|16792,16793
8|16794,16795
units|16796,16801
;|16801,16802
<EOL>|16802,16803
351|16803,16806
-|16806,16807
400|16807,16810
-|16811,16812
10|16813,16815
units|16816,16821
;|16821,16822
<EOL>|16822,16823
over|16823,16827
400|16828,16831
-|16832,16833
10|16834,16836
units|16837,16842
and|16843,16846
call|16847,16851
MD|16852,16854
.|16854,16855
<EOL>|16857,16858
8.|16858,16860
miconazole|16861,16871
nitrate|16872,16879
2|16880,16881
%|16882,16883
Powder|16884,16890
Sig|16891,16894
:|16894,16895
One|16896,16899
(|16900,16901
1|16901,16902
)|16902,16903
Appl|16904,16908
Topical|16909,16916
TID|16917,16920
<EOL>|16921,16922
(|16922,16923
3|16923,16924
times|16925,16930
a|16931,16932
day|16933,16936
)|16936,16937
as|16938,16940
needed|16941,16947
for|16948,16951
rash|16952,16956
.|16956,16957
<EOL>|16959,16960
9.|16960,16962
ondansetron|16963,16974
HCl|16975,16978
2|16979,16980
mg|16981,16983
/|16983,16984
mL|16984,16986
Solution|16987,16995
Sig|16996,16999
:|16999,17000
Four|17001,17005
(|17006,17007
4|17007,17008
)|17008,17009
mg|17010,17012
Intravenous|17013,17024
<EOL>|17025,17026
every|17026,17031
eight|17032,17037
(|17038,17039
8|17039,17040
)|17040,17041
hours|17042,17047
as|17048,17050
needed|17051,17057
for|17058,17061
nausea|17062,17068
.|17068,17069
<EOL>|17071,17072
10.|17072,17075
olanzapine|17076,17086
2.5|17087,17090
mg|17091,17093
Tablet|17094,17100
Sig|17101,17104
:|17104,17105
One|17106,17109
(|17110,17111
1|17111,17112
)|17112,17113
Tablet|17114,17120
PO|17121,17123
HS|17124,17126
(|17127,17128
at|17128,17130
<EOL>|17131,17132
bedtime|17132,17139
)|17139,17140
as|17141,17143
needed|17144,17150
for|17151,17154
anxiety|17155,17162
/|17162,17163
insomnia|17163,17171
.|17171,17172
<EOL>|17174,17175
11.|17175,17178
olanzapine|17179,17189
2.5|17190,17193
mg|17194,17196
Tablet|17197,17203
Sig|17204,17207
:|17207,17208
One|17209,17212
(|17213,17214
1|17214,17215
)|17215,17216
Tablet|17217,17223
PO|17224,17226
DAILY|17227,17232
<EOL>|17233,17234
(|17234,17235
Daily|17235,17240
)|17240,17241
as|17242,17244
needed|17245,17251
for|17252,17255
anxiety|17256,17263
.|17263,17264
<EOL>|17266,17267
12.|17267,17270
vancomycin|17271,17281
250|17282,17285
mg|17286,17288
Capsule|17289,17296
Sig|17297,17300
:|17300,17301
Two|17302,17305
(|17306,17307
2|17307,17308
)|17308,17309
Capsule|17310,17317
PO|17318,17320
Q6H|17321,17324
(|17325,17326
every|17326,17331
<EOL>|17332,17333
6|17333,17334
hours|17335,17340
)|17340,17341
for|17342,17345
12|17346,17348
days|17349,17353
:|17353,17354
Continue|17355,17363
through|17364,17371
_|17372,17373
_|17373,17374
_|17374,17375
.|17375,17376
<EOL>|17378,17379
<EOL>|17379,17380
<EOL>|17381,17382
Discharge|17382,17391
Disposition|17392,17403
:|17403,17404
<EOL>|17404,17405
Extended|17405,17413
Care|17414,17418
<EOL>|17418,17419
<EOL>|17420,17421
Facility|17421,17429
:|17429,17430
<EOL>|17430,17431
_|17431,17432
_|17432,17433
_|17433,17434
<EOL>|17434,17435
<EOL>|17436,17437
Discharge|17437,17446
Diagnosis|17447,17456
:|17456,17457
<EOL>|17457,17458
Primary|17458,17465
diagnoses|17466,17475
:|17475,17476
<EOL>|17476,17477
Clostridium|17477,17488
difficile|17489,17498
colitis|17499,17506
and|17507,17510
sepsis|17511,17517
<EOL>|17517,17518
Pleural|17518,17525
effusion|17526,17534
with|17535,17539
pigtail|17540,17547
catheter|17548,17556
placed|17557,17563
<EOL>|17563,17564
<EOL>|17564,17565
<EOL>|17566,17567
Discharge|17567,17576
Condition|17577,17586
:|17586,17587
<EOL>|17587,17588
Mental|17588,17594
Status|17595,17601
:|17601,17602
Confused|17603,17611
-|17612,17613
sometimes|17614,17623
.|17623,17624
<EOL>|17624,17625
Level|17625,17630
of|17631,17633
Consciousness|17634,17647
:|17647,17648
Lethargic|17649,17658
but|17659,17662
arousable|17663,17672
.|17672,17673
<EOL>|17673,17674
Activity|17674,17682
Status|17683,17689
:|17689,17690
Out|17691,17694
of|17695,17697
Bed|17698,17701
with|17702,17706
assistance|17707,17717
to|17718,17720
chair|17721,17726
or|17727,17729
<EOL>|17730,17731
wheelchair|17731,17741
.|17741,17742
<EOL>|17742,17743
<EOL>|17743,17744
<EOL>|17745,17746
Discharge|17746,17755
Instructions|17756,17768
:|17768,17769
<EOL>|17769,17770
Dear|17770,17774
Ms.|17775,17778
_|17779,17780
_|17780,17781
_|17781,17782
,|17782,17783
<EOL>|17783,17784
<EOL>|17784,17785
It|17785,17787
was|17788,17791
a|17792,17793
pleasure|17794,17802
taking|17803,17809
care|17810,17814
of|17815,17817
you|17818,17821
during|17822,17828
your|17829,17833
admission|17834,17843
to|17844,17846
<EOL>|17847,17848
_|17848,17849
_|17849,17850
_|17850,17851
for|17852,17855
abdominal|17856,17865
pain|17866,17870
.|17870,17871
You|17873,17876
were|17877,17881
found|17882,17887
to|17888,17890
have|17891,17895
an|17896,17898
infection|17899,17908
<EOL>|17909,17910
called|17910,17916
C.|17917,17919
diff|17920,17924
.|17924,17925
This|17927,17931
was|17932,17935
treated|17936,17943
with|17944,17948
antibiotics|17949,17960
which|17961,17966
you|17967,17970
<EOL>|17971,17972
will|17972,17976
continue|17977,17985
after|17986,17991
discharge|17992,18001
.|18001,18002
You|18004,18007
also|18008,18012
had|18013,18016
shortness|18017,18026
of|18027,18029
breath|18030,18036
<EOL>|18037,18038
and|18038,18041
were|18042,18046
found|18047,18052
to|18053,18055
have|18056,18060
a|18061,18062
large|18063,18068
collection|18069,18079
of|18080,18082
fluid|18083,18088
around|18089,18095
your|18096,18100
<EOL>|18101,18102
right|18102,18107
lung|18108,18112
and|18113,18116
a|18117,18118
catheter|18119,18127
was|18128,18131
placed|18132,18138
to|18139,18141
drain|18142,18147
this|18148,18152
fluid|18153,18158
.|18158,18159
This|18161,18165
<EOL>|18166,18167
catheter|18167,18175
will|18176,18180
remain|18181,18187
in|18188,18190
place|18191,18196
when|18197,18201
you|18202,18205
go|18206,18208
to|18209,18211
rehab|18212,18217
and|18218,18221
you|18222,18225
will|18226,18230
<EOL>|18231,18232
follow|18232,18238
-|18238,18239
up|18239,18241
with|18242,18246
the|18247,18250
lung|18251,18255
doctors|18256,18263
after|18264,18269
_|18270,18271
_|18271,18272
_|18272,18273
.|18273,18274
<EOL>|18274,18275
<EOL>|18275,18276
The|18276,18279
following|18280,18289
changes|18290,18297
have|18298,18302
been|18303,18307
made|18308,18312
to|18313,18315
your|18316,18320
medications|18321,18332
:|18332,18333
<EOL>|18333,18334
STOP|18334,18338
lisinopril|18339,18349
<EOL>|18349,18350
STOP|18350,18354
omeprazole|18355,18365
<EOL>|18365,18366
STOP|18366,18370
tiotropium|18371,18381
<EOL>|18381,18382
START|18382,18387
Zofran|18388,18394
4mg|18395,18398
IV|18399,18401
<EOL>|18402,18403
START|18403,18408
vancomycin|18409,18419
500mg|18420,18425
by|18426,18428
mouth|18429,18434
every|18435,18440
6|18441,18442
hours|18443,18448
through|18449,18456
_|18457,18458
_|18458,18459
_|18459,18460
<EOL>|18460,18461
START|18461,18466
olanzapine|18467,18477
2.5|18478,18481
mg|18481,18483
twice|18484,18489
daily|18490,18495
as|18496,18498
needed|18499,18505
for|18506,18509
anxiety|18510,18517
<EOL>|18517,18518
<EOL>|18519,18520
Followup|18520,18528
Instructions|18529,18541
:|18541,18542
<EOL>|18542,18543
_|18543,18544
_|18544,18545
_|18545,18546
<EOL>|18546,18547

