CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|true|false||Unit
null|Unit device|Device|true|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|true|false||Unit
null|Unit of Measure|LabModifier|true|false||Unit
null|Unit|LabModifier|true|false||Unit
null|Enzyme Unit|LabModifier|true|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Pharmaceutical Preparations|Drug|true|false||MEDICINEnull|Medicine|Title|true|false||MEDICINEnull|Known|Modifier|true|false||Knownnull|Hypersensitivity|Finding|true|false||Allergiesnull|null|Attribute|true|false||Allergiesnull|Adverse reaction to drug|Finding|true|false||Adverse Drug Reactionsnull|Adverse reaction to drug|Finding|true|false||Drug Reactionsnull|Pharmaceutical Preparations|Drug|true|false||Drug
null|Pharmacologic Substance|Drug|true|false||Drugnull|Drug problem|Finding|true|false||Drugnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|subjective (symptom)|Finding|false|false||subjectivenull|null|Attribute|false|false||subjectivenull|Subjective observation (qualifier value)|Modifier|false|false||subjectivenull|Fever|Finding|false|false||feversnull|Lethargy|Finding|false|false||lethargynull|Bloody|Finding|false|false||bloodynull|Hemorrhagic|Modifier|false|false||bloodynull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|system output|Finding|false|false||outputnull|Measurement of fluid output|Procedure|false|false||outputnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|LARGE1 wt Allele|Finding|false|false||large
null|LARGE1 gene|Finding|false|false||largenull|Large|LabModifier|false|false||largenull|Pelvis|Anatomy|false|false||pelvicnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Repositioning (procedure)|Procedure|false|false||repositioningnull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|Clinical act of insertion|Procedure|false|false||placement
null|Implantation procedure|Procedure|false|false||placement
null|null|Procedure|false|false||placementnull|Placement|Modifier|false|false||placementnull|Additional|Finding|false|false||additionalnull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|removal technique|Procedure|false|false||Removal
null|Excision|Procedure|false|false||Removal
null|Extraction|Procedure|false|false||Removalnull|Removing (action)|Event|false|false||Removalnull|More|LabModifier|false|false||morenull|Recent|Time|false|false||recentlynull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|PMH - past medical history|Finding|false|false||PMH
null|Medical History|Finding|false|false||PMHnull|Hypertensive disease|Disorder|false|false||hypertensionnull|Neoplasm of uncertain or unknown behavior of bladder|Disorder|false|false||bladder
null|Benign neoplasm of bladder|Disorder|false|false||bladder
null|Carcinoma in situ of bladder|Disorder|false|false||bladdernull|Procedures on bladder|Procedure|false|false||bladdernull|Urinary Bladder|Anatomy|false|false||bladdernull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Enneking High Surgical Grade|Finding|false|false||high grade
null|Severe (severity modifier)|Finding|false|false||high gradenull|Message Waiting Priority - High|Finding|false|false||high
null|high - ActExposureLevelCode|Finding|false|false||high
null|IPSS Risk Category High|Finding|false|false||high
null|IPSS-R Risk Category High|Finding|false|false||high
null|High (finding)|Finding|false|false||highnull|Observation Value - High|Modifier|false|false||high
null|High|Modifier|false|false||high
null|Abnormally high|Modifier|false|false||highnull|Histopathologic Grade|Finding|false|false||grade
null|Grade|Finding|false|false||grade
null|School Grade|Finding|false|false||gradenull|Invasive Urothelial Carcinoma|Disorder|false|false||invasive urothelial carcinomanull|Invasive|Modifier|false|false||invasivenull|Urothelial Carcinoma|Disorder|false|false||urothelial carcinoma
null|Carcinoma, Transitional Cell|Disorder|false|false||urothelial carcinomanull|Carcinoma|Disorder|false|false||carcinomanull|pT2b TNM Finding|Finding|false|false||pT2bnull|Total abdominal hysterectomy with bilateral salpingo-oophorectomy|Procedure|false|false||TAH/BSOnull|Total abdominal hysterectomy|Procedure|false|false||TAHnull|Tahitian language|Entity|false|false||TAHnull|Buthionine Sulfoximine|Drug|false|false||BSO
null|Buthionine Sulfoximine|Drug|false|false||BSO
null|Buthionine Sulfoximine|Drug|false|false||BSOnull|Complete cystectomy|Procedure|false|false||radical cystectomynull|Radicals (chemistry)|Drug|false|false||radicalnull|Radical (qualifier value)|Modifier|false|false||radicalnull|Cystectomy|Procedure|false|false||cystectomynull|Structure of ileal conduit|Disorder|false|false||ileal conduitnull|Ileal conduit procedure|Procedure|false|false||ileal conduitnull|ileum|Anatomy|false|false||ilealnull|Conduit implant|Device|false|false||conduitnull|Intraabdominal Route of Administration|Finding|false|false||intra-abdominalnull|Intra-abdominal|Modifier|false|false||intra-abdominalnull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|Pelvic fluid collection|Disorder|false|false||pelvic fluid collectionnull|Pelvis|Anatomy|false|false||pelvicnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Collection Object - UML Entity|Finding|false|false||collection
null|Item Collection|Finding|false|false||collection
null|Collections (publication)|Finding|false|false||collection
null|Collection (action)|Finding|false|false||collectionnull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|Clinical act of insertion|Procedure|false|false||placement
null|Implantation procedure|Procedure|false|false||placement
null|null|Procedure|false|false||placementnull|Placement|Modifier|false|false||placementnull|2 Days|Time|false|false||2 daysnull|day|Time|false|false||daysnull|Generalized|Modifier|false|false||generalizednull|Malaise|Finding|false|false||malaisenull|1 Day|Time|false|false||1 daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Fever|Finding|false|false||feversnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Drain placement|Procedure|false|false||drain placementnull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|null|Procedure|false|false||placement
null|Implantation procedure|Procedure|false|false||placement
null|Clinical act of insertion|Procedure|false|false||placementnull|Placement|Modifier|false|false||placementnull|Intra-abdominal fluid collection|Disorder|false|false||intra-abdominal fluid collectionnull|Intraabdominal Route of Administration|Finding|false|false||intra-abdominalnull|Intra-abdominal|Modifier|false|false||intra-abdominalnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Collection Object - UML Entity|Finding|false|false||collection
null|Item Collection|Finding|false|false||collection
null|Collections (publication)|Finding|false|false||collection
null|Collection (action)|Finding|false|false||collectionnull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|Thought|Finding|false|false||thought
null|null|Finding|false|false||thoughtnull|Recent|Time|false|false||recentnull|Total abdominal hysterectomy with bilateral salpingo-oophorectomy|Procedure|false|false||TAH/BSOnull|Total abdominal hysterectomy|Procedure|false|false||TAHnull|Tahitian language|Entity|false|false||TAHnull|Buthionine Sulfoximine|Drug|false|false||BSO
null|Buthionine Sulfoximine|Drug|false|false||BSO
null|Buthionine Sulfoximine|Drug|false|false||BSOnull|Complete cystectomy|Procedure|false|false||radical cystectomynull|Radicals (chemistry)|Drug|false|false||radicalnull|Radical (qualifier value)|Modifier|false|false||radicalnull|Cystectomy|Procedure|false|false||cystectomynull|Pelvis|Anatomy|false|false||pelvicnull|Biopsy of lymph node|Procedure|false|false||lymph node biopsynull|lymph nodes|Anatomy|false|false||lymph nodenull|Lymph|Finding|false|false||lymphnull|biopsy characteristics|Finding|false|false||biopsy
null|null|Finding|false|false||biopsynull|Biopsy Procedures on the Pharynx, Adenoids, and Tonsils|Procedure|false|false||biopsy
null|Biopsy|Procedure|false|false||biopsy
null|Consent Type - biopsy|Procedure|false|false||biopsynull|Procedure (set of actions)|Finding|false|false||procedurenull|Interventional procedure|Procedure|false|false||procedurenull|null|Attribute|false|false||procedurenull|Act Class - procedure|Event|false|false||procedurenull|Last 2 Days|Time|false|false||past 2 daysnull|2 Days|Time|false|false||2 daysnull|day|Time|false|false||daysnull|Generalized|Modifier|false|false||generalizednull|Malaise|Finding|false|false||malaisenull|1 Day|Time|false|false||1 daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Fever symptoms (finding)|Finding|false|false||fever
null|Fever|Finding|false|false||fevernull|Rigor - Temperature-associated observation|Finding|false|false||rigorsnull|Tmax|LabModifier|false|false||Tmaxnull|At home|Finding|false|false||at homenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Body Substance Discharge|Finding|false|false||drainage
null|Body Fluid Discharge|Finding|false|false||drainagenull|Drainage procedure|Procedure|false|false||drainagenull|Intraabdominal Route of Administration|Finding|false|false||intra-abdominalnull|Intra-abdominal|Modifier|false|false||intra-abdominalnull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|Urostomy procedure|Procedure|false|false||urostomynull|Urological stoma|Anatomy|false|false||urostomynull|system output|Finding|false|false||outputnull|Measurement of fluid output|Procedure|false|false||outputnull|null|Finding|false|false||unchangednull|About The Same|Modifier|false|false||unchangednull|Associated with|Modifier|false|false||associatednull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Left lower quadrant pain|Finding|false|false||LLQ painnull|Structure of left lower quadrant of abdomen|Anatomy|false|false||LLQnull|Left lower quadrant|Modifier|false|false||LLQnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|rectal discharge diarrhea (physical finding)|Finding|true|false||diarrhea
null|Diarrhea|Finding|true|false||diarrheanull|Hematochezia|Disorder|true|false||BRBPRnull|Eruption of skin (disorder)|Disorder|true|false||rashnull|Skin rash|Finding|true|false||rash
null|Eruptions|Finding|true|false||rash
null|Exanthema|Finding|true|false||rashnull|Cough (guaifenesin)|Drug|true|false||cough
null|Cough (guaifenesin)|Drug|true|false||coughnull|Coughing|Finding|true|false||coughnull|Headache|Finding|false|false||headachenull|Neck stiffness|Finding|false|false||neck stiffnessnull|Passive joint movement of neck (finding)|Finding|false|false||neck
null|Neck problem|Finding|false|false||necknull|dendritic spine neck|Anatomy|false|false||neck
null|Neck|Anatomy|false|false||necknull|Stiffness|Finding|false|false||stiffnessnull|Initially|Time|false|false||initiallynull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|Culture Dose Form|Drug|false|false||culturenull|Culture (Anthropological)|Finding|false|false||culture
null|Cultural aspects|Finding|false|false||culturenull|Microbial culture (procedure)|Procedure|false|false||culture
null|Laboratory culture|Procedure|false|false||culturenull|Zosyn|Drug|false|false||zosyn
null|Zosyn|Drug|false|false||zosynnull|vancomycin|Drug|false|false||vancomycin
null|vancomycin|Drug|false|false||vancomycinnull|Vancomycin measurement|Procedure|false|false||vancomycinnull|Acetaminophen [EPC]|Drug|false|false||acetaminophen
null|acetaminophen|Drug|false|false||acetaminophen
null|acetaminophen|Drug|false|false||acetaminophennull|Acetaminophen measurement|Procedure|false|false||acetaminophennull|Further|Modifier|false|false||furthernull|Disease Management|Procedure|false|false||managementnull|Management Occupations|Subject|false|false||managementnull|Management procedure|Event|false|false||management
null|Administration occupational activities|Event|false|false||managementnull|Hypertensive disease|Disorder|false|false||Hypertensionnull|ACP2 protein, human|Drug|false|false||lap
null|ACP2 protein, human|Drug|false|false||lapnull|Congenital laryngeal adductor palsy|Disorder|false|false||lapnull|Left atrial pressure|Finding|false|false||lap
null|ACP2 gene|Finding|false|false||lap
null|PICALM wt Allele|Finding|false|false||lap
null|LAP3 wt Allele|Finding|false|false||lap
null|ACP2 wt Allele|Finding|false|false||lap
null|LAP3 gene|Finding|false|false||lap
null|CENPJ gene|Finding|false|false||lap
null|CEBPB wt Allele|Finding|false|false||lap
null|PICALM gene|Finding|false|false||lap
null|CEBPB gene|Finding|false|false||lapnull|Laparoscopy|Procedure|false|false||lapnull|Lap - unit|LabModifier|false|false||lapnull|Structure of left knee region|Anatomy|false|false||left knee
null|Structure of left knee|Anatomy|false|false||left kneenull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Knee Replacement Arthroplasty|Procedure|false|false||knee replacementnull|null|Attribute|false|false||knee replacementnull|Examination of knee joint|Procedure|false|false||kneenull|Knee region structure|Anatomy|false|false||knee
null|Knee|Anatomy|false|false||knee
null|Lower extremity>Knee|Anatomy|false|false||knee
null|Knee joint|Anatomy|false|false||kneenull|Replacement|Finding|false|false||replacementnull|Replacement - supply|Procedure|false|false||replacement
null|Surgical Replantation|Procedure|false|false||replacementnull|Laminectomy|Procedure|false|false||laminectomynull|Glycation End Products, Advanced|Drug|false|false||age
null|Glycation End Products, Advanced|Drug|false|false||agenull|null|Attribute|false|false||agenull|Age|Subject|false|false||agenull|Malignant neoplasm of urinary bladder|Disorder|false|false||Bladder Cancer
null|Carcinoma of bladder|Disorder|false|false||Bladder Cancer
null|Bladder Neoplasm|Disorder|false|false||Bladder Cancernull|Carcinoma in situ of bladder|Disorder|false|false||Bladder
null|Benign neoplasm of bladder|Disorder|false|false||Bladder
null|Neoplasm of uncertain or unknown behavior of bladder|Disorder|false|false||Bladdernull|Procedures on bladder|Procedure|false|false||Bladdernull|Urinary Bladder|Anatomy|false|false||Bladdernull|Malignant Neoplasms|Disorder|false|false||Cancernull|Specialty Type - cancer|Title|false|false||Cancernull|Cancer <Cancridae>|Entity|false|false||Cancernull|Enneking High Surgical Grade|Finding|false|false||high grade
null|Severe (severity modifier)|Finding|false|false||high gradenull|Message Waiting Priority - High|Finding|false|false||high
null|high - ActExposureLevelCode|Finding|false|false||high
null|IPSS Risk Category High|Finding|false|false||high
null|IPSS-R Risk Category High|Finding|false|false||high
null|High (finding)|Finding|false|false||highnull|Observation Value - High|Modifier|false|false||high
null|High|Modifier|false|false||high
null|Abnormally high|Modifier|false|false||highnull|Histopathologic Grade|Finding|false|false||grade
null|Grade|Finding|false|false||grade
null|School Grade|Finding|false|false||gradenull|Membrane Attack Complex|Drug|false|false||TCC
null|triclocarban|Drug|false|false||TCC
null|triclocarban|Drug|false|false||TCC
null|Membrane Attack Complex|Drug|false|false||TCCnull|TARSAL-CARPAL COALITION SYNDROME|Disorder|false|false||TCCnull|membrane attack complex location|Anatomy|false|false||TCCnull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|Magnetic Resonance Imaging (MRI) of Pelvis|Procedure|false|false||pelvic MRInull|Pelvis|Anatomy|false|false||pelvicnull|CYREN gene|Finding|false|false||MRInull|Magnetic resonance imaging service|Procedure|false|false||MRI
null|Magnetic Resonance Imaging|Procedure|false|false||MRInull|Maori Language|Entity|false|false||MRInull|Tumor Cell Invasion|Disorder|false|false||invasionnull|Cell Invasion|Finding|false|false||invasionnull|Into urinary bladder|Modifier|false|false||into bladdernull|Wall of bladder|Anatomy|false|false||bladder wallnull|Neoplasm of uncertain or unknown behavior of bladder|Disorder|false|false||bladder
null|Benign neoplasm of bladder|Disorder|false|false||bladder
null|Carcinoma in situ of bladder|Disorder|false|false||bladdernull|Procedures on bladder|Procedure|false|false||bladdernull|Urinary Bladder|Anatomy|false|false||bladdernull|Walls of a building|Device|false|false||wallnull|Neck+Chest>Soft tissue|Anatomy|false|false||soft tissue
null|soft tissue|Anatomy|false|false||soft tissuenull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||softnull|Soft|Modifier|false|false||softnull|Tissue Specimen Code|Finding|false|false||tissuenull|Body tissue|Anatomy|false|false||tissuenull|Adenohypophyseal Diseases|Disorder|false|false||anteriornull|Anterior|Modifier|false|false||anteriornull|Vaginal wall|Anatomy|false|false||vaginal wallnull|Vaginal Dosage Form|Drug|false|false||vaginalnull|Vaginal Route of Administration|Finding|false|false||vaginal
null|Vaginal (intended site)|Finding|false|false||vaginalnull|Vagina|Anatomy|false|false||vaginalnull|Vaginal|Modifier|false|false||vaginalnull|Walls of a building|Device|false|false||wallnull|With staging|Finding|false|false||stagingnull|Consent Type - Hysterectomy|Finding|false|false||hysterectomynull|Hysterectomy|Procedure|false|false||hysterectomynull|Bilateral oophorectomy|Procedure|false|false||bilateral oophorectomynull|Bilateral|Modifier|false|false||bilateralnull|Ovariectomy|Procedure|false|false||oophorectomynull|Enlarged uterus|Finding|false|false||large uterusnull|LARGE1 wt Allele|Finding|false|false||large
null|LARGE1 gene|Finding|false|false||largenull|Large|LabModifier|false|false||largenull|Neoplasm of uncertain or unknown behavior of uterus|Disorder|false|false||uterus
null|Uterine Diseases|Disorder|false|false||uterusnull|examination of uterus|Procedure|false|false||uterusnull|Pelvis>Uterus|Anatomy|false|false||uterus
null|Mouse Uterus|Anatomy|false|false||uterus
null|Uterus|Anatomy|false|false||uterusnull|Fibroid Tumor|Disorder|false|false||fibroidnull|Pelvic lymph node group|Anatomy|false|false||pelvic lymph nodenull|Pelvis|Anatomy|false|false||pelvicnull|lymph nodes|Anatomy|false|false||lymph nodenull|Lymph|Finding|false|false||lymphnull|removal technique|Procedure|false|false||resection
null|Excision|Procedure|false|false||resectionnull|Complete cystectomy|Procedure|false|false||radical cystectomynull|Radicals (chemistry)|Drug|false|false||radicalnull|Radical (qualifier value)|Modifier|false|false||radicalnull|Cystectomy|Procedure|false|false||cystectomynull|Adenohypophyseal Diseases|Disorder|false|false||anteriornull|Anterior|Modifier|false|false||anteriornull|Vaginectomy|Procedure|false|false||vaginectomynull|Vaginal Dosage Form|Drug|false|false||vaginalnull|Vaginal Route of Administration|Finding|false|false||vaginal
null|Vaginal (intended site)|Finding|false|false||vaginalnull|Vagina|Anatomy|false|false||vaginalnull|Vaginal|Modifier|false|false||vaginalnull|Optical Image Reconstruction|Procedure|false|false||reconstruction
null|Reconstructive Surgical Procedures|Procedure|false|false||reconstructionnull|Structure of ileal conduit|Disorder|false|false||ileal conduitnull|Ileal conduit procedure|Procedure|false|false||ileal conduitnull|ileum|Anatomy|false|false||ilealnull|Conduit implant|Device|false|false||conduitnull|Surgical construction|Procedure|false|false||creationnull|Creation|Event|false|false||creationnull|Course|Time|false|false||coursenull|Bacteremia|Finding|false|false||bacteremianull|Growth and Development function|Finding|true|false||development
null|development aspects|Finding|true|false||development
null|biological development|Finding|true|false||development
null|Development|Finding|true|false||developmentnull|Intraabdominal Route of Administration|Finding|true|false||intra-abdominalnull|Intra-abdominal|Modifier|true|false||intra-abdominalnull|fluid - substance|Drug|true|false||fluid
null|Liquid substance|Drug|true|false||fluidnull|Fluid Specimen Code|Finding|true|false||fluidnull|Fluid behavior|Modifier|true|false||fluidnull|Collection Object - UML Entity|Finding|true|false||collection
null|Item Collection|Finding|true|false||collection
null|Collections (publication)|Finding|true|false||collection
null|Collection (action)|Finding|true|false||collectionnull|Drain placement|Procedure|true|false||drain placementnull|Drain - SpecimenType|Drug|true|false||drainnull|Drain Specimen Code|Finding|true|false||drainnull|Drain device|Device|true|false||drainnull|null|Procedure|true|false||placement
null|Implantation procedure|Procedure|true|false||placement
null|Clinical act of insertion|Procedure|true|false||placementnull|Placement|Modifier|true|false||placementnull|Deep thrombophlebitis|Disorder|false|false||DVT
null|Deep Vein Thrombosis|Disorder|false|false||DVTnull|area DVT|Anatomy|false|false||DVTnull|null|Attribute|false|false||DVTnull|Lovenox|Drug|false|false||lovenox
null|Lovenox|Drug|false|false||lovenoxnull|Negative|Finding|false|false||Negative fornull|Rh Negative Blood Group|Finding|false|false||Negative
null|Negative|Finding|false|false||Negative
null|Negative Finding|Finding|false|false||Negativenull|Expression Negative|Lab|false|false||Negativenull|Negative - qualifier|Modifier|false|false||Negative
null|Negative Charge|Modifier|false|false||Negativenull|Negative Number|LabModifier|false|false||Negativenull|Malignant neoplasm of urinary bladder|Disorder|true|false||bladder CAnull|Neoplasm of uncertain or unknown behavior of bladder|Disorder|true|false||bladder
null|Benign neoplasm of bladder|Disorder|true|false||bladder
null|Carcinoma in situ of bladder|Disorder|true|false||bladdernull|Procedures on bladder|Procedure|true|false||bladdernull|Urinary Bladder|Anatomy|true|false||bladdernull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|Exam|Finding|false|false||EXAMnull|Medical Examination|Procedure|false|false||EXAMnull|Taking vital signs|Procedure|false|false||Vital Signsnull|null|Attribute|false|false||Vital Signs
null|Vital signs|Attribute|false|false||Vital Signsnull|Vital High Nitrogen Enteral Nutrition|Drug|false|false||Vitalnull|Vital (qualifier value)|Modifier|false|false||Vitalnull|Aspects of signs|Finding|false|false||Signs
null|Physical findings|Finding|false|false||Signsnull|Manufactured sign|Device|false|false||Signsnull|Telling untruths|Finding|false|false||Lyingnull|Supine Position|Modifier|false|false||Lyingnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||Generalnull|General medical service|Procedure|false|false||Generalnull|Generalized|Modifier|false|false||Generalnull|Alert brand of caffeine|Drug|true|false||Alert
null|Alert brand of caffeine|Drug|true|false||Alertnull|Mentally alert|Finding|true|false||Alert
null|Consciousness clear|Finding|true|false||Alert
null|Alert note|Finding|true|false||Alert
null|Alert|Finding|true|false||Alertnull|null|Attribute|true|false||Alertnull|Admission Level of Care Code - Acute|Finding|true|false||acute
null|Acute - Triage Code|Finding|true|false||acutenull|acute|Time|true|false||acutenull|Emotional distress|Finding|true|false||distress
null|Distress|Finding|true|false||distressnull|HEENT|Anatomy|true|false||HEENTnull|Anicteric|Finding|false|false||anictericnull|Myelofibrosis|Disorder|false|false||MMMnull|Medial part of medial mammillary nucleus|Anatomy|false|false||MMMnull|Oropharyngeal|Anatomy|false|false||oropharynxnull|Remote control command - Clear|Finding|false|false||clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|Systolic Murmurs|Finding|true|false||systolic murmurnull|Systole|Finding|true|false||systolicnull|Heart murmur|Finding|true|false||murmurnull|Pericardial friction rub|Finding|true|false||RUBSnull|Pericardial friction rub|Finding|true|false||rubsnull|Lung|Anatomy|true|false||Lungsnull|Remote control command - Clear|Finding|true|false||Clearnull|Clear|Modifier|true|false||Clear
null|Transparent (qualitative concept)|Modifier|true|false||Clearnull|Auscultation|Procedure|true|false||auscultationnull|Wheezing|Finding|true|false||wheezesnull|Basilar Rales|Finding|true|false||rales
null|Rales|Finding|true|false||ralesnull|Rhonchi|Finding|true|false||rhonchinull|Malignant neoplasm of abdomen|Disorder|false|false||Abdomennull|Abdomen problem|Finding|false|false||Abdomennull|Abdomen|Anatomy|false|false||Abdomen
null|Abdominal Cavity|Anatomy|false|false||Abdomennull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||Softnull|Soft|Modifier|false|false||Softnull|Bowel sounds|Finding|false|false||bowel soundsnull|Intestines|Anatomy|false|false||bowelnull|null|Device|false|false||soundsnull|null|Phenomenon|false|false||soundsnull|Present|Finding|false|false||present
null|Presentation|Finding|false|false||presentnull|Structure of ileal conduit|Disorder|false|false||ileal conduitnull|Ileal conduit procedure|Procedure|false|false||ileal conduitnull|ileum|Anatomy|false|false||ilealnull|Conduit implant|Device|false|false||conduitnull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|Structure of right lower quadrant of abdomen|Anatomy|false|false||RLQnull|Right lower quadrant|Modifier|false|false||RLQnull|Pigtail Drain|Device|false|false||pigtail drainnull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|Structure of left lower quadrant of abdomen|Anatomy|false|false||LLQnull|Left lower quadrant|Modifier|false|false||LLQnull|Dark color|Modifier|false|false||darknull|GNAS-AS1 gene|Finding|false|false||sangnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Hereditary Multiple Exostoses|Disorder|true|false||Extnull|EXT1 wt Allele|Finding|true|false||Ext
null|EXT1 gene|Finding|true|false||Extnull|Feels warm|Finding|false|false||Warmnull|warming process|Phenomenon|false|false||Warmnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Neurology speciality|Title|false|false||Neuronull|Neurologic (qualifier value)|Modifier|false|false||Neuronull|CNDP2 gene|Finding|false|false||CN2null|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|All extremities|Anatomy|false|false||all extremitiesnull|All extremities|Anatomy|false|false||extremities
null|Limb structure|Anatomy|false|false||extremitiesnull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|Exam|Finding|false|false||EXAMnull|Medical Examination|Procedure|false|false||EXAMnull|Taking vital signs|Procedure|false|false||Vital signsnull|null|Attribute|false|false||Vital signs
null|Vital signs|Attribute|false|false||Vital signsnull|Vital High Nitrogen Enteral Nutrition|Drug|false|false||Vitalnull|Vital (qualifier value)|Modifier|false|false||Vitalnull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||Generalnull|General medical service|Procedure|false|false||Generalnull|Generalized|Modifier|false|false||Generalnull|HEENT|Anatomy|false|false||HEENTnull|Scleral Diseases|Disorder|false|false||Scleranull|examination of sclera|Procedure|false|false||Scleranull|Sclera|Anatomy|false|false||Scleranull|Anicteric|Finding|false|false||anictericnull|Passive joint movement of neck (finding)|Finding|false|false||Neck
null|Neck problem|Finding|false|false||Necknull|dendritic spine neck|Anatomy|false|false||Neck
null|Neck|Anatomy|false|false||Necknull|Supple|Finding|false|false||supplenull|Lung|Anatomy|false|false||Lungsnull|Remote control command - Clear|Finding|true|false||Clearnull|Clear|Modifier|true|false||Clear
null|Transparent (qualitative concept)|Modifier|true|false||Clearnull|Auscultation|Procedure|true|false||auscultationnull|Wheezing|Finding|true|false||wheezesnull|Basilar Rales|Finding|true|false||rales
null|Rales|Finding|true|false||ralesnull|Rhonchi|Finding|true|false||rhonchinull|Adenohypophyseal Diseases|Disorder|false|false||anteriornull|Anterior|Modifier|false|false||anteriornull|Auscultation|Procedure|false|false||auscultationnull|Regular|Modifier|false|false||Regularnull|Amount type - Rate|Finding|false|false||ratenull|Rating (action)|Event|false|false||ratenull|Rate|LabModifier|false|false||ratenull|Rhythm|Finding|false|false||rhythm
null|rhythmic process (biological)|Finding|false|false||rhythmnull|SYSTOLIC EJECTION MURMUR|Finding|false|false||SEMnull|Microscopes, Electron, Scanning|Device|false|false||SEMnull|Standard Error|LabModifier|false|false||SEMnull|Malignant neoplasm of abdomen|Disorder|false|false||Abdomennull|Abdomen problem|Finding|false|false||Abdomennull|Abdomen|Anatomy|false|false||Abdomen
null|Abdominal Cavity|Anatomy|false|false||Abdomennull|Structure of ileal conduit|Disorder|false|false||ileal conduitnull|Ileal conduit procedure|Procedure|false|false||ileal conduitnull|ileum|Anatomy|false|false||ilealnull|Conduit implant|Device|false|false||conduitnull|Clear Yellow|Modifier|false|false||clear yellownull|Remote control command - Clear|Finding|false|false||clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|Yellow color|Modifier|false|false||yellownull|Portion of urine|Finding|false|false||urine
null|null|Finding|false|false||urine
null|Urine|Finding|false|false||urine
null|In Urine|Finding|false|false||urine
null|Urine specimen|Finding|false|false||urinenull|Structure of left lower quadrant of abdomen|Anatomy|false|false||LLQnull|Left lower quadrant|Modifier|false|false||LLQnull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|Place - dosing instruction imperative|Finding|false|false||placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|Serosanguinous fluid|Finding|false|false||serosanguinous fluidnull|Serosanguineous|Modifier|false|false||serosanguinousnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Hereditary Multiple Exostoses|Disorder|false|false||Extnull|EXT1 wt Allele|Finding|false|false||Ext
null|EXT1 gene|Finding|false|false||Extnull|Feels warm|Finding|false|false||Warmnull|warming process|Phenomenon|false|false||Warmnull|Well (answer to question)|Finding|true|false||wellnull|Well (container)|Device|true|false||wellnull|Microplate Well|Modifier|true|false||well
null|Good|Modifier|true|false||well
null|Healthy|Modifier|true|false||wellnull|null|Drug|true|false||pulsesnull|Physiologic pulse|Finding|true|false||pulsesnull|Pulse taking|Procedure|true|false||pulsesnull|Clubbing|Disorder|true|false||clubbingnull|Cyanosis|Finding|true|false||cyanosisnull|Edema|Finding|true|false||edemanull|null|Attribute|true|false||edemanull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|Laboratory test finding|Lab|false|false||LABSnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Lymph|Finding|false|false||Lymphsnull|Monos|Drug|false|false||Monos
null|Mono-S|Drug|false|false||Monos
null|Monos|Drug|false|false||Monosnull|SARCOIDOSIS, EARLY-ONSET|Disorder|false|false||Eos
null|Familial eosinophilia|Disorder|false|false||Eosnull|PRSS33 gene|Finding|false|false||Eos
null|IKZF4 gene|Finding|false|false||Eosnull|Eos <Loriini>|Entity|false|false||Eosnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|RET protein, human|Drug|false|false||Retnull|RET protein, human|Finding|false|false||Ret
null|RET gene|Finding|false|false||Ret
null|Oncogene RET|Finding|false|false||Ret
null|RET wt Allele|Finding|false|false||Retnull|ret unit of radiation dose|LabModifier|false|false||Retnull|CONSTRICTING BANDS, CONGENITAL|Disorder|false|false||Abs
null|Amniotic Band Syndrome|Disorder|false|false||Absnull|DDX41 wt Allele|Finding|false|false||Abs
null|DDX41 gene|Finding|false|false||Absnull|RET protein, human|Drug|false|false||Retnull|RET protein, human|Finding|false|false||Ret
null|RET gene|Finding|false|false||Ret
null|Oncogene RET|Finding|false|false||Ret
null|RET wt Allele|Finding|false|false||Retnull|ret unit of radiation dose|LabModifier|false|false||Retnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Alanine Transaminase|Drug|false|false||ALT
null|Alanine Transaminase|Drug|false|false||ALTnull|Liposarcoma, well differentiated|Disorder|false|false||ALT
null|Atypical Lipoma|Disorder|false|false||ALTnull|null|Finding|false|false||ALT
null|Alternative Billing Concepts|Finding|false|false||ALT
null|GPT gene|Finding|false|false||ALTnull|Antibiotic Lock Therapy|Procedure|false|false||ALTnull|Southern Altai Language|Entity|false|false||ALTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||ASTnull|Atypical Spitz Nevus|Disorder|false|false||ASTnull|SLC17A5 wt Allele|Finding|false|false||AST
null|SLC17A5 gene|Finding|false|false||AST
null|GOT1 gene|Finding|false|false||ASTnull|Asterion|Anatomy|false|false||ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|Alkaline Phosphatase|Drug|false|false||AlkPhos
null|Alkaline Phosphatase|Drug|false|false||AlkPhosnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|lipase|Drug|false|false||Lipase
null|lipase|Drug|false|false||Lipase
null|lipase|Drug|false|false||Lipasenull|Lipase measurement|Procedure|false|false||Lipasenull|Blood albumin|Procedure|false|false||BLOOD Albuminnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Albumin|Drug|false|false||Albumin
null|Albumins|Drug|false|false||Albumin
null|Albumins|Drug|false|false||Albumin
null|Albumin|Drug|false|false||Albuminnull|Albumin metabolic function|Finding|false|false||Albumin
null|ALB gene|Finding|false|false||Albuminnull|Albumin measurement|Procedure|false|false||Albuminnull|Iron Drug Class|Drug|false|false||Iron
null|iron|Drug|false|false||Iron
null|iron|Drug|false|false||Iron
null|iron|Drug|false|false||Iron
null|Ferrum metallicum, Homeopathic preparation|Drug|false|false||Ironnull|Iron measurement|Procedure|false|false||Ironnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Thyrotropin-Releasing Hormone, human|Drug|false|false||TRF
null|IL5 protein, human|Drug|false|false||TRF
null|IL5 protein, human|Drug|false|false||TRF
null|thyrotropin-releasing hormone|Drug|false|false||TRF
null|thyrotropin-releasing hormone|Drug|false|false||TRF
null|thyrotropin-releasing hormone|Drug|false|false||TRF
null|Tocotrienol-rich Fraction|Drug|false|false||TRF
null|Thyrotropin-Releasing Hormone, human|Drug|false|false||TRFnull|TERF1 wt Allele|Finding|false|false||TRF
null|TERF1 gene|Finding|false|false||TRF
null|IL5 gene|Finding|false|false||TRFnull|lactate in blood (lab test)|Procedure|false|false||BLOOD Lactatenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|lactate|Drug|false|false||Lactate
null|lactate|Drug|false|false||Lactate
null|Lactates|Drug|false|false||Lactatenull|Lactic acid measurement|Procedure|false|false||Lactatenull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|Laboratory test finding|Lab|false|false||LABSnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood calcium measurement|Procedure|false|false||BLOOD Calciumnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Microbiology Diagnostic Service Section ID|Finding|false|false||MICROBIOLOGY
null|Microbiological|Finding|false|false||MICROBIOLOGY
null|Microbiology - Laboratory Class|Finding|false|false||MICROBIOLOGYnull|Microbiology procedure|Procedure|false|false||MICROBIOLOGYnull|Science of Microbiology|Title|false|false||MICROBIOLOGYnull|Blood culture|Procedure|false|false||Blood culturesnull|Blood and lymphatic system disorders|Disorder|false|false||Bloodnull|peripheral blood|Finding|false|false||Blood
null|Blood|Finding|false|false||Blood
null|In Blood|Finding|false|false||Bloodnull|Culture (Anthropological)|Finding|false|false||culturesnull|Pending - Allergy Clinical Status|Finding|false|false||pending
null|Pending - referral status|Finding|false|false||pendingnull|Pending - status|Time|false|false||pendingnull|pending - ManagedParticipationStatus|Modifier|false|false||pending
null|pending - RoleStatus|Modifier|false|false||pending
null|Pending - Day type|Modifier|false|false||pendingnull|Pelvis|Anatomy|false|false||pelvicnull|Respiratory Aspiration|Disorder|false|false||aspirationnull|Aspiration into respiratory tract|Finding|false|false||aspiration
null|Endotracheal aspiration|Finding|false|false||aspiration
null|Pulmonary aspiration|Finding|false|false||aspirationnull|null|Procedure|false|false||aspirationnull|Gram's stain|Drug|false|false||GRAM STAIN
null|Gram's stain|Drug|false|false||GRAM STAINnull|Bacterial stain, routine|Procedure|false|false||GRAM STAINnull|gram|LabModifier|false|false||GRAMnull|Stains|Drug|false|false||STAINnull|Staining method|Procedure|false|false||STAINnull|Diagnosis Type - Final|Finding|false|false||Finalnull|Final|Time|false|false||Finalnull|End-stage|Modifier|false|false||Finalnull|Knowledge Field|Finding|false|false||FIELD
null|Force Field|Finding|false|false||FIELD
null|Field|Finding|false|false||FIELDnull|field - patient encounter|Procedure|false|false||FIELDnull|Specimen Type - Leukocytes|Finding|false|false||LEUKOCYTES
null|null|Finding|false|false||LEUKOCYTESnull|Leukocytes|Anatomy|false|false||LEUKOCYTESnull|Microorganisms seen|Finding|true|false||MICROORGANISMS SEENnull|Microorganism|Entity|true|false||MICROORGANISMSnull|fluid - substance|Drug|false|false||FLUID
null|Liquid substance|Drug|false|false||FLUIDnull|Fluid Specimen Code|Finding|false|false||FLUIDnull|Fluid behavior|Modifier|false|false||FLUIDnull|Culture Dose Form|Drug|false|false||CULTUREnull|Culture (Anthropological)|Finding|false|false||CULTURE
null|Cultural aspects|Finding|false|false||CULTUREnull|Microbial culture (procedure)|Procedure|false|false||CULTURE
null|Laboratory culture|Procedure|false|false||CULTUREnull|Diagnosis Type - Final|Finding|false|false||Finalnull|Final|Time|false|false||Finalnull|End-stage|Modifier|false|false||Finalnull|Growth & development aspects|Finding|true|false||GROWTH
null|Tissue Growth|Finding|true|false||GROWTH
null|Growth|Finding|true|false||GROWTH
null|growth aspects|Finding|true|false||GROWTHnull|Growth action|Phenomenon|true|false||GROWTHnull|Anaerobic microbial culture|Procedure|false|false||ANAEROBIC CULTUREnull|Anaerobic|Modifier|false|false||ANAEROBICnull|Culture Dose Form|Drug|false|false||CULTUREnull|Culture (Anthropological)|Finding|false|false||CULTURE
null|Cultural aspects|Finding|false|false||CULTUREnull|Microbial culture (procedure)|Procedure|false|false||CULTURE
null|Laboratory culture|Procedure|false|false||CULTUREnull|Preliminary|Time|false|false||Preliminarynull|Growth & development aspects|Finding|true|false||GROWTH
null|Tissue Growth|Finding|true|false||GROWTH
null|Growth|Finding|true|false||GROWTH
null|growth aspects|Finding|true|false||GROWTHnull|Growth action|Phenomenon|true|false||GROWTHnull|Imaging problem|Finding|false|false||IMAGINGnull|Diagnostic Imaging|Procedure|false|false||IMAGING
null|Imaging Techniques|Procedure|false|false||IMAGINGnull|Imaging Technology|Title|false|false||IMAGINGnull|null|Attribute|false|false||CT ABDnull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false||ABDnull|ABD (body structure)|Anatomy|false|false||ABD
null|Abdomen|Anatomy|false|false||ABDnull|Pel crisis|Disorder|false|false||PEL
null|Primary Effusion Lymphoma|Disorder|false|false||PEL
null|Pure Erythroid Leukemia|Disorder|false|false||PELnull|PEL (body structure)|Anatomy|false|false||PELnull|Contrast Media|Drug|false|false||CONTRASTnull|Contrast|Modifier|false|false||CONTRASTnull|Parameterized Data Type - Interval|Finding|false|false||Intervalnull|Interval|Time|false|false||Intervalnull|Reduced|Finding|false|false||decreasenull|Decrease|LabModifier|false|false||decreasenull|size|Modifier|false|false||sizenull|size - solid dosage form|LabModifier|false|false||sizenull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Collection Object - UML Entity|Finding|false|false||collection
null|Item Collection|Finding|false|false||collection
null|Collections (publication)|Finding|false|false||collection
null|Collection (action)|Finding|false|false||collectionnull|Anterior approach|Modifier|false|false||anterior approachnull|Adenohypophyseal Diseases|Disorder|false|false||anteriornull|Anterior|Modifier|false|false||anteriornull|Approach (contact)|Finding|false|false||approachnull|Approach (spatial)|Modifier|false|false||approachnull|null|Device|false|false||pigtail catheternull|null|Finding|false|false||catheternull|catheter device|Device|false|false||catheter
null|XXX>Catheter|Device|false|false||catheternull|null|Finding|false|false||unchangednull|About The Same|Modifier|false|false||unchangednull|Position of phenotypic abnormality|Modifier|false|false||position
null|Positioning (attribute)|Modifier|false|false||positionnull|Collection Object - UML Entity|Finding|false|false||collection
null|Item Collection|Finding|false|false||collection
null|Collections (publication)|Finding|false|false||collection
null|Collection (action)|Finding|false|false||collectionnull|Walls of a building|Device|false|false||wallnull|Parameterized Data Type - Interval|Finding|false|false||Intervalnull|Interval|Time|false|false||Intervalnull|increase in size|Finding|false|false||increase in sizenull|Increase|Finding|false|false||increasenull|size|Modifier|false|false||sizenull|size - solid dosage form|LabModifier|false|false||sizenull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Pelvis|Anatomy|false|false||pelvicnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Collection Object - UML Entity|Finding|false|false||collection
null|Item Collection|Finding|false|false||collection
null|Collections (publication)|Finding|false|false||collection
null|Collection (action)|Finding|false|false||collectionnull|Peripheral|Modifier|false|false||peripheralnull|Refractive surgery enhancement|Procedure|false|false||enhancementnull|Enhance (action)|Event|false|false||enhancementnull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|Query Status Code - new|Finding|true|false||new
null|Act Status - new|Finding|true|false||newnull|Newar Language|Entity|true|false||newnull|New|Modifier|true|false||newnull|fluid - substance|Drug|true|false||fluid
null|Liquid substance|Drug|true|false||fluidnull|Fluid Specimen Code|Finding|true|false||fluidnull|Fluid behavior|Modifier|true|false||fluidnull|Collection Object - UML Entity|Finding|true|false||collection
null|Item Collection|Finding|true|false||collection
null|Collections (publication)|Finding|true|false||collection
null|Collection (action)|Finding|true|false||collectionnull|Cancer/Testis Antigen|Drug|false|false||CTAnull|PCYT1A wt Allele|Finding|false|false||CTA
null|CERNA3 gene|Finding|false|false||CTAnull|Cardiac Computerized Tomographic Angiography|Procedure|false|false||CTAnull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false||ABDnull|ABD (body structure)|Anatomy|false|false||ABD
null|Abdomen|Anatomy|false|false||ABDnull|Malignant neoplasm of pelvis|Disorder|false|false||PELVISnull|Pelvis problem|Finding|false|false||PELVISnull|Pelvis+|Anatomy|false|false||PELVIS
null|Pelvic cavity structure|Anatomy|false|false||PELVIS
null|Pelvis|Anatomy|false|false||PELVISnull|Reduced|Finding|false|false||Decreasenull|Decrease|LabModifier|false|false||Decreasenull|size|Modifier|false|false||sizenull|size - solid dosage form|LabModifier|false|false||sizenull|Structure of right lower quadrant of abdomen|Anatomy|false|false||right lower quadrantnull|Right lower quadrant|Modifier|false|false||right lower quadrantnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Quadrant|Modifier|false|false||quadrantnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Collection Object - UML Entity|Finding|false|false||collection
null|Item Collection|Finding|false|false||collection
null|Collections (publication)|Finding|false|false||collection
null|Collection (action)|Finding|false|false||collectionnull|Percutaneous Route of Drug Administration|Finding|false|false||percutaneousnull|Percutaneous|Modifier|false|false||percutaneousnull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|Areas <Spilosomini>|Entity|false|false||areasnull|Area|Modifier|false|false||areasnull|Message Waiting Priority - High|Finding|false|false||high
null|high - ActExposureLevelCode|Finding|false|false||high
null|IPSS Risk Category High|Finding|false|false||high
null|IPSS-R Risk Category High|Finding|false|false||high
null|High (finding)|Finding|false|false||highnull|Observation Value - High|Modifier|false|false||high
null|High|Modifier|false|false||high
null|Abnormally high|Modifier|false|false||highnull|Attenuation|Event|false|false||attenuationnull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Consistent with|Finding|false|false||consistent withnull|Compatible|Modifier|false|false||consistent withnull|Consistent with|Finding|false|false||consistentnull|Blood product|Drug|false|false||blood productsnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Associated with|Modifier|false|false||associatednull|Hyperemia|Disorder|false|false||hyperemianull|Likely Inflammatory Activity|Finding|false|false||likely inflammatorynull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Inflammatory|Finding|false|false||inflammatorynull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Contrast Media|Drug|true|false||contrastnull|Contrast|Modifier|true|false||contrastnull|Extravasation of Diagnostic and Therapeutic Materials|Disorder|true|false||extravasationnull|Extravasation|Finding|true|false||extravasationnull|LARGE1 wt Allele|Finding|false|false||large
null|LARGE1 gene|Finding|false|false||largenull|Large|LabModifier|false|false||largenull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Collection Object - UML Entity|Finding|false|false||collection
null|Item Collection|Finding|false|false||collection
null|Collections (publication)|Finding|false|false||collection
null|Collection (action)|Finding|false|false||collectionnull|IPSS-R Risk Category Low|Finding|false|false||low
null|IPSS Risk Category Low|Finding|false|false||low
null|low confidentiality|Finding|false|false||lownull|Low - MessageWaitingPriority|Modifier|false|false||low
null|low|Modifier|false|false||low
null|low exposure|Modifier|false|false||lownull|null|LabModifier|false|false||lownull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Malignant neoplasm of abdomen|Disorder|false|false||abdomennull|Abdomen problem|Finding|false|false||abdomennull|Abdomen|Anatomy|false|false||abdomen
null|Abdominal Cavity|Anatomy|false|false||abdomennull|Malignant neoplasm of pelvis|Disorder|false|false||pelvisnull|Pelvis problem|Finding|false|false||pelvisnull|Pelvis+|Anatomy|false|false||pelvis
null|Pelvic cavity structure|Anatomy|false|false||pelvis
null|Pelvis|Anatomy|false|false||pelvisnull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Linear|Modifier|true|false||linearnull|Peripheral|Modifier|true|false||peripheralnull|Refractive surgery enhancement|Procedure|true|false||enhancementnull|Enhance (action)|Event|true|false||enhancementnull|Communicable Diseases|Disorder|true|false||infectionnull|Infection|Finding|true|false||infectionnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Moderate to severe|Modifier|false|false||moderate to severenull|Moderate - Severity of Illness Code|Finding|false|false||moderate
null|Moderate|Finding|false|false||moderatenull|Moderate (severity modifier)|Modifier|false|false||moderate
null|Moderate - Allergy Severity|Modifier|false|false||moderate
null|Moderation|Modifier|false|false||moderatenull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Hydroureteronephrosis|Disorder|false|false||hydroureteronephrosisnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Mass Effect|Finding|false|false||Mass effectnull|Morphology, Attenuation, Size, and Structure Criteria|Finding|false|false||Mass
null|null|Finding|false|false||Mass
null|FBN1 wt Allele|Finding|false|false||Mass
null|FBN1 gene|Finding|false|false||Mass
null|Mass of body region|Finding|false|false||Mass
null|Mass of body structure|Finding|false|false||Massnull|Mass, a measure of quantity of matter|LabModifier|false|false||Mass
null|Molecular Mass|LabModifier|false|false||Massnull|Effect, Appearance|Modifier|false|false||effect
null|Effect|Modifier|false|false||effectnull|Anastomosis|Disorder|false|false||anastomosisnull|null|Procedure|false|false||anastomosisnull|Anatomical anastomosis|Anatomy|false|false||anastomosisnull|Distal Resection Margin|Attribute|false|false||distalnull|Distal (qualifier value)|Modifier|false|false||distalnull|Ureter|Anatomy|false|false||uretersnull|Neobladder|Anatomy|false|false||neobladdernull|Hydronephrosis|Disorder|false|false||hydronephrosisnull|Residual|Modifier|false|false||residualnull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Alternative|Modifier|true|false||alternativenull|Etiology aspects|Finding|true|false||etiologiesnull|Stenosis|Finding|true|false||stenosisnull|Stenosis <Pimeliinae>|Entity|true|false||stenosisnull|Stenosis Morphology|Modifier|true|false||stenosisnull|Neoplasms|Disorder|false|false||tumornull|Tumor Mass|Finding|false|false||tumor
null|null|Finding|false|false||tumornull|Infiltration Route of Administration|Finding|false|false||infiltration
null|Infiltration|Finding|false|false||infiltration
null|Spread by direct extension|Finding|false|false||infiltrationnull|Infiltration (procedure)|Procedure|false|false||infiltrationnull|Lesion of liver|Finding|false|false||hepatic lesionnull|Hepatic|Anatomy|false|false||hepaticnull|Lesion|Finding|false|false||lesion
null|null|Finding|false|false||lesionnull|Anatomical segmentation|Modifier|false|false||segmentnull|Attention - G-code|Finding|false|false||attention
null|Attention|Finding|false|false||attentionnull|Academic Research Enhancement Awards|Event|false|false||areanull|Geographic Locations|Entity|false|false||areanull|Area|Modifier|false|false||areanull|Following|Time|false|false||subsequentnull|Interventional procedure|Procedure|false|false||INTERVENTIONAL PROCEDUREnull|Interventional procedure|Procedure|false|false||INTERVENTIONAL
null|interventional (invasive) radiology|Procedure|false|false||INTERVENTIONALnull|Procedure (set of actions)|Finding|false|false||PROCEDUREnull|Interventional procedure|Procedure|false|false||PROCEDUREnull|null|Attribute|false|false||PROCEDUREnull|Act Class - procedure|Event|false|false||PROCEDUREnull|Complete, Multiple Vitamins with Iron|Drug|false|false||Complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||Complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||Completenull|Completion Status for valid values - Complete|Finding|false|false||Complete
null|Data operation - complete|Finding|false|false||Complete
null|Finish - dosing instruction imperative|Finding|false|false||Completenull|Complete|Modifier|false|false||Completenull|Collapse (finding)|Finding|false|false||collapse
null|Shock|Finding|false|false||collapse
null|null|Finding|false|false||collapsenull|Collapse (morphologic abnormality)|Phenomenon|false|false||collapsenull|Has patient|Finding|false|false||patient hasnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Recent|Time|false|false||recentlynull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Quadrant|Modifier|false|false||quadrantnull|Collection Object - UML Entity|Finding|false|false||collection
null|Item Collection|Finding|false|false||collection
null|Collections (publication)|Finding|false|false||collection
null|Collection (action)|Finding|false|false||collectionnull|null|Finding|false|false||catheternull|catheter device|Device|false|false||catheter
null|XXX>Catheter|Device|false|false||catheternull|Collection Object - UML Entity|Finding|false|false||collection
null|Item Collection|Finding|false|false||collection
null|Collections (publication)|Finding|false|false||collection
null|Collection (action)|Finding|false|false||collectionnull|Near complete|Finding|false|false||Near completenull|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||completenull|Completion Status for valid values - Complete|Finding|false|false||complete
null|Data operation - complete|Finding|false|false||complete
null|Finish - dosing instruction imperative|Finding|false|false||completenull|Complete|Modifier|false|false||completenull|Collapse (finding)|Finding|false|false||collapse
null|Shock|Finding|false|false||collapse
null|null|Finding|false|false||collapsenull|Collapse (morphologic abnormality)|Phenomenon|false|false||collapsenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Collection Object - UML Entity|Finding|false|false||collection
null|Item Collection|Finding|false|false||collection
null|Collections (publication)|Finding|false|false||collection
null|Collection (action)|Finding|false|false||collectionnull|Middle|Modifier|false|false||midnull|Malignant neoplasm of pelvis|Disorder|false|false||pelvisnull|Pelvis problem|Finding|false|false||pelvisnull|Pelvis+|Anatomy|false|false||pelvis
null|Pelvic cavity structure|Anatomy|false|false||pelvis
null|Pelvis|Anatomy|false|false||pelvisnull|null|Device|false|false||pigtail catheternull|null|Finding|false|false||catheternull|catheter device|Device|false|false||catheter
null|XXX>Catheter|Device|false|false||catheternull|Place - dosing instruction imperative|Finding|false|false||placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|Structure of left lower quadrant of abdomen|Anatomy|false|false||Left lower quadrantnull|Left lower quadrant|Modifier|false|false||Left lower quadrantnull|Table Cell Horizontal Align - left|Finding|false|false||Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Quadrant|Modifier|false|false||quadrantnull|Deep Resection Margin|Attribute|false|false||deepnull|Deep (qualifier value)|Modifier|false|false||deepnull|Pelvis|Anatomy|false|false||pelvicnull|Table Frame - above|Finding|false|false||abovenull|Upper|Modifier|false|false||abovenull|findings aspects|Finding|false|false||findingsnull|null|Attribute|false|false||findingsnull|Team|Subject|false|false||teamnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Clinical status|Attribute|false|false||clinical status
null|null|Attribute|false|false||clinical statusnull|Clinical NEC (not elsewhere classified in LNC)|Finding|false|false||clinicalnull|Clinical|Modifier|false|false||clinicalnull|What subject filter - Status|Finding|false|false||statusnull|null|Attribute|false|false||statusnull|Social status|Modifier|false|false||status
null|Status|Modifier|false|false||statusnull|Decision|Finding|true|false||decisionnull|Further|Modifier|true|false||furthernull|Collection Object - UML Entity|Finding|true|false||collection
null|Item Collection|Finding|true|false||collection
null|Collections (publication)|Finding|true|false||collection
null|Collection (action)|Finding|true|false||collectionnull|Body Substance Discharge|Finding|true|false||drainage
null|Body Fluid Discharge|Finding|true|false||drainagenull|Drainage procedure|Procedure|true|false||drainagenull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|true|false||time
null|Time (foundation metadata concept)|Finding|true|false||time
null|Value type - Time|Finding|true|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|true|false||time
null|Data types - Time|Finding|true|false||time
null|null|Finding|true|false||timenull|Time|Time|true|false||timenull|Severe - Severity of Illness Code|Finding|false|false||Severe
null|Intensity and Distress 5|Finding|false|false||Severe
null|Severe - Triage Code|Finding|false|false||Severe
null|Severe (severity modifier)|Finding|false|false||Severe
null|Allergy Severity - Severe|Finding|false|false||Severenull|Bilateral hydronephrosis|Disorder|false|false||bilateral hydronephrosisnull|Bilateral|Modifier|false|false||bilateralnull|Hydronephrosis|Disorder|false|false||hydronephrosisnull|null|Time|false|false||priornull|Physical Examination|Procedure|false|false||examinationsnull|Recommendation|Finding|false|false||RECOMMENDATIONnull|Persistence|Finding|false|false||persistencenull|Severe hydronephrosis|Disorder|false|false||severe hydronephrosisnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Hydronephrosis|Disorder|false|false||hydronephrosisnull|Percutaneous Route of Drug Administration|Finding|false|false||percutaneousnull|Percutaneous|Modifier|false|false||percutaneousnull|Nephrostomy tube|Device|false|false||nephrostomy tubesnull|Has nephrostomy|Finding|false|false||nephrostomynull|Nephrostomy (procedure)|Procedure|false|false||nephrostomynull|null|Finding|false|false||tubesnull|biomedical tube device|Device|false|false||tubesnull|Tube Dosing Unit|LabModifier|false|false||tubesnull|BRIEF Health Literacy Screening Tool|Finding|false|false||BRIEF
null|Behavior Rating Inventory of Executive Function|Finding|false|false||BRIEFnull|Brief|Time|false|false||BRIEFnull|Shortened|Modifier|false|false||BRIEFnull|summary - ActRelationshipSubset|Finding|false|false||SUMMARY
null|Summary (document)|Finding|false|false||SUMMARYnull|Transaction counts and value totals - year|Finding|false|false||year
null|Precision - year|Finding|false|false||yearnull|year|Time|false|false||yearnull|Old|Time|false|false||oldnull|Woman|Subject|false|false||womennull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Malignant neoplasm of urinary bladder|Disorder|false|false||bladder cancer
null|Carcinoma of bladder|Disorder|false|false||bladder cancer
null|Bladder Neoplasm|Disorder|false|false||bladder cancernull|Neoplasm of uncertain or unknown behavior of bladder|Disorder|false|false||bladder
null|Benign neoplasm of bladder|Disorder|false|false||bladder
null|Carcinoma in situ of bladder|Disorder|false|false||bladdernull|Procedures on bladder|Procedure|false|false||bladdernull|Urinary Bladder|Anatomy|false|false||bladdernull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Cystectomy|Procedure|false|false||cystectomynull|Consent Type - Hysterectomy|Finding|false|false||hysterectomynull|Hysterectomy|Procedure|false|false||hysterectomynull|Buthionine Sulfoximine|Drug|false|false||BSO
null|Buthionine Sulfoximine|Drug|false|false||BSO
null|Buthionine Sulfoximine|Drug|false|false||BSOnull|Structure of ileal conduit|Disorder|false|false||ileal conduitnull|Ileal conduit procedure|Procedure|false|false||ileal conduitnull|ileum|Anatomy|false|false||ilealnull|Conduit implant|Device|false|false||conduitnull|post operative (finding)|Finding|false|false||post operativenull|Operative|Time|false|false||operativenull|Course|Time|false|false||coursenull|Deep thrombophlebitis|Disorder|false|false||DVT
null|Deep Vein Thrombosis|Disorder|false|false||DVTnull|area DVT|Anatomy|false|false||DVTnull|null|Attribute|false|false||DVTnull|Intestinal obstruction co-occurrent and due to decreased peristalsis|Disorder|false|false||ileus
null|Ileus|Disorder|false|false||ileusnull|Pelvis|Anatomy|false|false||pelvicnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Structure of left lower quadrant of abdomen|Anatomy|false|false||LLQnull|Left lower quadrant|Modifier|false|false||LLQnull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|subjective (symptom)|Finding|false|false||subjectivenull|null|Attribute|false|false||subjectivenull|Subjective observation (qualifier value)|Modifier|false|false||subjectivenull|Fever|Finding|false|false||feversnull|Lethargy|Finding|false|false||lethargynull|Bloody|Finding|false|false||bloodynull|Hemorrhagic|Modifier|false|false||bloodynull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|system output|Finding|false|false||outputnull|Measurement of fluid output|Procedure|false|false||outputnull|Patient Outcome - Worsening|Finding|false|false||worseningnull|Worsening (qualifier value)|Modifier|false|false||worseningnull|Anemia|Disorder|false|false||anemianull|Anemia <Anemiaceae>|Entity|false|false||anemianull|Unit of Measure|LabModifier|false|false||units
null|Unit - NCI Thesaurus Property|LabModifier|false|false||units
null|Unit|LabModifier|false|false||unitsnull|Appropriate|Modifier|false|false||appropriatenull|Increase|Finding|false|false||increasenull|Hemoglobin|Drug|false|false||hemoglobin
null|chrysarobin|Drug|false|false||hemoglobin
null|chrysarobin|Drug|false|false||hemoglobin
null|Hemoglobin|Drug|false|false||hemoglobinnull|Hemoglobin finding|Finding|false|false||hemoglobinnull|Hemoglobin measurement|Procedure|false|false||hemoglobinnull|Imaging problem|Finding|false|false||imagingnull|Diagnostic Imaging|Procedure|false|false||imaging
null|Imaging Techniques|Procedure|false|false||imagingnull|Imaging Technology|Title|false|false||imagingnull|Parameterized Data Type - Interval|Finding|false|false||intervalnull|Interval|Time|false|false||intervalnull|increase in size|Finding|false|false||increase in sizenull|Increase|Finding|false|false||increasenull|size|Modifier|false|false||sizenull|size - solid dosage form|LabModifier|false|false||sizenull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Abdominal Fluid|Finding|false|false||abdominal fluidnull|Abdomen|Anatomy|false|false||abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Collection Object - UML Entity|Finding|false|false||collection
null|Item Collection|Finding|false|false||collection
null|Collections (publication)|Finding|false|false||collection
null|Collection (action)|Finding|false|false||collectionnull|Decision|Finding|false|false||Decisionnull|Place - dosing instruction imperative|Finding|false|false||placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|fluid - substance|Drug|false|false||Fluid
null|Liquid substance|Drug|false|false||Fluidnull|Fluid Specimen Code|Finding|false|false||Fluidnull|Fluid behavior|Modifier|false|false||Fluidnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Culture (Anthropological)|Finding|true|false||culturesnull|Rh Negative Blood Group|Finding|true|false||negative
null|Negative|Finding|true|false||negative
null|Negative Finding|Finding|true|false||negativenull|Expression Negative|Lab|true|false||negativenull|Negative - qualifier|Modifier|true|false||negative
null|Negative Charge|Modifier|true|false||negativenull|Negative Number|LabModifier|true|false||negativenull|Tumor cells, malignant|Anatomy|true|false||malignant cellsnull|Malignant (qualifier value)|Modifier|true|false||malignantnull|Cells|Anatomy|true|false||cellsnull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Lymphatic problem|Finding|true|false||lymphaticnull|Lymphatic vessel|Anatomy|true|false||lymphaticnull|Lymphatic|Modifier|true|false||lymphaticnull|Urinary tract|Anatomy|true|false||urinarynull|urinary|Modifier|true|false||urinarynull|fluid - substance|Drug|true|false||fluid
null|Liquid substance|Drug|true|false||fluidnull|Fluid Specimen Code|Finding|true|false||fluidnull|Fluid behavior|Modifier|true|false||fluidnull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Collection Object - UML Entity|Finding|false|false||collection
null|Item Collection|Finding|false|false||collection
null|Collections (publication)|Finding|false|false||collection
null|Collection (action)|Finding|false|false||collectionnull|Completely - dosing instruction fragment|Finding|false|false||completelynull|Complete|Modifier|false|false||completelynull|null|Time|false|false||priornull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|Still|Disorder|false|false||stillnull|Serosanguinous fluid|Finding|false|false||serosanguinous fluidnull|Serosanguineous|Modifier|false|false||serosanguinousnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Fever|Finding|false|false||feversnull|Leukocytosis|Disorder|false|false||leukocytosisnull|Blood leukocyte number above reference range|Finding|false|false||leukocytosisnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE|Drug|false|false||antibiotics
null|Antibiotics|Drug|false|false||antibiotics
null|Antibiotics, ophthalmologic|Drug|false|false||antibiotics
null|Antibiotics, Gynecological|Drug|false|false||antibiotics
null|antibiotics, intestinal|Drug|false|false||antibiotics
null|Antibiotic throat preparations|Drug|false|false||antibiotics
null|Antibiotics, Antitubercular|Drug|false|false||antibiotics
null|Antibiotics for systemic use|Drug|false|false||antibiotics
null|Antifungal Antibiotics, Topical|Drug|false|false||antibioticsnull|Widening|Modifier|false|false||broadnull|Spectrum|Finding|false|false||spectrumnull|Electromagnetic Spectrum|LabModifier|false|false||spectrumnull|ertapenem|Drug|false|false||ertapenem
null|ertapenem|Drug|false|false||ertapenemnull|At discharge|Time|false|false||at dischargenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Numerous|LabModifier|false|false||multiplenull|Follow - dosing instruction imperative|Finding|false|false||follow
null|Follow|Finding|false|false||follownull|Followed by|Time|false|false||follownull|Malignant Fibrous Histiocytoma|Disorder|false|false||upsnull|HMBS gene|Finding|false|false||upsnull|United Parcel Service|Entity|false|false||upsnull|Imaging problem|Finding|false|false||imagingnull|Diagnostic Imaging|Procedure|false|false||imaging
null|Imaging Techniques|Procedure|false|false||imagingnull|Imaging Technology|Title|false|false||imagingnull|Marketing basis - Transitional|Finding|false|false||transitionalnull|Transitional cell morphology|Modifier|false|false||transitionalnull|Admission Level of Care Code - Acute|Finding|false|false||ACUTE
null|Acute - Triage Code|Finding|false|false||ACUTEnull|acute|Time|false|false||ACUTEnull|Pelvis|Anatomy|false|false||Pelvicnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Adenohypophyseal Diseases|Disorder|false|false||anteriornull|Anterior|Modifier|false|false||anteriornull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|Serosanguinous fluid|Finding|false|false||serosanguinous fluidnull|Serosanguineous|Modifier|false|false||serosanguinousnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|CT of abdomen|Procedure|false|false||CT abdomennull|null|Attribute|false|false||CT abdomennull|Malignant neoplasm of abdomen|Disorder|false|false||abdomennull|Abdomen problem|Finding|false|false||abdomennull|Abdomen|Anatomy|false|false||abdomen
null|Abdominal Cavity|Anatomy|false|false||abdomennull|Malignant neoplasm of pelvis|Disorder|false|false||pelvisnull|Pelvis problem|Finding|false|false||pelvisnull|Pelvis+|Anatomy|false|false||pelvis
null|Pelvic cavity structure|Anatomy|false|false||pelvis
null|Pelvis|Anatomy|false|false||pelvisnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Collection Object - UML Entity|Finding|false|false||collection
null|Item Collection|Finding|false|false||collection
null|Collections (publication)|Finding|false|false||collection
null|Collection (action)|Finding|false|false||collectionnull|Decision|Finding|false|false||decisionnull|Place - dosing instruction imperative|Finding|false|false||placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|fluid - substance|Drug|true|false||fluid
null|Liquid substance|Drug|true|false||fluidnull|Fluid Specimen Code|Finding|true|false||fluidnull|Fluid behavior|Modifier|true|false||fluidnull|Negative|Finding|false|false||negative fornull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Malignant (qualifier value)|Modifier|true|false||malignantnull|Cells|Anatomy|true|false||cellsnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Triglycerides|Drug|false|false||triglycerides
null|Triglycerides|Drug|false|false||triglyceridesnull|Triglycerides metabolic function|Finding|false|false||triglyceridesnull|Triglycerides measurement|Procedure|false|false||triglyceridesnull|fluid - substance|Drug|true|false||fluid
null|Liquid substance|Drug|true|false||fluidnull|Fluid Specimen Code|Finding|true|false||fluidnull|Fluid behavior|Modifier|true|false||fluidnull|Collection Object - UML Entity|Finding|true|false||collection
null|Item Collection|Finding|true|false||collection
null|Collections (publication)|Finding|true|false||collection
null|Collection (action)|Finding|true|false||collectionnull|Portion of urine|Finding|true|false||urine
null|null|Finding|true|false||urine
null|Urine|Finding|true|false||urine
null|In Urine|Finding|true|false||urine
null|Urine specimen|Finding|true|false||urinenull|Lymphatic problem|Finding|true|false||lymphaticnull|Lymphatic vessel|Anatomy|true|false||lymphaticnull|Lymphatic|Modifier|true|false||lymphaticnull|fluid - substance|Drug|true|false||fluid
null|Liquid substance|Drug|true|false||fluidnull|Fluid Specimen Code|Finding|true|false||fluidnull|Fluid behavior|Modifier|true|false||fluidnull|fluid - substance|Drug|true|false||Fluid
null|Liquid substance|Drug|true|false||Fluidnull|Fluid Specimen Code|Finding|true|false||Fluidnull|Fluid behavior|Modifier|true|false||Fluidnull|Culture Dose Form|Drug|true|false||culturenull|Culture (Anthropological)|Finding|true|false||culture
null|Cultural aspects|Finding|true|false||culturenull|Microbial culture (procedure)|Procedure|true|false||culture
null|Laboratory culture|Procedure|true|false||culturenull|Negative|Finding|false|false||negative fornull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|bacteria aspects|Finding|true|false||bacterianull|Bacteria <walking sticks>|Entity|true|false||bacteria
null|Bacteria|Entity|true|false||bacterianull|Parameterized Data Type - Interval|Finding|false|false||intervalnull|Interval|Time|false|false||intervalnull|Imaging problem|Finding|false|false||imagingnull|Diagnostic Imaging|Procedure|false|false||imaging
null|Imaging Techniques|Procedure|false|false||imagingnull|Imaging Technology|Title|false|false||imagingnull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Collection Object - UML Entity|Finding|false|false||collection
null|Item Collection|Finding|false|false||collection
null|Collections (publication)|Finding|false|false||collection
null|Collection (action)|Finding|false|false||collectionnull|Completely - dosing instruction fragment|Finding|false|false||completelynull|Complete|Modifier|false|false||completelynull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Collection Object - UML Entity|Finding|false|false||collection
null|Item Collection|Finding|false|false||collection
null|Collections (publication)|Finding|false|false||collection
null|Collection (action)|Finding|false|false||collectionnull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|Serosanguinous fluid|Finding|false|false||serosanguinous fluidnull|Serosanguineous|Modifier|false|false||serosanguinousnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Serosanguinous fluid|Finding|false|false||serosanguinous fluidnull|Serosanguineous|Modifier|false|false||serosanguinousnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Amount type - Rate|Finding|false|false||ratenull|Rating (action)|Event|false|false||ratenull|Rate|LabModifier|false|false||ratenull|null|Time|false|false||prior tonull|null|Time|false|false||priornull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Place - dosing instruction imperative|Finding|false|false||placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|fluid - substance|Drug|true|false||fluid
null|Liquid substance|Drug|true|false||fluidnull|Fluid Specimen Code|Finding|true|false||fluidnull|Fluid behavior|Modifier|true|false||fluidnull|Collection Object - UML Entity|Finding|true|false||collection
null|Item Collection|Finding|true|false||collection
null|Collections (publication)|Finding|true|false||collection
null|Collection (action)|Finding|true|false||collectionnull|Imaging problem|Finding|true|false||imagingnull|Diagnostic Imaging|Procedure|true|false||imaging
null|Imaging Techniques|Procedure|true|false||imagingnull|Imaging Technology|Title|true|false||imagingnull|Completely - dosing instruction fragment|Finding|true|false||completelynull|Complete|Modifier|true|false||completelynull|Collapsed|Finding|true|false||collapsed
null|Collapse (finding)|Finding|true|false||collapsednull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Culture (Anthropological)|Finding|false|false||culturesnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Collection Object - UML Entity|Finding|false|false||collection
null|Item Collection|Finding|false|false||collection
null|Collections (publication)|Finding|false|false||collection
null|Collection (action)|Finding|false|false||collectionnull|Positive|Finding|false|false||positive fornull|BRAF Gene Rearrangement|Disorder|false|false||positivenull|Rh Positive Blood Group|Finding|false|false||positive
null|Positive Finding|Finding|false|false||positive
null|Positive|Finding|false|false||positivenull|Positive Charge|Modifier|false|false||positivenull|Positive Number|LabModifier|false|false||positivenull|Encounter due to being carrier or suspected carrier of Methicillin susceptible Staphylococcus aureus|Finding|false|false||MSSAnull|Methicillin susceptible Staphylococcus aureus|Entity|false|false||MSSAnull|Ruta graveolens preparation|Drug|true|false||rue
null|Ruta graveolens preparation|Drug|true|false||ruenull|Ruta graveolens|Entity|true|false||rue
null|Ruta|Entity|true|false||ruenull|Abdominal Infection|Disorder|true|false||intra-abdominal infectionnull|Intraabdominal Route of Administration|Finding|true|false||intra-abdominalnull|Intra-abdominal|Modifier|true|false||intra-abdominalnull|Communicable Diseases|Disorder|true|false||infectionnull|Infection|Finding|true|false||infectionnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Fever symptoms (finding)|Finding|false|false||fever
null|Fever|Finding|false|false||fevernull|Leukocytosis|Disorder|false|false||leukocytosisnull|Blood leukocyte number above reference range|Finding|false|false||leukocytosisnull|Widening|Modifier|false|false||broadnull|Spectrum|Finding|false|false||spectrumnull|Electromagnetic Spectrum|LabModifier|false|false||spectrumnull|Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE|Drug|false|false||antibiotics
null|Antibiotics|Drug|false|false||antibiotics
null|Antibiotics, ophthalmologic|Drug|false|false||antibiotics
null|Antibiotics, Gynecological|Drug|false|false||antibiotics
null|antibiotics, intestinal|Drug|false|false||antibiotics
null|Antibiotic throat preparations|Drug|false|false||antibiotics
null|Antibiotics, Antitubercular|Drug|false|false||antibiotics
null|Antibiotics for systemic use|Drug|false|false||antibiotics
null|Antifungal Antibiotics, Topical|Drug|false|false||antibioticsnull|Flagyl|Drug|false|false||flagyl
null|Flagyl|Drug|false|false||flagylnull|Team|Subject|false|false||teamnull|Zosyn|Drug|false|false||zosyn
null|Zosyn|Drug|false|false||zosynnull|On discharge|Time|false|false||On dischargenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|ertapenem|Drug|false|false||ertapenem
null|ertapenem|Drug|false|false||ertapenemnull|Approximate|Modifier|false|false||approximatelynull|4 Weeks|Time|false|false||4 weeksnull|week|Time|false|false||weeksnull|Diagnosis Type - Final|Finding|false|false||finalnull|Final|Time|false|false||finalnull|End-stage|Modifier|false|false||finalnull|Length|LabModifier|false|false||lengthnull|Biomaterial Treatment|Finding|false|false||treatment
null|Treating|Finding|false|false||treatment
null|therapeutic aspects|Finding|false|false||treatmentnull|treatment - ActInformationManagementReason|Procedure|false|false||treatment
null|Administration (procedure)|Procedure|false|false||treatment
null|Therapeutic procedure|Procedure|false|false||treatmentnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Collection Object - UML Entity|Finding|false|false||collection
null|Item Collection|Finding|false|false||collection
null|Collections (publication)|Finding|false|false||collection
null|Collection (action)|Finding|false|false||collectionnull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|Repeat Object|Finding|false|false||repeat
null|Repeat|Finding|false|false||repeatnull|Repeat Pattern|Time|false|false||repeatnull|Imaging problem|Finding|false|false||imagingnull|Diagnostic Imaging|Procedure|false|false||imaging
null|Imaging Techniques|Procedure|false|false||imagingnull|Imaging Technology|Title|false|false||imagingnull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|Basis|Drug|false|false||basisnull|Basis - conceptual entity|Finding|false|false||basisnull|Apyrexial|Finding|false|false||afebrilenull|Leukocytosis|Disorder|false|false||leukocytosisnull|Blood leukocyte number above reference range|Finding|false|false||leukocytosisnull|Pulmonary Embolism|Finding|false|false||Pulmonary embolismnull|Pulmonary (intended site)|Finding|false|false||Pulmonarynull|Lung|Anatomy|false|false||Pulmonarynull|null|Attribute|false|false||Pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||Pulmonarynull|Embolism|Finding|false|false||embolism
null|Embolus|Finding|false|false||embolismnull|Probable diagnosis|Finding|false|false||Likely
null|Probably|Finding|false|false||Likelynull|contextual factors|Finding|false|false||settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|Deep thrombophlebitis|Disorder|false|false||DVT
null|Deep Vein Thrombosis|Disorder|false|false||DVTnull|area DVT|Anatomy|false|false||DVTnull|null|Attribute|false|false||DVTnull|Lovenox|Drug|false|false||lovenox
null|Lovenox|Drug|false|false||lovenoxnull|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparinnull|Gamma-glutamyl transferase|Drug|false|false||ggt
null|Gamma-glutamyl transferase|Drug|false|false||ggtnull|GGT2P gene|Finding|false|false||ggt
null|GGT1 gene|Finding|false|false||ggtnull|Gamma glutamyl transferase measurement|Procedure|false|false||ggtnull|Procedure (set of actions)|Finding|false|false||procedures
null|Methods aspects|Finding|false|false||proceduresnull|Interventional procedure|Procedure|false|false||proceduresnull|Lovenox|Drug|false|false||lovenox
null|Lovenox|Drug|false|false||lovenoxnull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|infant weight for previous delivery (history)|Finding|false|false||weight
null|Weight symptom (finding)|Finding|false|false||weightnull|Weighing patient|Procedure|false|false||weightnull|null|Attribute|false|false||weightnull|Body Weight|Subject|false|false||weightnull|Importance Weight|Modifier|false|false||weightnull|Weight|LabModifier|false|false||weightnull|Every twelve hours|Time|false|false||q12Hnull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Acute kidney injury|Disorder|false|false||Acute renal injurynull|Admission Level of Care Code - Acute|Finding|false|false||Acute
null|Acute - Triage Code|Finding|false|false||Acutenull|acute|Time|false|false||Acutenull|Injury of kidney|Disorder|false|false||renal injurynull|Urologic Diseases|Disorder|false|false||renalnull|Kidney|Anatomy|false|false||renalnull|Traumatic AND/OR non-traumatic injury|Disorder|false|false||injury
null|Traumatic injury|Disorder|false|false||injurynull|Solitary Cutaneous Reticulohistiocytosis|Disorder|false|false||SCrnull|Stringent Complete Response|Finding|false|false||SCr
null|FBXL20 gene|Finding|false|false||SCrnull|BaseLine dental cement|Drug|false|false||baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Urologic Diseases|Disorder|false|false||uropathynull|LARGE1 wt Allele|Finding|false|false||large
null|LARGE1 gene|Finding|false|false||largenull|Large|LabModifier|false|false||largenull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Course|Time|false|false||coursenull|Hospital Stay|Time|false|false||hospital staynull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Diagnosis Type - Final|Finding|false|false||finalnull|Final|Time|false|false||finalnull|End-stage|Modifier|false|false||finalnull|Hydronephrosis|Disorder|false|false||Hydronephrosisnull|Bilateral|Modifier|false|false||bilateralnull|Parameterized Data Type - Interval|Finding|false|false||intervalnull|Interval|Time|false|false||intervalnull|Imaging problem|Finding|false|false||imagingnull|Diagnostic Imaging|Procedure|false|false||imaging
null|Imaging Techniques|Procedure|false|false||imagingnull|Imaging Technology|Title|false|false||imagingnull|null|Time|false|false||priornull|Scientific Study|Procedure|false|false||studiesnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Glycation End Products, Advanced|Drug|false|false||age
null|Glycation End Products, Advanced|Drug|false|false||agenull|null|Attribute|false|false||agenull|Age|Subject|false|false||agenull|Adequate|Modifier|false|false||adequate
null|Sufficient|Modifier|false|false||adequatenull|Urinary tract|Anatomy|false|false||urinarynull|urinary|Modifier|false|false||urinarynull|system output|Finding|true|false||outputnull|Measurement of fluid output|Procedure|true|false||outputnull|Adequate|Modifier|true|false||adequate
null|Sufficient|Modifier|true|false||adequatenull|Creatinine renal clearance measurement|Procedure|true|false||creatinine clearancenull|Creatinine clearance|Phenomenon|true|false||creatinine clearancenull|creatinine|Drug|true|false||creatinine
null|creatinine|Drug|true|false||creatininenull|Creatinine metabolic function|Finding|true|false||creatininenull|Creatinine measurement|Procedure|true|false||creatininenull|Clearance procedure|Procedure|true|false||clearancenull|Clearance of substance|Attribute|true|false||clearancenull|Clearance [PK]|Phenomenon|true|false||clearancenull|Clearance|Modifier|true|false||clearancenull|Significant|Finding|true|false||significantnull|Event Seriousness - Significant|Modifier|true|false||significantnull|Electrolyte [EPC]|Drug|true|false||electrolyte
null|Electrolytes|Drug|true|false||electrolyte
null|Electrolytes|Drug|true|false||electrolytenull|Congenital Abnormality|Disorder|true|false||abnormalitiesnull|teratologic|Finding|true|false||abnormalitiesnull|Relationship modifier - Patient|Finding|true|false||patient
null|Specimen Type - Patient|Finding|true|false||patient
null|Mail Claim Party - Patient|Finding|true|false||patient
null|Report source - Patient|Finding|true|false||patient
null|null|Finding|true|false||patient
null|Disabled Person Code - Patient|Finding|true|false||patientnull|Patients|Subject|true|false||patientnull|Veterinary Patient|Entity|true|false||patientnull|Probable diagnosis|Finding|true|false||likely
null|Probably|Finding|true|false||likelynull|Intervention regimes|Procedure|true|false||intervention
null|Nursing interventions|Procedure|true|false||intervention
null|Interventional procedure|Procedure|true|false||interventionnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|PROGRESSIVE ENCEPHALOMYELITIS WITH RIGIDITY|Disorder|false|false||Pernull|Per - dosing instruction fragment|Finding|false|false||Per
null|PER1 gene|Finding|false|false||Per
null|Follow|Finding|false|false||Per
null|PER1 wt Allele|Finding|false|false||Pernull|PER (body structure)|Anatomy|false|false||Pernull|Per (qualifier)|Modifier|false|false||Pernull|Urology|Title|false|false||urologynull|Consultation|Procedure|false|false||consultnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Recommendation|Finding|false|false||recommendednull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|Urology|Title|false|false||urologynull|follow-up|Procedure|false|false||followupnull|Anemia|Disorder|false|false||Anemianull|Anemia <Anemiaceae>|Entity|false|false||Anemianull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|combination - answer to question|Finding|false|false||combinationnull|combination of objects|Entity|false|false||combinationnull|Combined|Modifier|false|false||combinationnull|Anemia of chronic disease|Disorder|false|false||anemia of chronic inflammationnull|Anemia|Disorder|false|false||anemianull|Anemia <Anemiaceae>|Entity|false|false||anemianull|Chronic inflammation|Finding|false|false||chronic inflammationnull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Inflammation|Finding|false|false||inflammationnull|Acute hemorrhage|Finding|false|false||acute blood lossnull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Blood Loss|Finding|false|false||blood loss
null|Hemorrhage|Finding|false|false||blood lossnull|Actual blood loss|LabModifier|false|false||blood lossnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Loss (adaptation)|Finding|false|false||lossnull|Loss (quantitative)|LabModifier|false|false||lossnull|Adenohypophyseal Diseases|Disorder|false|false||anteriornull|Anterior|Modifier|false|false||anteriornull|abdominal drain in place|Finding|false|false||abdominal drainnull|Abdominal drain (physical object)|Device|false|false||abdominal drainnull|Abdomen|Anatomy|false|false||abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|Serosanguinous fluid|Finding|false|false||serosanguinous fluidnull|Serosanguineous|Modifier|false|false||serosanguinousnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Laboratory test finding|Lab|true|false||Labsnull|Consistent with|Finding|true|false||consistent withnull|Compatible|Modifier|true|false||consistent withnull|Consistent with|Finding|true|false||consistentnull|Hemolysis (biological function)|Finding|true|false||hemolysis
null|null|Finding|true|false||hemolysis
null|Hemolysis (finding)|Finding|true|false||hemolysis
null|Hemolysis (disorder)|Finding|true|false||hemolysisnull|Specimen Reject Reason - Hemolysis|Modifier|true|false||hemolysisnull|Unit of Measure|LabModifier|false|false||units
null|Unit - NCI Thesaurus Property|LabModifier|false|false||units
null|Unit|LabModifier|false|false||unitsnull|Appropriate|Modifier|false|false||appropriatenull|Communication Response|Finding|false|false||response
null|Disease Response|Finding|false|false||response
null|Answer (statement)|Finding|false|false||responsenull|Response process|Subject|false|false||responsenull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemorrhage|Finding|false|false||hemnull|altretamine/etoposide/methotrexate protocol|Procedure|false|false||hemnull|Assistant Secretary for Technology Policy/Office of the National Coordinator for Health Information Technology|Entity|false|false||oncnull|Recommendation|Finding|false|false||recommendationnull|Threshold|Modifier|false|false||thresholdnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Observation Interpretation - better|Finding|false|false||betternull|Better|Modifier|false|false||betternull|High|Modifier|false|false||highernull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|counts|LabModifier|false|false||countsnull|Hypokalemia|Finding|false|false||Hypokalemianull|Oral Dosage Form|Drug|false|false||oralnull|Oral Route of Administration|Finding|false|false||oral
null|Oral (intended site)|Finding|false|false||oralnull|Oral cavity|Anatomy|false|false||oralnull|Oral|Modifier|false|false||oralnull|potassium chloride|Drug|false|false||KCl
null|potassium chloride|Drug|false|false||KClnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Chronic - Admission Level of Care Code|Finding|false|false||CHRONICnull|Provision of recurring care for chronic illness|Procedure|false|false||CHRONICnull|chronic|Time|false|false||CHRONICnull|Invasive|Modifier|false|false||Invasivenull|Urothelial Carcinoma, High Grade|Disorder|false|false||high-grade urothelial carcinomanull|Message Waiting Priority - High|Finding|false|false||high
null|high - ActExposureLevelCode|Finding|false|false||high
null|IPSS Risk Category High|Finding|false|false||high
null|IPSS-R Risk Category High|Finding|false|false||high
null|High (finding)|Finding|false|false||highnull|Observation Value - High|Modifier|false|false||high
null|High|Modifier|false|false||high
null|Abnormally high|Modifier|false|false||highnull|Histopathologic Grade|Finding|false|false||grade
null|Grade|Finding|false|false||grade
null|School Grade|Finding|false|false||gradenull|Urothelial Carcinoma|Disorder|false|false||urothelial carcinoma
null|Carcinoma, Transitional Cell|Disorder|false|false||urothelial carcinomanull|Carcinoma|Disorder|false|false||carcinomanull|Deep Resection Margin|Attribute|false|false||deepnull|Deep (qualifier value)|Modifier|false|false||deepnull|Bladder Detrusor Muscle|Anatomy|false|false||muscularis proprianull|Bladder Detrusor Muscle|Anatomy|false|false||muscularis
null|Muscle layer|Anatomy|false|false||muscularisnull|Cystectomy|Procedure|false|false||cystectomynull|Consent Type - Hysterectomy|Finding|false|false||hysterectomynull|Hysterectomy|Procedure|false|false||hysterectomynull|Buthionine Sulfoximine|Drug|false|false||BSO
null|Buthionine Sulfoximine|Drug|false|false||BSO
null|Buthionine Sulfoximine|Drug|false|false||BSOnull|Structure of ileal conduit|Disorder|false|false||ileal conduitnull|Ileal conduit procedure|Procedure|false|false||ileal conduitnull|ileum|Anatomy|false|false||ilealnull|Conduit implant|Device|false|false||conduitnull|post operative (finding)|Finding|false|false||post operativenull|Operative|Time|false|false||operativenull|Course|Time|false|false||coursenull|Deep thrombophlebitis|Disorder|false|false||DVT
null|Deep Vein Thrombosis|Disorder|false|false||DVTnull|area DVT|Anatomy|false|false||DVTnull|null|Attribute|false|false||DVTnull|Intestinal obstruction co-occurrent and due to decreased peristalsis|Disorder|false|false||ileus
null|Ileus|Disorder|false|false||ileusnull|Pelvis|Anatomy|false|false||pelvicnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Relationship modifier - Patient|Finding|true|false||Patient
null|Specimen Type - Patient|Finding|true|false||Patient
null|Mail Claim Party - Patient|Finding|true|false||Patient
null|Report source - Patient|Finding|true|false||Patient
null|null|Finding|true|false||Patient
null|Disabled Person Code - Patient|Finding|true|false||Patientnull|Patients|Subject|true|false||Patientnull|Veterinary Patient|Entity|true|false||Patientnull|Infantile Neuroaxonal Dystrophy|Disorder|true|false||plannull|Treatment Plan|Finding|true|false||plan
null|Planned|Finding|true|false||plan
null|null|Finding|true|false||plannull|Chemotherapy Regimen|Procedure|true|false||chemo
null|Chemotherapy|Procedure|true|false||chemonull|Radiation Ionizing Radiotherapy|Procedure|true|false||radiation
null|Radiotherapy Research|Procedure|true|false||radiation
null|Radiation therapy (procedure)|Procedure|true|false||radiationnull|Electromagnetic Radiation|Phenomenon|true|false||radiation
null|Radiation|Phenomenon|true|false||radiationnull|Unit of radiation dose|LabModifier|true|false||radiationnull|Positron-Emission Tomography|Procedure|false|false||PET scannull|Tomography, Emission-Computed|Procedure|false|false||PET
null|Positron-Emission Tomography|Procedure|false|false||PETnull|Pet Animal|Entity|false|false||PETnull|Radionuclide Imaging|Procedure|false|false||scan
null|Scanning|Procedure|false|false||scannull|Focal|Modifier|false|false||foci ofnull|Foci|Finding|false|false||focinull|Focal|Modifier|false|false||focinull|Metastatic malignant neoplasm|Disorder|false|false||metastatic disease
null|Metastatic Neoplasm|Disorder|false|false||metastatic disease
null|Neoplasm Metastasis|Disorder|false|false||metastatic diseasenull|Metastatic Lesion|Finding|false|false||metastatic diseasenull|metastatic qualifier|Finding|false|false||metastatic
null|Metastatic to|Finding|false|false||metastaticnull|Disease|Disorder|false|false||diseasenull|Lung diseases|Disorder|false|false||lungnull|Lung Problem|Finding|false|false||lungnull|Chest>Lung|Anatomy|false|false||lung
null|Lung|Anatomy|false|false||lungnull|Neoplasm of uncertain or unknown behavior of peritoneum|Disorder|false|false||peritoneum
null|Benign neoplasm of peritoneum|Disorder|false|false||peritoneumnull|Serous layer of peritoneum|Anatomy|false|false||peritoneum
null|Peritoneum|Anatomy|false|false||peritoneum
null|Abdomen>Peritoneum|Anatomy|false|false||peritoneumnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|SON gene|Finding|false|false||sonnull|Son (person)|Subject|false|false||sonnull|Songhay Languages|Entity|false|false||sonnull|Doctor - Title|Finding|false|false||doctornull|Physicians|Subject|false|false||doctornull|Work-up|Procedure|false|false||work upnull|Work|Event|false|false||worknull|Lung mass|Finding|false|false||lung massnull|Lung diseases|Disorder|false|false||lungnull|Lung Problem|Finding|false|false||lungnull|Chest>Lung|Anatomy|false|false||lung
null|Lung|Anatomy|false|false||lungnull|Mass of body structure|Finding|false|false||mass
null|Morphology, Attenuation, Size, and Structure Criteria|Finding|false|false||mass
null|null|Finding|false|false||mass
null|FBN1 wt Allele|Finding|false|false||mass
null|FBN1 gene|Finding|false|false||mass
null|Mass of body region|Finding|false|false||massnull|Mass, a measure of quantity of matter|LabModifier|false|false||mass
null|Molecular Mass|LabModifier|false|false||massnull|Continuous|Finding|false|false||ongoingnull|Discussion (communication)|Finding|false|false||discussionnull|Discussion (procedure)|Procedure|false|false||discussionnull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|Hemorrhage|Finding|false|false||hemnull|altretamine/etoposide/methotrexate protocol|Procedure|false|false||hemnull|Assistant Secretary for Technology Policy/Office of the National Coordinator for Health Information Technology|Entity|false|false||oncnull|Vitelliform Macular Dystrophy|Disorder|false|false||bestnull|BEST1 wt Allele|Finding|false|false||best
null|BEST1 gene|Finding|false|false||bestnull|best (quality)|Modifier|false|false||bestnull|Lesion|Finding|false|false||lesionsnull|Mass in breast|Finding|false|false||Breast massnull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false||Breastnull|Breast problem|Finding|false|false||Breastnull|Procedures on breast|Procedure|false|false||Breastnull|Breast|Anatomy|false|false||Breastnull|Mass of body structure|Finding|false|false||mass
null|Morphology, Attenuation, Size, and Structure Criteria|Finding|false|false||mass
null|null|Finding|false|false||mass
null|FBN1 wt Allele|Finding|false|false||mass
null|FBN1 gene|Finding|false|false||mass
null|Mass of body region|Finding|false|false||massnull|Mass, a measure of quantity of matter|LabModifier|false|false||mass
null|Molecular Mass|LabModifier|false|false||massnull|Encounter due to Screening for malignant neoplasm of breast|Finding|false|false||mammogramnull|Mammography|Procedure|false|false||mammogramnull|Breast Imaging-Reporting and Data System Assessment Category 5|Finding|false|false||BI-RADS 5null|Breast Imaging Reporting and Data System|Finding|false|false||BI-RADSnull|Solid Dose Form|Drug|false|false||Solid
null|solid substance|Drug|false|false||Solidnull|Solid|Modifier|false|false||Solidnull|Mass of body structure|Finding|false|false||mass
null|Morphology, Attenuation, Size, and Structure Criteria|Finding|false|false||mass
null|null|Finding|false|false||mass
null|FBN1 wt Allele|Finding|false|false||mass
null|FBN1 gene|Finding|false|false||mass
null|Mass of body region|Finding|false|false||massnull|Mass, a measure of quantity of matter|LabModifier|false|false||mass
null|Molecular Mass|LabModifier|false|false||massnull|3 o'clock|Time|false|false||3 o'clocknull|CLOCK protein, human|Drug|false|false||clock
null|CLOCK protein, human|Drug|false|false||clocknull|CLOCK gene|Finding|false|false||clocknull|Clock Device|Device|false|false||clocknull|Left breast|Anatomy|false|false||left breastnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false||breastnull|Breast problem|Finding|false|false||breastnull|Procedures on breast|Procedure|false|false||breastnull|Breast|Anatomy|false|false||breastnull|High|Modifier|false|false||highlynull|Suspicious for Malignancy|Finding|false|false||suspicious for malignancynull|Suspicious|Modifier|false|false||suspiciousnull|Primary malignant neoplasm|Disorder|false|false||malignancy
null|Malignant Neoplasms|Disorder|false|false||malignancynull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|SON gene|Finding|false|false||sonnull|Son (person)|Subject|false|false||sonnull|Songhay Languages|Entity|false|false||sonnull|Doctor - Title|Finding|false|false||doctornull|Physicians|Subject|false|false||doctornull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|Mass in breast|Finding|false|false||breast massnull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false||breastnull|Breast problem|Finding|false|false||breastnull|Procedures on breast|Procedure|false|false||breastnull|Breast|Anatomy|false|false||breastnull|Mass of body structure|Finding|false|false||mass
null|Morphology, Attenuation, Size, and Structure Criteria|Finding|false|false||mass
null|null|Finding|false|false||mass
null|FBN1 wt Allele|Finding|false|false||mass
null|FBN1 gene|Finding|false|false||mass
null|Mass of body region|Finding|false|false||massnull|Mass, a measure of quantity of matter|LabModifier|false|false||mass
null|Molecular Mass|LabModifier|false|false||massnull|Continuous|Finding|false|false||ongoingnull|Discussion (communication)|Finding|false|false||discussionnull|Discussion (procedure)|Procedure|false|false||discussionnull|Doctor - Title|Finding|false|false||doctornull|Physicians|Subject|false|false||doctornull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|Assistant Secretary for Technology Policy/Office of the National Coordinator for Health Information Technology|Entity|false|false||oncnull|Infantile Neuroaxonal Dystrophy|Disorder|false|false||plannull|Treatment Plan|Finding|false|false||plan
null|Planned|Finding|false|false||plan
null|null|Finding|false|false||plannull|atorvastatin|Drug|true|false||atorvastatin
null|atorvastatin|Drug|true|false||atorvastatinnull|Changing|Finding|true|false||changesnull|Changed status|LabModifier|true|false||changesnull|consider|Finding|false|false||Considernull|Processing type - Evaluation|Finding|false|false||evaluationnull|Evaluation procedure|Procedure|false|false||evaluation
null|Evaluation|Procedure|false|false||evaluationnull|Stop brand of fluoride|Drug|false|false||stopping
null|Stop brand of fluoride|Drug|false|false||stoppingnull|atorvastatin|Drug|false|false||atorvastatin
null|atorvastatin|Drug|false|false||atorvastatinnull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|Basis|Drug|false|false||basisnull|Basis - conceptual entity|Finding|false|false||basisnull|Hypothyroidism|Disorder|false|false||Hypothyroidismnull|Synthetic Levothyroxine|Drug|true|false||levothyroxine
null|Synthetic Levothyroxine|Drug|true|false||levothyroxine
null|levothyroxine|Drug|true|false||levothyroxine
null|levothyroxine|Drug|true|false||levothyroxine
null|levothyroxine|Drug|true|false||levothyroxinenull|Changing|Finding|true|false||changesnull|Changed status|LabModifier|true|false||changesnull|Hereditary Coproporphyria|Disorder|false|false||HCPnull|PTPN6 wt Allele|Finding|false|false||HCP
null|CPOX gene|Finding|false|false||HCP
null|AMBP wt Allele|Finding|false|false||HCP
null|PTPN6 gene|Finding|false|false||HCP
null|AMBP gene|Finding|false|false||HCPnull|SON gene|Finding|false|false||sonnull|Son (person)|Subject|false|false||sonnull|Songhay Languages|Entity|false|false||sonnull|null|Attribute|false|false||physiciannull|Physicians|Subject|false|false||physiciannull|CODE STATUS|Procedure|false|false||Code statusnull|MDF Attribute Type - Code|Finding|false|false||Code
null|A Codes|Finding|false|false||Code
null|Code|Finding|false|false||Codenull|Coding|Event|false|false||Codenull|What subject filter - Status|Finding|false|false||statusnull|null|Attribute|false|false||statusnull|Social status|Modifier|false|false||status
null|Status|Modifier|false|false||statusnull|Full|Modifier|false|false||fullnull|MDF Attribute Type - Code|Finding|false|false||code
null|A Codes|Finding|false|false||code
null|Code|Finding|false|false||codenull|Coding|Event|false|false||codenull|Disabled Person Code - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|Relationship modifier - Patient|Finding|false|false||patient
null|null|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Marketing basis - Transitional|Finding|false|false||TRANSITIONALnull|Transitional cell morphology|Modifier|false|false||TRANSITIONALnull|Communicable Diseases|Disorder|false|false||infectious diseasenull|Infectious Disease Medicine|Title|false|false||infectious diseasenull|Communicable Diseases|Disorder|false|false||infectiousnull|infectious - Entity Risk|Modifier|false|false||infectiousnull|Disease|Disorder|false|false||diseasenull|Follow-up status|Finding|false|false||follow upnull|follow-up|Procedure|false|false||follow upnull|Follow - dosing instruction imperative|Finding|false|false||follow
null|Follow|Finding|false|false||follownull|Followed by|Time|false|false||follownull|Preparation|Event|false|false||set upnull|SET protein, human|Drug|false|false||set
null|SET protein, human|Drug|false|false||setnull|Parameterized Data Type - Set|Finding|false|false||set
null|Set scale|Finding|false|false||set
null|Set (Psychology)|Finding|false|false||set
null|SET gene|Finding|false|false||set
null|set (group)|Finding|false|false||setnull|Appointments|Event|false|false||appointmentnull|Appointments|Event|false|false||appointmentnull|CT of abdomen|Procedure|false|false||CT abdomennull|null|Attribute|false|false||CT abdomennull|Malignant neoplasm of abdomen|Disorder|false|false||abdomennull|Abdomen problem|Finding|false|false||abdomennull|Abdomen|Anatomy|false|false||abdomen
null|Abdominal Cavity|Anatomy|false|false||abdomennull|Malignant neoplasm of pelvis|Disorder|false|false||pelvisnull|Pelvis problem|Finding|false|false||pelvisnull|Pelvis+|Anatomy|false|false||pelvis
null|Pelvic cavity structure|Anatomy|false|false||pelvis
null|Pelvis|Anatomy|false|false||pelvisnull|Assure|Device|false|false||Assurenull|CT of abdomen|Procedure|false|false||CT abdomennull|null|Attribute|false|false||CT abdomennull|Malignant neoplasm of abdomen|Disorder|false|false||abdomennull|Abdomen problem|Finding|false|false||abdomennull|Abdomen|Anatomy|false|false||abdomen
null|Abdominal Cavity|Anatomy|false|false||abdomennull|Malignant neoplasm of pelvis|Disorder|false|false||pelvisnull|Pelvis problem|Finding|false|false||pelvisnull|Pelvis+|Anatomy|false|false||pelvis
null|Pelvic cavity structure|Anatomy|false|false||pelvis
null|Pelvis|Anatomy|false|false||pelvisnull|Contrast Media|Drug|false|false||contrastnull|Contrast|Modifier|false|false||contrastnull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|Weekly|Time|false|false||weeklynull|AML Lab Table|Finding|false|false||lab
null|LAT2 gene|Finding|false|false||lab
null|EWS Lab Table|Finding|false|false||labnull|Laboratory|Device|false|false||labnull|Labrador retriever|Entity|false|false||lab
null|Laboratory|Entity|false|false||labnull|Following|Time|false|false||following
null|Status post|Time|false|false||followingnull|Complete Blood Count|Procedure|false|false||CBCnull|Nuclear cap binding complex location|Anatomy|false|false||CBCnull|Amount type - Differential|Finding|false|false||differentialnull|Differential (qualifier value)|Modifier|false|false||differential
null|Different|Modifier|false|false||differential
null|Differential - view|Modifier|false|false||differentialnull|Blood Urea Nitrogen|Drug|false|false||BUN
null|Blood Urea Nitrogen|Drug|false|false||BUNnull|Blood urea nitrogen measurement|Procedure|false|false||BUNnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||ASTnull|Atypical Spitz Nevus|Disorder|false|false||ASTnull|SLC17A5 wt Allele|Finding|false|false||AST
null|SLC17A5 gene|Finding|false|false||AST
null|GOT1 gene|Finding|false|false||ASTnull|Asterion|Anatomy|false|false||ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|Alanine Transaminase|Drug|false|false||ALT
null|Alanine Transaminase|Drug|false|false||ALTnull|Liposarcoma, well differentiated|Disorder|false|false||ALT
null|Atypical Lipoma|Disorder|false|false||ALTnull|null|Finding|false|false||ALT
null|Alternative Billing Concepts|Finding|false|false||ALT
null|GPT gene|Finding|false|false||ALTnull|Antibiotic Lock Therapy|Procedure|false|false||ALTnull|Southern Altai Language|Entity|false|false||ALTnull|Alkaline Phosphatase|Drug|false|false||ALK PHOS
null|Alkaline Phosphatase|Drug|false|false||ALK PHOSnull|Alkaline phosphatase measurement|Procedure|false|false||ALK PHOSnull|ALK protein, human|Drug|false|false||ALK
null|ALK protein, human|Drug|false|false||ALKnull|ALK protein, human|Finding|false|false||ALK
null|ALK gene|Finding|false|false||ALK
null|ALK wt Allele|Finding|false|false||ALKnull|Phos <Photinae>|Entity|false|false||PHOSnull|AML Lab Table|Finding|false|false||LAB
null|LAT2 gene|Finding|false|false||LAB
null|EWS Lab Table|Finding|false|false||LABnull|Laboratory|Device|false|false||LABnull|Labrador retriever|Entity|false|false||LAB
null|Laboratory|Entity|false|false||LABnull|null|Event|false|false||REQUESTSnull|Annotated - ParameterizedDataType|Finding|false|false||ANNOTATEDnull|Clinic|Device|false|false||CLINIC
null|Ambulatory Care Facilities|Device|false|false||CLINICnull|Clinic|Entity|false|false||CLINIC
null|Ambulatory Care Facilities|Entity|false|false||CLINICnull|Patient location type - Clinic|Modifier|false|false||CLINIC
null|Person location type - Clinic|Modifier|false|false||CLINICnull|Authorization Mode - Fax|Finding|false|false||FAX
null|Fax Number|Finding|false|false||FAXnull|Facsimile Machine|Device|false|false||FAX
null|Telefacsimile|Device|false|false||FAXnull|Possible|Finding|false|false||possiblenull|Possible diagnosis|Modifier|false|false||possible
null|Possibly Related to Intervention|Modifier|false|false||possiblenull|ertapenem|Drug|false|false||ertapenem
null|ertapenem|Drug|false|false||ertapenemnull|Night time|Time|true|false||at nightnull|Night time|Time|true|false||nightnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|true|false||time
null|Time (foundation metadata concept)|Finding|true|false||time
null|Value type - Time|Finding|true|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|true|false||time
null|Data types - Time|Finding|true|false||time
null|null|Finding|true|false||timenull|Time|Time|true|false||timenull|daily activities|Finding|true|false||daily activitiesnull|Daily|Time|true|false||dailynull|activities (history)|Finding|true|false||activitiesnull|Activities|Event|true|false||activitiesnull|ertapenem|Drug|false|false||ertapenem
null|ertapenem|Drug|false|false||ertapenemnull|week|Time|false|false||weeksnull|Diagnosis Type - Final|Finding|false|false||finalnull|Final|Time|false|false||finalnull|End-stage|Modifier|false|false||finalnull|Biomaterial Treatment|Finding|false|false||treatment
null|Treating|Finding|false|false||treatment
null|therapeutic aspects|Finding|false|false||treatmentnull|treatment - ActInformationManagementReason|Procedure|false|false||treatment
null|Administration (procedure)|Procedure|false|false||treatment
null|Therapeutic procedure|Procedure|false|false||treatmentnull|Length|LabModifier|false|false||lengthnull|Communicable Diseases|Disorder|false|false||infectious diseasenull|Infectious Disease Medicine|Title|false|false||infectious diseasenull|Communicable Diseases|Disorder|false|false||infectiousnull|infectious - Entity Risk|Modifier|false|false||infectiousnull|Disease|Disorder|false|false||diseasenull|Team|Subject|false|false||teamnull|Continuous|Finding|false|false||ongoingnull|Discussion (communication)|Finding|false|false||discussionnull|Discussion (procedure)|Procedure|false|false||discussionnull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|Hemorrhage|Finding|false|false||hemnull|altretamine/etoposide/methotrexate protocol|Procedure|false|false||hemnull|Assistant Secretary for Technology Policy/Office of the National Coordinator for Health Information Technology|Entity|false|false||oncnull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|Lesion of breast|Finding|false|false||breast lesionnull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false||breastnull|Breast problem|Finding|false|false||breastnull|Procedures on breast|Procedure|false|false||breastnull|Breast|Anatomy|false|false||breastnull|Lesion|Finding|false|false||lesion
null|null|Finding|false|false||lesionnull|Lung diseases|Disorder|false|false||lungnull|Lung Problem|Finding|false|false||lungnull|Chest>Lung|Anatomy|false|false||lung
null|Lung|Anatomy|false|false||lungnull|Neoplasm of uncertain or unknown behavior of peritoneum|Disorder|false|false||peritoneum
null|Benign neoplasm of peritoneum|Disorder|false|false||peritoneumnull|Serous layer of peritoneum|Anatomy|false|false||peritoneum
null|Peritoneum|Anatomy|false|false||peritoneum
null|Abdomen>Peritoneum|Anatomy|false|false||peritoneumnull|Lesion|Finding|false|false||lesionsnull|Patient need for (contextual qualifier)|Finding|false|false||need fornull|Patient need for (contextual qualifier)|Finding|false|false||neednull|Needs|Modifier|false|false||neednull|atorvastatin|Drug|false|false||atorvastatin
null|atorvastatin|Drug|false|false||atorvastatinnull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|Urology|Title|false|false||urologynull|Team|Subject|false|false||teamnull|Patient Outcome - Worsening|Finding|false|false||worseningnull|Worsening (qualifier value)|Modifier|false|false||worseningnull|Hydronephrosis|Disorder|false|false||hydronephrosisnull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|MEDICATION LIST|Finding|false|false||Medication listnull|Pharmaceutical Preparations|Drug|false|false||Medicationnull|medication - HL7 publishing domain|Finding|false|false||Medication
null|Medications|Finding|false|false||Medicationnull|List|Finding|false|false||list
null|Sequence Data Type|Finding|false|false||listnull|Accurate (qualifier value)|Modifier|false|false||accuratenull|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||completenull|Completion Status for valid values - Complete|Finding|false|false||complete
null|Data operation - complete|Finding|false|false||complete
null|Finish - dosing instruction imperative|Finding|false|false||completenull|Complete|Modifier|false|false||completenull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Every six hours|Time|false|false||Q6Hnull|atorvastatin|Drug|false|false||Atorvastatin
null|atorvastatin|Drug|false|false||Atorvastatinnull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|enoxaparin sodium|Drug|false|false||Enoxaparin Sodium
null|enoxaparin sodium|Drug|false|false||Enoxaparin Sodiumnull|enoxaparin|Drug|false|false||Enoxaparin
null|enoxaparin|Drug|false|false||Enoxaparinnull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|Every twelve hours|Time|false|false||Q12Hnull|Firstly|Modifier|false|false||Firstnull|First (number)|LabModifier|false|false||Firstnull|Unit dose|LabModifier|false|false||Dose
null|Dosage|LabModifier|false|false||Dosenull|next - HtmlLinkType|Finding|false|false||Nextnull|Following|Time|false|false||Next
null|Then|Time|false|false||Nextnull|Adjacent|Modifier|false|false||Nextnull|Extended Priority Codes - Routine|Finding|false|false||Routine
null|Report priority - Routine|Finding|false|false||Routine
null|Admission Type - Routine|Finding|false|false||Routine
null|Level of Care - Routine|Finding|false|false||Routine
null|Processing priority - Routine|Finding|false|false||Routine
null|Referral priority - Routine|Finding|false|false||Routinenull|Routine coag|Procedure|false|false||Routinenull|Priority - Routine|Time|false|false||Routinenull|Routine|Modifier|false|false||Routinenull|Administration (procedure)|Procedure|false|false||Administrationnull|Administration occupational activities|Event|false|false||Administrationnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||Time
null|Time (foundation metadata concept)|Finding|false|false||Time
null|Value type - Time|Finding|false|false||Time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||Time
null|Data types - Time|Finding|false|false||Time
null|null|Finding|false|false||Timenull|Time|Time|false|false||Timenull|levothyroxine sodium|Drug|false|false||Levothyroxine Sodium
null|levothyroxine sodium|Drug|false|false||Levothyroxine Sodium
null|levothyroxine sodium|Drug|false|false||Levothyroxine Sodiumnull|Synthetic Levothyroxine|Drug|false|false||Levothyroxine
null|Synthetic Levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxinenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|microgram|LabModifier|false|false||mcgnull|Daily|Time|false|false||DAILYnull|lorazepam|Drug|false|false||LORazepam
null|lorazepam|Drug|false|false||LORazepamnull|Daily|Time|false|false||DAILYnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Anxiety Disorders|Disorder|false|false||anxiety
null|Anxiety|Disorder|false|false||anxietynull|Anxiety symptoms|Finding|false|false||anxietynull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|ertapenem sodium|Drug|false|false||Ertapenem Sodium
null|ertapenem sodium|Drug|false|false||Ertapenem Sodiumnull|ertapenem|Drug|false|false||Ertapenem
null|ertapenem|Drug|false|false||Ertapenemnull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|Duration brand of oxymetazoline|Drug|false|false||Durationnull|Duration (temporal concept)|Time|false|false||Durationnull|Unit dose|LabModifier|false|false||Dose
null|Dosage|LabModifier|false|false||Dosenull|ertapenem|Drug|true|false||ertapenem
null|ertapenem|Drug|true|false||ertapenemnull|Daily|Time|true|false||dailynull|Interferes with|Finding|true|false||interferenull|daily activities|Finding|true|false||daily activitiesnull|Daily|Time|true|false||dailynull|activities (history)|Finding|true|false||activitiesnull|Activities|Event|true|false||activitiesnull|Milk of Magnesia (Brand Name)|Drug|false|false||Milk of Magnesia
null|Milk of Magnesia (Brand Name)|Drug|false|false||Milk of Magnesia
null|magnesium hydroxide Oral Suspension|Drug|false|false||Milk of Magnesianull|cow milk allergenic extract|Drug|false|false||Milk
null|Milk antigen|Drug|false|false||Milk
null|Milk Beverage|Drug|false|false||Milk
null|Plant-Based Milk|Drug|false|false||Milk
null|cow milk allergenic extract|Drug|false|false||Milk
null|Milk Specimen|Drug|false|false||Milk
null|Cow's milk|Drug|false|false||Milk
null|null|Drug|false|false||Milknull|Milk (body substance)|Finding|false|false||Milk
null|Milk Specimen Code|Finding|false|false||Milknull|magnesium oxide|Drug|false|false||Magnesia
null|magnesium oxide|Drug|false|false||Magnesianull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Constipation|Finding|false|false||constipationnull|enoxaparin sodium|Drug|false|false||Enoxaparin Sodium
null|enoxaparin sodium|Drug|false|false||Enoxaparin Sodiumnull|enoxaparin|Drug|false|false||Enoxaparin
null|enoxaparin|Drug|false|false||Enoxaparinnull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|Every twelve hours|Time|false|false||Q12Hnull|Firstly|Modifier|false|false||Firstnull|First (number)|LabModifier|false|false||Firstnull|Unit dose|LabModifier|false|false||Dose
null|Dosage|LabModifier|false|false||Dosenull|next - HtmlLinkType|Finding|false|false||Nextnull|Following|Time|false|false||Next
null|Then|Time|false|false||Nextnull|Adjacent|Modifier|false|false||Nextnull|Extended Priority Codes - Routine|Finding|false|false||Routine
null|Report priority - Routine|Finding|false|false||Routine
null|Admission Type - Routine|Finding|false|false||Routine
null|Level of Care - Routine|Finding|false|false||Routine
null|Processing priority - Routine|Finding|false|false||Routine
null|Referral priority - Routine|Finding|false|false||Routinenull|Routine coag|Procedure|false|false||Routinenull|Priority - Routine|Time|false|false||Routinenull|Routine|Modifier|false|false||Routinenull|Administration (procedure)|Procedure|false|false||Administrationnull|Administration occupational activities|Event|false|false||Administrationnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||Time
null|Time (foundation metadata concept)|Finding|false|false||Time
null|Value type - Time|Finding|false|false||Time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||Time
null|Data types - Time|Finding|false|false||Time
null|null|Finding|false|false||Timenull|Time|Time|false|false||Timenull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Every six hours|Time|false|false||Q6Hnull|atorvastatin|Drug|false|false||Atorvastatin
null|atorvastatin|Drug|false|false||Atorvastatinnull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|levothyroxine sodium|Drug|false|false||Levothyroxine Sodium
null|levothyroxine sodium|Drug|false|false||Levothyroxine Sodium
null|levothyroxine sodium|Drug|false|false||Levothyroxine Sodiumnull|Synthetic Levothyroxine|Drug|false|false||Levothyroxine
null|Synthetic Levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxinenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|microgram|LabModifier|false|false||mcgnull|Daily|Time|false|false||DAILYnull|lorazepam|Drug|false|false||LORazepam
null|lorazepam|Drug|false|false||LORazepamnull|Daily|Time|false|false||DAILYnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Anxiety Disorders|Disorder|false|false||anxiety
null|Anxiety|Disorder|false|false||anxietynull|Anxiety symptoms|Finding|false|false||anxietynull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|long-term care|Procedure|false|false||Extended Carenull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|In care (finding)|Finding|false|false||Care
null|Continuity Assessment Record and Evaluation|Finding|false|false||Carenull|care activity|Event|false|false||Carenull|ADMIN.FACILITY|Finding|false|false||Facilitynull|Facility (object)|Device|false|false||Facilitynull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|null|Attribute|false|false||Primary diagnosisnull|Principal diagnosis|Modifier|false|false||Primary diagnosisnull|True primary (qualifier value)|Time|false|false||Primarynull|Primary|Modifier|false|false||Primarynull|Diagnosis Classification - Diagnosis|Finding|false|false||diagnosis
null|diagnosis aspects|Finding|false|false||diagnosisnull|Diagnosis|Procedure|false|false||diagnosisnull|null|Attribute|false|false||diagnosisnull|Pelvic fluid collection|Disorder|false|false||Pelvic fluid collectionnull|Pelvis|Anatomy|false|false||Pelvicnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Collection Object - UML Entity|Finding|false|false||collection
null|Item Collection|Finding|false|false||collection
null|Collections (publication)|Finding|false|false||collection
null|Collection (action)|Finding|false|false||collectionnull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Iron deficiency anemia secondary to chronic blood loss|Disorder|false|false||blood loss anemia
null|Anemia due to blood loss|Disorder|false|false||blood loss anemia
null|Acute posthaemorrhagic anaemia|Disorder|false|false||blood loss anemianull|Blood Loss|Finding|false|false||blood loss
null|Hemorrhage|Finding|false|false||blood lossnull|Actual blood loss|LabModifier|false|false||blood lossnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Loss (adaptation)|Finding|false|false||lossnull|Loss (quantitative)|LabModifier|false|false||lossnull|Anemia|Disorder|false|false||anemianull|Anemia <Anemiaceae>|Entity|false|false||anemianull|Secondary diagnosis|Finding|false|false||Secondary diagnosisnull|null|Attribute|false|false||Secondary diagnosisnull|Neoplasm Metastasis|Disorder|false|false||Secondarynull|metastatic qualifier|Finding|false|false||Secondarynull|Secondary to|Modifier|false|false||Secondarynull|second (number)|LabModifier|false|false||Secondarynull|Diagnosis Classification - Diagnosis|Finding|false|false||diagnosis
null|diagnosis aspects|Finding|false|false||diagnosisnull|Diagnosis|Procedure|false|false||diagnosisnull|null|Attribute|false|false||diagnosisnull|Kidney Failure, Acute|Disorder|false|false||acute renal failurenull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Kidney Failure, Acute|Disorder|false|false||renal failure, acutenull|Kidney Failure|Disorder|false|false||renal failurenull|Urologic Diseases|Disorder|false|false||renalnull|Kidney|Anatomy|false|false||renalnull|Failure (biologic function)|Finding|false|false||failure
null|Failure|Finding|false|false||failure
null|Personal failure|Finding|false|false||failurenull|Acute-on-chronic|Time|false|false||acute on chronicnull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Anemia|Disorder|false|false||anemianull|Anemia <Anemiaceae>|Entity|false|false||anemianull|Recent|Time|false|false||recentnull|Pulmonary Embolism|Finding|false|false||pulmonary embolismnull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Embolism|Finding|false|false||embolism
null|Embolus|Finding|false|false||embolismnull|Invasive|Modifier|false|false||invasivenull|Message Waiting Priority - High|Finding|false|false||high
null|high - ActExposureLevelCode|Finding|false|false||high
null|IPSS Risk Category High|Finding|false|false||high
null|IPSS-R Risk Category High|Finding|false|false||high
null|High (finding)|Finding|false|false||highnull|Observation Value - High|Modifier|false|false||high
null|High|Modifier|false|false||high
null|Abnormally high|Modifier|false|false||highnull|Histopathologic Grade|Finding|false|false||grade
null|Grade|Finding|false|false||grade
null|School Grade|Finding|false|false||gradenull|Urothelial Carcinoma|Disorder|false|false||urothelial carcinoma
null|Carcinoma, Transitional Cell|Disorder|false|false||urothelial carcinomanull|Carcinoma|Disorder|false|false||carcinomanull|Left breast|Anatomy|false|false||left breastnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Mass in breast|Finding|false|false||breast massnull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false||breastnull|Breast problem|Finding|false|false||breastnull|Procedures on breast|Procedure|false|false||breastnull|Breast|Anatomy|false|false||breastnull|Mass of body structure|Finding|false|false||mass
null|Morphology, Attenuation, Size, and Structure Criteria|Finding|false|false||mass
null|null|Finding|false|false||mass
null|FBN1 wt Allele|Finding|false|false||mass
null|FBN1 gene|Finding|false|false||mass
null|Mass of body region|Finding|false|false||massnull|Mass, a measure of quantity of matter|LabModifier|false|false||mass
null|Molecular Mass|LabModifier|false|false||massnull|Breast Imaging Reporting and Data System|Finding|false|false||BIRADSnull|Hypothyroidism|Disorder|false|false||hypothyroidismnull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Helping Behavior|Finding|false|false||assistancenull|Assisted (qualifier value)|Modifier|false|false||assistancenull|AICDA protein, human|Drug|false|false||aid
null|AICDA protein, human|Drug|false|false||aidnull|AICDA wt Allele|Finding|false|false||aid
null|AICDA gene|Finding|false|false||aidnull|AID - Artificial insemination by donor|Procedure|false|false||aid
null|dacarbazine/doxorubicin/ifosfamide protocol|Procedure|false|false||aidnull|Aid (attribute)|Modifier|false|false||aid
null|Assisted (qualifier value)|Modifier|false|false||aidnull|Walkers|Device|false|false||walkernull|CANE, INCLUDES CANES OF ALL MATERIALS, ADJUSTABLE OR FIXED, WITH TIP|Device|false|false||canenull|Cane - plant part|Entity|false|false||canenull|FBXW7-AS1 gene|Finding|false|false||Dearnull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Feeling tired|Finding|false|false||feeling tirednull|Feeling tired|Finding|false|false||tired
null|Feel Tired question|Finding|false|false||tired
null|Fatigue|Finding|false|false||tirednull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|system output|Finding|false|false||outputnull|Measurement of fluid output|Procedure|false|false||outputnull|Bloody|Finding|false|false||bloodynull|Hemorrhagic|Modifier|false|false||bloodynull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|X-Ray Computed Tomography|Procedure|false|false||CT scannull|Radionuclide Imaging|Procedure|false|false||scan
null|Scanning|Procedure|false|false||scannull|Very large|Finding|false|false||very largenull|Very|Modifier|false|false||verynull|LARGE1 wt Allele|Finding|false|false||large
null|LARGE1 gene|Finding|false|false||largenull|Large|LabModifier|false|false||largenull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Malignant neoplasm of pelvis|Disorder|false|false||pelvisnull|Pelvis problem|Finding|false|false||pelvisnull|Pelvis+|Anatomy|false|false||pelvis
null|Pelvic cavity structure|Anatomy|false|false||pelvis
null|Pelvis|Anatomy|false|false||pelvisnull|radiologist|Subject|false|false||radiologistsnull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|LARGE1 wt Allele|Finding|false|false||large
null|LARGE1 gene|Finding|false|false||largenull|Large|LabModifier|false|false||largenull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Collection Object - UML Entity|Finding|false|false||collection
null|Item Collection|Finding|false|false||collection
null|Collections (publication)|Finding|false|false||collection
null|Collection (action)|Finding|false|false||collectionnull|Blood Transfusion|Procedure|false|false||blood transfusionnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|null|Finding|false|false||transfusionnull|Blood Transfusion|Procedure|false|false||transfusion
null|Transfusion (procedure)|Procedure|false|false||transfusionnull|Peripherally Inserted Central Catheter Line Insertion|Procedure|false|false||PICCnull|Peripherally inserted central catheter (physical object)|Device|false|false||PICCnull|Long Variable|Modifier|false|false||long
null|Long|Modifier|false|false||longnull|Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE|Drug|false|false||antibiotics
null|Antibiotics|Drug|false|false||antibiotics
null|Antibiotics, ophthalmologic|Drug|false|false||antibiotics
null|Antibiotics, Gynecological|Drug|false|false||antibiotics
null|antibiotics, intestinal|Drug|false|false||antibiotics
null|Antibiotic throat preparations|Drug|false|false||antibiotics
null|Antibiotics, Antitubercular|Drug|false|false||antibiotics
null|Antibiotics for systemic use|Drug|false|false||antibiotics
null|Antifungal Antibiotics, Topical|Drug|false|false||antibioticsnull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Physicians|Subject|false|false||doctorsnull|Lung diseases|Disorder|false|false||lungnull|Lung Problem|Finding|false|false||lungnull|Chest>Lung|Anatomy|false|false||lung
null|Lung|Anatomy|false|false||lungnull|Lesion of breast|Finding|false|false||breast lesionsnull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false||breastnull|Breast problem|Finding|false|false||breastnull|Procedures on breast|Procedure|false|false||breastnull|Breast|Anatomy|false|false||breastnull|Lesion|Finding|false|false||lesionsnull|Recommendation|Finding|false|false||recommendationsnull|Continuous|Finding|false|false||Continuenull|Lovenox|Drug|false|false||Lovenox
null|Lovenox|Drug|false|false||Lovenoxnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Blood Clot|Finding|false|false||blood clot
null|Thrombus|Finding|false|false||blood clotnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|In Blood|Finding|false|false||blood
null|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||bloodnull|clotrimazole|Drug|false|false||clot
null|clotrimazole|Drug|false|false||clotnull|Blood Clot|Finding|false|false||clotnull|Lung diseases|Disorder|false|false||lungnull|Lung Problem|Finding|false|false||lungnull|Chest>Lung|Anatomy|false|false||lung
null|Lung|Anatomy|false|false||lungnull|Communicable Diseases|Disorder|true|false||infectious diseasenull|Infectious Disease Medicine|Title|true|false||infectious diseasenull|Communicable Diseases|Disorder|true|false||infectiousnull|infectious - Entity Risk|Modifier|true|false||infectiousnull|Disease|Disorder|true|false||diseasenull|Doctor - Title|Finding|true|false||doctornull|Physicians|Subject|true|false||doctornull|Following|Time|false|false||following
null|Status post|Time|false|false||followingnull|MDF AttributeType - Number|Finding|false|false||numbernull|Count of entities|LabModifier|false|false||number
null|Numbers|LabModifier|false|false||numbernull|Appointments|Event|false|false||appointmentnull|SURE Test|Finding|false|false||surenull|Certain (qualifier value)|Modifier|false|false||surenull|Repeat Object|Finding|false|false||repeat
null|Repeat|Finding|false|false||repeatnull|Repeat Pattern|Time|false|false||repeatnull|X-Ray Computed Tomography|Procedure|false|false||CT scannull|Radionuclide Imaging|Procedure|false|false||scan
null|Scanning|Procedure|false|false||scannull|Appointments|Event|false|false||appointmentnull|Communicable Diseases|Disorder|false|false||infectious diseasenull|Infectious Disease Medicine|Title|false|false||infectious diseasenull|Communicable Diseases|Disorder|false|false||infectiousnull|infectious - Entity Risk|Modifier|false|false||infectiousnull|Disease|Disorder|false|false||diseasenull|Doctor - Title|Finding|false|false||doctornull|Physicians|Subject|false|false||doctornull|Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE|Drug|false|false||antibiotics
null|Antibiotics|Drug|false|false||antibiotics
null|Antibiotics, ophthalmologic|Drug|false|false||antibiotics
null|Antibiotics, Gynecological|Drug|false|false||antibiotics
null|antibiotics, intestinal|Drug|false|false||antibiotics
null|Antibiotic throat preparations|Drug|false|false||antibiotics
null|Antibiotics, Antitubercular|Drug|false|false||antibiotics
null|Antibiotics for systemic use|Drug|false|false||antibiotics
null|Antifungal Antibiotics, Topical|Drug|false|false||antibioticsnull|Several|LabModifier|false|false||severalnull|week|Time|false|false||weeksnull|Communicable Diseases|Disorder|false|false||infectious diseasenull|Infectious Disease Medicine|Title|false|false||infectious diseasenull|Communicable Diseases|Disorder|false|false||infectiousnull|infectious - Entity Risk|Modifier|false|false||infectiousnull|Disease|Disorder|false|false||diseasenull|Doctor - Title|Finding|false|false||doctornull|Physicians|Subject|false|false||doctornull|Long Variable|Modifier|false|false||long
null|Long|Modifier|false|false||longnull|Production Class Code - Pleasure|Finding|false|false||pleasure
null|pleasurable emotion|Finding|false|false||pleasurenull|Pleasure - Animals raised for recreation|Entity|false|false||pleasurenull|care of - AddressPartType|Finding|false|false||care ofnull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Team|Subject|false|false||teamnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions