 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|28,32
No|33,35
:|35,36
_|39,40
_|40,41
_|41,42
<EOL>|42,43
<EOL>|44,45
Admission|45,54
Date|55,59
:|59,60
_|62,63
_|63,64
_|64,65
Discharge|79,88
Date|89,93
:|93,94
_|97,98
_|98,99
_|99,100
<EOL>|100,101
<EOL>|102,103
Date|103,107
of|108,110
Birth|111,116
:|116,117
_|119,120
_|120,121
_|121,122
Sex|135,138
:|138,139
F|142,143
<EOL>|143,144
<EOL>|145,146
Service|146,153
:|153,154
MEDICINE|155,163
<EOL>|163,164
<EOL>|165,166
Allergies|166,175
:|175,176
<EOL>|177,178
Codeine|178,185
/|186,187
Augmentin|188,197
/|198,199
Topamax|200,207
<EOL>|207,208
<EOL>|209,210
Attending|210,219
:|219,220
_|221,222
_|222,223
_|223,224
.|224,225
<EOL>|225,226
<EOL>|227,228
Chief|228,233
Complaint|234,243
:|243,244
<EOL>|244,245
Shortness|245,254
of|255,257
Breath|258,264
<EOL>|264,265
<EOL>|266,267
Major|267,272
Surgical|273,281
or|282,284
Invasive|285,293
Procedure|294,303
:|303,304
<EOL>|304,305
None|305,309
<EOL>|309,310
<EOL>|310,311
<EOL>|312,313
History|313,320
of|321,323
Present|324,331
Illness|332,339
:|339,340
<EOL>|340,341
Ms.|341,344
_|345,346
_|346,347
_|347,348
is|349,351
a|352,353
_|354,355
_|355,356
_|356,357
with|358,362
history|363,370
of|371,373
cerebral|374,382
aneurysm|383,391
,|391,392
<EOL>|393,394
presenting|394,404
with|405,409
shortness|410,419
of|420,422
breath|423,429
,|429,430
found|431,436
to|437,439
have|440,444
PE|445,447
at|448,450
OSH|451,454
,|454,455
<EOL>|456,457
and|457,460
transferred|461,472
here|473,477
for|478,481
further|482,489
management|490,500
.|500,501
Earlier|502,509
in|510,512
the|513,516
<EOL>|517,518
month|518,523
,|523,524
pt|525,527
developed|528,537
swelling|538,546
in|547,549
RLE|550,553
with|554,558
warmth|559,565
and|566,569
erythema|570,578
<EOL>|579,580
consistent|580,590
with|591,595
cellulitis|596,606
.|606,607
LENIs|608,613
at|614,616
this|617,621
time|622,626
did|627,630
not|631,634
<EOL>|635,636
demontrate|636,646
any|647,650
DVT|651,654
.|654,655
She|656,659
was|660,663
treated|664,671
with|672,676
a|677,678
course|679,685
of|686,688
cephalexin|689,699
<EOL>|700,701
with|701,705
improvement|706,717
in|718,720
erythema|721,729
and|730,733
pain|734,738
.|738,739
Additionally|740,752
swelling|753,761
<EOL>|762,763
went|763,767
down|768,772
substantially|773,786
.|786,787
However|788,795
,|795,796
2|797,798
days|799,803
ago|804,807
,|807,808
she|809,812
begn|813,817
<EOL>|818,819
developing|819,829
worsening|830,839
dyspnea|840,847
on|848,850
exertion|851,859
.|859,860
Promotes|861,869
chest|870,875
<EOL>|876,877
heaviness|877,886
but|887,890
no|891,893
pain|894,898
.|898,899
Denies|900,906
other|907,912
URI|913,916
symptoms|917,925
.|925,926
No|927,929
prior|930,935
hx|936,938
of|939,941
<EOL>|942,943
DVT|943,946
.|946,947
The|947,950
patient|951,958
denies|959,965
any|966,969
fever|970,975
,|975,976
chills|977,983
,|983,984
abdominal|985,994
pain|995,999
,|999,1000
bowel|1001,1006
<EOL>|1007,1008
or|1008,1010
bladder|1011,1018
changes|1019,1026
.|1026,1027
Up|1028,1030
to|1031,1033
date|1034,1038
on|1039,1041
all|1042,1045
age|1046,1049
appropriate|1050,1061
cancer|1062,1068
<EOL>|1069,1070
screening|1070,1079
.|1079,1080
No|1081,1083
recent|1084,1090
weight|1091,1097
loss|1098,1102
.|1102,1103
<EOL>|1105,1106
<EOL>|1106,1107
She|1107,1110
was|1111,1114
transferred|1115,1126
from|1127,1131
the|1132,1135
_|1136,1137
_|1137,1138
_|1138,1139
the|1140,1143
patient|1144,1151
has|1152,1155
a|1156,1157
known|1158,1163
<EOL>|1164,1165
history|1165,1172
of|1173,1175
a|1176,1177
brain|1178,1183
aneurysm|1184,1192
and|1193,1196
the|1197,1200
inpatient|1201,1210
team|1211,1215
at|1216,1218
the|1219,1222
<EOL>|1223,1224
_|1224,1225
_|1225,1226
_|1226,1227
was|1228,1231
uncomfortable|1232,1245
admitting|1246,1255
her|1256,1259
in|1260,1262
case|1263,1267
thrombolytics|1268,1281
<EOL>|1282,1283
were|1283,1287
used|1288,1292
.|1292,1293
She|1294,1297
was|1298,1301
placed|1302,1308
on|1309,1311
a|1312,1313
heparin|1314,1321
drip|1322,1326
prior|1327,1332
to|1333,1335
transfer|1336,1344
.|1344,1345
<EOL>|1347,1348
<EOL>|1348,1349
In|1349,1351
the|1352,1355
ED|1356,1358
,|1358,1359
initial|1360,1367
vital|1368,1373
signs|1374,1379
were|1380,1384
:|1384,1385
98.4|1386,1390
82|1391,1393
150|1394,1397
/|1397,1398
70|1398,1400
18|1401,1403
95|1404,1406
%|1406,1407
<EOL>|1409,1410
Exam|1410,1414
was|1415,1418
reportedly|1419,1429
unremarkable|1430,1442
.|1442,1443
A|1444,1445
bedside|1446,1453
echo|1454,1458
showed|1459,1465
no|1466,1468
<EOL>|1469,1470
obvious|1470,1477
signs|1478,1483
of|1484,1486
right|1487,1492
heart|1493,1498
strain|1499,1505
.|1505,1506
Patient|1507,1514
was|1515,1518
given|1519,1524
nothing|1525,1532
<EOL>|1533,1534
other|1534,1539
than|1540,1544
heparin|1545,1552
gtt|1553,1556
continued|1557,1566
from|1567,1571
_|1572,1573
_|1573,1574
_|1574,1575
with|1576,1580
lab|1581,1584
notable|1585,1592
<EOL>|1593,1594
for|1594,1597
PTT|1598,1601
128|1602,1605
.|1605,1606
<EOL>|1607,1608
<EOL>|1609,1610
On|1610,1612
Transfer|1613,1621
Vitals|1622,1628
were|1629,1633
:|1633,1634
97.9|1635,1639
77|1640,1642
119|1643,1646
/|1646,1647
74|1647,1649
16|1650,1652
97|1653,1655
%|1655,1656
Nasal|1657,1662
Cannula|1663,1670
.|1670,1671
<EOL>|1672,1673
Her|1673,1676
breathing|1677,1686
is|1687,1689
greatly|1690,1697
improved|1698,1706
.|1706,1707
She|1708,1711
denies|1712,1718
any|1719,1722
chest|1723,1728
pain|1729,1733
.|1733,1734
<EOL>|1736,1737
<EOL>|1737,1738
<EOL>|1739,1740
Past|1740,1744
Medical|1745,1752
History|1753,1760
:|1760,1761
<EOL>|1761,1762
CEREBRAL|1762,1770
ANEURYSM|1771,1779
<EOL>|1781,1782
incidental|1782,1792
finding|1793,1800
_|1801,1802
_|1802,1803
_|1803,1804
when|1805,1809
she|1810,1813
was|1814,1817
hospialized|1818,1829
at|1830,1832
_|1833,1834
_|1834,1835
_|1835,1836
<EOL>|1838,1839
_|1839,1840
_|1840,1841
_|1841,1842
with|1843,1847
severe|1848,1854
HA|1855,1857
,|1857,1858
dizziness|1859,1868
.|1868,1869
Head|1870,1874
CT|1875,1877
also|1878,1882
<EOL>|1883,1884
showed|1884,1890
<EOL>|1892,1893
tiny|1893,1897
lacunar|1898,1905
infarcts|1906,1914
in|1915,1917
both|1918,1922
basal|1923,1928
ganglia|1929,1936
.|1936,1937
<EOL>|1939,1940
most|1940,1944
recent|1945,1951
_|1952,1953
_|1953,1954
_|1954,1955
of|1956,1958
_|1959,1960
_|1960,1961
_|1961,1962
without|1963,1970
contrast|1971,1979
:|1979,1980
<EOL>|1982,1983
stable|1983,1989
3|1990,1991
mm|1992,1994
protuberance|1995,2007
off|2008,2011
the|2012,2015
genu|2016,2020
of|2021,2023
the|2024,2027
left|2028,2032
internal|2033,2041
<EOL>|2043,2044
carotid|2044,2051
artery|2052,2058
.|2058,2059
<EOL>|2061,2062
Followed|2062,2070
by|2071,2073
Dr.|2074,2077
_|2078,2079
_|2079,2080
_|2080,2081
at|2082,2084
_|2085,2086
_|2086,2087
_|2087,2088
.|2088,2089
<EOL>|2091,2092
MRA|2092,2095
q|2096,2097
_|2098,2099
_|2099,2100
_|2100,2101
years|2102,2107
advised|2108,2115
.|2115,2116
<EOL>|2118,2119
BRCA1|2119,2124
GENE|2125,2129
MUTATION|2130,2138
<EOL>|2140,2141
CHRONIC|2141,2148
OBSTRUCTIVE|2149,2160
PULMONARY|2161,2170
DISEASE|2171,2178
<EOL>|2180,2181
SLEEP|2181,2186
APNEA|2187,2192
<EOL>|2194,2195
COLONIC|2195,2202
POLYPS|2203,2209
<EOL>|2211,2212
GASTROESOPHAGEAL|2212,2228
REFLUX|2229,2235
<EOL>|2237,2238
DEPRESSION|2238,2248
<EOL>|2250,2251
PRE-DIABETES|2251,2263
<EOL>|2265,2266
hx|2266,2268
HEMATURIA|2269,2278
<EOL>|2280,2281
LOW|2281,2284
BACK|2285,2289
PAIN|2290,2294
VARICOSE|2295,2303
VEINS|2304,2309
R|2310,2311
>|2311,2312
L|2312,2313
<EOL>|2315,2316
SCABIES|2316,2323
<EOL>|2325,2326
HYPERLIPIDEMIA|2326,2340
<EOL>|2342,2343
ROTATOR|2343,2350
CUFF|2351,2355
TEAR|2356,2360
<EOL>|2362,2363
syncope|2363,2370
vs|2371,2373
TIA|2374,2377
carotid|2378,2385
US|2386,2388
_|2389,2390
_|2390,2391
_|2391,2392
no|2393,2395
hemodynamically|2396,2411
significant|2412,2423
<EOL>|2425,2426
<EOL>|2426,2427
stenosis|2427,2435
,|2435,2436
ECHO|2437,2441
nl|2442,2444
.|2444,2445
<EOL>|2447,2448
TAH|2448,2451
/|2451,2452
BSO|2452,2455
<EOL>|2457,2458
CHOLECYSTECTOMY|2458,2473
<EOL>|2475,2476
<EOL>|2476,2477
<EOL>|2478,2479
Social|2479,2485
History|2486,2493
:|2493,2494
<EOL>|2494,2495
_|2495,2496
_|2496,2497
_|2497,2498
<EOL>|2498,2499
Family|2499,2505
History|2506,2513
:|2513,2514
<EOL>|2514,2515
No|2515,2517
family|2518,2524
hx|2525,2527
of|2528,2530
DVT|2531,2534
or|2535,2537
PE|2538,2540
,|2540,2541
two|2542,2545
sisters|2546,2553
have|2554,2558
atrial|2559,2565
fibrillation|2566,2578
<EOL>|2580,2581
<EOL>|2581,2582
<EOL>|2582,2583
<EOL>|2584,2585
Physical|2585,2593
Exam|2594,2598
:|2598,2599
<EOL>|2599,2600
ON|2600,2602
ADMISSION|2603,2612
:|2612,2613
<EOL>|2613,2614
<EOL>|2614,2615
VS|2615,2617
:|2617,2618
98.9|2619,2623
105|2624,2627
/|2627,2628
54|2628,2630
65|2631,2633
18|2634,2636
96|2637,2639
%|2639,2640
on|2641,2643
RA|2644,2646
<EOL>|2646,2647
GENERAL|2647,2654
:|2654,2655
NAD|2656,2659
,|2659,2660
obese|2661,2666
<EOL>|2668,2669
HEENT|2669,2674
:|2674,2675
AT|2676,2678
/|2678,2679
NC|2679,2681
,|2681,2682
EOMI|2683,2687
,|2687,2688
PERRL|2689,2694
,|2694,2695
anicteric|2696,2705
sclera|2706,2712
,|2712,2713
pink|2714,2718
conjunctiva|2719,2730
,|2730,2731
<EOL>|2732,2733
MMM|2733,2736
,|2736,2737
good|2738,2742
dentition|2743,2752
<EOL>|2754,2755
NECK|2755,2759
:|2759,2760
nontender|2761,2770
supple|2771,2777
neck|2778,2782
,|2782,2783
no|2784,2786
LAD|2787,2790
,|2790,2791
no|2792,2794
JVD|2795,2798
<EOL>|2800,2801
CARDIAC|2801,2808
:|2808,2809
RRR|2810,2813
,|2813,2814
S1|2815,2817
/|2817,2818
S2|2818,2820
,|2820,2821
no|2822,2824
murmurs|2825,2832
,|2832,2833
gallops|2834,2841
,|2841,2842
or|2843,2845
rubs|2846,2850
<EOL>|2852,2853
LUNG|2853,2857
:|2857,2858
CTAB|2859,2863
,|2863,2864
no|2865,2867
wheezes|2868,2875
,|2875,2876
rales|2877,2882
,|2882,2883
rhonchi|2884,2891
,|2891,2892
breathing|2893,2902
comfortably|2903,2914
<EOL>|2915,2916
without|2916,2923
use|2924,2927
of|2928,2930
accessory|2931,2940
muscles|2941,2948
<EOL>|2950,2951
ABDOMEN|2951,2958
:|2958,2959
nondistended|2960,2972
,|2972,2973
+|2974,2975
BS|2975,2977
,|2977,2978
nontender|2979,2988
in|2989,2991
all|2992,2995
quadrants|2996,3005
,|3005,3006
no|3007,3009
<EOL>|3010,3011
rebound|3011,3018
/|3018,3019
guarding|3019,3027
,|3027,3028
no|3029,3031
hepatosplenomegaly|3032,3050
<EOL>|3052,3053
EXTREMITIES|3053,3064
:|3064,3065
no|3066,3068
appreciable|3069,3080
lower|3081,3086
exam|3087,3091
swelling|3092,3100
althught|3101,3109
R|3110,3111
calf|3112,3116
<EOL>|3117,3118
is|3118,3120
tender|3121,3127
to|3128,3130
palpation|3131,3140
<EOL>|3140,3141
PULSES|3141,3147
:|3147,3148
2|3149,3150
+|3150,3151
DP|3152,3154
pulses|3155,3161
bilaterally|3162,3173
<EOL>|3175,3176
NEURO|3176,3181
:|3181,3182
CN|3183,3185
II|3186,3188
-|3188,3189
XII|3189,3192
intact|3193,3199
,|3199,3200
no|3201,3203
focal|3204,3209
deficits|3210,3218
<EOL>|3220,3221
SKIN|3221,3225
:|3225,3226
warm|3227,3231
and|3232,3235
well|3236,3240
perfused|3241,3249
,|3249,3250
no|3251,3253
excoriations|3254,3266
or|3267,3269
lesions|3270,3277
,|3277,3278
no|3279,3281
<EOL>|3282,3283
rashes|3283,3289
<EOL>|3289,3290
<EOL>|3292,3293
<EOL>|3293,3294
ON|3294,3296
DISCHARGE|3297,3306
:|3306,3307
<EOL>|3307,3308
VS|3308,3310
:|3310,3311
98.5|3312,3316
124|3317,3320
/|3320,3321
61|3321,3323
77|3324,3326
18|3327,3329
98|3330,3332
%|3332,3333
on|3334,3336
RA|3337,3339
<EOL>|3339,3340
GENERAL|3340,3347
:|3347,3348
NAD|3349,3352
,|3352,3353
obese|3354,3359
<EOL>|3361,3362
HEENT|3362,3367
:|3367,3368
AT|3369,3371
/|3371,3372
NC|3372,3374
,|3374,3375
EOMI|3376,3380
,|3380,3381
PERRL|3382,3387
,|3387,3388
anicteric|3389,3398
sclera|3399,3405
,|3405,3406
pink|3407,3411
conjunctiva|3412,3423
,|3423,3424
<EOL>|3425,3426
MMM|3426,3429
,|3429,3430
good|3431,3435
dentition|3436,3445
<EOL>|3447,3448
NECK|3448,3452
:|3452,3453
nontender|3454,3463
supple|3464,3470
neck|3471,3475
,|3475,3476
no|3477,3479
LAD|3480,3483
,|3483,3484
no|3485,3487
JVD|3488,3491
<EOL>|3493,3494
CARDIAC|3494,3501
:|3501,3502
RRR|3503,3506
,|3506,3507
S1|3508,3510
/|3510,3511
S2|3511,3513
,|3513,3514
no|3515,3517
murmurs|3518,3525
,|3525,3526
gallops|3527,3534
,|3534,3535
or|3536,3538
rubs|3539,3543
<EOL>|3545,3546
LUNG|3546,3550
:|3550,3551
CTAB|3552,3556
,|3556,3557
no|3558,3560
wheezes|3561,3568
,|3568,3569
rales|3570,3575
,|3575,3576
rhonchi|3577,3584
,|3584,3585
breathing|3586,3595
comfortably|3596,3607
<EOL>|3608,3609
without|3609,3616
use|3617,3620
of|3621,3623
accessory|3624,3633
muscles|3634,3641
<EOL>|3643,3644
ABDOMEN|3644,3651
:|3651,3652
nondistended|3653,3665
,|3665,3666
+|3667,3668
BS|3668,3670
,|3670,3671
nontender|3672,3681
in|3682,3684
all|3685,3688
quadrants|3689,3698
,|3698,3699
no|3700,3702
<EOL>|3703,3704
rebound|3704,3711
/|3711,3712
guarding|3712,3720
,|3720,3721
no|3722,3724
hepatosplenomegaly|3725,3743
<EOL>|3745,3746
EXTREMITIES|3746,3757
:|3757,3758
no|3759,3761
appreciable|3762,3773
lower|3774,3779
exam|3780,3784
swelling|3785,3793
althught|3794,3802
R|3803,3804
calf|3805,3809
<EOL>|3810,3811
is|3811,3813
tender|3814,3820
to|3821,3823
palpation|3824,3833
<EOL>|3833,3834
PULSES|3834,3840
:|3840,3841
2|3842,3843
+|3843,3844
DP|3845,3847
pulses|3848,3854
bilaterally|3855,3866
<EOL>|3868,3869
NEURO|3869,3874
:|3874,3875
CN|3876,3878
II|3879,3881
-|3881,3882
XII|3882,3885
intact|3886,3892
,|3892,3893
no|3894,3896
focal|3897,3902
deficits|3903,3911
<EOL>|3913,3914
SKIN|3914,3918
:|3918,3919
warm|3920,3924
and|3925,3928
well|3929,3933
perfused|3934,3942
,|3942,3943
no|3944,3946
excoriations|3947,3959
or|3960,3962
lesions|3963,3970
,|3970,3971
no|3972,3974
<EOL>|3975,3976
rashes|3976,3982
<EOL>|3982,3983
<EOL>|3983,3984
ON|3984,3986
DISCHARGE|3987,3996
:|3996,3997
<EOL>|3997,3998
<EOL>|3999,4000
Pertinent|4000,4009
Results|4010,4017
:|4017,4018
<EOL>|4018,4019
_|4019,4020
_|4020,4021
_|4021,4022
04|4023,4025
:|4025,4026
52PM|4026,4030
_|4033,4034
_|4034,4035
_|4035,4036
PTT|4037,4040
-|4040,4041
128|4041,4044
.|4044,4045
0|4045,4046
*|4046,4047
_|4048,4049
_|4049,4050
_|4050,4051
<EOL>|4051,4052
_|4052,4053
_|4053,4054
_|4054,4055
04|4056,4058
:|4058,4059
52PM|4059,4063
PLT|4066,4069
COUNT|4070,4075
-|4075,4076
150|4076,4079
<EOL>|4079,4080
_|4080,4081
_|4081,4082
_|4082,4083
04|4084,4086
:|4086,4087
52PM|4087,4091
NEUTS|4094,4099
-|4099,4100
56.6|4100,4104
_|4105,4106
_|4106,4107
_|4107,4108
MONOS|4109,4114
-|4114,4115
6.0|4115,4118
EOS|4119,4122
-|4122,4123
1.6|4123,4126
<EOL>|4127,4128
BASOS|4128,4133
-|4133,4134
0.7|4134,4137
<EOL>|4137,4138
_|4138,4139
_|4139,4140
_|4140,4141
04|4142,4144
:|4144,4145
52PM|4145,4149
GLUCOSE|4152,4159
-|4159,4160
130|4160,4163
*|4163,4164
UREA|4165,4169
N|4170,4171
-|4171,4172
16|4172,4174
CREAT|4175,4180
-|4180,4181
0.9|4181,4184
SODIUM|4185,4191
-|4191,4192
140|4192,4195
<EOL>|4196,4197
POTASSIUM|4197,4206
-|4206,4207
3.8|4207,4210
CHLORIDE|4211,4219
-|4219,4220
101|4220,4223
TOTAL|4224,4229
CO2|4230,4233
-|4233,4234
27|4234,4236
ANION|4237,4242
GAP|4243,4246
-|4246,4247
16|4247,4249
<EOL>|4249,4250
_|4250,4251
_|4251,4252
_|4252,4253
04|4254,4256
:|4256,4257
52PM|4257,4261
_|4264,4265
_|4265,4266
_|4266,4267
PTT|4268,4271
-|4271,4272
128|4272,4275
.|4275,4276
0|4276,4277
*|4277,4278
_|4279,4280
_|4280,4281
_|4281,4282
history|4283,4290
of|4291,4293
cerebral|4294,4302
aneurysm|4303,4311
,|4311,4312
recent|4313,4319
treatment|4320,4329
for|4330,4333
RLE|4334,4337
<EOL>|4338,4339
swelling|4339,4347
and|4348,4351
erythema|4352,4360
with|4361,4365
keflex|4366,4372
x|4373,4374
5|4375,4376
days|4377,4381
s|4382,4383
/|4383,4384
p|4384,4385
negative|4386,4394
RLE|4395,4398
U|4399,4400
/|4400,4401
S|4401,4402
<EOL>|4403,4404
now|4404,4407
presenting|4408,4418
with|4419,4423
shortness|4424,4433
of|4434,4436
breath|4437,4443
,|4443,4444
found|4445,4450
to|4451,4453
have|4454,4458
PE|4459,4461
.|4461,4462
<EOL>|4463,4464
<EOL>|4464,4465
#|4465,4466
Pulmonary|4467,4476
embolism|4477,4485
-|4485,4486
Treated|4486,4493
with|4494,4498
lovenox|4499,4506
while|4507,4512
hospitalized|4513,4525
,|4525,4526
<EOL>|4527,4528
transitioned|4528,4540
to|4541,4543
warfarin|4544,4552
at|4553,4555
discharge|4556,4565
.|4565,4566
Shortness|4567,4576
of|4577,4579
breath|4580,4586
<EOL>|4587,4588
resolved|4588,4596
while|4597,4602
hospitalized|4603,4615
without|4616,4623
the|4624,4627
need|4628,4632
for|4633,4636
supplemental|4637,4649
<EOL>|4650,4651
oxygen|4651,4657
.|4657,4658
<EOL>|4658,4659
<EOL>|4659,4660
#|4660,4661
History|4662,4669
of|4670,4672
cerebral|4673,4681
aneurysm|4682,4690
-|4690,4691
Per|4691,4694
Dr.|4695,4698
_|4699,4700
_|4700,4701
_|4701,4702
who|4703,4706
<EOL>|4707,4708
follows|4708,4715
the|4716,4719
patient|4720,4727
's|4727,4729
aneurysm|4730,4738
)|4738,4739
she|4740,4743
should|4744,4750
have|4751,4755
another|4756,4763
follow|4764,4770
<EOL>|4771,4772
up|4772,4774
MRI|4775,4778
(|4779,4780
last|4780,4784
was|4785,4788
_|4789,4790
_|4790,4791
_|4791,4792
to|4793,4795
assess|4796,4802
the|4803,4806
size|4807,4811
of|4812,4814
the|4815,4818
aneurysm|4819,4827
.|4827,4828
<EOL>|4829,4830
Careful|4830,4837
consideration|4838,4851
was|4852,4855
given|4856,4861
to|4862,4864
continuing|4865,4875
the|4876,4879
aspirin|4880,4887
which|4888,4893
<EOL>|4894,4895
she|4895,4898
takes|4899,4904
for|4905,4908
her|4909,4912
aneurysm|4913,4921
and|4922,4925
what|4926,4930
the|4931,4934
_|4935,4936
_|4936,4937
_|4937,4938
anti-coagulant|4939,4953
<EOL>|4954,4955
would|4955,4960
be|4961,4963
in|4964,4966
light|4967,4972
of|4973,4975
the|4976,4979
aneurysm|4980,4988
to|4989,4991
minimize|4992,5000
her|5001,5004
risk|5005,5009
of|5010,5012
<EOL>|5013,5014
bleeding|5014,5022
.|5022,5023
After|5024,5029
discussion|5030,5040
with|5041,5045
Dr.|5046,5049
_|5050,5051
_|5051,5052
_|5052,5053
Dr.|5054,5057
_|5058,5059
_|5059,5060
_|5060,5061
<EOL>|5062,5063
decision|5063,5071
was|5072,5075
made|5076,5080
to|5081,5083
bridge|5084,5090
to|5091,5093
Coumadin|5094,5102
with|5103,5107
lovenox|5108,5115
and|5116,5119
hold|5120,5124
<EOL>|5125,5126
the|5126,5129
aspirin|5130,5137
.|5137,5138
Her|5139,5142
MRA|5143,5146
which|5147,5152
was|5153,5156
performed|5157,5166
to|5167,5169
assess|5170,5176
the|5177,5180
size|5181,5185
of|5186,5188
<EOL>|5189,5190
the|5190,5193
aneurysm|5194,5202
while|5203,5208
the|5209,5212
patient|5213,5220
was|5221,5224
admitted|5225,5233
showed|5234,5240
stable|5241,5247
size|5248,5252
<EOL>|5253,5254
of|5254,5256
the|5257,5260
aneurysm|5261,5269
(|5270,5271
4mm|5271,5274
)|5274,5275
with|5276,5280
no|5281,5283
change|5284,5290
since|5291,5296
_|5297,5298
_|5298,5299
_|5299,5300
.|5300,5301
<EOL>|5301,5302
<EOL>|5302,5303
#|5303,5304
Hyperlipidemia|5304,5318
:|5318,5319
continued|5320,5329
atorvastatin|5330,5342
20|5343,5345
<EOL>|5346,5347
<EOL>|5348,5349
#|5349,5350
Depression|5350,5360
:|5360,5361
continued|5362,5371
home|5372,5376
sertaline|5377,5386
<EOL>|5388,5389
<EOL>|5389,5390
#|5390,5391
GERD|5391,5395
:|5395,5396
continued|5397,5406
home|5407,5411
omeprazole|5412,5422
<EOL>|5424,5425
<EOL>|5425,5426
#|5426,5427
Asthma|5427,5433
:|5433,5434
no|5435,5437
evidence|5438,5446
of|5447,5449
reactive|5450,5458
airway|5459,5465
disease|5466,5473
on|5474,5476
exam|5477,5481
,|5481,5482
<EOL>|5483,5484
continued|5484,5493
albuterol|5494,5503
inhaler|5504,5511
as|5512,5514
needed|5515,5521
.|5521,5522
<EOL>|5524,5525
<EOL>|5525,5526
Transitional|5526,5538
Issues|5539,5545
<EOL>|5545,5546
<EOL>|5546,5547
#|5547,5548
Anti-coagulation|5549,5565
:|5565,5566
Please|5567,5573
assess|5574,5580
optimal|5581,5588
length|5589,5595
of|5596,5598
treatment|5599,5608
<EOL>|5609,5610
for|5610,5613
the|5614,5617
patient|5618,5625
.|5625,5626
<EOL>|5626,5627
<EOL>|5627,5628
#|5628,5629
Cigarette|5630,5639
smoking|5640,5647
:|5647,5648
The|5649,5652
patient|5653,5660
quit|5661,5665
smoking|5666,5673
on|5674,5676
admission|5677,5686
to|5687,5689
<EOL>|5690,5691
the|5691,5694
ER|5695,5697
_|5698,5699
_|5699,5700
_|5700,5701
,|5701,5702
please|5703,5709
provide|5710,5717
encouragement|5718,5731
and|5732,5735
resources|5736,5745
<EOL>|5746,5747
regarding|5747,5756
smoking|5757,5764
cessation|5765,5774
.|5774,5775
<EOL>|5775,5776
<EOL>|5776,5777
<EOL>|5778,5779
Medications|5779,5790
on|5791,5793
Admission|5794,5803
:|5803,5804
<EOL>|5804,5805
The|5805,5808
Preadmission|5809,5821
Medication|5822,5832
list|5833,5837
is|5838,5840
accurate|5841,5849
and|5850,5853
complete|5854,5862
.|5862,5863
<EOL>|5863,5864
1.|5864,5866
Lovastatin|5867,5877
40|5878,5880
mg|5881,5883
oral|5884,5888
daily|5889,5894
<EOL>|5895,5896
2.|5896,5898
Sertraline|5899,5909
100|5910,5913
mg|5914,5916
PO|5917,5919
DAILY|5920,5925
<EOL>|5926,5927
3.|5927,5929
Aspirin|5930,5937
325|5938,5941
mg|5942,5944
PO|5945,5947
DAILY|5948,5953
<EOL>|5954,5955
4.|5955,5957
Omeprazole|5958,5968
20|5969,5971
mg|5972,5974
PO|5975,5977
BID|5978,5981
<EOL>|5982,5983
5.|5983,5985
albuterol|5986,5995
sulfate|5996,6003
90|6004,6006
mcg|6007,6010
/|6010,6011
actuation|6011,6020
inhalation|6021,6031
q4hrs|6032,6037
prn|6038,6041
<EOL>|6042,6043
wheezing|6043,6051
<EOL>|6052,6053
6.|6053,6055
Vitamin|6056,6063
D|6064,6065
_|6066,6067
_|6067,6068
_|6068,6069
UNIT|6070,6074
PO|6075,6077
DAILY|6078,6083
<EOL>|6084,6085
7.|6085,6087
Multivitamins|6088,6101
W|6102,6103
/|6103,6104
minerals|6104,6112
1|6113,6114
TAB|6115,6118
PO|6119,6121
DAILY|6122,6127
<EOL>|6128,6129
<EOL>|6129,6130
<EOL>|6131,6132
Discharge|6132,6141
Medications|6142,6153
:|6153,6154
<EOL>|6154,6155
1.|6155,6157
Lovastatin|6158,6168
40|6169,6171
mg|6172,6174
oral|6175,6179
daily|6180,6185
<EOL>|6186,6187
2.|6187,6189
Multivitamins|6190,6203
W|6204,6205
/|6205,6206
minerals|6206,6214
1|6215,6216
TAB|6217,6220
PO|6221,6223
DAILY|6224,6229
<EOL>|6230,6231
3.|6231,6233
Omeprazole|6234,6244
20|6245,6247
mg|6248,6250
PO|6251,6253
BID|6254,6257
<EOL>|6258,6259
4.|6259,6261
Sertraline|6262,6272
100|6273,6276
mg|6277,6279
PO|6280,6282
DAILY|6283,6288
<EOL>|6289,6290
5.|6290,6292
Vitamin|6293,6300
D|6301,6302
_|6303,6304
_|6304,6305
_|6305,6306
UNIT|6307,6311
PO|6312,6314
DAILY|6315,6320
<EOL>|6321,6322
6.|6322,6324
Enoxaparin|6325,6335
Sodium|6336,6342
110|6343,6346
mg|6347,6349
SC|6350,6352
Q12H|6353,6357
<EOL>|6358,6359
Start|6359,6364
:|6364,6365
Today|6366,6371
-|6372,6373
_|6374,6375
_|6375,6376
_|6376,6377
,|6377,6378
First|6379,6384
Dose|6385,6389
:|6389,6390
Next|6391,6395
Routine|6396,6403
Administration|6404,6418
<EOL>|6419,6420
Time|6420,6424
<EOL>|6425,6426
RX|6426,6428
*|6429,6430
enoxaparin|6430,6440
120|6441,6444
mg|6445,6447
/|6447,6448
0.8|6448,6451
mL|6452,6454
110|6455,6458
mg|6459,6461
Q12H|6462,6466
SQ|6467,6469
every|6470,6475
twelve|6476,6482
(|6483,6484
12|6484,6486
)|6486,6487
<EOL>|6488,6489
hours|6489,6494
Disp|6495,6499
#|6500,6501
*|6501,6502
12|6502,6504
Syringe|6505,6512
Refills|6513,6520
:|6520,6521
*|6521,6522
0|6522,6523
<EOL>|6523,6524
7.|6524,6526
Nicotine|6527,6535
Patch|6536,6541
14|6542,6544
mg|6545,6547
TD|6548,6550
DAILY|6551,6556
<EOL>|6557,6558
RX|6558,6560
*|6561,6562
nicotine|6562,6570
[|6571,6572
Nicoderm|6572,6580
CQ|6581,6583
]|6583,6584
14|6585,6587
mg|6588,6590
/|6590,6591
24|6591,6593
hour|6594,6598
Apply|6599,6604
one|6605,6608
patch|6609,6614
daily|6615,6620
<EOL>|6621,6622
Disp|6622,6626
#|6627,6628
*|6628,6629
30|6629,6631
Patch|6632,6637
Refills|6638,6645
:|6645,6646
*|6646,6647
0|6647,6648
<EOL>|6648,6649
8.|6649,6651
Warfarin|6652,6660
5|6661,6662
mg|6663,6665
PO|6666,6668
DAILY16|6669,6676
<EOL>|6677,6678
RX|6678,6680
*|6681,6682
warfarin|6682,6690
[|6691,6692
Coumadin|6692,6700
]|6700,6701
5|6702,6703
mg|6704,6706
1|6707,6708
tablet|6709,6715
(|6715,6716
s|6716,6717
)|6717,6718
by|6719,6721
mouth|6722,6727
qdaily|6728,6734
Disp|6735,6739
<EOL>|6740,6741
#|6741,6742
*|6742,6743
30|6743,6745
Tablet|6746,6752
Refills|6753,6760
:|6760,6761
*|6761,6762
0|6762,6763
<EOL>|6763,6764
9.|6764,6766
albuterol|6767,6776
sulfate|6777,6784
90|6785,6787
mcg|6788,6791
/|6791,6792
actuation|6792,6801
inhalation|6802,6812
q4hrs|6813,6818
prn|6819,6822
<EOL>|6823,6824
wheezing|6824,6832
<EOL>|6833,6834
10.|6834,6837
Outpatient|6838,6848
Lab|6849,6852
Work|6853,6857
<EOL>|6857,6858
Please|6858,6864
check|6865,6870
INR|6871,6874
on|6875,6877
_|6878,6879
_|6879,6880
_|6880,6881
.|6881,6882
<EOL>|6882,6883
<EOL>|6883,6884
ICD|6884,6887
-|6887,6888
9|6888,6889
:|6889,6890
415.1|6891,6896
<EOL>|6897,6898
<EOL>|6898,6899
Please|6899,6905
fax|6906,6909
result|6910,6916
to|6917,6919
Dr.|6920,6923
_|6924,6925
_|6925,6926
_|6926,6927
at|6928,6930
_|6931,6932
_|6932,6933
_|6933,6934
<EOL>|6934,6935
<EOL>|6935,6936
<EOL>|6937,6938
Discharge|6938,6947
Disposition|6948,6959
:|6959,6960
<EOL>|6960,6961
Home|6961,6965
<EOL>|6965,6966
<EOL>|6967,6968
Discharge|6968,6977
Diagnosis|6978,6987
:|6987,6988
<EOL>|6988,6989
Primary|6989,6996
Diagnosis|6997,7006
:|7006,7007
Pulmonary|7008,7017
embolism|7018,7026
<EOL>|7026,7027
<EOL>|7027,7028
Secondary|7028,7037
Diagnosis|7038,7047
:|7047,7048
Superficial|7049,7060
thrombophlebitis|7061,7077
<EOL>|7077,7078
<EOL>|7078,7079
Primary|7079,7086
Diagnosis|7087,7096
:|7096,7097
Pulmonary|7098,7107
embolism|7108,7116
<EOL>|7116,7117
<EOL>|7117,7118
Secondary|7118,7127
Diagnosis|7128,7137
:|7137,7138
Superficial|7139,7150
thrombophlebitis|7151,7167
<EOL>|7167,7168
<EOL>|7168,7169
<EOL>|7170,7171
Discharge|7171,7180
Condition|7181,7190
:|7190,7191
<EOL>|7191,7192
Mental|7192,7198
Status|7199,7205
:|7205,7206
Clear|7207,7212
and|7213,7216
coherent|7217,7225
.|7225,7226
<EOL>|7226,7227
Level|7227,7232
of|7233,7235
Consciousness|7236,7249
:|7249,7250
Alert|7251,7256
and|7257,7260
interactive|7261,7272
.|7272,7273
<EOL>|7273,7274
Activity|7274,7282
Status|7283,7289
:|7289,7290
Ambulatory|7291,7301
-|7302,7303
Independent|7304,7315
.|7315,7316
<EOL>|7316,7317
<EOL>|7317,7318
<EOL>|7319,7320
Discharge|7320,7329
Instructions|7330,7342
:|7342,7343
<EOL>|7343,7344
Dear|7344,7348
Ms.|7349,7352
_|7353,7354
_|7354,7355
_|7355,7356
,|7356,7357
<EOL>|7357,7358
<EOL>|7358,7359
It|7359,7361
was|7362,7365
a|7366,7367
pleasure|7368,7376
caring|7377,7383
for|7384,7387
you|7388,7391
at|7392,7394
the|7395,7398
_|7399,7400
_|7400,7401
_|7401,7402
<EOL>|7403,7404
_|7404,7405
_|7405,7406
_|7406,7407
.|7407,7408
You|7409,7412
were|7413,7417
admitted|7418,7426
because|7427,7434
of|7435,7437
a|7438,7439
pulmonary|7440,7449
<EOL>|7450,7451
embolism|7451,7459
(|7460,7461
blood|7461,7466
clot|7467,7471
in|7472,7474
the|7475,7478
lungs|7479,7484
)|7484,7485
.|7485,7486
We|7487,7489
treated|7490,7497
this|7498,7502
blood|7503,7508
clot|7509,7513
<EOL>|7514,7515
by|7515,7517
giving|7518,7524
you|7525,7528
anti-coagulation|7529,7545
medicine|7546,7554
which|7555,7560
you|7561,7564
will|7565,7569
continue|7570,7578
<EOL>|7579,7580
to|7580,7582
take|7583,7587
as|7588,7590
an|7591,7593
outpatient|7594,7604
.|7604,7605
You|7606,7609
should|7610,7616
continue|7617,7625
taking|7626,7632
this|7633,7637
<EOL>|7638,7639
medication|7639,7649
until|7650,7655
your|7656,7660
primary|7661,7668
care|7669,7673
doctor|7674,7680
(|7681,7682
_|7682,7683
_|7683,7684
_|7684,7685
)|7685,7686
says|7687,7691
it|7692,7694
<EOL>|7695,7696
is|7696,7698
okay|7699,7703
to|7704,7706
stop|7707,7711
(|7712,7713
likely|7713,7719
_|7720,7721
_|7721,7722
_|7722,7723
months|7724,7730
)|7730,7731
.|7731,7732
We|7733,7735
spoke|7736,7741
with|7742,7746
your|7747,7751
<EOL>|7752,7753
neurosurgeon|7753,7765
(|7766,7767
Dr|7767,7769
.|7769,7770
_|7771,7772
_|7772,7773
_|7773,7774
who|7775,7778
follows|7779,7786
your|7787,7791
aneurysm|7792,7800
and|7801,7804
he|7805,7807
<EOL>|7808,7809
recommended|7809,7820
that|7821,7825
you|7826,7829
get|7830,7833
a|7834,7835
repeat|7836,7842
MRI|7843,7846
of|7847,7849
your|7850,7854
brain|7855,7860
while|7861,7866
you|7867,7870
<EOL>|7871,7872
were|7872,7876
admitted|7877,7885
.|7885,7886
This|7887,7891
MRI|7892,7895
showed|7896,7902
that|7903,7907
the|7908,7911
anuerysm|7912,7920
has|7921,7924
not|7925,7928
changed|7929,7936
<EOL>|7937,7938
in|7938,7940
size|7941,7945
since|7946,7951
_|7952,7953
_|7953,7954
_|7954,7955
,|7955,7956
it|7957,7959
is|7960,7962
still|7963,7968
4mm|7969,7972
in|7973,7975
size|7976,7980
.|7980,7981
We|7982,7984
wish|7985,7989
you|7990,7993
all|7994,7997
the|7998,8001
<EOL>|8002,8003
_|8003,8004
_|8004,8005
_|8005,8006
in|8007,8009
your|8010,8014
continued|8015,8024
recovery|8025,8033
.|8033,8034
<EOL>|8034,8035
<EOL>|8035,8036
Sincerely|8036,8045
,|8045,8046
<EOL>|8046,8047
<EOL>|8047,8048
Your|8048,8052
_|8053,8054
_|8054,8055
_|8055,8056
Team|8057,8061
<EOL>|8061,8062
<EOL>|8063,8064
Followup|8064,8072
Instructions|8073,8085
:|8085,8086
<EOL>|8086,8087
_|8087,8088
_|8088,8089
_|8089,8090
<EOL>|8090,8091

