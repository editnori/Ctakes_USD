 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|29,33
No|34,36
:|36,37
_|40,41
_|41,42
_|42,43
<EOL>|43,44
<EOL>|45,46
Admission|46,55
Date|56,60
:|60,61
_|63,64
_|64,65
_|65,66
Discharge|80,89
Date|90,94
:|94,95
_|98,99
_|99,100
_|100,101
<EOL>|101,102
<EOL>|103,104
Date|104,108
of|109,111
Birth|112,117
:|117,118
_|120,121
_|121,122
_|122,123
Sex|136,139
:|139,140
F|143,144
<EOL>|144,145
<EOL>|146,147
Service|147,154
:|154,155
MEDICINE|156,164
<EOL>|164,165
<EOL>|166,167
lisinopril|179,189
<EOL>|189,190
<EOL>|191,192
Attending|192,201
:|201,202
_|203,204
_|204,205
_|205,206
.|206,207
<EOL>|207,208
<EOL>|209,210
Left|227,231
diabetic|232,240
foot|241,245
ulcer|246,251
<EOL>|251,252
<EOL>|253,254
Major|254,259
Surgical|260,268
or|269,271
Invasive|272,280
Procedure|281,290
:|290,291
<EOL>|291,292
Left|292,296
partial|297,304
hallux|305,311
amputation|312,322
<EOL>|322,323
<EOL>|323,324
<EOL>|325,326
_|354,355
_|355,356
_|356,357
with|358,362
poorly|363,369
controlled|370,380
diabetes|381,389
(|390,391
complicated|391,402
by|403,405
retinopathy|406,417
,|417,418
<EOL>|418,419
neuropathy|419,429
,|429,430
PAD|431,434
,|434,435
foot|436,440
ulcer|441,446
L|447,448
hallux|449,455
)|455,456
,|456,457
CAD|458,461
with|462,466
_|467,468
_|468,469
_|469,470
s|471,472
/|472,473
p|473,474
<EOL>|475,476
CABG|476,480
,|480,481
<EOL>|481,482
and|482,485
narcotics|486,495
agreement|496,505
,|505,506
presenting|507,517
with|518,522
3|523,524
days|525,529
subjective|530,540
<EOL>|541,542
fever|542,547
,|547,548
<EOL>|548,549
chills|549,555
,|555,556
increased|557,566
pain|567,571
in|572,574
L|575,576
great|577,582
toe|583,586
.|586,587
Pt|588,590
recently|591,599
had|600,603
ulcer|604,609
<EOL>|609,610
debrided|610,618
by|619,621
podiatry|622,630
on|631,633
_|634,635
_|635,636
_|636,637
,|637,638
ulcer|639,644
had|645,648
healed|649,655
to|656,658
the|659,662
size|663,667
of|668,670
a|671,672
<EOL>|672,673
pin|673,676
,|676,677
but|678,681
within|682,688
the|689,692
span|693,697
of|698,700
a|701,702
week|703,707
enlarged|708,716
to|717,719
size|720,724
of|725,727
a|728,729
tennis|730,736
<EOL>|736,737
ball|737,741
.|741,742
Presented|743,752
to|753,755
_|756,757
_|757,758
_|758,759
urgent|760,766
care|767,771
in|772,774
_|775,776
_|776,777
_|777,778
,|778,779
found|780,785
to|786,788
be|789,791
<EOL>|791,792
febrile|792,799
to|800,802
_|803,804
_|804,805
_|805,806
,|806,807
given|808,813
Tylenol|814,821
,|821,822
sent|823,827
to|828,830
ER|831,833
and|834,837
was|838,841
afebrile|842,850
and|851,854
<EOL>|854,855
normotensive|855,867
upon|868,872
arrival|873,880
,|880,881
though|882,888
sustained|889,898
tachycardia|899,910
to|911,913
low|914,917
<EOL>|917,918
100s|918,922
.|922,923
Podiatry|924,932
consulted|933,942
in|943,945
ER|946,948
,|948,949
wound|950,955
to|956,958
left|959,963
medial|964,970
hallux|971,977
<EOL>|977,978
probes|978,984
to|985,987
bone|988,992
w|993,994
/|994,995
high|996,1000
c|1001,1002
/|1002,1003
f|1003,1004
osteomyelitis|1005,1018
.|1018,1019
X-rays|1020,1026
show|1027,1031
bony|1032,1036
<EOL>|1036,1037
erosion|1037,1044
but|1045,1048
no|1049,1051
subcutaneous|1052,1064
gas|1065,1068
.|1068,1069
Plan|1070,1074
for|1075,1078
IV|1079,1081
antibiotics|1082,1093
and|1094,1097
<EOL>|1097,1098
partial|1098,1105
amputation|1106,1116
of|1117,1119
left|1120,1124
great|1125,1130
toe|1131,1134
tomorrow|1135,1143
(|1144,1145
_|1145,1146
_|1146,1147
_|1147,1148
)|1148,1149
.|1149,1150
_|1151,1152
_|1152,1153
_|1153,1154
n|1155,1156
/|1156,1157
v|1157,1158
,|1158,1159
<EOL>|1159,1160
abd|1160,1163
pain|1164,1168
,|1168,1169
diarrhea|1170,1178
,|1178,1179
excessive|1180,1189
urination|1190,1199
,|1199,1200
orthostasis|1201,1212
,|1212,1213
dyspnea|1214,1221
,|1221,1222
<EOL>|1222,1223
chest|1223,1228
pain|1229,1233
.|1233,1234
<EOL>|1234,1235
<EOL>|1235,1236
In|1236,1238
the|1239,1242
ED|1243,1245
:|1245,1246
<EOL>|1246,1247
<EOL>|1247,1248
Initial|1248,1255
vital|1256,1261
signs|1262,1267
were|1268,1272
notable|1273,1280
for|1281,1284
:|1284,1285
afebrile|1286,1294
,|1294,1295
tachycardia|1296,1307
to|1308,1310
<EOL>|1310,1311
118|1311,1314
,|1314,1315
normotensive|1316,1328
<EOL>|1328,1329
<EOL>|1329,1330
Exam|1330,1334
notable|1335,1342
for|1343,1346
:|1346,1347
<EOL>|1347,1348
PE|1348,1350
:|1350,1351
warm|1352,1356
,|1356,1357
slightly|1358,1366
diaphoretic|1367,1378
<EOL>|1378,1379
CV|1379,1381
:|1381,1382
RRR|1383,1386
,|1386,1387
+|1388,1389
S1|1389,1391
/|1391,1392
S2|1392,1394
<EOL>|1394,1395
Resp|1395,1399
:|1400,1401
lungs|1401,1406
clear|1407,1412
b|1413,1414
/|1414,1415
l|1415,1416
<EOL>|1416,1417
MSK|1417,1420
:|1420,1421
erythema|1422,1430
involving|1431,1440
L|1441,1442
big|1443,1446
toe|1447,1450
,|1450,1451
tracking|1452,1460
along|1461,1466
inferior|1467,1475
base|1476,1480
.|1480,1481
<EOL>|1481,1482
Tenderness|1482,1492
tracking|1493,1501
along|1502,1507
path|1508,1512
of|1513,1515
great|1516,1521
saphenous|1522,1531
on|1532,1534
L|1535,1536
calf|1537,1541
.|1541,1542
<EOL>|1542,1543
Limited|1543,1550
dorsiflexion|1551,1563
and|1564,1567
plantar|1568,1575
flexion|1576,1583
.|1583,1584
Limited|1585,1592
ROM|1593,1596
of|1597,1599
ankle|1600,1605
<EOL>|1605,1606
and|1606,1609
toe|1610,1613
.|1613,1614
<EOL>|1614,1615
Mental|1615,1621
Status|1622,1628
:|1628,1629
A|1630,1631
&|1631,1632
ox4|1632,1635
<EOL>|1635,1636
Lines|1636,1641
&|1642,1643
Drains|1644,1650
:|1650,1651
20g|1652,1655
L|1656,1657
hand|1658,1662
<EOL>|1662,1663
<EOL>|1663,1664
Labs|1664,1668
were|1669,1673
notable|1674,1681
for|1682,1685
:|1685,1686
<EOL>|1686,1687
<EOL>|1687,1688
136|1688,1691
98|1693,1695
26|1697,1699
*|1699,1700
AGap|1705,1709
=|1709,1710
20|1710,1712
<EOL>|1713,1714
-|1714,1715
-|1715,1716
-|1716,1717
-|1717,1718
-|1718,1719
-|1719,1720
-|1720,1721
-|1721,1722
-|1722,1723
-|1723,1724
-|1724,1725
-|1725,1726
<|1726,1727
266|1727,1730
*|1730,1731
<EOL>|1732,1733
4.2|1733,1736
18|1738,1740
*|1740,1741
1.6|1742,1745
*|1745,1746
<EOL>|1748,1749
<EOL>|1749,1750
Lactate|1750,1757
elevated|1758,1766
:|1766,1767
2.4|1768,1771
<EOL>|1771,1772
Whites|1772,1778
elevated|1779,1787
:|1787,1788
23.4|1789,1793
,|1793,1794
neut|1795,1799
predominance|1800,1812
<EOL>|1812,1813
<EOL>|1813,1814
Studies|1814,1821
performed|1822,1831
include|1832,1839
:|1839,1840
<EOL>|1840,1841
<EOL>|1841,1842
Xray|1842,1846
Foot|1847,1851
Ap|1852,1854
,|1854,1855
Lat|1855,1858
&|1859,1860
Obl|1861,1864
Left|1865,1869
(|1870,1871
prelim|1871,1877
read|1878,1882
)|1882,1883
:|1883,1884
Re-demonstration|1885,1901
of|1902,1904
<EOL>|1904,1905
ulceration|1905,1915
along|1916,1921
the|1922,1925
medial|1926,1932
distal|1933,1939
aspect|1940,1946
of|1947,1949
the|1950,1953
great|1954,1959
toe|1960,1963
and|1964,1967
<EOL>|1967,1968
erosion|1968,1975
along|1976,1981
the|1982,1985
medial|1986,1992
base|1993,1997
of|1998,2000
the|2001,2004
distal|2005,2011
phalanx|2012,2019
of|2020,2022
the|2023,2026
great|2027,2032
<EOL>|2032,2033
toe|2033,2036
perhaps|2037,2044
slightly|2045,2053
progressed|2054,2064
in|2065,2067
the|2068,2071
interval|2072,2080
.|2080,2081
Findings|2082,2090
again|2091,2096
<EOL>|2096,2097
remain|2097,2103
concerning|2104,2114
<EOL>|2115,2116
for|2116,2119
osteomyelitis|2120,2133
and|2134,2137
MRI|2138,2141
with|2142,2146
contrast|2147,2155
could|2156,2161
be|2162,2164
obtained|2165,2173
for|2174,2177
<EOL>|2177,2178
further|2178,2185
<EOL>|2186,2187
assessment|2187,2197
.|2197,2198
<EOL>|2199,2200
<EOL>|2200,2201
Patient|2201,2208
was|2209,2212
given|2213,2218
:|2218,2219
<EOL>|2219,2220
Piperacillin|2220,2232
-|2232,2233
Tazobactam|2233,2243
<EOL>|2245,2246
Vancomycin|2246,2256
<EOL>|2256,2257
<EOL>|2257,2258
Consults|2258,2266
:|2266,2267
Podiatry|2268,2276
<EOL>|2276,2277
<EOL>|2277,2278
Vitals|2278,2284
on|2285,2287
transfer|2288,2296
:|2296,2297
T100|2298,2302
.5|2302,2304
,|2304,2305
BP|2306,2308
154|2309,2312
/|2312,2313
80|2313,2315
,|2315,2316
HR117|2317,2322
,|2322,2323
RR18|2324,2328
,|2328,2329
99|2330,2332
Ra|2333,2335
<EOL>|2336,2337
<EOL>|2337,2338
Upon|2338,2342
arrival|2343,2350
to|2351,2353
the|2354,2357
floor|2358,2363
,|2363,2364
patient|2365,2372
resting|2373,2380
comfortably|2381,2392
in|2393,2395
bed|2396,2399
,|2399,2400
<EOL>|2400,2401
complains|2401,2410
of|2411,2413
chills|2414,2420
,|2420,2421
which|2422,2427
resolve|2428,2435
with|2436,2440
blankets|2441,2449
.|2449,2450
Left|2451,2455
foot|2456,2460
<EOL>|2460,2461
wrapped|2461,2468
in|2469,2471
gauze|2472,2477
dressing|2478,2486
,|2486,2487
very|2488,2492
tender|2493,2499
up|2500,2502
to|2503,2505
midcalf|2506,2513
.|2513,2514
<EOL>|2514,2515
<EOL>|2515,2516
REVIEW|2516,2522
OF|2523,2525
SYSTEMS|2526,2533
:|2533,2534
<EOL>|2534,2535
<EOL>|2535,2536
Complete|2536,2544
ROS|2545,2548
obtained|2549,2557
and|2558,2561
is|2562,2564
otherwise|2565,2574
negative|2575,2583
<EOL>|2583,2584
<EOL>|2585,2586
-|2608,2609
COPD|2609,2613
<EOL>|2613,2614
-|2614,2615
CAD|2615,2618
s|2619,2620
/|2620,2621
p|2621,2622
BMS|2623,2626
proximal|2627,2635
-|2635,2636
LAD|2636,2639
_|2640,2641
_|2641,2642
_|2642,2643
,|2643,2644
DES|2645,2648
to|2649,2651
mid|2652,2655
LAD|2656,2659
_|2660,2661
_|2661,2662
_|2662,2663
,|2663,2664
DES|2665,2668
to|2669,2671
edge|2672,2676
<EOL>|2677,2678
ISR|2678,2681
of|2682,2684
mid|2685,2688
LAD|2689,2692
DES|2693,2696
and|2697,2700
stenosis|2701,2709
distal|2710,2716
to|2717,2719
stent|2720,2725
_|2726,2727
_|2727,2728
_|2728,2729
,|2729,2730
DES|2731,2734
to|2735,2737
OM1|2738,2741
<EOL>|2742,2743
_|2743,2744
_|2744,2745
_|2745,2746
,|2746,2747
s|2748,2749
/|2749,2750
p|2750,2751
3|2752,2753
v|2754,2755
CABG|2756,2760
LIMA|2761,2765
-|2765,2766
LAD|2766,2769
,|2769,2770
SVG|2771,2774
-|2774,2775
OM1|2775,2778
,|2778,2779
<EOL>|2780,2781
_|2781,2782
_|2782,2783
_|2783,2784
<EOL>|2785,2786
-|2786,2787
HFpEF|2787,2792
<EOL>|2792,2793
-|2793,2794
Depression|2794,2804
<EOL>|2806,2807
-|2807,2808
DM|2808,2810
<EOL>|2812,2813
-|2813,2814
GERD|2814,2818
<EOL>|2820,2821
-|2821,2822
Hypertension|2822,2834
<EOL>|2834,2835
-|2835,2836
Migraines|2836,2845
<EOL>|2845,2846
-|2846,2847
Chronic|2847,2854
shoulder|2855,2863
pain|2864,2868
on|2869,2871
narcotics|2872,2881
<EOL>|2881,2882
-|2882,2883
OSA|2883,2886
<EOL>|2886,2887
-|2887,2888
Peripheral|2888,2898
neuropathy|2899,2909
<EOL>|2909,2910
-|2910,2911
Restless|2911,2919
leg|2920,2923
<EOL>|2923,2924
<EOL>|2925,2926
:|2940,2941
<EOL>|2941,2942
_|2942,2943
_|2943,2944
_|2944,2945
<EOL>|2945,2946
:|2960,2961
<EOL>|2961,2962
Patient|2962,2969
was|2970,2973
ward|2974,2978
of|2979,2981
the|2982,2985
_|2986,2987
_|2987,2988
_|2988,2989
,|2989,2990
does|2991,2995
n't|2995,2998
know|2999,3003
full|3004,3008
details|3009,3016
of|3017,3019
<EOL>|3020,3021
.|3035,3036
Mother|3037,3043
with|3044,3048
possible|3049,3057
alcohol|3058,3065
abuse|3066,3071
.|3071,3072
Father|3073,3079
<EOL>|3080,3081
deceased|3081,3089
at|3090,3092
_|3093,3094
_|3094,3095
_|3095,3096
from|3097,3101
Hodgkin|3102,3109
's|3109,3111
Disease|3112,3119
per|3120,3123
old|3124,3127
records|3128,3135
.|3135,3136
<EOL>|3136,3137
<EOL>|3138,3139
ADMISSION|3154,3163
EXAM|3164,3168
<EOL>|3168,3169
=|3169,3170
=|3170,3171
=|3171,3172
=|3172,3173
=|3173,3174
=|3174,3175
=|3175,3176
=|3176,3177
=|3177,3178
=|3178,3179
=|3179,3180
=|3180,3181
=|3181,3182
=|3182,3183
<EOL>|3183,3184
VITALS|3184,3190
:|3190,3191
T100|3192,3196
.5|3196,3198
,|3198,3199
BP|3200,3202
154|3203,3206
/|3206,3207
80|3207,3209
,|3209,3210
HR117|3211,3216
,|3216,3217
RR18|3218,3222
,|3222,3223
99|3224,3226
Ra|3227,3229
<EOL>|3230,3231
GENERAL|3231,3238
:|3238,3239
Alert|3240,3245
and|3246,3249
interactive|3250,3261
.|3261,3262
In|3263,3265
no|3266,3268
acute|3269,3274
distress|3275,3283
.|3283,3284
<EOL>|3284,3285
HEENT|3285,3290
:|3290,3291
NCAT|3292,3296
.|3296,3297
MMM|3298,3301
.|3301,3302
<EOL>|3302,3303
CARDIAC|3303,3310
:|3310,3311
RRR|3312,3315
,|3315,3316
no|3317,3319
MRG|3320,3323
<EOL>|3323,3324
LUNGS|3324,3329
:|3329,3330
Normal|3331,3337
WOB|3338,3341
,|3341,3342
CTA|3343,3346
B|3347,3348
/|3348,3349
L|3349,3350
<EOL>|3350,3351
ABDOMEN|3351,3358
:|3358,3359
Soft|3360,3364
,|3364,3365
nontender|3366,3375
to|3376,3378
deep|3379,3383
palpation|3384,3393
,|3393,3394
nondistended|3395,3407
,|3407,3408
<EOL>|3408,3409
normoactive|3409,3420
bowel|3421,3426
sounds|3427,3433
.|3433,3434
<EOL>|3434,3435
EXTREMITIES|3435,3446
:|3446,3447
left|3448,3452
foot|3453,3457
wrapped|3458,3465
in|3466,3468
gauze|3469,3474
dressing|3475,3483
,|3483,3484
mildly|3485,3491
<EOL>|3491,3492
erythematous|3492,3504
and|3505,3508
very|3509,3513
tender|3514,3520
up|3521,3523
to|3524,3526
lower|3527,3532
calf|3533,3537
,|3537,3538
RLE|3539,3542
no|3543,3545
edema|3546,3551
,|3551,3552
<EOL>|3552,3553
thready|3553,3560
DP|3561,3563
pulses|3564,3570
<EOL>|3570,3571
NEUROLOGIC|3571,3581
:|3581,3582
Sensory|3583,3590
and|3591,3594
motor|3595,3600
function|3601,3609
grossly|3610,3617
intact|3618,3624
.|3624,3625
<EOL>|3625,3626
<EOL>|3626,3627
DISCHARGE|3627,3636
EXAM|3637,3641
<EOL>|3641,3642
=|3642,3643
=|3643,3644
=|3644,3645
=|3645,3646
=|3646,3647
=|3647,3648
=|3648,3649
=|3649,3650
=|3650,3651
=|3651,3652
=|3652,3653
=|3653,3654
=|3654,3655
=|3655,3656
<EOL>|3656,3657
VS|3657,3659
:|3659,3660
98.5|3661,3665
,|3665,3666
134|3667,3670
/|3671,3672
75|3673,3675
,|3675,3676
75|3676,3678
,|3678,3679
18|3680,3682
,|3682,3683
97|3684,3686
%|3686,3687
RA|3688,3690
<EOL>|3690,3691
General|3691,3698
Appearance|3699,3709
:|3709,3710
Well|3711,3715
-|3715,3716
groomed|3716,3723
,|3723,3724
in|3725,3727
NAD|3728,3731
.|3731,3732
<EOL>|3732,3733
HEENT|3733,3738
:|3738,3739
Atraumatic|3740,3750
,|3750,3751
normocephalic|3752,3765
.|3765,3766
Sclera|3767,3773
anicteric|3774,3783
b|3784,3785
/|3785,3786
l|3786,3787
.|3787,3788
MMM|3789,3792
.|3792,3793
No|3794,3796
<EOL>|3796,3797
oropharyngeal|3797,3810
lesions|3811,3818
.|3818,3819
No|3820,3822
LAD|3823,3826
.|3826,3827
<EOL>|3827,3828
Lungs|3828,3833
:|3833,3834
Equal|3835,3840
chest|3841,3846
rise|3847,3851
.|3851,3852
Good|3853,3857
air|3858,3861
movement|3862,3870
.|3870,3871
No|3872,3874
increased|3875,3884
work|3885,3889
of|3890,3892
<EOL>|3892,3893
breathing|3893,3902
.|3902,3903
Decreased|3904,3913
breath|3914,3920
sounds|3921,3927
in|3928,3930
LLL|3931,3934
.|3934,3935
Rales|3936,3941
in|3942,3944
left|3945,3949
base|3950,3954
.|3954,3955
<EOL>|3956,3957
No|3957,3959
<EOL>|3959,3960
wheezes|3960,3967
or|3968,3970
rhonchi|3971,3978
.|3978,3979
<EOL>|3979,3980
CV|3980,3982
:|3982,3983
RRR|3984,3987
.|3987,3988
Normal|3989,3995
S1|3996,3998
,|3998,3999
S2|4000,4002
.|4002,4003
No|4004,4006
murmurs|4007,4014
,|4014,4015
gallops|4016,4023
,|4023,4024
or|4025,4027
rubs|4028,4032
.|4032,4033
No|4034,4036
carotid|4037,4044
<EOL>|4044,4045
bruits|4045,4051
b|4052,4053
/|4053,4054
l|4054,4055
.|4055,4056
+|4057,4058
2|4058,4059
carotid|4060,4067
pulses|4068,4074
b|4075,4076
/|4076,4077
l|4077,4078
,|4078,4079
+|4080,4081
2|4081,4082
radial|4083,4089
pulses|4090,4096
b|4097,4098
/|4098,4099
l|4099,4100
,|4100,4101
+|4102,4103
1|4103,4104
<EOL>|4104,4105
dorsalis|4105,4113
pedis|4114,4119
pulse|4120,4125
on|4126,4128
right|4129,4134
,|4134,4135
unable|4136,4142
to|4143,4145
palpate|4146,4153
on|4154,4156
left|4157,4161
due|4162,4165
to|4166,4168
<EOL>|4168,4169
surgical|4169,4177
bandage|4178,4185
.|4185,4186
<EOL>|4186,4187
Abdomen|4187,4194
:|4194,4195
Non-distended|4196,4209
.|4209,4210
Bowel|4211,4216
sounds|4217,4223
present|4224,4231
.|4231,4232
Soft|4233,4237
,|4237,4238
non-tender|4239,4249
<EOL>|4250,4251
to|4251,4253
<EOL>|4253,4254
palpation|4254,4263
throughout|4264,4274
.|4274,4275
<EOL>|4276,4277
Extremities|4277,4288
:|4288,4289
No|4290,4292
clubbing|4293,4301
or|4302,4304
cyanosis|4305,4313
.|4313,4314
Left|4315,4319
foot|4320,4324
dressing|4325,4333
clean|4334,4339
<EOL>|4339,4340
today|4340,4345
.|4345,4346
Erythema|4347,4355
and|4356,4359
edema|4360,4365
around|4366,4372
margin|4373,4379
of|4380,4382
surgical|4383,4391
site|4392,4396
is|4397,4399
<EOL>|4399,4400
improved|4400,4408
today|4409,4414
.|4414,4415
Suture|4416,4422
site|4423,4427
is|4428,4430
clean|4431,4436
with|4437,4441
no|4442,4444
pus|4445,4448
.|4448,4449
<EOL>|4449,4450
Skin|4450,4454
:|4454,4455
No|4456,4458
rashes|4459,4465
or|4466,4468
lesions|4469,4476
besides|4477,4484
surgical|4485,4493
site|4494,4498
.|4498,4499
<EOL>|4499,4500
Neuro|4500,4505
:|4505,4506
A|4507,4508
+|4508,4509
O|4509,4510
to|4511,4513
person|4514,4520
,|4520,4521
place|4522,4527
,|4527,4528
and|4529,4532
time|4533,4537
.|4537,4538
CN|4539,4541
III|4542,4545
-|4545,4546
XII|4546,4549
grossly|4550,4557
<EOL>|4558,4559
intact|4559,4565
.|4565,4566
<EOL>|4566,4567
<EOL>|4568,4569
Pertinent|4569,4578
Results|4579,4586
:|4586,4587
<EOL>|4587,4588
ADMISSION|4588,4597
LABS|4598,4602
<EOL>|4602,4603
=|4603,4604
=|4604,4605
=|4605,4606
=|4606,4607
=|4607,4608
=|4608,4609
=|4609,4610
=|4610,4611
=|4611,4612
=|4612,4613
=|4613,4614
=|4614,4615
=|4615,4616
=|4616,4617
<EOL>|4617,4618
_|4618,4619
_|4619,4620
_|4620,4621
05|4622,4624
:|4624,4625
50PM|4625,4629
BLOOD|4630,4635
WBC|4636,4639
-|4639,4640
23|4640,4642
.|4642,4643
4|4643,4644
*|4644,4645
RBC|4646,4649
-|4649,4650
4|4650,4651
.|4651,4652
01|4652,4654
Hgb|4655,4658
-|4658,4659
13.3|4659,4663
Hct|4664,4667
-|4667,4668
37.9|4668,4672
<EOL>|4673,4674
MCV|4674,4677
-|4677,4678
95|4678,4680
MCH|4681,4684
-|4684,4685
33|4685,4687
.|4687,4688
2|4688,4689
*|4689,4690
MCHC|4691,4695
-|4695,4696
35.1|4696,4700
RDW|4701,4704
-|4704,4705
12.0|4705,4709
RDWSD|4710,4715
-|4715,4716
42.1|4716,4720
Plt|4721,4724
_|4725,4726
_|4726,4727
_|4727,4728
<EOL>|4728,4729
_|4729,4730
_|4730,4731
_|4731,4732
05|4733,4735
:|4735,4736
50PM|4736,4740
BLOOD|4741,4746
Neuts|4747,4752
-|4752,4753
81|4753,4755
.|4755,4756
4|4756,4757
*|4757,4758
Lymphs|4759,4765
-|4765,4766
10|4766,4768
.|4768,4769
5|4769,4770
*|4770,4771
Monos|4772,4777
-|4777,4778
7.1|4778,4781
<EOL>|4782,4783
Eos|4783,4786
-|4786,4787
0|4787,4788
.|4788,4789
0|4789,4790
*|4790,4791
Baso|4792,4796
-|4796,4797
0.3|4797,4800
Im|4801,4803
_|4804,4805
_|4805,4806
_|4806,4807
AbsNeut|4808,4815
-|4815,4816
19|4816,4818
.|4818,4819
09|4819,4821
*|4821,4822
AbsLymp|4823,4830
-|4830,4831
2|4831,4832
.|4832,4833
47|4833,4835
<EOL>|4836,4837
AbsMono|4837,4844
-|4844,4845
1|4845,4846
.|4846,4847
66|4847,4849
*|4849,4850
AbsEos|4851,4857
-|4857,4858
0|4858,4859
.|4859,4860
00|4860,4862
*|4862,4863
AbsBaso|4864,4871
-|4871,4872
0.06|4872,4876
<EOL>|4876,4877
_|4877,4878
_|4878,4879
_|4879,4880
05|4881,4883
:|4883,4884
50PM|4884,4888
BLOOD|4889,4894
Glucose|4895,4902
-|4902,4903
266|4903,4906
*|4906,4907
UreaN|4908,4913
-|4913,4914
26|4914,4916
*|4916,4917
Creat|4918,4923
-|4923,4924
1|4924,4925
.|4925,4926
6|4926,4927
*|4927,4928
Na|4929,4931
-|4931,4932
136|4932,4935
<EOL>|4936,4937
K|4937,4938
-|4938,4939
4.2|4939,4942
Cl|4943,4945
-|4945,4946
98|4946,4948
HCO3|4949,4953
-|4953,4954
18|4954,4956
*|4956,4957
AnGap|4958,4963
-|4963,4964
20|4964,4966
*|4966,4967
<EOL>|4967,4968
_|4968,4969
_|4969,4970
_|4970,4971
05|4972,4974
:|4974,4975
50PM|4975,4979
BLOOD|4980,4985
CRP|4986,4989
-|4989,4990
180|4990,4993
.|4993,4994
1|4994,4995
*|4995,4996
<EOL>|4996,4997
_|4997,4998
_|4998,4999
_|4999,5000
07|5001,5003
:|5003,5004
45PM|5004,5008
BLOOD|5009,5014
_|5015,5016
_|5016,5017
_|5017,5018
pO2|5019,5022
-|5022,5023
22|5023,5025
*|5025,5026
pCO2|5027,5031
-|5031,5032
44|5032,5034
pH|5035,5037
-|5037,5038
7|5038,5039
.|5039,5040
32|5040,5042
*|5042,5043
<EOL>|5044,5045
calTCO2|5045,5052
-|5052,5053
24|5053,5055
Base|5056,5060
XS|5061,5063
-|5063,5064
-|5064,5065
4|5065,5066
<EOL>|5066,5067
_|5067,5068
_|5068,5069
_|5069,5070
05|5071,5073
:|5073,5074
50PM|5074,5078
BLOOD|5079,5084
Lactate|5085,5092
-|5092,5093
2|5093,5094
.|5094,5095
4|5095,5096
*|5096,5097
<EOL>|5097,5098
_|5098,5099
_|5099,5100
_|5100,5101
07|5102,5104
:|5104,5105
40PM|5105,5109
URINE|5110,5115
Color|5116,5121
-|5121,5122
Straw|5122,5127
Appear|5128,5134
-|5134,5135
Clear|5135,5140
Sp|5141,5143
_|5144,5145
_|5145,5146
_|5146,5147
<EOL>|5147,5148
_|5148,5149
_|5149,5150
_|5150,5151
07|5152,5154
:|5154,5155
40PM|5155,5159
URINE|5160,5165
Blood|5166,5171
-|5171,5172
NEG|5172,5175
Nitrite|5176,5183
-|5183,5184
NEG|5184,5187
Protein|5188,5195
-|5195,5196
TR|5196,5198
*|5198,5199
<EOL>|5200,5201
Glucose|5201,5208
-|5208,5209
1000|5209,5213
*|5213,5214
Ketone|5215,5221
-|5221,5222
TR|5222,5224
*|5224,5225
Bilirub|5226,5233
-|5233,5234
NEG|5234,5237
Urobiln|5238,5245
-|5245,5246
NEG|5246,5249
pH|5250,5252
-|5252,5253
6.0|5253,5256
<EOL>|5257,5258
Leuks|5258,5263
-|5263,5264
SM|5264,5266
*|5266,5267
<EOL>|5267,5268
_|5268,5269
_|5269,5270
_|5270,5271
07|5272,5274
:|5274,5275
40PM|5275,5279
URINE|5280,5285
RBC|5286,5289
-|5289,5290
4|5290,5291
*|5291,5292
WBC|5293,5296
-|5296,5297
7|5297,5298
*|5298,5299
Bacteri|5300,5307
-|5307,5308
FEW|5308,5311
*|5311,5312
Yeast|5313,5318
-|5318,5319
NONE|5319,5323
<EOL>|5324,5325
Epi|5325,5328
-|5328,5329
1|5329,5330
TransE|5331,5337
-|5337,5338
<|5338,5339
1|5339,5340
<EOL>|5340,5341
_|5341,5342
_|5342,5343
_|5343,5344
07|5345,5347
:|5347,5348
40PM|5348,5352
URINE|5353,5358
Mucous|5359,5365
-|5365,5366
RARE|5366,5370
*|5370,5371
<EOL>|5371,5372
<EOL>|5372,5373
PERTINENT|5373,5382
INTERVAL|5383,5391
LABS|5392,5396
<EOL>|5396,5397
=|5397,5398
=|5398,5399
=|5399,5400
=|5400,5401
=|5401,5402
=|5402,5403
=|5403,5404
=|5404,5405
=|5405,5406
=|5406,5407
=|5407,5408
=|5408,5409
=|5409,5410
=|5410,5411
=|5411,5412
=|5412,5413
=|5413,5414
=|5414,5415
=|5415,5416
=|5416,5417
=|5417,5418
=|5418,5419
=|5419,5420
<EOL>|5420,5421
_|5421,5422
_|5422,5423
_|5423,5424
09|5425,5427
:|5427,5428
48AM|5428,5432
BLOOD|5433,5438
ALT|5439,5442
-|5442,5443
25|5443,5445
AST|5446,5449
-|5449,5450
29|5450,5452
LD|5453,5455
(|5455,5456
LDH|5456,5459
)|5459,5460
-|5460,5461
210|5461,5464
AlkPhos|5465,5472
-|5472,5473
130|5473,5476
*|5476,5477
<EOL>|5478,5479
TotBili|5479,5486
-|5486,5487
0.8|5487,5490
<EOL>|5490,5491
<EOL>|5491,5492
DISCHARGE|5492,5501
LABS|5502,5506
<EOL>|5506,5507
=|5507,5508
=|5508,5509
=|5509,5510
=|5510,5511
=|5511,5512
=|5512,5513
=|5513,5514
=|5514,5515
=|5515,5516
=|5516,5517
=|5517,5518
=|5518,5519
=|5519,5520
=|5520,5521
<EOL>|5521,5522
_|5522,5523
_|5523,5524
_|5524,5525
07|5526,5528
:|5528,5529
17AM|5529,5533
BLOOD|5534,5539
WBC|5540,5543
-|5543,5544
9.9|5544,5547
RBC|5548,5551
-|5551,5552
3|5552,5553
.|5553,5554
07|5554,5556
*|5556,5557
Hgb|5558,5561
-|5561,5562
9|5562,5563
.|5563,5564
8|5564,5565
*|5565,5566
Hct|5567,5570
-|5570,5571
30|5571,5573
.|5573,5574
4|5574,5575
*|5575,5576
<EOL>|5577,5578
MCV|5578,5581
-|5581,5582
99|5582,5584
*|5584,5585
MCH|5586,5589
-|5589,5590
31.9|5590,5594
MCHC|5595,5599
-|5599,5600
32.2|5600,5604
RDW|5605,5608
-|5608,5609
12.3|5609,5613
RDWSD|5614,5619
-|5619,5620
44.2|5620,5624
Plt|5625,5628
_|5629,5630
_|5630,5631
_|5631,5632
<EOL>|5632,5633
_|5633,5634
_|5634,5635
_|5635,5636
07|5637,5639
:|5639,5640
29AM|5640,5644
BLOOD|5645,5650
Glucose|5651,5658
-|5658,5659
109|5659,5662
*|5662,5663
UreaN|5664,5669
-|5669,5670
18|5670,5672
Creat|5673,5678
-|5678,5679
1|5679,5680
.|5680,5681
2|5681,5682
*|5682,5683
Na|5684,5686
-|5686,5687
140|5687,5690
<EOL>|5691,5692
K|5692,5693
-|5693,5694
4.0|5694,5697
Cl|5698,5700
-|5700,5701
100|5701,5704
HCO3|5705,5709
-|5709,5710
25|5710,5712
AnGap|5713,5718
-|5718,5719
15|5719,5721
<EOL>|5721,5722
_|5722,5723
_|5723,5724
_|5724,5725
07|5726,5728
:|5728,5729
29AM|5729,5733
BLOOD|5734,5739
Calcium|5740,5747
-|5747,5748
8.8|5748,5751
Phos|5752,5756
-|5756,5757
4.3|5757,5760
Mg|5761,5763
-|5763,5764
1.8|5764,5767
<EOL>|5767,5768
_|5768,5769
_|5769,5770
_|5770,5771
07|5772,5774
:|5774,5775
29AM|5775,5779
BLOOD|5780,5785
CRP|5786,5789
-|5789,5790
44|5790,5792
.|5792,5793
6|5793,5794
*|5794,5795
<EOL>|5795,5796
<EOL>|5796,5797
IMAGING|5797,5804
<EOL>|5804,5805
=|5805,5806
=|5806,5807
=|5807,5808
=|5808,5809
=|5809,5810
=|5810,5811
=|5811,5812
<EOL>|5812,5813
LEFT|5813,5817
FOOT|5818,5822
XRAY|5823,5827
(|5828,5829
_|5829,5830
_|5830,5831
_|5831,5832
)|5832,5833
<EOL>|5833,5834
Re-demonstration|5849,5865
of|5866,5868
ulceration|5869,5879
along|5880,5885
the|5886,5889
medial|5890,5896
distal|5897,5903
aspect|5904,5910
of|5911,5913
<EOL>|5914,5915
the|5915,5918
great|5919,5924
toe|5925,5928
<EOL>|5928,5929
and|5929,5932
erosion|5933,5940
along|5941,5946
the|5947,5950
medial|5951,5957
base|5958,5962
of|5963,5965
the|5966,5969
distal|5970,5976
phalanx|5977,5984
of|5985,5987
the|5988,5991
<EOL>|5992,5993
great|5993,5998
toe|5999,6002
,|6002,6003
the|6004,6007
<EOL>|6007,6008
latter|6008,6014
of|6015,6017
which|6018,6023
is|6024,6026
perhaps|6027,6034
slightly|6035,6043
progressed|6044,6054
in|6055,6057
the|6058,6061
interval|6062,6070
.|6070,6071
<EOL>|6072,6073
again|6082,6087
<EOL>|6087,6088
remain|6088,6094
concerning|6095,6105
for|6106,6109
osteomyelitis|6110,6123
and|6124,6127
MRI|6128,6131
with|6132,6136
contrast|6137,6145
could|6146,6151
<EOL>|6152,6153
be|6153,6155
obtained|6156,6164
<EOL>|6164,6165
for|6165,6168
further|6169,6176
assessment|6177,6187
.|6187,6188
<EOL>|6188,6189
<EOL>|6189,6190
NIAS|6190,6194
(|6195,6196
_|6196,6197
_|6197,6198
_|6198,6199
)|6199,6200
<EOL>|6200,6201
-|6201,6202
-|6202,6203
-|6203,6204
-|6204,6205
-|6205,6206
-|6206,6207
-|6207,6208
-|6208,6209
-|6209,6210
-|6210,6211
-|6211,6212
-|6212,6213
-|6213,6214
-|6214,6215
-|6215,6216
<EOL>|6216,6217
:|6225,6226
<EOL>|6227,6228
<EOL>|6229,6230
On|6230,6232
the|6233,6236
right|6237,6242
side|6243,6247
,|6247,6248
triphasic|6249,6258
Doppler|6259,6266
waveforms|6267,6276
are|6277,6280
seen|6281,6285
in|6286,6288
the|6289,6292
<EOL>|6293,6294
right|6294,6299
femoral|6300,6307
,|6307,6308
<EOL>|6308,6309
popliteal|6309,6318
,|6318,6319
and|6320,6323
dorsalis|6324,6332
pedis|6333,6338
arteries|6339,6347
.|6347,6348
Absent|6350,6356
waveform|6357,6365
in|6366,6368
the|6369,6372
<EOL>|6373,6374
posterior|6374,6383
<EOL>|6383,6384
tibial|6384,6390
artery|6391,6397
.|6397,6398
<EOL>|6398,6399
The|6399,6402
right|6403,6408
ABI|6409,6412
was|6413,6416
1.6|6417,6420
,|6420,6421
artifactually|6422,6435
elevated|6436,6444
due|6445,6448
to|6449,6451
<EOL>|6452,6453
noncompressible|6453,6468
vessels|6469,6476
.|6476,6477
<EOL>|6477,6478
<EOL>|6479,6480
On|6480,6482
the|6483,6486
left|6487,6491
side|6492,6496
,|6496,6497
triphasic|6498,6507
Doppler|6508,6515
waveforms|6516,6525
are|6526,6529
seen|6530,6534
at|6535,6537
the|6538,6541
<EOL>|6542,6543
left|6543,6547
femoral|6548,6555
and|6556,6559
<EOL>|6559,6560
popliteal|6560,6569
arteries|6570,6578
.|6578,6579
Monophasic|6581,6591
waveforms|6592,6601
are|6602,6605
seen|6606,6610
in|6611,6613
the|6614,6617
<EOL>|6618,6619
posterior|6619,6628
tibial|6629,6635
and|6636,6639
<EOL>|6639,6640
dorsalis|6640,6648
pedis|6649,6654
arteries|6655,6663
.|6663,6664
<EOL>|6664,6665
The|6665,6668
left|6669,6673
ABI|6674,6677
could|6678,6683
not|6684,6687
be|6688,6690
calculated|6691,6701
<EOL>|6701,6702
<EOL>|6703,6704
Pulse|6704,6709
volume|6710,6716
recordings|6717,6727
showed|6728,6734
decreased|6735,6744
amplitudes|6745,6755
at|6756,6758
the|6759,6762
level|6763,6768
<EOL>|6769,6770
the|6770,6773
right|6774,6779
<EOL>|6779,6780
calf|6780,6784
,|6784,6785
ankle|6786,6791
and|6792,6795
metatarsal|6796,6806
.|6806,6807
<EOL>|6807,6808
<EOL>|6809,6810
Significant|6825,6836
bilateral|6837,6846
tibial|6847,6853
arterial|6854,6862
insufficiency|6863,6876
to|6877,6879
the|6880,6883
lower|6884,6889
<EOL>|6890,6891
extremities|6891,6902
<EOL>|6902,6903
at|6903,6905
rest|6906,6910
,|6910,6911
more|6912,6916
significant|6917,6928
on|6929,6931
the|6932,6935
right|6936,6941
side|6942,6946
.|6946,6947
<EOL>|6947,6948
<EOL>|6948,6949
CXR|6949,6952
(|6953,6954
_|6954,6955
_|6955,6956
_|6956,6957
)|6957,6958
<EOL>|6958,6959
-|6959,6960
-|6960,6961
-|6961,6962
-|6962,6963
-|6963,6964
-|6964,6965
-|6965,6966
-|6966,6967
-|6967,6968
-|6968,6969
-|6969,6970
-|6970,6971
-|6971,6972
-|6972,6973
<EOL>|6973,6974
Comparison|6989,6999
to|7000,7002
_|7003,7004
_|7004,7005
_|7005,7006
.|7006,7007
No|7009,7011
relevant|7012,7020
change|7021,7027
is|7028,7030
noted|7031,7036
.|7036,7037
<EOL>|7039,7040
Alignment|7040,7049
of|7050,7052
the|7053,7056
<EOL>|7056,7057
sternal|7057,7064
wires|7065,7070
is|7071,7073
unremarkable|7074,7086
.|7086,7087
Mild|7089,7093
elongation|7094,7104
of|7105,7107
the|7108,7111
<EOL>|7112,7113
descending|7113,7123
aorta|7124,7129
.|7129,7130
<EOL>|7131,7132
Borderline|7132,7142
size|7143,7147
of|7148,7150
the|7151,7154
heart|7155,7160
.|7160,7161
No|7163,7165
pleural|7166,7173
effusions|7174,7183
.|7183,7184
No|7186,7188
<EOL>|7189,7190
pneumonia|7190,7199
,|7199,7200
no|7201,7203
<EOL>|7203,7204
pulmonary|7204,7213
edema|7214,7219
.|7219,7220
<EOL>|7220,7221
<EOL>|7221,7222
MRI|7222,7225
LEFT|7226,7230
FOOT|7231,7235
(|7236,7237
_|7237,7238
_|7238,7239
_|7239,7240
)|7240,7241
<EOL>|7241,7242
1.|7258,7260
Nonenhancing|7261,7273
stump|7274,7279
soft|7280,7284
tissue|7285,7291
and|7292,7295
the|7296,7299
plantar|7300,7307
fat|7308,7311
pad|7312,7315
under|7316,7321
<EOL>|7322,7323
the|7323,7326
middle|7327,7333
<EOL>|7333,7334
phalanges|7334,7343
,|7343,7344
concerning|7345,7355
for|7356,7359
devitalized|7360,7371
tissue|7372,7378
.|7378,7379
No|7381,7383
evidence|7384,7392
of|7393,7395
<EOL>|7396,7397
drainable|7397,7406
<EOL>|7406,7407
abscess|7407,7414
.|7414,7415
<EOL>|7415,7416
2.|7416,7418
4|7419,7420
mm|7421,7423
focus|7424,7429
of|7430,7432
low|7433,7436
T1|7437,7439
signal|7440,7446
with|7447,7451
edema|7452,7457
at|7458,7460
the|7461,7464
most|7465,7469
distal|7470,7476
<EOL>|7477,7478
cortex|7478,7484
of|7485,7487
the|7488,7491
<EOL>|7491,7492
first|7492,7497
metatarsal|7498,7508
.|7508,7509
This|7511,7515
is|7516,7518
nonspecific|7519,7530
as|7531,7533
there|7534,7539
was|7540,7543
no|7544,7546
<EOL>|7547,7548
comparison|7548,7558
study|7559,7564
and|7565,7568
<EOL>|7568,7569
focus|7569,7574
of|7575,7577
osteomyelitis|7578,7591
can|7592,7595
not|7595,7598
be|7599,7601
excluded|7602,7610
.|7610,7611
<EOL>|7611,7612
3.|7612,7614
2|7615,7616
sinus|7617,7622
tracts|7623,7629
medial|7630,7636
to|7637,7639
the|7640,7643
head|7644,7648
of|7649,7651
the|7652,7655
first|7656,7661
metatarsal|7662,7672
,|7672,7673
<EOL>|7674,7675
status|7675,7681
post|7682,7686
<EOL>|7686,7687
amputation|7687,7697
at|7698,7700
the|7701,7704
first|7705,7710
MTP|7711,7714
with|7715,7719
postsurgical|7720,7732
changes|7733,7740
.|7740,7741
<EOL>|7741,7742
4.|7742,7744
Dorsal|7745,7751
swelling|7752,7760
and|7761,7764
diffuse|7765,7772
skin|7773,7777
edema|7778,7783
.|7783,7784
<EOL>|7784,7785
<EOL>|7785,7786
CXR|7786,7789
PICC|7790,7794
PLACEMENT|7795,7804
(|7805,7806
_|7806,7807
_|7807,7808
_|7808,7809
)|7809,7810
<EOL>|7810,7811
New|7826,7829
right|7830,7835
PICC|7836,7840
with|7841,7845
tip|7846,7849
projecting|7850,7860
over|7861,7865
the|7866,7869
junction|7870,7878
of|7879,7881
the|7882,7885
<EOL>|7886,7887
superior|7887,7895
vena|7896,7900
cava|7901,7905
<EOL>|7905,7906
and|7906,7909
right|7910,7915
atrium|7916,7922
.|7922,7923
No|7925,7927
pneumothorax|7928,7940
.|7940,7941
Clear|7943,7948
lungs|7949,7954
.|7954,7955
<EOL>|7955,7956
<EOL>|7956,7957
PATHOLOGY|7957,7966
<EOL>|7966,7967
=|7967,7968
=|7968,7969
=|7969,7970
=|7970,7971
=|7971,7972
=|7972,7973
=|7973,7974
=|7974,7975
=|7975,7976
=|7976,7977
<EOL>|7977,7978
SURGICAL|7978,7986
TISSUE|7987,7993
(|7994,7995
_|7995,7996
_|7996,7997
_|7997,7998
)|7998,7999
<EOL>|7999,8000
-|8000,8001
Bone|8002,8006
with|8007,8011
reparative|8012,8022
changes|8023,8030
,|8030,8031
consistent|8032,8042
with|8043,8047
chronic|8048,8055
<EOL>|8056,8057
osteomyelitis|8057,8070
.|8070,8071
<EOL>|8071,8072
-|8072,8073
There|8074,8079
is|8080,8082
no|8083,8085
evidence|8086,8094
of|8095,8097
acute|8098,8103
osteomyelitis|8104,8117
.|8117,8118
<EOL>|8119,8120
<EOL>|8120,8121
SURGICAL|8121,8129
TISSUE|8130,8136
(|8137,8138
_|8138,8139
_|8139,8140
_|8140,8141
)|8141,8142
<EOL>|8142,8143
1.|8143,8145
LEFT|8146,8150
GREAT|8151,8156
TOE|8157,8160
,|8160,8161
EXCISION|8162,8170
:|8170,8171
<EOL>|8171,8172
-|8172,8173
Acute|8174,8179
osteomyelitis|8180,8193
,|8193,8194
focal|8195,8200
.|8200,8201
<EOL>|8201,8202
-|8202,8203
Bone|8204,8208
with|8209,8213
reparative|8214,8224
changes|8225,8232
.|8232,8233
<EOL>|8233,8234
-|8234,8235
Skin|8236,8240
and|8241,8244
subcutis|8245,8253
with|8254,8258
ulceration|8259,8269
and|8270,8273
acute|8274,8279
inflammation|8280,8292
.|8292,8293
<EOL>|8293,8294
-|8294,8295
Atherosclerosis|8296,8311
,|8311,8312
severe|8313,8319
.|8319,8320
<EOL>|8320,8321
2.|8321,8323
PROXIMAL|8324,8332
PHALANX|8333,8340
BASE|8341,8345
MARGIN|8346,8352
,|8352,8353
LEFT|8354,8358
,|8358,8359
EXCISION|8360,8368
:|8368,8369
<EOL>|8369,8370
-|8370,8371
Bone|8372,8376
with|8377,8381
reparative|8382,8392
changes|8393,8400
.|8400,8401
<EOL>|8401,8402
-|8402,8403
There|8404,8409
is|8410,8412
no|8413,8415
evidence|8416,8424
of|8425,8427
acute|8428,8433
osteomyelitis|8434,8447
.|8447,8448
<EOL>|8448,8449
3.|8449,8451
PROXIMAL|8452,8460
PHALANX|8461,8468
,|8468,8469
LEFT|8470,8474
,|8474,8475
EXCISION|8476,8484
:|8484,8485
<EOL>|8485,8486
-|8486,8487
Bone|8488,8492
with|8493,8497
reparative|8498,8508
changes|8509,8516
.|8516,8517
<EOL>|8517,8518
-|8518,8519
There|8520,8525
is|8526,8528
no|8529,8531
evidence|8532,8540
of|8541,8543
acute|8544,8549
osteomyelitis|8550,8563
.|8563,8564
<EOL>|8564,8565
<EOL>|8565,8566
MICROBIOLOGY|8566,8578
<EOL>|8578,8579
=|8579,8580
=|8580,8581
=|8581,8582
=|8582,8583
=|8583,8584
=|8584,8585
=|8585,8586
=|8586,8587
=|8587,8588
=|8588,8589
=|8589,8590
=|8590,8591
<EOL>|8591,8592
_|8592,8593
_|8593,8594
_|8594,8595
10|8596,8598
:|8598,8599
00|8599,8601
am|8602,8604
TISSUE|8605,8611
PROXIMAL|8617,8625
PHALYNX|8626,8633
.|8633,8634
<EOL>|8635,8636
<EOL>|8636,8637
GRAM|8640,8644
STAIN|8645,8650
(|8651,8652
Final|8652,8657
_|8658,8659
_|8659,8660
_|8660,8661
:|8661,8662
<EOL>|8663,8664
2|8670,8671
+|8671,8672
_|8675,8676
_|8676,8677
_|8677,8678
per|8679,8682
1000X|8683,8688
FIELD|8689,8694
)|8694,8695
:|8695,8696
POLYMORPHONUCLEAR|8699,8716
<EOL>|8717,8718
LEUKOCYTES|8718,8728
.|8728,8729
<EOL>|8730,8731
2|8737,8738
+|8738,8739
_|8742,8743
_|8743,8744
_|8744,8745
per|8746,8749
1000X|8750,8755
FIELD|8756,8761
)|8761,8762
:|8762,8763
GRAM|8766,8770
POSITIVE|8771,8779
COCCI|8780,8785
IN|8786,8788
<EOL>|8789,8790
PAIRS|8790,8795
.|8795,8796
<EOL>|8797,8798
Reported|8804,8812
to|8813,8815
and|8816,8819
read|8820,8824
back|8825,8829
by|8830,8832
_|8833,8834
_|8834,8835
_|8835,8836
(|8837,8838
_|8838,8839
_|8839,8840
_|8840,8841
)|8841,8842
ON|8843,8845
<EOL>|8846,8847
_|8847,8848
_|8848,8849
_|8849,8850
AT|8851,8853
<EOL>|8853,8854
1|8860,8861
:|8861,8862
20PM|8862,8866
.|8866,8867
<EOL>|8868,8869
<EOL>|8869,8870
TISSUE|8873,8879
(|8880,8881
Final|8881,8886
_|8887,8888
_|8888,8889
_|8889,8890
:|8890,8891
<EOL>|8892,8893
STAPH|8899,8904
AUREUS|8905,8911
COAG|8912,8916
+|8917,8918
.|8918,8919
SPARSE|8923,8929
GROWTH|8930,8936
.|8936,8937
<EOL>|8938,8939
Susceptibility|8948,8962
testing|8963,8970
performed|8971,8980
on|8981,8983
culture|8984,8991
#|8992,8993
_|8994,8995
_|8995,8996
_|8996,8997
<EOL>|8998,8999
_|8999,9000
_|9000,9001
_|9001,9002
.|9002,9003
<EOL>|9004,9005
<EOL>|9005,9006
ANAEROBIC|9009,9018
CULTURE|9019,9026
(|9027,9028
Final|9028,9033
_|9034,9035
_|9035,9036
_|9036,9037
:|9037,9038
NO|9042,9044
ANAEROBES|9045,9054
ISOLATED|9055,9063
.|9063,9064
<EOL>|9065,9066
<EOL>|9066,9067
<EOL>|9067,9068
ACID|9071,9075
FAST|9076,9080
SMEAR|9081,9086
(|9087,9088
Final|9088,9093
_|9094,9095
_|9095,9096
_|9096,9097
:|9097,9098
<EOL>|9099,9100
NO|9106,9108
ACID|9109,9113
FAST|9114,9118
BACILLI|9119,9126
SEEN|9127,9131
ON|9132,9134
DIRECT|9135,9141
SMEAR|9142,9147
.|9147,9148
<EOL>|9149,9150
<EOL>|9150,9151
ACID|9154,9158
FAST|9159,9163
CULTURE|9164,9171
(|9172,9173
Preliminary|9173,9184
)|9184,9185
:|9185,9186
<EOL>|9187,9188
_|9188,9189
_|9189,9190
_|9190,9191
_|9191,9192
_|9192,9193
_|9193,9194
_|9194,9195
_|9195,9196
_|9196,9197
_|9197,9198
_|9198,9199
_|9199,9200
_|9200,9201
_|9201,9202
_|9202,9203
_|9203,9204
_|9204,9205
_|9205,9206
_|9206,9207
_|9207,9208
_|9208,9209
_|9209,9210
_|9210,9211
_|9211,9212
_|9212,9213
_|9213,9214
_|9214,9215
_|9215,9216
_|9216,9217
_|9217,9218
_|9218,9219
_|9219,9220
_|9220,9221
_|9221,9222
_|9222,9223
_|9223,9224
_|9224,9225
_|9225,9226
_|9226,9227
_|9227,9228
_|9228,9229
_|9229,9230
_|9230,9231
_|9231,9232
_|9232,9233
_|9233,9234
_|9234,9235
_|9235,9236
_|9236,9237
_|9237,9238
_|9238,9239
_|9239,9240
_|9240,9241
_|9241,9242
_|9242,9243
_|9243,9244
_|9244,9245
_|9245,9246
<EOL>|9246,9247
_|9247,9248
_|9248,9249
_|9249,9250
7|9251,9252
:|9252,9253
00|9253,9255
pm|9256,9258
BLOOD|9259,9264
CULTURE|9265,9272
<EOL>|9272,9273
<EOL>|9273,9274
*|9302,9303
*|9303,9304
FINAL|9304,9309
REPORT|9310,9316
_|9317,9318
_|9318,9319
_|9319,9320
<EOL>|9320,9321
<EOL>|9321,9322
Blood|9325,9330
Culture|9331,9338
,|9338,9339
Routine|9340,9347
(|9348,9349
Final|9349,9354
_|9355,9356
_|9356,9357
_|9357,9358
:|9358,9359
NO|9363,9365
GROWTH|9366,9372
.|9372,9373
<EOL>|9374,9375
_|9375,9376
_|9376,9377
_|9377,9378
_|9378,9379
_|9379,9380
_|9380,9381
_|9381,9382
_|9382,9383
_|9383,9384
_|9384,9385
_|9385,9386
_|9386,9387
_|9387,9388
_|9388,9389
_|9389,9390
_|9390,9391
_|9391,9392
_|9392,9393
_|9393,9394
_|9394,9395
_|9395,9396
_|9396,9397
_|9397,9398
_|9398,9399
_|9399,9400
_|9400,9401
_|9401,9402
_|9402,9403
_|9403,9404
_|9404,9405
_|9405,9406
_|9406,9407
_|9407,9408
_|9408,9409
_|9409,9410
_|9410,9411
_|9411,9412
_|9412,9413
_|9413,9414
_|9414,9415
_|9415,9416
_|9416,9417
_|9417,9418
_|9418,9419
_|9419,9420
_|9420,9421
_|9421,9422
_|9422,9423
_|9423,9424
_|9424,9425
_|9425,9426
_|9426,9427
_|9427,9428
_|9428,9429
_|9429,9430
_|9430,9431
_|9431,9432
_|9432,9433
<EOL>|9433,9434
_|9434,9435
_|9435,9436
_|9436,9437
5|9438,9439
:|9439,9440
38|9440,9442
pm|9443,9445
BLOOD|9446,9451
CULTURE|9452,9459
<EOL>|9459,9460
<EOL>|9460,9461
*|9489,9490
*|9490,9491
FINAL|9491,9496
REPORT|9497,9503
_|9504,9505
_|9505,9506
_|9506,9507
<EOL>|9507,9508
<EOL>|9508,9509
Blood|9512,9517
Culture|9518,9525
,|9525,9526
Routine|9527,9534
(|9535,9536
Final|9536,9541
_|9542,9543
_|9543,9544
_|9544,9545
:|9545,9546
NO|9550,9552
GROWTH|9553,9559
.|9559,9560
<EOL>|9561,9562
_|9562,9563
_|9563,9564
_|9564,9565
_|9565,9566
_|9566,9567
_|9567,9568
_|9568,9569
_|9569,9570
_|9570,9571
_|9571,9572
_|9572,9573
_|9573,9574
_|9574,9575
_|9575,9576
_|9576,9577
_|9577,9578
_|9578,9579
_|9579,9580
_|9580,9581
_|9581,9582
_|9582,9583
_|9583,9584
_|9584,9585
_|9585,9586
_|9586,9587
_|9587,9588
_|9588,9589
_|9589,9590
_|9590,9591
_|9591,9592
_|9592,9593
_|9593,9594
_|9594,9595
_|9595,9596
_|9596,9597
_|9597,9598
_|9598,9599
_|9599,9600
_|9600,9601
_|9601,9602
_|9602,9603
_|9603,9604
_|9604,9605
_|9605,9606
_|9606,9607
_|9607,9608
_|9608,9609
_|9609,9610
_|9610,9611
_|9611,9612
_|9612,9613
_|9613,9614
_|9614,9615
_|9615,9616
_|9616,9617
_|9617,9618
_|9618,9619
_|9619,9620
<EOL>|9620,9621
_|9621,9622
_|9622,9623
_|9623,9624
12|9625,9627
:|9627,9628
34|9628,9630
am|9631,9633
BLOOD|9634,9639
CULTURE|9640,9647
<EOL>|9647,9648
<EOL>|9648,9649
*|9677,9678
*|9678,9679
FINAL|9679,9684
REPORT|9685,9691
_|9692,9693
_|9693,9694
_|9694,9695
<EOL>|9695,9696
<EOL>|9696,9697
Blood|9700,9705
Culture|9706,9713
,|9713,9714
Routine|9715,9722
(|9723,9724
Final|9724,9729
_|9730,9731
_|9731,9732
_|9732,9733
:|9733,9734
NO|9738,9740
GROWTH|9741,9747
.|9747,9748
<EOL>|9749,9750
_|9750,9751
_|9751,9752
_|9752,9753
_|9753,9754
_|9754,9755
_|9755,9756
_|9756,9757
_|9757,9758
_|9758,9759
_|9759,9760
_|9760,9761
_|9761,9762
_|9762,9763
_|9763,9764
_|9764,9765
_|9765,9766
_|9766,9767
_|9767,9768
_|9768,9769
_|9769,9770
_|9770,9771
_|9771,9772
_|9772,9773
_|9773,9774
_|9774,9775
_|9775,9776
_|9776,9777
_|9777,9778
_|9778,9779
_|9779,9780
_|9780,9781
_|9781,9782
_|9782,9783
_|9783,9784
_|9784,9785
_|9785,9786
_|9786,9787
_|9787,9788
_|9788,9789
_|9789,9790
_|9790,9791
_|9791,9792
_|9792,9793
_|9793,9794
_|9794,9795
_|9795,9796
_|9796,9797
_|9797,9798
_|9798,9799
_|9799,9800
_|9800,9801
_|9801,9802
_|9802,9803
_|9803,9804
_|9804,9805
_|9805,9806
_|9806,9807
_|9807,9808
<EOL>|9808,9809
_|9809,9810
_|9810,9811
_|9811,9812
11|9813,9815
:|9815,9816
00|9816,9818
pm|9819,9821
BLOOD|9822,9827
CULTURE|9828,9835
<EOL>|9835,9836
<EOL>|9836,9837
*|9865,9866
*|9866,9867
FINAL|9867,9872
REPORT|9873,9879
_|9880,9881
_|9881,9882
_|9882,9883
<EOL>|9883,9884
<EOL>|9884,9885
Blood|9888,9893
Culture|9894,9901
,|9901,9902
Routine|9903,9910
(|9911,9912
Final|9912,9917
_|9918,9919
_|9919,9920
_|9920,9921
:|9921,9922
NO|9926,9928
GROWTH|9929,9935
.|9935,9936
<EOL>|9937,9938
_|9938,9939
_|9939,9940
_|9940,9941
_|9941,9942
_|9942,9943
_|9943,9944
_|9944,9945
_|9945,9946
_|9946,9947
_|9947,9948
_|9948,9949
_|9949,9950
_|9950,9951
_|9951,9952
_|9952,9953
_|9953,9954
_|9954,9955
_|9955,9956
_|9956,9957
_|9957,9958
_|9958,9959
_|9959,9960
_|9960,9961
_|9961,9962
_|9962,9963
_|9963,9964
_|9964,9965
_|9965,9966
_|9966,9967
_|9967,9968
_|9968,9969
_|9969,9970
_|9970,9971
_|9971,9972
_|9972,9973
_|9973,9974
_|9974,9975
_|9975,9976
_|9976,9977
_|9977,9978
_|9978,9979
_|9979,9980
_|9980,9981
_|9981,9982
_|9982,9983
_|9983,9984
_|9984,9985
_|9985,9986
_|9986,9987
_|9987,9988
_|9988,9989
_|9989,9990
_|9990,9991
_|9991,9992
_|9992,9993
_|9993,9994
_|9994,9995
_|9995,9996
<EOL>|9996,9997
_|9997,9998
_|9998,9999
_|9999,10000
12|10001,10003
:|10003,10004
18|10004,10006
am|10007,10009
BLOOD|10010,10015
CULTURE|10016,10023
<EOL>|10023,10024
<EOL>|10024,10025
*|10053,10054
*|10054,10055
FINAL|10055,10060
REPORT|10061,10067
_|10068,10069
_|10069,10070
_|10070,10071
<EOL>|10071,10072
<EOL>|10072,10073
Blood|10076,10081
Culture|10082,10089
,|10089,10090
Routine|10091,10098
(|10099,10100
Final|10100,10105
_|10106,10107
_|10107,10108
_|10108,10109
:|10109,10110
NO|10114,10116
GROWTH|10117,10123
.|10123,10124
<EOL>|10125,10126
_|10126,10127
_|10127,10128
_|10128,10129
_|10129,10130
_|10130,10131
_|10131,10132
_|10132,10133
_|10133,10134
_|10134,10135
_|10135,10136
_|10136,10137
_|10137,10138
_|10138,10139
_|10139,10140
_|10140,10141
_|10141,10142
_|10142,10143
_|10143,10144
_|10144,10145
_|10145,10146
_|10146,10147
_|10147,10148
_|10148,10149
_|10149,10150
_|10150,10151
_|10151,10152
_|10152,10153
_|10153,10154
_|10154,10155
_|10155,10156
_|10156,10157
_|10157,10158
_|10158,10159
_|10159,10160
_|10160,10161
_|10161,10162
_|10162,10163
_|10163,10164
_|10164,10165
_|10165,10166
_|10166,10167
_|10167,10168
_|10168,10169
_|10169,10170
_|10170,10171
_|10171,10172
_|10172,10173
_|10173,10174
_|10174,10175
_|10175,10176
_|10176,10177
_|10177,10178
_|10178,10179
_|10179,10180
_|10180,10181
_|10181,10182
_|10182,10183
_|10183,10184
<EOL>|10184,10185
_|10185,10186
_|10186,10187
_|10187,10188
10|10189,10191
:|10191,10192
53|10192,10194
pm|10195,10197
BLOOD|10198,10203
CULTURE|10204,10211
<EOL>|10211,10212
<EOL>|10212,10213
*|10241,10242
*|10242,10243
FINAL|10243,10248
REPORT|10249,10255
_|10256,10257
_|10257,10258
_|10258,10259
<EOL>|10259,10260
<EOL>|10260,10261
Blood|10264,10269
Culture|10270,10277
,|10277,10278
Routine|10279,10286
(|10287,10288
Final|10288,10293
_|10294,10295
_|10295,10296
_|10296,10297
:|10297,10298
NO|10302,10304
GROWTH|10305,10311
.|10311,10312
<EOL>|10313,10314
<EOL>|10314,10315
<EOL>|10316,10317
=|10340,10341
=|10341,10342
=|10342,10343
=|10343,10344
=|10344,10345
=|10345,10346
=|10346,10347
=|10347,10348
=|10348,10349
=|10349,10350
=|10350,10351
=|10351,10352
=|10352,10353
<EOL>|10353,10354
SUMMARY|10354,10361
<EOL>|10361,10362
=|10362,10363
=|10363,10364
=|10364,10365
=|10365,10366
=|10366,10367
=|10367,10368
=|10368,10369
=|10369,10370
=|10370,10371
=|10371,10372
=|10372,10373
=|10373,10374
=|10374,10375
<EOL>|10375,10376
<EOL>|10376,10377
_|10377,10378
_|10378,10379
_|10379,10380
yo|10381,10383
F|10384,10385
with|10386,10390
hx|10391,10393
of|10394,10396
DMII|10397,10401
,|10401,10402
HTN|10403,10406
who|10407,10410
presented|10411,10420
with|10421,10425
diabetic|10426,10434
foot|10435,10439
<EOL>|10440,10441
ulcer|10441,10446
on|10447,10449
her|10450,10453
left|10454,10458
hallux|10459,10465
complicated|10466,10477
by|10478,10480
osteomyelitis|10481,10494
.|10494,10495
She|10496,10499
<EOL>|10500,10501
underwent|10501,10510
surgical|10511,10519
debridement|10520,10531
and|10532,10535
partial|10536,10543
tissue|10544,10550
and|10551,10554
bone|10555,10559
<EOL>|10560,10561
removal|10561,10568
on|10569,10571
_|10572,10573
_|10573,10574
_|10574,10575
.|10575,10576
However|10577,10584
the|10585,10588
infection|10589,10598
persisted|10599,10608
,|10608,10609
and|10610,10613
she|10614,10617
<EOL>|10618,10619
underwent|10619,10628
left|10629,10633
hallux|10634,10640
amputation|10641,10651
on|10652,10654
_|10655,10656
_|10656,10657
_|10657,10658
.|10658,10659
She|10660,10663
was|10664,10667
started|10668,10675
<EOL>|10676,10677
on|10677,10679
IV|10680,10682
nafcillin|10683,10692
for|10693,10696
MSSA|10697,10701
infection|10702,10711
with|10712,10716
plan|10717,10721
to|10722,10724
continue|10725,10733
home|10734,10738
<EOL>|10739,10740
infusions|10740,10749
of|10750,10752
nafcillin|10753,10762
until|10763,10768
at|10769,10771
least|10772,10777
_|10778,10779
_|10779,10780
_|10780,10781
<EOL>|10781,10782
<EOL>|10782,10783
ACTIVE|10783,10789
ISSUES|10790,10796
<EOL>|10796,10797
=|10797,10798
=|10798,10799
=|10799,10800
=|10800,10801
=|10801,10802
=|10802,10803
=|10803,10804
=|10804,10805
=|10805,10806
=|10806,10807
=|10807,10808
=|10808,10809
=|10809,10810
<EOL>|10810,10811
#|10811,10812
Osteomyelitis|10812,10825
of|10826,10828
left|10829,10833
hallux|10834,10840
:|10840,10841
Due|10842,10845
to|10846,10848
diabetic|10849,10857
ulcer|10858,10863
of|10864,10866
left|10867,10871
<EOL>|10872,10873
hallux|10873,10879
.|10879,10880
Patient|10881,10888
underwent|10889,10898
partial|10899,10906
left|10907,10911
hallux|10912,10918
amputation|10919,10929
on|10930,10932
_|10933,10934
_|10934,10935
_|10935,10936
<EOL>|10937,10938
by|10938,10940
podiatry|10941,10949
.|10949,10950
She|10951,10954
was|10955,10958
initially|10959,10968
placed|10969,10975
on|10976,10978
IV|10979,10981
Vancomycin|10982,10992
,|10992,10993
Flagyl|10994,11000
,|11000,11001
<EOL>|11002,11003
and|11003,11006
cefepime|11007,11015
.|11015,11016
Initial|11017,11024
surgical|11025,11033
cultures|11034,11042
came|11043,11047
back|11048,11052
positive|11053,11061
for|11062,11065
<EOL>|11066,11067
MSSA|11067,11071
,|11071,11072
so|11073,11075
was|11076,11079
changed|11080,11087
to|11088,11090
IV|11091,11093
nafcillin|11094,11103
.|11103,11104
Patient|11105,11112
continued|11113,11122
to|11123,11125
be|11126,11128
<EOL>|11129,11130
afebrile|11130,11138
,|11138,11139
but|11140,11143
her|11144,11147
left|11148,11152
foot|11153,11157
continued|11158,11167
to|11168,11170
have|11171,11175
erythema|11176,11184
,|11184,11185
edema|11186,11191
,|11191,11192
<EOL>|11193,11194
pain|11194,11198
,|11198,11199
and|11200,11203
the|11204,11207
ulcer|11208,11213
was|11214,11217
not|11218,11221
healing|11222,11229
well|11230,11234
.|11234,11235
There|11236,11241
was|11242,11245
concern|11246,11253
for|11254,11257
<EOL>|11258,11259
poor|11259,11263
arterial|11264,11272
blood|11273,11278
flow|11279,11283
and|11284,11287
therefore|11288,11297
underwent|11298,11307
noninvasive|11308,11319
<EOL>|11320,11321
arterial|11321,11329
studies|11330,11337
on|11338,11340
bilateral|11341,11350
lower|11351,11356
extremities|11357,11368
.|11368,11369
The|11370,11373
studies|11374,11381
<EOL>|11382,11383
showed|11383,11389
mild|11390,11394
atherosclerotic|11395,11410
disease|11411,11418
in|11419,11421
her|11422,11425
left|11426,11430
leg|11431,11434
and|11435,11438
foot|11439,11443
,|11443,11444
<EOL>|11445,11446
and|11446,11449
severe|11450,11456
atherosclerotic|11457,11472
disease|11473,11480
in|11481,11483
her|11484,11487
right|11488,11493
leg|11494,11497
and|11498,11501
foot|11502,11506
.|11506,11507
<EOL>|11508,11509
Vascular|11509,11517
surgery|11518,11525
was|11526,11529
consulted|11530,11539
for|11540,11543
potential|11544,11553
intervention|11554,11566
,|11566,11567
but|11568,11571
<EOL>|11572,11573
they|11573,11577
felt|11578,11582
that|11583,11587
no|11588,11590
further|11591,11598
vascular|11599,11607
intervention|11608,11620
was|11621,11624
warranted|11625,11634
<EOL>|11635,11636
prior|11636,11641
to|11642,11644
podiatric|11645,11654
surgery|11655,11662
.|11662,11663
The|11664,11667
patient|11668,11675
was|11676,11679
brought|11680,11687
back|11688,11692
to|11693,11695
the|11696,11699
<EOL>|11700,11701
OR|11701,11703
by|11704,11706
podiatry|11707,11715
on|11716,11718
_|11719,11720
_|11720,11721
_|11721,11722
for|11723,11726
total|11727,11732
left|11733,11737
hallux|11738,11744
amputation|11745,11755
<EOL>|11756,11757
given|11757,11762
lack|11763,11767
of|11768,11770
clinical|11771,11779
improvement|11780,11791
.|11791,11792
Her|11793,11796
_|11797,11798
_|11798,11799
_|11799,11800
blood|11801,11806
cell|11807,11811
count|11812,11817
<EOL>|11818,11819
continued|11819,11828
to|11829,11831
down|11832,11836
trend|11837,11842
.|11842,11843
The|11844,11847
pathology|11848,11857
report|11858,11864
showed|11865,11871
clean|11872,11877
<EOL>|11878,11879
margins|11879,11886
.|11886,11887
However|11888,11895
,|11895,11896
patient|11897,11904
was|11905,11908
continuing|11909,11919
to|11920,11922
have|11923,11927
pain|11928,11932
,|11932,11933
and|11934,11937
there|11938,11943
<EOL>|11944,11945
was|11945,11948
increased|11949,11958
erythema|11959,11967
and|11968,11971
swelling|11972,11980
around|11981,11987
surgical|11988,11996
site|11997,12001
.|12001,12002
An|12003,12005
MRI|12006,12009
<EOL>|12010,12011
of|12011,12013
the|12014,12017
left|12018,12022
foot|12023,12027
was|12028,12031
done|12032,12036
,|12036,12037
which|12038,12043
showed|12044,12050
devitalization|12051,12065
of|12066,12068
the|12069,12072
<EOL>|12073,12074
surgical|12074,12082
flap|12083,12087
,|12087,12088
some|12089,12093
edema|12094,12099
,|12099,12100
and|12101,12104
a|12105,12106
hyperintense|12107,12119
focal|12120,12125
spot|12126,12130
at|12131,12133
the|12134,12137
<EOL>|12138,12139
site|12139,12143
of|12144,12146
the|12147,12150
surgery|12151,12158
.|12158,12159
There|12160,12165
were|12166,12170
no|12171,12173
signs|12174,12179
of|12180,12182
abscess|12183,12190
or|12191,12193
fluid|12194,12199
<EOL>|12200,12201
collection|12201,12211
.|12211,12212
Podiatry|12213,12221
team|12222,12226
felt|12227,12231
patient|12232,12239
did|12240,12243
not|12244,12247
need|12248,12252
any|12253,12256
acute|12257,12262
<EOL>|12263,12264
surgical|12264,12272
intervention|12273,12285
and|12286,12289
will|12290,12294
have|12295,12299
close|12300,12305
follow|12306,12312
-|12312,12313
up|12313,12315
on|12316,12318
<EOL>|12319,12320
_|12320,12321
_|12321,12322
_|12322,12323
.|12323,12324
A|12325,12326
PICC|12327,12331
line|12332,12336
was|12337,12340
placed|12341,12347
in|12348,12350
the|12351,12354
right|12355,12360
arm|12361,12364
<EOL>|12365,12366
_|12366,12367
_|12367,12368
_|12368,12369
with|12370,12374
tentative|12375,12384
plan|12385,12389
to|12390,12392
complete|12393,12401
a|12402,12403
two|12404,12407
-|12407,12408
week|12408,12412
course|12413,12419
of|12420,12422
IV|12423,12425
<EOL>|12426,12427
nafcillin|12427,12436
on|12437,12439
_|12440,12441
_|12441,12442
_|12442,12443
.|12443,12444
For|12445,12448
the|12449,12452
wound|12453,12458
,|12458,12459
podiatry|12460,12468
recommends|12469,12479
daily|12480,12485
<EOL>|12486,12487
dressing|12487,12495
changes|12496,12503
to|12504,12506
left|12507,12511
foot|12512,12516
surgical|12517,12525
site|12526,12530
:|12530,12531
Betadine|12532,12540
moistened|12541,12550
<EOL>|12551,12552
gauze|12552,12557
,|12557,12558
4x4|12559,12562
gauze|12563,12568
,|12568,12569
and|12570,12573
kerlix|12574,12580
.|12580,12581
<EOL>|12581,12582
<EOL>|12582,12583
#|12583,12584
Cough|12584,12589
:|12589,12590
During|12591,12597
her|12598,12601
stay|12602,12606
the|12607,12610
patient|12611,12618
developed|12619,12628
cough|12629,12634
that|12635,12639
was|12640,12643
<EOL>|12644,12645
nonproductive|12645,12658
.|12658,12659
It|12660,12662
was|12663,12666
thought|12667,12674
to|12675,12677
be|12678,12680
due|12681,12684
to|12685,12687
atelectasis|12688,12699
after|12700,12705
<EOL>|12706,12707
surgery|12707,12714
,|12714,12715
especially|12716,12726
since|12727,12732
her|12733,12736
rales|12737,12742
on|12743,12745
exam|12746,12750
would|12751,12756
clear|12757,12762
with|12763,12767
<EOL>|12768,12769
coughing|12769,12777
.|12777,12778
A|12779,12780
repeat|12781,12787
chest|12788,12793
x-ray|12794,12799
was|12800,12803
negative|12804,12812
for|12813,12816
any|12817,12820
acute|12821,12826
<EOL>|12827,12828
cardiopulmonary|12828,12843
processes|12844,12853
and|12854,12857
on|12858,12860
comparison|12861,12871
to|12872,12874
previous|12875,12883
chest|12884,12889
<EOL>|12890,12891
x-ray|12891,12896
during|12897,12903
this|12904,12908
hospital|12909,12917
stay|12918,12922
there|12923,12928
were|12929,12933
no|12934,12936
changes|12937,12944
.|12944,12945
Will|12946,12950
<EOL>|12951,12952
restart|12952,12959
home|12960,12964
Lasix|12965,12970
at|12971,12973
discharge|12974,12983
.|12983,12984
<EOL>|12984,12985
<EOL>|12985,12986
#|12986,12987
Hypertension|12987,12999
:|12999,13000
Patient|13001,13008
's|13008,13010
antihypertensives|13011,13028
were|13029,13033
held|13034,13038
upon|13039,13043
<EOL>|13044,13045
admission|13045,13054
given|13055,13060
that|13061,13065
her|13066,13069
blood|13070,13075
pressures|13076,13085
were|13086,13090
low|13091,13094
with|13095,13099
systolic|13100,13108
<EOL>|13109,13110
blood|13110,13115
pressures|13116,13125
in|13126,13128
the|13129,13132
_|13133,13134
_|13134,13135
_|13135,13136
likely|13137,13143
due|13144,13147
to|13148,13150
sepsis|13151,13157
in|13158,13160
the|13161,13164
<EOL>|13165,13166
setting|13166,13173
of|13174,13176
her|13177,13180
osteomyelitis|13181,13194
from|13195,13199
her|13200,13203
diabetic|13204,13212
foot|13213,13217
ulcer|13218,13223
.|13223,13224
After|13225,13230
<EOL>|13231,13232
her|13232,13235
first|13236,13241
debridement|13242,13253
,|13253,13254
patient|13255,13262
's|13262,13264
blood|13265,13270
pressures|13271,13280
increase|13281,13289
to|13290,13292
<EOL>|13293,13294
160s|13294,13298
-|13298,13299
170s|13299,13303
so|13304,13306
we|13307,13309
restarted|13310,13319
her|13320,13323
losartan|13324,13332
and|13333,13336
furosemide|13337,13347
.|13347,13348
However|13349,13356
<EOL>|13357,13358
her|13358,13361
blood|13362,13367
pressure|13368,13376
dipped|13377,13383
back|13384,13388
down|13389,13393
again|13394,13399
to|13400,13402
the|13403,13406
_|13407,13408
_|13408,13409
_|13409,13410
systolic|13411,13419
<EOL>|13420,13421
and|13421,13424
her|13425,13428
creatinine|13429,13439
bumped|13440,13446
up|13447,13449
to|13450,13452
1.8|13453,13456
so|13457,13459
we|13460,13462
discontinued|13463,13475
her|13476,13479
<EOL>|13480,13481
losartan|13481,13489
and|13490,13493
furosemide|13494,13504
.|13504,13505
Her|13506,13509
metoprolol|13510,13520
was|13521,13524
continued|13525,13534
with|13535,13539
<EOL>|13540,13541
holding|13541,13548
parameters|13549,13559
,|13559,13560
and|13561,13564
it|13565,13567
was|13568,13571
held|13572,13576
when|13577,13581
her|13582,13585
systolic|13586,13594
blood|13595,13600
<EOL>|13601,13602
pressure|13602,13610
was|13611,13614
less|13615,13619
than|13620,13624
110|13625,13628
.|13628,13629
Her|13630,13633
_|13634,13635
_|13635,13636
_|13636,13637
resolved|13638,13646
,|13646,13647
and|13648,13651
she|13652,13655
became|13656,13662
<EOL>|13663,13664
hypertensive|13664,13676
again|13677,13682
,|13682,13683
so|13684,13686
we|13687,13689
restarted|13690,13699
her|13700,13703
losartan|13704,13712
while|13713,13718
in|13719,13721
the|13722,13725
<EOL>|13726,13727
hospital|13727,13735
and|13736,13739
instructed|13740,13750
the|13751,13754
patient|13755,13762
to|13763,13765
restart|13766,13773
her|13774,13777
Lasix|13778,13783
upon|13784,13788
<EOL>|13789,13790
discharge|13790,13799
from|13800,13804
the|13805,13808
hospital|13809,13817
.|13817,13818
<EOL>|13818,13819
<EOL>|13819,13820
#|13820,13821
Acute|13821,13826
Kidney|13827,13833
Injury|13834,13840
:|13840,13841
Her|13842,13845
baseline|13846,13854
creatinine|13855,13865
is|13866,13868
1.0|13869,13872
.|13872,13873
It|13874,13876
bumped|13877,13883
<EOL>|13884,13885
up|13885,13887
to|13888,13890
1.8|13891,13894
in|13895,13897
the|13898,13901
setting|13902,13909
of|13910,13912
sepsis|13913,13919
,|13919,13920
restarting|13921,13931
her|13932,13935
losartan|13936,13944
and|13945,13948
<EOL>|13949,13950
furosemide|13950,13960
,|13960,13961
and|13962,13965
hypotension|13966,13977
.|13977,13978
We|13979,13981
gave|13982,13986
her|13987,13990
IV|13991,13993
fluids|13994,14000
and|14001,14004
stopped|14005,14012
<EOL>|14013,14014
her|14014,14017
losartan|14018,14026
and|14027,14030
furosemide|14031,14041
.|14041,14042
Her|14043,14046
creatinine|14047,14057
continued|14058,14067
to|14068,14070
improve|14071,14078
<EOL>|14079,14080
with|14080,14084
these|14085,14090
measures|14091,14099
and|14100,14103
upon|14104,14108
discharge|14109,14118
it|14119,14121
was|14122,14125
1.1|14126,14129
-|14129,14130
1|14130,14131
.|14131,14132
2|14132,14133
,|14133,14134
which|14135,14140
is|14141,14143
<EOL>|14144,14145
around|14145,14151
her|14152,14155
baseline|14156,14164
.|14164,14165
<EOL>|14165,14166
<EOL>|14166,14167
CHRONIC|14167,14174
ISSUES|14175,14181
<EOL>|14181,14182
=|14182,14183
=|14183,14184
=|14184,14185
=|14185,14186
=|14186,14187
=|14187,14188
=|14188,14189
=|14189,14190
=|14190,14191
=|14191,14192
=|14192,14193
=|14193,14194
=|14194,14195
=|14195,14196
<EOL>|14196,14197
#|14197,14198
Diabetes|14198,14206
Mellitus|14207,14215
Type|14216,14220
2|14221,14222
:|14222,14223
Upon|14224,14228
admission|14229,14238
,|14238,14239
patient|14240,14247
was|14248,14251
started|14252,14259
<EOL>|14260,14261
on|14261,14263
80|14264,14266
%|14266,14267
of|14268,14270
home|14271,14275
insulin|14276,14283
doses|14284,14289
.|14289,14290
Her|14291,14294
Lantus|14295,14301
inpatient|14302,14311
dose|14312,14316
was|14317,14320
32|14321,14323
<EOL>|14324,14325
units|14325,14330
,|14330,14331
and|14332,14335
her|14336,14339
Humalog|14340,14347
inpatient|14348,14357
dose|14358,14362
was|14363,14366
12|14367,14369
units|14370,14375
3|14376,14377
times|14378,14383
<EOL>|14384,14385
daily|14385,14390
.|14390,14391
Patient|14392,14399
's|14399,14401
blood|14402,14407
sugars|14408,14414
were|14415,14419
hard|14420,14424
to|14425,14427
control|14428,14435
while|14436,14441
she|14442,14445
was|14446,14449
<EOL>|14450,14451
inpatient|14451,14460
.|14460,14461
Working|14462,14469
with|14470,14474
the|14475,14478
_|14479,14480
_|14480,14481
_|14481,14482
diabetes|14483,14491
consult|14492,14499
team|14500,14504
we|14505,14507
<EOL>|14508,14509
adjusted|14509,14517
her|14518,14521
insulin|14522,14529
doses|14530,14535
as|14536,14538
needed|14539,14545
.|14545,14546
_|14547,14548
_|14548,14549
_|14549,14550
recommended|14551,14562
<EOL>|14563,14564
discharging|14564,14575
the|14576,14579
patient|14580,14587
on|14588,14590
48|14591,14593
units|14594,14599
of|14600,14602
Toujeo|14603,14609
and|14610,14613
18|14614,14616
units|14617,14622
of|14623,14625
<EOL>|14626,14627
Novolog|14627,14634
with|14635,14639
meals|14640,14645
as|14646,14648
well|14649,14653
as|14654,14656
resuming|14657,14665
her|14666,14669
Trajenta|14670,14678
and|14679,14682
<EOL>|14683,14684
Jardiance|14684,14693
.|14693,14694
<EOL>|14694,14695
<EOL>|14695,14696
#|14696,14697
CODE|14697,14701
STATUS|14702,14708
:|14708,14709
Full|14710,14714
(|14715,14716
presumed|14716,14724
)|14724,14725
<EOL>|14725,14726
#|14726,14727
CONTACT|14727,14734
:|14734,14735
_|14736,14737
_|14737,14738
_|14738,14739
(|14740,14741
grandson|14741,14749
's|14749,14751
girlfriend|14752,14762
)|14762,14763
_|14764,14765
_|14765,14766
_|14766,14767
<EOL>|14767,14768
<EOL>|14768,14769
TRANSITIONAL|14769,14781
ISSUES|14782,14788
<EOL>|14788,14789
=|14789,14790
=|14790,14791
=|14791,14792
=|14792,14793
=|14793,14794
=|14794,14795
=|14795,14796
=|14796,14797
=|14797,14798
=|14798,14799
=|14799,14800
=|14800,14801
=|14801,14802
=|14802,14803
=|14803,14804
=|14804,14805
=|14805,14806
=|14806,14807
=|14807,14808
<EOL>|14808,14809
[|14809,14810
]|14811,14812
Patient|14813,14820
is|14821,14823
on|14824,14826
oxycodone|14827,14836
5|14837,14838
mg|14839,14841
Q8H|14842,14845
for|14846,14849
her|14850,14853
foot|14854,14858
pain|14859,14863
from|14864,14868
the|14869,14872
<EOL>|14873,14874
surgery|14874,14881
.|14881,14882
She|14883,14886
was|14887,14890
given|14891,14896
enough|14897,14903
to|14904,14906
get|14907,14910
her|14911,14914
to|14915,14917
her|14918,14921
PCP|14922,14925
appointment|14926,14937
,|14937,14938
<EOL>|14939,14940
which|14940,14945
is|14946,14948
_|14949,14950
_|14950,14951
_|14951,14952
.|14952,14953
Please|14954,14960
re-assess|14961,14970
pain|14971,14975
management|14976,14986
.|14986,14987
<EOL>|14987,14988
<EOL>|14988,14989
[|14989,14990
]|14991,14992
Osteomyelitis|14993,15006
,|15006,15007
infected|15008,15016
diabetic|15017,15025
foot|15026,15030
ulcer|15031,15036
:|15036,15037
Surgical|15038,15046
margin|15047,15053
<EOL>|15054,15055
from|15055,15059
total|15060,15065
left|15066,15070
hallux|15071,15077
amputation|15078,15088
on|15089,15091
_|15092,15093
_|15093,15094
_|15094,15095
was|15096,15099
negative|15100,15108
for|15109,15112
<EOL>|15113,15114
osteomyelitis|15114,15127
.|15127,15128
Patient|15129,15136
to|15137,15139
complete|15140,15148
a|15149,15150
2|15151,15152
week|15153,15157
course|15158,15164
of|15165,15167
nafcillin|15168,15177
<EOL>|15178,15179
for|15179,15182
ongoing|15183,15190
soft|15191,15195
tissue|15196,15202
infection|15203,15212
and|15213,15216
will|15217,15221
follow|15222,15228
up|15229,15231
with|15232,15236
ID|15237,15239
<EOL>|15240,15241
prior|15241,15246
to|15247,15249
completion|15250,15260
of|15261,15263
antibiotics|15264,15275
to|15276,15278
ensure|15279,15285
resolution|15286,15296
.|15296,15297
Will|15298,15302
be|15303,15305
<EOL>|15306,15307
discharged|15307,15317
on|15318,15320
q4|15321,15323
hour|15324,15328
nafcillin|15329,15338
to|15339,15341
be|15342,15344
infused|15345,15352
via|15353,15356
a|15357,15358
pump|15359,15363
.|15363,15364
Once|15365,15369
<EOL>|15370,15371
finished|15371,15379
an|15380,15382
antibiotic|15383,15393
should|15394,15400
also|15401,15405
have|15406,15410
right|15411,15416
arm|15417,15420
PICC|15421,15425
line|15426,15430
<EOL>|15431,15432
removed|15432,15439
.|15439,15440
For|15441,15444
the|15445,15448
wound|15449,15454
,|15454,15455
podiatry|15456,15464
recommends|15465,15475
daily|15476,15481
dressing|15482,15490
<EOL>|15491,15492
changes|15492,15499
to|15500,15502
left|15503,15507
foot|15508,15512
surgical|15513,15521
site|15522,15526
:|15526,15527
Betadine|15528,15536
moistened|15537,15546
gauze|15547,15552
,|15552,15553
<EOL>|15554,15555
4x4|15555,15558
gauze|15559,15564
,|15564,15565
and|15566,15569
kerlix|15570,15576
<EOL>|15576,15577
<EOL>|15577,15578
[|15578,15579
]|15580,15581
Diabetes|15582,15590
mellitus|15591,15599
type|15600,15604
2|15605,15606
:|15606,15607
Patient|15608,15615
's|15615,15617
blood|15618,15623
sugars|15624,15630
were|15631,15635
very|15636,15640
<EOL>|15641,15642
labile|15642,15648
.|15648,15649
Given|15650,15655
that|15656,15660
she|15661,15664
came|15665,15669
in|15670,15672
with|15673,15677
a|15678,15679
diabetic|15680,15688
foot|15689,15693
ulcer|15694,15699
<EOL>|15700,15701
suggesting|15701,15711
that|15712,15716
her|15717,15720
blood|15721,15726
sugars|15727,15733
are|15734,15737
not|15738,15741
well|15742,15746
-|15746,15747
controlled|15747,15757
at|15758,15760
<EOL>|15761,15762
home|15762,15766
,|15766,15767
she|15768,15771
needs|15772,15777
close|15778,15783
follow|15784,15790
-|15790,15791
up|15791,15793
to|15794,15796
optimize|15797,15805
her|15806,15809
diabetic|15810,15818
<EOL>|15819,15820
medication|15820,15830
regimen|15831,15838
.|15838,15839
She|15840,15843
is|15844,15846
being|15847,15852
discharged|15853,15863
on|15864,15866
reduced|15867,15874
dose|15875,15879
<EOL>|15880,15881
Toujeo|15881,15887
and|15888,15891
regular|15892,15899
home|15900,15904
Novolog|15905,15912
along|15913,15918
with|15919,15923
her|15924,15927
usual|15928,15933
Trajenta|15934,15942
<EOL>|15943,15944
and|15944,15947
Jardiance|15948,15957
with|15958,15962
close|15963,15968
follow|15969,15975
-|15975,15976
up|15976,15978
with|15979,15983
_|15984,15985
_|15985,15986
_|15986,15987
provider|15988,15996
on|15997,15999
<EOL>|16000,16001
_|16001,16002
_|16002,16003
_|16003,16004
,|16004,16005
_|16006,16007
_|16007,16008
_|16008,16009
at|16010,16012
1|16013,16014
_|16015,16016
_|16016,16017
_|16017,16018
.|16018,16019
Please|16020,16026
reassess|16027,16035
patient|16036,16043
's|16043,16045
need|16046,16050
for|16051,16054
<EOL>|16055,16056
Jardiance|16056,16065
given|16066,16071
history|16072,16079
of|16080,16082
recurrent|16083,16092
AKIs|16093,16097
<EOL>|16097,16098
<EOL>|16098,16099
[|16099,16100
]|16101,16102
Cough|16103,16108
:|16108,16109
Patient|16110,16117
developed|16118,16127
non-productive|16128,16142
cough|16143,16148
while|16149,16154
in|16155,16157
<EOL>|16158,16159
hospital|16159,16167
but|16168,16171
afebrile|16172,16180
,|16180,16181
no|16182,16184
leukocytosis|16185,16197
,|16197,16198
CXR|16199,16202
no|16203,16205
signs|16206,16211
of|16212,16214
pleural|16215,16222
<EOL>|16223,16224
effusion|16224,16232
or|16233,16235
consolidation|16236,16249
.|16249,16250
Suspect|16251,16258
due|16259,16262
to|16263,16265
atelectasis|16266,16277
in|16278,16280
post-op|16281,16288
<EOL>|16289,16290
period|16290,16296
after|16297,16302
foot|16303,16307
surgery|16308,16315
.|16315,16316
Will|16317,16321
discharge|16322,16331
on|16332,16334
incentive|16335,16344
<EOL>|16345,16346
spirometer|16346,16356
and|16357,16360
restarting|16361,16371
home|16372,16376
Lasix|16377,16382
as|16383,16385
outpatient|16386,16396
.|16396,16397
If|16398,16400
not|16401,16404
<EOL>|16405,16406
improved|16406,16414
once|16415,16419
back|16420,16424
on|16425,16427
outpatient|16428,16438
Lasix|16439,16444
,|16444,16445
would|16446,16451
consider|16452,16460
further|16461,16468
<EOL>|16469,16470
workup|16470,16476
.|16476,16477
<EOL>|16477,16478
<EOL>|16478,16479
[|16479,16480
]|16481,16482
Hypertension|16483,16495
:|16495,16496
Patient|16497,16504
was|16505,16508
discharged|16509,16519
on|16520,16522
her|16523,16526
regular|16527,16534
home|16535,16539
<EOL>|16540,16541
medications|16541,16552
.|16552,16553
While|16554,16559
she|16560,16563
was|16564,16567
an|16568,16570
inpatient|16571,16580
,|16580,16581
she|16582,16585
became|16586,16592
hypotensive|16593,16604
<EOL>|16605,16606
when|16606,16610
we|16611,16613
restarted|16614,16623
her|16624,16627
on|16628,16630
all|16631,16634
of|16635,16637
her|16638,16641
antihypertensives|16642,16659
.|16659,16660
Please|16661,16667
<EOL>|16668,16669
follow|16669,16675
her|16676,16679
blood|16680,16685
pressure|16686,16694
to|16695,16697
ensure|16698,16704
that|16705,16709
she|16710,16713
is|16714,16716
on|16717,16719
the|16720,16723
right|16724,16729
<EOL>|16730,16731
regimen|16731,16738
.|16738,16739
If|16740,16742
too|16743,16746
low|16747,16750
,|16750,16751
might|16752,16757
consider|16758,16766
removing|16767,16775
furosemide|16776,16786
.|16786,16787
<EOL>|16787,16788
<EOL>|16788,16789
[|16789,16790
]|16791,16792
_|16793,16794
_|16794,16795
_|16795,16796
:|16796,16797
Discharge|16798,16807
creatinine|16808,16818
1.2|16819,16822
on|16823,16825
_|16826,16827
_|16827,16828
_|16828,16829
.|16829,16830
Suspect|16831,16838
patient|16839,16846
will|16847,16851
<EOL>|16852,16853
have|16853,16857
a|16858,16859
slight|16860,16866
bump|16867,16871
in|16872,16874
creatinine|16875,16885
after|16886,16891
restarting|16892,16902
losartan|16903,16911
on|16912,16914
<EOL>|16915,16916
_|16916,16917
_|16917,16918
_|16918,16919
.|16919,16920
Patient|16921,16928
had|16929,16932
weekly|16933,16939
labs|16940,16944
checked|16945,16952
with|16953,16957
IV|16958,16960
antibiotic|16961,16971
<EOL>|16972,16973
infusions|16973,16982
.|16982,16983
If|16984,16986
continues|16987,16996
to|16997,16999
rise|17000,17004
,|17004,17005
may|17006,17009
be|17010,17012
due|17013,17016
to|17017,17019
nafcillin|17020,17029
and|17030,17033
<EOL>|17034,17035
would|17035,17040
consider|17041,17049
switching|17050,17059
antibiotic|17060,17070
to|17071,17073
cefazolin|17074,17083
.|17083,17084
<EOL>|17084,17085
<EOL>|17085,17086
#|17086,17087
CODE|17087,17091
STATUS|17092,17098
:|17098,17099
Full|17100,17104
(|17105,17106
presumed|17106,17114
)|17114,17115
<EOL>|17115,17116
#|17116,17117
CONTACT|17117,17124
:|17124,17125
_|17126,17127
_|17127,17128
_|17128,17129
(|17130,17131
grandson|17131,17139
's|17139,17141
girlfriend|17142,17152
)|17152,17153
_|17154,17155
_|17155,17156
_|17156,17157
<EOL>|17157,17158
<EOL>|17158,17159
>|17159,17160
30|17160,17162
minutes|17163,17170
spent|17171,17176
on|17177,17179
complex|17180,17187
discharge|17188,17197
<EOL>|17198,17199
<EOL>|17200,17201
Medications|17201,17212
on|17213,17215
Admission|17216,17225
:|17225,17226
<EOL>|17226,17227
The|17227,17230
Preadmission|17231,17243
Medication|17244,17254
list|17255,17259
is|17260,17262
accurate|17263,17271
and|17272,17275
complete|17276,17284
.|17284,17285
<EOL>|17285,17286
1.|17286,17288
canagliflozin|17289,17302
100|17303,17306
mg|17307,17309
oral|17310,17314
DAILY|17315,17320
<EOL>|17321,17322
2.|17322,17324
Nitroglycerin|17325,17338
SL|17339,17341
0.4|17342,17345
mg|17346,17348
SL|17349,17351
Q5MIN|17352,17357
:|17357,17358
PRN|17358,17361
angina|17362,17368
<EOL>|17369,17370
3.|17370,17372
rOPINIRole|17373,17383
0.5|17384,17387
mg|17388,17390
PO|17391,17393
QHS|17394,17397
restless|17398,17406
leg|17407,17410
syndrome|17411,17419
<EOL>|17420,17421
4.|17421,17423
TraZODone|17424,17433
50|17434,17436
mg|17437,17439
PO|17440,17442
QHS|17443,17446
:|17446,17447
PRN|17447,17450
insomnia|17451,17459
<EOL>|17460,17461
5.|17461,17463
Pantoprazole|17464,17476
40|17477,17479
mg|17480,17482
PO|17483,17485
BID|17486,17489
<EOL>|17490,17491
6.|17491,17493
Gabapentin|17494,17504
400|17505,17508
mg|17509,17511
PO|17512,17514
QHS|17515,17518
:|17518,17519
PRN|17519,17522
Neuropathic|17523,17534
pain|17535,17539
<EOL>|17540,17541
7.|17541,17543
Atorvastatin|17544,17556
80|17557,17559
mg|17560,17562
PO|17563,17565
QPM|17566,17569
<EOL>|17570,17571
8.|17571,17573
Fluticasone|17574,17585
Propionate|17586,17596
110mcg|17597,17603
2|17604,17605
PUFF|17606,17610
IH|17611,17613
BID|17614,17617
<EOL>|17618,17619
9.|17619,17621
linaGLIPtin|17622,17633
5|17634,17635
mg|17636,17638
oral|17639,17643
DAILY|17644,17649
<EOL>|17650,17651
10.|17651,17654
Losartan|17655,17663
Potassium|17664,17673
25|17674,17676
mg|17677,17679
PO|17680,17682
DAILY|17683,17688
<EOL>|17689,17690
11.|17690,17693
OxyCODONE|17694,17703
-|17703,17704
-|17704,17705
Acetaminophen|17705,17718
(|17719,17720
5mg|17720,17723
-|17723,17724
325mg|17724,17729
)|17729,17730
1|17731,17732
TAB|17733,17736
PO|17737,17739
TID|17740,17743
:|17743,17744
PRN|17744,17747
Pain|17748,17752
-|17753,17754
<EOL>|17755,17756
Severe|17756,17762
<EOL>|17763,17764
12.|17764,17767
Lidocaine|17768,17777
5|17778,17779
%|17779,17780
Patch|17781,17786
1|17787,17788
PTCH|17789,17793
TD|17794,17796
QPM|17797,17800
<EOL>|17801,17802
13.|17802,17805
Furosemide|17806,17816
20|17817,17819
mg|17820,17822
PO|17823,17825
DAILY|17826,17831
<EOL>|17832,17833
14.|17833,17836
Metoprolol|17837,17847
Succinate|17848,17857
XL|17858,17860
150|17861,17864
mg|17865,17867
PO|17868,17870
DAILY|17871,17876
<EOL>|17877,17878
15.|17878,17881
albuterol|17882,17891
sulfate|17892,17899
90|17900,17902
mcg|17903,17906
/|17906,17907
actuation|17907,17916
inhalation|17917,17927
Q4H|17928,17931
:|17931,17932
PRN|17932,17935
<EOL>|17936,17937
16|17937,17939
.|17939,17940
Aspirin|17941,17948
EC|17949,17951
325|17952,17955
mg|17956,17958
PO|17959,17961
DAILY|17962,17967
<EOL>|17968,17969
17.|17969,17972
MetronidAZOLE|17973,17986
Topical|17987,17994
1|17995,17996
%|17997,17998
Gel|17999,18002
1|18003,18004
Appl|18005,18009
TP|18010,18012
DAILY|18013,18018
Rosacea|18019,18026
<EOL>|18027,18028
18.|18028,18031
nystatin|18032,18040
100,000|18041,18048
unit|18049,18053
/|18053,18054
gram|18054,18058
topical|18059,18066
DAILY|18067,18072
:|18072,18073
PRN|18073,18076
<EOL>|18077,18078
<EOL>|18078,18079
<EOL>|18080,18081
Discharge|18081,18090
Medications|18091,18102
:|18102,18103
<EOL>|18103,18104
1.|18104,18106
Acetaminophen|18108,18121
1000|18122,18126
mg|18127,18129
PO|18130,18132
Q8H|18133,18136
<EOL>|18137,18138
RX|18138,18140
*|18141,18142
acetaminophen|18142,18155
500|18156,18159
mg|18160,18162
2|18163,18164
tablet|18165,18171
(|18171,18172
s|18172,18173
)|18173,18174
by|18175,18177
mouth|18178,18183
Every|18184,18189
8|18190,18191
hours|18192,18197
for|18198,18201
<EOL>|18202,18203
foot|18203,18207
pain|18208,18212
Disp|18213,18217
#|18218,18219
*|18219,18220
60|18220,18222
Tablet|18223,18229
Refills|18230,18237
:|18237,18238
*|18238,18239
0|18239,18240
<EOL>|18241,18242
2.|18242,18244
Bisacodyl|18246,18255
10|18256,18258
mg|18259,18261
PO|18262,18264
DAILY|18265,18270
:|18270,18271
PRN|18271,18274
Constipation|18275,18287
-|18288,18289
Second|18290,18296
Line|18297,18301
<EOL>|18302,18303
RX|18303,18305
*|18306,18307
bisacodyl|18307,18316
5|18317,18318
mg|18319,18321
2|18322,18323
tablet|18324,18330
(|18330,18331
s|18331,18332
)|18332,18333
by|18334,18336
mouth|18337,18342
Once|18343,18347
a|18348,18349
day|18350,18353
as|18354,18356
needed|18357,18363
for|18364,18367
<EOL>|18368,18369
constipation|18369,18381
Disp|18382,18386
#|18387,18388
*|18388,18389
60|18389,18391
Tablet|18392,18398
Refills|18399,18406
:|18406,18407
*|18407,18408
0|18408,18409
<EOL>|18410,18411
3.|18411,18413
Docusate|18415,18423
Sodium|18424,18430
100|18431,18434
mg|18435,18437
PO|18438,18440
BID|18441,18444
<EOL>|18445,18446
RX|18446,18448
*|18449,18450
docusate|18450,18458
sodium|18459,18465
100|18466,18469
mg|18470,18472
1|18473,18474
capsule|18475,18482
(|18482,18483
s|18483,18484
)|18484,18485
by|18486,18488
mouth|18489,18494
Twice|18495,18500
a|18501,18502
day|18503,18506
<EOL>|18507,18508
Disp|18508,18512
#|18513,18514
*|18514,18515
30|18515,18517
Capsule|18518,18525
Refills|18526,18533
:|18533,18534
*|18534,18535
0|18535,18536
<EOL>|18537,18538
4.|18538,18540
Nafcillin|18542,18551
2|18552,18553
g|18554,18555
IV|18556,18558
Q4H|18559,18562
<EOL>|18563,18564
RX|18564,18566
*|18567,18568
nafcillin|18568,18577
in|18578,18580
dextrose|18581,18589
iso|18590,18593
-|18593,18594
osm|18594,18597
2|18598,18599
gram|18600,18604
/|18604,18605
100|18605,18608
mL|18609,18611
2|18612,18613
g|18614,18615
IV|18616,18618
Every|18619,18624
<EOL>|18625,18626
four|18626,18630
hours|18631,18636
Disp|18637,18641
#|18642,18643
*|18643,18644
84|18644,18646
Intravenous|18647,18658
Bag|18659,18662
Refills|18663,18670
:|18670,18671
*|18671,18672
0|18672,18673
<EOL>|18674,18675
5.|18675,18677
OxyCODONE|18679,18688
(|18689,18690
Immediate|18690,18699
Release|18700,18707
)|18707,18708
5|18709,18710
mg|18711,18713
PO|18714,18716
Q8H|18717,18720
:|18720,18721
PRN|18721,18724
Pain|18725,18729
-|18730,18731
<EOL>|18732,18733
Moderate|18733,18741
<EOL>|18742,18743
RX|18743,18745
*|18746,18747
oxycodone|18747,18756
5|18757,18758
mg|18759,18761
1|18762,18763
capsule|18764,18771
(|18771,18772
s|18772,18773
)|18773,18774
by|18775,18777
mouth|18778,18783
Once|18784,18788
every|18789,18794
8|18795,18796
hours|18797,18802
as|18803,18805
<EOL>|18806,18807
needed|18807,18813
for|18814,18817
severe|18818,18824
foot|18825,18829
pain|18830,18834
.|18834,18835
Disp|18836,18840
#|18841,18842
*|18842,18843
15|18843,18845
Capsule|18846,18853
Refills|18854,18861
:|18861,18862
*|18862,18863
0|18863,18864
<EOL>|18865,18866
6.|18866,18868
Senna|18870,18875
8.6|18876,18879
mg|18880,18882
PO|18883,18885
BID|18886,18889
:|18889,18890
PRN|18890,18893
Constipation|18894,18906
-|18907,18908
First|18909,18914
Line|18915,18919
<EOL>|18920,18921
RX|18921,18923
*|18924,18925
sennosides|18925,18935
[|18936,18937
senna|18937,18942
]|18942,18943
8.6|18944,18947
mg|18948,18950
1|18951,18952
tablet|18953,18959
by|18960,18962
mouth|18963,18968
Twice|18969,18974
a|18975,18976
day|18977,18980
as|18981,18983
<EOL>|18984,18985
needed|18985,18991
for|18992,18995
constipation|18996,19008
Disp|19009,19013
#|19014,19015
*|19015,19016
30|19016,19018
Tablet|19019,19025
Refills|19026,19033
:|19033,19034
*|19034,19035
0|19035,19036
<EOL>|19037,19038
7.|19038,19040
Novolog|19042,19049
18|19050,19052
Units|19053,19058
Breakfast|19059,19068
<EOL>|19068,19069
Novolog|19069,19076
18|19077,19079
Units|19080,19085
Lunch|19086,19091
<EOL>|19091,19092
Novolog|19092,19099
18|19100,19102
Units|19103,19108
Dinner|19109,19115
<EOL>|19116,19117
8.|19117,19119
albuterol|19121,19130
sulfate|19131,19138
90|19139,19141
mcg|19142,19145
/|19145,19146
actuation|19146,19155
inhalation|19156,19166
Q4H|19167,19170
:|19170,19171
PRN|19171,19174
<EOL>|19176,19177
9.|19177,19179
Aspirin|19181,19188
EC|19189,19191
325|19192,19195
mg|19196,19198
PO|19199,19201
DAILY|19202,19207
<EOL>|19209,19210
10.|19210,19213
Atorvastatin|19215,19227
80|19228,19230
mg|19231,19233
PO|19234,19236
QPM|19237,19240
<EOL>|19242,19243
11.|19243,19246
canagliflozin|19248,19261
100|19262,19265
mg|19266,19268
oral|19269,19273
DAILY|19274,19279
<EOL>|19281,19282
12.|19282,19285
Fluticasone|19287,19298
Propionate|19299,19309
110mcg|19310,19316
2|19317,19318
PUFF|19319,19323
IH|19324,19326
BID|19327,19330
<EOL>|19332,19333
13.|19333,19336
Furosemide|19338,19348
20|19349,19351
mg|19352,19354
PO|19355,19357
DAILY|19358,19363
<EOL>|19365,19366
14.|19366,19369
Gabapentin|19371,19381
400|19382,19385
mg|19386,19388
PO|19389,19391
QHS|19392,19395
:|19395,19396
PRN|19396,19399
Neuropathic|19400,19411
pain|19412,19416
<EOL>|19418,19419
15|19419,19421
.|19421,19422
Lidocaine|19424,19433
5|19434,19435
%|19435,19436
Patch|19437,19442
1|19443,19444
PTCH|19445,19449
TD|19450,19452
QPM|19453,19456
<EOL>|19458,19459
16.|19459,19462
linaGLIPtin|19464,19475
5|19476,19477
mg|19478,19480
oral|19481,19485
DAILY|19486,19491
<EOL>|19493,19494
17.|19494,19497
Losartan|19499,19507
Potassium|19508,19517
25|19518,19520
mg|19521,19523
PO|19524,19526
DAILY|19527,19532
<EOL>|19534,19535
18.|19535,19538
Metoprolol|19540,19550
Succinate|19551,19560
XL|19561,19563
150|19564,19567
mg|19568,19570
PO|19571,19573
DAILY|19574,19579
<EOL>|19581,19582
19|19582,19584
.|19584,19585
MetronidAZOLE|19587,19600
Topical|19601,19608
1|19609,19610
%|19611,19612
Gel|19613,19616
1|19617,19618
Appl|19619,19623
TP|19624,19626
DAILY|19627,19632
Rosacea|19633,19640
<EOL>|19642,19643
20|19643,19645
.|19645,19646
Nitroglycerin|19648,19661
SL|19662,19664
0.4|19665,19668
mg|19669,19671
SL|19672,19674
Q5MIN|19675,19680
:|19680,19681
PRN|19681,19684
angina|19685,19691
<EOL>|19693,19694
21.|19694,19697
nystatin|19699,19707
100,000|19708,19715
unit|19716,19720
/|19720,19721
gram|19721,19725
topical|19726,19733
DAILY|19734,19739
:|19739,19740
PRN|19740,19743
<EOL>|19745,19746
22.|19746,19749
OxyCODONE|19751,19760
-|19760,19761
-|19761,19762
Acetaminophen|19762,19775
(|19776,19777
5mg|19777,19780
-|19780,19781
325mg|19781,19786
)|19786,19787
1|19788,19789
TAB|19790,19793
PO|19794,19796
TID|19797,19800
:|19800,19801
PRN|19801,19804
Pain|19805,19809
<EOL>|19810,19811
-|19811,19812
Severe|19813,19819
<EOL>|19821,19822
23|19822,19824
.|19824,19825
Pantoprazole|19827,19839
40|19840,19842
mg|19843,19845
PO|19846,19848
BID|19849,19852
<EOL>|19854,19855
24.|19855,19858
rOPINIRole|19860,19870
0.5|19871,19874
mg|19875,19877
PO|19878,19880
QHS|19881,19884
restless|19885,19893
leg|19894,19897
syndrome|19898,19906
<EOL>|19908,19909
25.|19909,19912
_|19914,19915
_|19915,19916
_|19916,19917
SoloStar|19918,19926
U-300|19927,19932
Insulin|19933,19940
(|19941,19942
insulin|19942,19949
glargine|19950,19958
)|19958,19959
300|19960,19963
<EOL>|19964,19965
unit|19965,19969
/|19969,19970
mL|19970,19972
(|19973,19974
1.5|19974,19977
mL|19978,19980
)|19980,19981
subcutaneous|19982,19994
QHS|19995,19998
<EOL>|19999,20000
Inject|20000,20006
48U|20007,20010
QHS|20011,20014
<EOL>|20016,20017
26|20017,20019
.|20019,20020
TraZODone|20022,20031
50|20032,20034
mg|20035,20037
PO|20038,20040
QHS|20041,20044
:|20044,20045
PRN|20045,20048
insomnia|20049,20057
<EOL>|20059,20060
27.|20060,20063
Outpatient|20063,20073
Lab|20074,20077
Work|20078,20082
<EOL>|20082,20083
ICD|20083,20086
-|20086,20087
10|20087,20089
:|20089,20090
E11|20091,20094
.|20094,20095
621|20095,20098
<EOL>|20099,20100
DATE|20100,20104
:|20104,20105
weekly|20106,20112
:|20112,20113
draw|20114,20118
on|20119,20121
_|20122,20123
_|20123,20124
_|20124,20125
and|20126,20129
_|20130,20131
_|20131,20132
_|20132,20133
<EOL>|20133,20134
LAB|20134,20137
TEST|20138,20142
:|20142,20143
CBC|20144,20147
with|20148,20152
differential|20153,20165
,|20165,20166
BUN|20167,20170
,|20170,20171
Cr|20172,20174
,|20174,20175
AST|20176,20179
,|20179,20180
ALT|20181,20184
,|20184,20185
Total|20186,20191
<EOL>|20191,20192
Bili|20192,20196
,|20196,20197
ALK|20198,20201
PHOS|20202,20206
,|20206,20207
ESR|20208,20211
,|20211,20212
CRP|20213,20216
<EOL>|20216,20217
PLEASE|20217,20223
FAX|20224,20227
RESULTS|20228,20235
TO|20236,20238
:|20238,20239
ATTN|20240,20244
:|20244,20245
_|20246,20247
_|20247,20248
_|20248,20249
CLINIC|20250,20256
-|20257,20258
FAX|20259,20262
:|20262,20263
<EOL>|20264,20265
_|20265,20266
_|20266,20267
_|20267,20268
<EOL>|20268,20269
28.|20269,20272
Rolling|20272,20279
Walker|20280,20286
<EOL>|20286,20287
EQUIPMENT|20287,20296
:|20296,20297
Rolling|20298,20305
Walker|20306,20312
<EOL>|20312,20313
DIAGNOSIS|20313,20322
:|20322,20323
Left|20324,20328
hallux|20329,20335
amputation|20336,20346
<EOL>|20346,20347
ICD|20347,20350
-|20350,20351
10|20351,20353
:|20353,20354
_|20355,20356
_|20356,20357
_|20357,20358
<EOL>|20359,20360
PX|20360,20362
:|20362,20363
Good|20364,20368
<EOL>|20368,20369
_|20369,20370
_|20370,20371
_|20371,20372
:|20372,20373
13|20374,20376
months|20377,20383
<EOL>|20383,20384
<EOL>|20384,20385
<EOL>|20386,20387
Discharge|20387,20396
Disposition|20397,20408
:|20408,20409
<EOL>|20409,20410
Home|20410,20414
With|20415,20419
Service|20420,20427
<EOL>|20427,20428
<EOL>|20429,20430
Facility|20430,20438
:|20438,20439
<EOL>|20439,20440
_|20440,20441
_|20441,20442
_|20442,20443
<EOL>|20443,20444
<EOL>|20445,20446
Discharge|20446,20455
Diagnosis|20456,20465
:|20465,20466
<EOL>|20466,20467
=|20485,20486
=|20486,20487
=|20487,20488
=|20488,20489
=|20489,20490
=|20490,20491
=|20491,20492
=|20492,20493
=|20493,20494
=|20494,20495
=|20495,20496
=|20496,20497
=|20497,20498
=|20498,20499
=|20499,20500
=|20500,20501
=|20501,20502
<EOL>|20502,20503
Osteomyelitis|20503,20516
of|20517,20519
left|20520,20524
hallux|20525,20531
<EOL>|20531,20532
<EOL>|20532,20533
SECONDARY|20533,20542
DIAGNOSES|20543,20552
<EOL>|20552,20553
=|20553,20554
=|20554,20555
=|20555,20556
=|20556,20557
=|20557,20558
=|20558,20559
=|20559,20560
=|20560,20561
=|20561,20562
=|20562,20563
=|20563,20564
=|20564,20565
=|20565,20566
=|20566,20567
=|20567,20568
=|20568,20569
=|20569,20570
=|20570,20571
=|20571,20572
<EOL>|20572,20573
Hypertension|20573,20585
<EOL>|20585,20586
Type|20586,20590
2|20591,20592
Diabetes|20593,20601
Mellitus|20602,20610
<EOL>|20610,20611
<EOL>|20611,20612
<EOL>|20613,20614
Mental|20635,20641
Status|20642,20648
:|20648,20649
Clear|20650,20655
and|20656,20659
coherent|20660,20668
.|20668,20669
<EOL>|20669,20670
Level|20670,20675
of|20676,20678
Consciousness|20679,20692
:|20692,20693
Alert|20694,20699
and|20700,20703
interactive|20704,20715
.|20715,20716
<EOL>|20716,20717
Activity|20717,20725
Status|20726,20732
:|20732,20733
Ambulatory|20734,20744
-|20745,20746
Independent|20747,20758
.|20758,20759
<EOL>|20759,20760
<EOL>|20760,20761
<EOL>|20762,20763
Dear|20787,20791
Ms.|20792,20795
_|20796,20797
_|20797,20798
_|20798,20799
,|20799,20800
<EOL>|20800,20801
<EOL>|20801,20802
It|20802,20804
was|20805,20808
a|20809,20810
pleasure|20811,20819
taking|20820,20826
care|20827,20831
of|20832,20834
you|20835,20838
.|20838,20839
<EOL>|20839,20840
<EOL>|20840,20841
WHY|20841,20844
WAS|20845,20848
I|20849,20850
ADMITTED|20851,20859
TO|20860,20862
THE|20863,20866
HOSPITAL|20867,20875
?|20875,20876
<EOL>|20876,20877
You|20877,20880
had|20881,20884
a|20885,20886
diabetic|20887,20895
foot|20896,20900
ulcer|20901,20906
on|20907,20909
your|20910,20914
left|20915,20919
toe|20920,20923
that|20924,20928
was|20929,20932
very|20933,20937
<EOL>|20938,20939
infected|20939,20947
and|20948,20951
had|20952,20955
caused|20956,20962
an|20963,20965
infection|20966,20975
in|20976,20978
your|20979,20983
bone|20984,20988
.|20988,20989
<EOL>|20989,20990
<EOL>|20990,20991
WHAT|20991,20995
WAS|20996,20999
DONE|21000,21004
WHILE|21005,21010
I|21011,21012
WAS|21013,21016
HERE|21017,21021
?|21021,21022
<EOL>|21022,21023
Your|21023,21027
big|21028,21031
left|21032,21036
toe|21037,21040
was|21041,21044
removed|21045,21052
because|21053,21060
you|21061,21064
had|21065,21068
a|21069,21070
bad|21071,21074
bone|21075,21079
<EOL>|21080,21081
infection|21081,21090
.|21090,21091
You|21092,21095
were|21096,21100
treated|21101,21108
with|21109,21113
antibiotics|21114,21125
to|21126,21128
fight|21129,21134
the|21135,21138
<EOL>|21139,21140
infection|21140,21149
and|21150,21153
will|21154,21158
need|21159,21163
to|21164,21166
go|21167,21169
home|21170,21174
on|21175,21177
IV|21178,21180
antibiotics|21181,21192
.|21192,21193
<EOL>|21193,21194
<EOL>|21194,21195
WHAT|21195,21199
DO|21200,21202
I|21203,21204
NEED|21205,21209
TO|21210,21212
DO|21213,21215
WHEN|21216,21220
I|21221,21222
LEAVE|21223,21228
?|21228,21229
<EOL>|21229,21230
Please|21230,21236
continue|21237,21245
to|21246,21248
take|21249,21253
your|21254,21258
medications|21259,21270
as|21271,21273
directed|21274,21282
.|21282,21283
You|21285,21288
will|21289,21293
<EOL>|21294,21295
go|21295,21297
home|21298,21302
with|21303,21307
an|21308,21310
antibiotic|21311,21321
infusion|21322,21330
pump|21331,21335
and|21336,21339
will|21340,21344
have|21345,21349
a|21350,21351
<EOL>|21352,21353
visiting|21353,21361
nurse|21362,21367
come|21368,21372
to|21373,21375
your|21376,21380
house|21381,21386
to|21387,21389
teach|21390,21395
you|21396,21399
how|21400,21403
to|21404,21406
use|21407,21410
it|21411,21413
.|21413,21414
<EOL>|21416,21417
You|21417,21420
will|21421,21425
need|21426,21430
to|21431,21433
administer|21434,21444
antibiotics|21445,21456
through|21457,21464
the|21465,21468
pump|21469,21473
every|21474,21479
4|21480,21481
<EOL>|21482,21483
hours|21483,21488
.|21488,21489
We|21491,21493
changed|21494,21501
your|21502,21506
diabetic|21507,21515
medication|21516,21526
regimen|21527,21534
,|21534,21535
so|21536,21538
please|21539,21545
<EOL>|21546,21547
follow|21547,21553
along|21554,21559
as|21560,21562
instructed|21563,21573
below|21574,21579
and|21580,21583
keep|21584,21588
close|21589,21594
track|21595,21600
of|21601,21603
your|21604,21608
<EOL>|21609,21610
sugars|21610,21616
at|21617,21619
home|21620,21624
.|21624,21625
Check|21626,21631
your|21632,21636
sugars|21637,21643
4|21644,21645
times|21646,21651
a|21652,21653
day|21654,21657
and|21658,21661
log|21662,21665
the|21666,21669
<EOL>|21670,21671
results|21671,21678
.|21678,21679
Bring|21680,21685
the|21686,21689
results|21690,21697
in|21698,21700
with|21701,21705
you|21706,21709
to|21710,21712
your|21713,21717
_|21718,21719
_|21719,21720
_|21720,21721
<EOL>|21722,21723
appointment|21723,21734
on|21735,21737
_|21738,21739
_|21739,21740
_|21740,21741
at|21742,21744
1|21745,21746
:|21746,21747
00|21747,21749
pm|21750,21752
so|21753,21755
that|21756,21760
they|21761,21765
can|21766,21769
<EOL>|21770,21771
adjust|21771,21777
your|21778,21782
medication|21783,21793
regimen|21794,21801
appropriately|21802,21815
.|21815,21816
Please|21817,21823
follow|21824,21830
-|21830,21831
up|21831,21833
<EOL>|21834,21835
with|21835,21839
Dr.|21840,21843
_|21844,21845
_|21845,21846
_|21846,21847
team|21848,21852
on|21853,21855
_|21856,21857
_|21857,21858
_|21858,21859
at|21860,21862
11|21863,21865
:|21865,21866
00|21866,21868
am|21869,21871
.|21871,21872
Please|21873,21879
<EOL>|21880,21881
follow|21881,21887
up|21888,21890
with|21891,21895
Dr.|21896,21899
_|21900,21901
_|21901,21902
_|21902,21903
your|21904,21908
antibiotic|21909,21919
regimen|21920,21927
on|21928,21930
<EOL>|21931,21932
_|21932,21933
_|21933,21934
_|21934,21935
at|21936,21938
10|21939,21941
:|21941,21942
30|21942,21944
am|21945,21947
.|21947,21948
Please|21949,21955
follow|21956,21962
-|21962,21963
up|21963,21965
with|21966,21970
Dr.|21971,21974
_|21975,21976
_|21976,21977
_|21977,21978
<EOL>|21979,21980
in|21980,21982
_|21983,21984
_|21984,21985
_|21985,21986
_|21987,21988
_|21988,21989
_|21989,21990
on|21991,21993
_|21994,21995
_|21995,21996
_|21996,21997
at|21998,22000
1|22001,22002
:|22002,22003
00|22003,22005
pm|22006,22008
.|22008,22009
<EOL>|22009,22010
<EOL>|22010,22011
Be|22011,22013
well|22014,22018
,|22018,22019
<EOL>|22019,22020
<EOL>|22020,22021
Your|22021,22025
_|22026,22027
_|22027,22028
_|22028,22029
Care|22030,22034
Team|22035,22039
<EOL>|22039,22040
<EOL>|22041,22042
Followup|22042,22050
Instructions|22051,22063
:|22063,22064
<EOL>|22064,22065
_|22065,22066
_|22066,22067
_|22067,22068
<EOL>|22068,22069

