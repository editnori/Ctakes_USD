 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|29,33
No|34,36
:|36,37
_|40,41
_|41,42
_|42,43
<EOL>|43,44
<EOL>|45,46
Admission|46,55
Date|56,60
:|60,61
_|63,64
_|64,65
_|65,66
Discharge|80,89
Date|90,94
:|94,95
_|98,99
_|99,100
_|100,101
<EOL>|101,102
<EOL>|103,104
Date|104,108
of|109,111
Birth|112,117
:|117,118
_|120,121
_|121,122
_|122,123
Sex|136,139
:|139,140
F|143,144
<EOL>|144,145
<EOL>|146,147
Service|147,154
:|154,155
MEDICINE|156,164
<EOL>|164,165
<EOL>|166,167
omeprazole|179,189
<EOL>|189,190
<EOL>|191,192
Attending|192,201
:|201,202
_|203,204
_|204,205
_|205,206
.|206,207
<EOL>|207,208
<EOL>|209,210
dysphagia|227,236
<EOL>|237,238
<EOL>|239,240
Major|240,245
Surgical|246,254
or|255,257
Invasive|258,266
Procedure|267,276
:|276,277
<EOL>|277,278
Upper|278,283
endoscopy|284,293
_|294,295
_|295,296
_|296,297
<EOL>|297,298
<EOL>|298,299
<EOL>|300,301
_|330,331
_|331,332
_|332,333
w|334,335
/|335,336
anxiety|337,344
and|345,348
several|349,356
years|357,362
of|363,365
dysphagia|366,375
who|376,379
p|380,381
/|381,382
w|382,383
worsened|384,392
<EOL>|393,394
foreign|394,401
body|402,406
sensation|407,416
.|416,417
<EOL>|418,419
<EOL>|419,420
She|420,423
describes|424,433
feeling|434,441
as|442,444
though|445,451
food|452,456
gets|457,461
stuck|462,467
in|468,470
her|471,474
neck|475,479
when|480,484
<EOL>|485,486
she|486,489
eats|490,494
.|494,495
She|496,499
put|500,503
herself|504,511
on|512,514
a|515,516
pureed|517,523
diet|524,528
to|529,531
address|532,539
this|540,544
over|545,549
<EOL>|550,551
the|551,554
last|555,559
10|560,562
days|563,567
.|567,568
When|569,573
she|574,577
has|578,581
food|582,586
stuck|587,592
in|593,595
the|596,599
throat|600,606
,|606,607
she|608,611
<EOL>|612,613
almost|613,619
feels|620,625
as|626,628
though|629,635
she|636,639
can|640,643
not|643,646
breath|647,653
,|653,654
but|655,658
she|659,662
denies|663,669
trouble|670,677
<EOL>|678,679
breathing|679,688
at|689,691
any|692,695
other|696,701
time|702,706
.|706,707
She|708,711
does|712,716
not|717,720
have|721,725
any|726,729
history|730,737
of|738,740
<EOL>|741,742
food|742,746
allergies|747,756
or|757,759
skin|760,764
rashes|765,771
.|771,772
<EOL>|773,774
<EOL>|775,776
In|776,778
the|779,782
ED|783,785
,|785,786
initial|787,794
vitals|795,801
:|801,802
97.6|804,808
81|810,812
148|814,817
/|817,818
83|818,820
16|822,824
100|826,829
%|829,830
RA|831,833
<EOL>|834,835
Imaging|835,842
showed|843,849
:|849,850
CXR|851,854
showed|855,861
a|862,863
prominent|864,873
esophagus|874,883
<EOL>|883,884
Consults|884,892
:|892,893
GI|894,896
was|897,900
consulted|901,910
.|910,911
<EOL>|911,912
<EOL>|912,913
Pt|913,915
underwent|916,925
EGD|926,929
which|930,935
showed|936,942
a|943,944
normal|945,951
appearing|952,961
esophagus|962,971
.|971,972
<EOL>|973,974
Biopsies|974,982
were|983,987
taken|988,993
.|993,994
<EOL>|994,995
<EOL>|995,996
Currently|996,1005
,|1005,1006
she|1007,1010
endorses|1011,1019
anxiety|1020,1027
about|1028,1033
eating|1034,1040
.|1040,1041
She|1042,1045
would|1046,1051
like|1052,1056
to|1057,1059
<EOL>|1060,1061
try|1061,1064
eating|1065,1071
here|1072,1076
prior|1077,1082
to|1083,1085
leaving|1086,1093
the|1094,1097
hospital|1098,1106
.|1106,1107
<EOL>|1108,1109
<EOL>|1109,1110
<EOL>|1111,1112
-|1134,1135
GERD|1136,1140
<EOL>|1142,1143
-|1144,1145
Hypercholesterolemia|1146,1166
<EOL>|1168,1169
-|1170,1171
Kidney|1172,1178
stones|1179,1185
<EOL>|1187,1188
-|1189,1190
Mitral|1191,1197
valve|1198,1203
prolapse|1204,1212
<EOL>|1214,1215
-|1216,1217
Uterine|1218,1225
fibroids|1226,1234
<EOL>|1236,1237
-|1238,1239
Osteoporosis|1240,1252
<EOL>|1254,1255
-|1256,1257
Migraine|1258,1266
headaches|1267,1276
<EOL>|1277,1278
<EOL>|1279,1280
:|1294,1295
<EOL>|1295,1296
_|1296,1297
_|1297,1298
_|1298,1299
<EOL>|1299,1300
:|1314,1315
<EOL>|1315,1316
+|1316,1317
HTN|1318,1321
-|1322,1323
father|1324,1330
<EOL>|1332,1333
+|1333,1334
Dementia|1335,1343
-|1344,1345
father|1346,1352
<EOL>|1354,1355
<EOL>|1356,1357
<EOL>|1358,1359
=|1374,1375
=|1375,1376
=|1376,1377
=|1377,1378
=|1378,1379
=|1379,1380
=|1380,1381
=|1381,1382
=|1382,1383
=|1383,1384
=|1384,1385
=|1385,1386
=|1386,1387
=|1387,1388
=|1388,1389
=|1389,1390
=|1390,1391
<EOL>|1391,1392
ADMISSION|1392,1401
/|1401,1402
DISCHARGE|1402,1411
EXAM|1412,1416
<EOL>|1416,1417
=|1417,1418
=|1418,1419
=|1419,1420
=|1420,1421
=|1421,1422
=|1422,1423
=|1423,1424
=|1424,1425
=|1425,1426
=|1426,1427
=|1427,1428
=|1428,1429
=|1429,1430
=|1430,1431
=|1431,1432
=|1432,1433
=|1433,1434
<EOL>|1434,1435
VS|1435,1437
:|1437,1438
97.9|1440,1444
PO|1446,1448
109|1449,1452
/|1453,1454
71|1455,1457
70|1458,1460
16|1461,1463
97|1464,1466
ra|1467,1469
<EOL>|1470,1471
GEN|1471,1474
:|1474,1475
Thin|1476,1480
anxious|1481,1488
woman|1489,1494
,|1494,1495
lying|1496,1501
in|1502,1504
bed|1505,1508
,|1508,1509
no|1510,1512
acute|1513,1518
distress|1519,1527
<EOL>|1529,1530
HEENT|1530,1535
:|1535,1536
Moist|1537,1542
MM|1543,1545
,|1545,1546
anicteric|1547,1556
sclerae|1557,1564
,|1564,1565
NCAT|1566,1570
,|1570,1571
PERRL|1572,1577
,|1577,1578
EOMI|1579,1583
<EOL>|1585,1586
NECK|1586,1590
:|1590,1591
Supple|1592,1598
without|1599,1606
LAD|1607,1610
,|1610,1611
no|1612,1614
JVD|1615,1618
<EOL>|1620,1621
PULM|1621,1625
:|1625,1626
CTABL|1627,1632
no|1633,1635
w|1636,1637
/|1637,1638
c|1638,1639
/|1639,1640
r|1640,1641
<EOL>|1641,1642
COR|1642,1645
:|1645,1646
RRR|1647,1650
(|1651,1652
+|1652,1653
)|1653,1654
S1|1654,1656
/|1656,1657
S2|1657,1659
no|1660,1662
m|1663,1664
/|1664,1665
r|1665,1666
/|1666,1667
g|1667,1668
<EOL>|1670,1671
ABD|1671,1674
:|1674,1675
Soft|1676,1680
,|1680,1681
non-tender|1682,1692
,|1692,1693
non-distended|1694,1707
,|1707,1708
+|1709,1710
BS|1710,1712
,|1712,1713
no|1714,1716
HSM|1717,1720
<EOL>|1722,1723
EXTREM|1723,1729
:|1729,1730
Warm|1731,1735
,|1735,1736
well|1737,1741
-|1741,1742
perfused|1742,1750
,|1750,1751
no|1752,1754
_|1755,1756
_|1756,1757
_|1757,1758
edema|1759,1764
<EOL>|1766,1767
NEURO|1767,1772
:|1772,1773
CN|1774,1776
II|1777,1779
-|1779,1780
XII|1780,1783
grossly|1784,1791
intact|1792,1798
,|1798,1799
motor|1800,1805
function|1806,1814
grossly|1815,1822
normal|1823,1829
,|1829,1830
<EOL>|1831,1832
sensation|1832,1841
grossly|1842,1849
intact|1850,1856
<EOL>|1858,1859
<EOL>|1860,1861
Pertinent|1861,1870
Results|1871,1878
:|1878,1879
<EOL>|1879,1880
=|1880,1881
=|1881,1882
=|1882,1883
=|1883,1884
=|1884,1885
=|1885,1886
=|1886,1887
=|1887,1888
=|1888,1889
=|1889,1890
=|1890,1891
=|1891,1892
=|1892,1893
<EOL>|1893,1894
ADMISSION|1894,1903
LABS|1904,1908
<EOL>|1908,1909
=|1909,1910
=|1910,1911
=|1911,1912
=|1912,1913
=|1913,1914
=|1914,1915
=|1915,1916
=|1916,1917
=|1917,1918
=|1918,1919
=|1919,1920
=|1920,1921
=|1921,1922
<EOL>|1922,1923
<EOL>|1923,1924
_|1924,1925
_|1925,1926
_|1926,1927
08|1928,1930
:|1930,1931
27AM|1931,1935
BLOOD|1936,1941
WBC|1942,1945
-|1945,1946
5.0|1946,1949
RBC|1950,1953
-|1953,1954
4|1954,1955
.|1955,1956
82|1956,1958
Hgb|1959,1962
-|1962,1963
14.9|1963,1967
Hct|1968,1971
-|1971,1972
44.4|1972,1976
MCV|1977,1980
-|1980,1981
92|1981,1983
<EOL>|1984,1985
MCH|1985,1988
-|1988,1989
30.9|1989,1993
MCHC|1994,1998
-|1998,1999
33.6|1999,2003
RDW|2004,2007
-|2007,2008
12.1|2008,2012
RDWSD|2013,2018
-|2018,2019
41.3|2019,2023
Plt|2024,2027
_|2028,2029
_|2029,2030
_|2030,2031
<EOL>|2031,2032
_|2032,2033
_|2033,2034
_|2034,2035
08|2036,2038
:|2038,2039
27AM|2039,2043
BLOOD|2044,2049
_|2050,2051
_|2051,2052
_|2052,2053
PTT|2054,2057
-|2057,2058
28.6|2058,2062
_|2063,2064
_|2064,2065
_|2065,2066
<EOL>|2066,2067
_|2067,2068
_|2068,2069
_|2069,2070
08|2071,2073
:|2073,2074
27AM|2074,2078
BLOOD|2079,2084
Glucose|2085,2092
-|2092,2093
85|2093,2095
UreaN|2096,2101
-|2101,2102
8|2102,2103
Creat|2104,2109
-|2109,2110
0.9|2110,2113
Na|2114,2116
-|2116,2117
142|2117,2120
K|2121,2122
-|2122,2123
3.6|2123,2126
<EOL>|2127,2128
Cl|2128,2130
-|2130,2131
104|2131,2134
HCO3|2135,2139
-|2139,2140
22|2140,2142
AnGap|2143,2148
-|2148,2149
20|2149,2151
<EOL>|2151,2152
_|2152,2153
_|2153,2154
_|2154,2155
08|2156,2158
:|2158,2159
27AM|2159,2163
BLOOD|2164,2169
ALT|2170,2173
-|2173,2174
11|2174,2176
AST|2177,2180
-|2180,2181
16|2181,2183
LD|2184,2186
(|2186,2187
LDH|2187,2190
)|2190,2191
-|2191,2192
154|2192,2195
AlkPhos|2196,2203
-|2203,2204
63|2204,2206
<EOL>|2207,2208
TotBili|2208,2215
-|2215,2216
1.0|2216,2219
<EOL>|2219,2220
_|2220,2221
_|2221,2222
_|2222,2223
08|2224,2226
:|2226,2227
27AM|2227,2231
BLOOD|2232,2237
Albumin|2238,2245
-|2245,2246
4.8|2246,2249
<EOL>|2249,2250
=|2250,2251
=|2251,2252
=|2252,2253
=|2253,2254
=|2254,2255
=|2255,2256
=|2256,2257
=|2257,2258
=|2258,2259
=|2259,2260
=|2260,2261
=|2261,2262
=|2262,2263
<EOL>|2263,2264
IMAGING|2264,2271
<EOL>|2271,2272
=|2272,2273
=|2273,2274
=|2274,2275
=|2275,2276
=|2276,2277
=|2277,2278
=|2278,2279
=|2279,2280
=|2280,2281
=|2281,2282
=|2282,2283
=|2283,2284
=|2284,2285
<EOL>|2285,2286
<EOL>|2286,2287
CXR|2287,2290
_|2291,2292
_|2292,2293
_|2293,2294
:|2294,2295
<EOL>|2296,2297
Prominent|2314,2323
esophagus|2324,2333
on|2334,2336
lateral|2337,2344
view|2345,2349
,|2349,2350
without|2351,2358
air|2359,2362
-|2362,2363
fluid|2363,2368
level|2369,2374
.|2374,2375
<EOL>|2376,2377
Given|2377,2382
the|2383,2386
patient|2387,2394
's|2394,2396
history|2397,2404
and|2405,2408
radiographic|2409,2421
appearance|2422,2432
,|2432,2433
barium|2434,2440
<EOL>|2441,2442
swallow|2442,2449
is|2450,2452
indicated|2453,2462
either|2463,2469
now|2470,2473
or|2474,2476
electively|2477,2487
.|2487,2488
<EOL>|2489,2490
<EOL>|2492,2493
NECK|2493,2497
X-ray|2498,2503
_|2504,2505
_|2505,2506
_|2506,2507
:|2507,2508
<EOL>|2508,2509
Within|2526,2532
the|2533,2536
limitation|2537,2547
of|2548,2550
plain|2551,2556
radiography|2557,2568
,|2568,2569
no|2570,2572
evidence|2573,2581
of|2582,2584
<EOL>|2585,2586
prevertebral|2586,2598
soft|2599,2603
tissue|2604,2610
swelling|2611,2619
or|2620,2622
soft|2623,2627
tissue|2628,2634
mass|2635,2639
in|2640,2642
the|2643,2646
<EOL>|2647,2648
neck|2648,2652
.|2652,2653
<EOL>|2654,2655
<EOL>|2656,2657
<EOL>|2657,2658
EGD|2658,2661
:|2661,2662
_|2663,2664
_|2664,2665
_|2665,2666
<EOL>|2666,2667
Impression|2668,2678
:|2678,2679
Hiatal|2680,2686
hernia|2687,2693
<EOL>|2693,2694
Angioectasia|2694,2706
in|2707,2709
the|2710,2713
stomach|2714,2721
<EOL>|2721,2722
Angioectasia|2722,2734
in|2735,2737
the|2738,2741
duodenum|2742,2750
<EOL>|2750,2751
(|2752,2753
biopsy|2753,2759
,|2759,2760
biopsy|2761,2767
)|2767,2768
<EOL>|2768,2769
Otherwise|2769,2778
normal|2779,2785
EGD|2786,2789
to|2790,2792
third|2793,2798
part|2799,2803
of|2804,2806
the|2807,2810
duodenum|2811,2819
<EOL>|2820,2821
<EOL>|2821,2822
Recommendations|2822,2837
:|2837,2838
-|2839,2840
no|2841,2843
obvious|2844,2851
anatomic|2852,2860
cause|2861,2866
for|2867,2870
the|2871,2874
patient|2875,2882
's|2882,2884
<EOL>|2885,2886
symptoms|2886,2894
<EOL>|2894,2895
-|2895,2896
follow|2897,2903
-|2903,2904
up|2904,2906
biopsy|2907,2913
results|2914,2921
to|2922,2924
rule|2925,2929
out|2930,2933
eosinophilic|2934,2946
esophagitis|2947,2958
<EOL>|2958,2959
-|2959,2960
follow|2961,2967
-|2967,2968
up|2968,2970
with|2971,2975
Dr.|2976,2979
_|2980,2981
_|2981,2982
_|2982,2983
if|2984,2986
biopsies|2987,2995
show|2996,3000
eosinophilic|3001,3013
<EOL>|3014,3015
esophagitis|3015,3026
<EOL>|3027,3028
<EOL>|3028,3029
<EOL>|3030,3031
Ms.|3054,3057
_|3058,3059
_|3059,3060
_|3060,3061
is|3062,3064
a|3065,3066
_|3067,3068
_|3068,3069
_|3069,3070
with|3071,3075
history|3076,3083
of|3084,3086
GERD|3087,3091
who|3092,3095
presents|3096,3104
with|3105,3109
<EOL>|3110,3111
subacute|3111,3119
worsening|3120,3129
of|3130,3132
dysphagia|3133,3142
and|3143,3146
foreign|3147,3154
body|3155,3159
sensation|3160,3169
.|3169,3170
This|3171,3175
<EOL>|3176,3177
had|3177,3180
worsened|3181,3189
to|3190,3192
the|3193,3196
point|3197,3202
where|3203,3208
she|3209,3212
placed|3213,3219
herself|3220,3227
on|3228,3230
a|3231,3232
pureed|3233,3239
<EOL>|3240,3241
diet|3241,3245
for|3246,3249
the|3250,3253
last|3254,3258
10|3259,3261
days|3262,3266
.|3266,3267
She|3268,3271
underwent|3272,3281
CXR|3282,3285
which|3286,3291
showed|3292,3298
a|3299,3300
<EOL>|3301,3302
prominent|3302,3311
esophagus|3312,3321
but|3322,3325
was|3326,3329
otherwise|3330,3339
normal|3340,3346
.|3346,3347
She|3348,3351
was|3352,3355
evaluated|3356,3365
<EOL>|3366,3367
by|3367,3369
Gastroenterology|3370,3386
and|3387,3390
underwent|3391,3400
an|3401,3403
upper|3404,3409
endoscopy|3410,3419
on|3420,3422
_|3423,3424
_|3424,3425
_|3425,3426
.|3426,3427
<EOL>|3428,3429
This|3429,3433
showed|3434,3440
a|3441,3442
normal|3443,3449
appearing|3450,3459
esophagus|3460,3469
.|3469,3470
Biopsies|3471,3479
were|3480,3484
taken|3485,3490
.|3490,3491
<EOL>|3492,3493
<EOL>|3493,3494
TRANSITIONAL|3494,3506
ISSUES|3507,3513
:|3513,3514
<EOL>|3514,3515
-|3515,3516
f|3516,3517
/|3517,3518
u|3518,3519
biopsies|3520,3528
from|3529,3533
EGD|3534,3537
<EOL>|3537,3538
-|3538,3539
if|3539,3541
results|3542,3549
show|3550,3554
eosinophilic|3555,3567
esophagitis|3568,3579
,|3579,3580
follow|3581,3587
-|3587,3588
up|3588,3590
with|3591,3595
Dr.|3596,3599
_|3600,3601
_|3601,3602
_|3602,3603
.|3603,3604
<EOL>|3605,3606
_|3606,3607
_|3607,3608
_|3608,3609
for|3610,3613
management|3614,3624
<EOL>|3624,3625
-|3625,3626
pt|3626,3628
should|3629,3635
undergo|3636,3643
barium|3644,3650
swallow|3651,3658
as|3659,3661
an|3662,3664
outpatient|3665,3675
for|3676,3679
further|3680,3687
<EOL>|3688,3689
workup|3689,3695
of|3696,3698
her|3699,3702
dysphagia|3703,3712
<EOL>|3712,3713
-|3713,3714
f|3714,3715
/|3715,3716
u|3716,3717
with|3718,3722
ENT|3723,3726
as|3727,3729
planned|3730,3737
<EOL>|3737,3738
#|3738,3739
Code|3739,3743
:|3743,3744
Full|3745,3749
(|3750,3751
presumed|3751,3759
)|3759,3760
<EOL>|3761,3762
<EOL>|3763,3764
Medications|3764,3775
on|3776,3778
Admission|3779,3788
:|3788,3789
<EOL>|3789,3790
The|3790,3793
Preadmission|3794,3806
Medication|3807,3817
list|3818,3822
is|3823,3825
accurate|3826,3834
and|3835,3838
complete|3839,3847
.|3847,3848
<EOL>|3848,3849
1.|3849,3851
Omeprazole|3852,3862
20|3863,3865
mg|3866,3868
PO|3869,3871
BID|3872,3875
<EOL>|3876,3877
<EOL>|3877,3878
<EOL>|3879,3880
Discharge|3880,3889
Medications|3890,3901
:|3901,3902
<EOL>|3902,3903
1.|3903,3905
Omeprazole|3907,3917
20|3918,3920
mg|3921,3923
PO|3924,3926
BID|3927,3930
<EOL>|3932,3933
<EOL>|3933,3934
<EOL>|3935,3936
Discharge|3936,3945
Disposition|3946,3957
:|3957,3958
<EOL>|3958,3959
Home|3959,3963
<EOL>|3963,3964
<EOL>|3965,3966
Discharge|3966,3975
Diagnosis|3976,3985
:|3985,3986
<EOL>|3986,3987
-|4006,4007
dysphagia|4007,4016
and|4017,4020
foreign|4021,4028
body|4029,4033
sensation|4034,4043
<EOL>|4043,4044
<EOL>|4044,4045
SECONDARY|4045,4054
DIAGNOSIS|4055,4064
:|4064,4065
<EOL>|4065,4066
-|4066,4067
GERD|4067,4071
<EOL>|4072,4073
<EOL>|4073,4074
<EOL>|4075,4076
Mental|4097,4103
Status|4104,4110
:|4110,4111
Clear|4112,4117
and|4118,4121
coherent|4122,4130
.|4130,4131
<EOL>|4131,4132
Level|4132,4137
of|4138,4140
Consciousness|4141,4154
:|4154,4155
Alert|4156,4161
and|4162,4165
interactive|4166,4177
.|4177,4178
<EOL>|4178,4179
Activity|4179,4187
Status|4188,4194
:|4194,4195
Ambulatory|4196,4206
-|4207,4208
Independent|4209,4220
.|4220,4221
<EOL>|4221,4222
<EOL>|4222,4223
<EOL>|4224,4225
Dear|4249,4253
Ms.|4254,4257
_|4258,4259
_|4259,4260
_|4260,4261
,|4261,4262
<EOL>|4262,4263
<EOL>|4263,4264
You|4264,4267
were|4268,4272
hospitalized|4273,4285
at|4286,4288
_|4289,4290
_|4290,4291
_|4291,4292
.|4292,4293
<EOL>|4293,4294
<EOL>|4294,4295
You|4295,4298
came|4299,4303
in|4304,4306
due|4307,4310
to|4311,4313
difficulty|4314,4324
swallowing|4325,4335
.|4335,4336
You|4337,4340
had|4341,4344
an|4345,4347
endoscopy|4348,4357
<EOL>|4358,4359
to|4359,4361
look|4362,4366
for|4367,4370
any|4371,4374
abnormalities|4375,4388
in|4389,4391
the|4392,4395
esophagus|4396,4405
.|4405,4406
Thankfully|4407,4417
,|4417,4418
this|4419,4423
<EOL>|4424,4425
was|4425,4428
normal|4429,4435
.|4435,4436
They|4437,4441
took|4442,4446
biopsies|4447,4455
,|4455,4456
and|4457,4460
you|4461,4464
will|4465,4469
be|4470,4472
called|4473,4479
with|4480,4484
the|4485,4488
<EOL>|4489,4490
results|4490,4497
.|4497,4498
You|4499,4502
should|4503,4509
have|4510,4514
a|4515,4516
test|4517,4521
called|4522,4528
a|4529,4530
barium|4531,4537
swallow|4538,4545
as|4546,4548
an|4549,4551
<EOL>|4552,4553
outpatient|4553,4563
.|4563,4564
<EOL>|4564,4565
<EOL>|4565,4566
We|4566,4568
wish|4569,4573
you|4574,4577
all|4578,4581
the|4582,4585
best|4586,4590
!|4590,4591
<EOL>|4591,4592
-|4592,4593
Your|4593,4597
_|4598,4599
_|4599,4600
_|4600,4601
Team|4602,4606
<EOL>|4607,4608
<EOL>|4609,4610
Followup|4610,4618
Instructions|4619,4631
:|4631,4632
<EOL>|4632,4633
_|4633,4634
_|4634,4635
_|4635,4636
<EOL>|4636,4637

