 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Procedure|Health Care Activity|SIMPLE_SEGMENT|40,49|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|40,54|false|false|false|C2598112||Admission Date
Finding|Body Substance|SIMPLE_SEGMENT|74,83|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|74,83|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|74,83|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|74,83|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|74,88|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|106,111|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|106,111|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|106,111|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|130,133|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|130,133|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|130,133|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|130,133|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|130,133|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|141,148|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|141,148|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|150,158|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Finding|Body Substance|Allergies|173,180|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Allergies|173,180|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Allergies|173,180|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Attribute|Clinical Attribute|Allergies|209,218|true|false|false|C1717415||Allergies
Finding|Pathologic Function|Allergies|209,218|true|false|false|C0020517|Hypersensitivity|Allergies
Drug|Pharmacologic Substance|Allergies|222,227|false|false|false|C0013227|Pharmaceutical Preparations|Drugs
Procedure|Therapeutic or Preventive Procedure|Allergies|222,227|false|false|false|C3687832|Drugs - dental services|Drugs
Finding|Functional Concept|Allergies|230,239|false|false|false|C1999232|Attending (action)|Attending
Anatomy|Body Location or Region|Chief Complaint|264,273|false|false|false|C0000726|Abdomen|Abdominal
Finding|Finding|Chief Complaint|264,284|false|false|false|C0000731|Abdomen distended|Abdominal distention
Finding|Finding|Chief Complaint|274,284|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distention
Finding|Pathologic Function|Chief Complaint|274,284|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distention
Finding|Classification|Chief Complaint|288,293|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|294,302|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|294,302|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|306,324|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|315,324|false|false|false|C0945766||Procedure
Event|Occupational Activity|Chief Complaint|315,324|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|315,324|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|315,324|false|false|false|C0184661|Interventional procedure|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|326,338|false|false|false|C0034115|Paracentesis|Paracentesis
Drug|Antibiotic|History of Present Illness|385,389|false|false|false|C4087029|Nitroglycerin/Sodium Citrate/Ethanol Solution|nice
Drug|Organic Chemical|History of Present Illness|385,389|false|false|false|C4087029|Nitroglycerin/Sodium Citrate/Ethanol Solution|nice
Drug|Organic Chemical|History of Present Illness|405,409|false|false|false|C0001962|ethanol|ETOH
Drug|Pharmacologic Substance|History of Present Illness|405,409|false|false|false|C0001962|ethanol|ETOH
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|405,415|false|false|false|C0085762|Alcohol abuse|ETOH abuse
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|410,415|false|false|false|C0013146|Drug abuse|abuse
Event|Event|History of Present Illness|410,415|false|false|false|C1546935|Abuse|abuse
Finding|Finding|History of Present Illness|410,415|false|false|false|C0562381|Victim of abuse (finding)|abuse
Finding|Sign or Symptom|History of Present Illness|435,447|false|false|false|C0009806|Constipation|constipation
Anatomy|Body Location or Region|History of Present Illness|449,458|false|false|false|C0000726|Abdomen|abdominal
Finding|Finding|History of Present Illness|449,469|false|false|false|C0000731|Abdomen distended|abdominal distention
Finding|Finding|History of Present Illness|459,469|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distention
Finding|Pathologic Function|History of Present Illness|459,469|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distention
Finding|Body Substance|History of Present Illness|483,490|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|483,490|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|483,490|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Food|History of Present Illness|519,523|false|false|false|C0043188|Wine|wine
Finding|Idea or Concept|History of Present Illness|551,556|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Intellectual Product|History of Present Illness|551,556|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Sign or Symptom|History of Present Illness|557,562|false|false|false|C5551396|Binge eating behavior|binge
Finding|Individual Behavior|History of Present Illness|557,571|false|false|false|C0556346|Binge Drinking|binge drinking
Finding|Idea or Concept|History of Present Illness|576,579|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|History of Present Illness|576,579|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Idea or Concept|History of Present Illness|601,606|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Intellectual Product|History of Present Illness|601,606|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Gene or Genome|History of Present Illness|607,610|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Anatomy|Body Location or Region|History of Present Illness|624,633|false|false|false|C0000726|Abdomen|abdominal
Finding|Finding|History of Present Illness|624,644|false|false|false|C0000731|Abdomen distended|abdominal distension
Finding|Finding|History of Present Illness|634,644|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distension
Finding|Pathologic Function|History of Present Illness|634,644|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distension
Finding|Functional Concept|History of Present Illness|645,656|false|false|false|C0205329|Progressive|progressive
Finding|Intellectual Product|History of Present Illness|671,675|false|false|false|C1561540|Transaction counts and value totals - week|week
Drug|Biomedical or Dental Material|History of Present Illness|700,705|false|false|false|C0302909;C1378566|Solid Dose Form;solid substance|solid
Drug|Substance|History of Present Illness|700,705|false|false|false|C0302909;C1378566|Solid Dose Form;solid substance|solid
Finding|Body Substance|History of Present Illness|706,711|false|false|false|C0015733|Feces|stool
Finding|Sign or Symptom|History of Present Illness|750,753|false|false|false|C0013404|Dyspnea|SOB
Finding|Sign or Symptom|History of Present Illness|754,757|false|false|false|C0231807|Dyspnea on exertion|DOE
Finding|Finding|History of Present Illness|761,769|false|false|false|C0392756|Reduced|decrease
Finding|Finding|History of Present Illness|787,796|false|false|false|C0013220;C0020963;C0220929;C0231197|Drug Tolerance;Immune Tolerance;Mental tolerance;Physiologic tolerance|tolerance
Finding|Mental Process|History of Present Illness|787,796|false|false|false|C0013220;C0020963;C0220929;C0231197|Drug Tolerance;Immune Tolerance;Mental tolerance;Physiologic tolerance|tolerance
Finding|Pathologic Function|History of Present Illness|787,796|false|false|false|C0013220;C0020963;C0220929;C0231197|Drug Tolerance;Immune Tolerance;Mental tolerance;Physiologic tolerance|tolerance
Finding|Physiologic Function|History of Present Illness|787,796|false|false|false|C0013220;C0020963;C0220929;C0231197|Drug Tolerance;Immune Tolerance;Mental tolerance;Physiologic tolerance|tolerance
Finding|Daily or Recreational Activity|History of Present Illness|810,816|false|false|false|C0040802|travel|travel
Procedure|Health Care Activity|History of Present Illness|810,816|false|false|false|C1555670|travel charge|travel
Drug|Pharmacologic Substance|History of Present Illness|866,872|true|false|false|C0003211;C0358845|Analgesics and non-steroidal anti-inflammatory drugs;Anti-Inflammatory Agents, Non-Steroidal|NSAIDs
Drug|Organic Chemical|History of Present Illness|874,881|true|false|false|C0699142|Tylenol|Tylenol
Drug|Pharmacologic Substance|History of Present Illness|874,881|true|false|false|C0699142|Tylenol|Tylenol
Drug|Pharmacologic Substance|History of Present Illness|885,888|false|false|false|C0013231|Drugs, Non-Prescription|OTC
Finding|Gene or Genome|History of Present Illness|885,888|false|false|false|C1418193|OTC gene|OTC
Attribute|Clinical Attribute|History of Present Illness|889,900|true|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|History of Present Illness|889,900|true|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|History of Present Illness|889,900|true|false|false|C4284232|Medications|medications
Drug|Pharmacologic Substance|History of Present Illness|889,906|true|false|false|C1115771||medications other
Finding|Organism Function|History of Present Illness|982,989|false|false|false|C0025344|Menstruation|periods
Disorder|Disease or Syndrome|History of Present Illness|1017,1024|false|false|false|C0003962|Ascites|ascites
Finding|Pathologic Function|History of Present Illness|1017,1024|false|false|false|C5441966|Peritoneal Effusion|ascites
Disorder|Disease or Syndrome|History of Present Illness|1035,1046|false|false|false|C0015695;C2711227|Fatty Liver;Steatohepatitis|fatty liver
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1041,1046|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|History of Present Illness|1041,1046|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|History of Present Illness|1041,1046|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|History of Present Illness|1041,1046|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|History of Present Illness|1041,1046|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|History of Present Illness|1041,1046|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Finding|Finding|History of Present Illness|1041,1046|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|History of Present Illness|1041,1046|false|false|false|C0872387|Procedures on liver|liver
Finding|Idea or Concept|History of Present Illness|1048,1052|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Anatomy|Body Location or Region|History of Present Illness|1054,1060|false|false|false|C0205054|Hepatic|portal
Phenomenon|Natural Phenomenon or Process|History of Present Illness|1061,1065|false|false|false|C0806140|Flow|flow
Finding|Body Substance|History of Present Illness|1068,1075|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|1068,1075|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|1068,1075|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Organic Chemical|History of Present Illness|1106,1112|false|false|false|C0699187|Valium|valium
Drug|Pharmacologic Substance|History of Present Illness|1106,1112|false|false|false|C0699187|Valium|valium
Anatomy|Body Space or Junction|History of Present Illness|1123,1126|false|false|false|C0016520|Structure of interventricular foramen|IVF
Disorder|Disease or Syndrome|History of Present Illness|1123,1126|false|false|false|C2751898|Ventricular Fibrillation, Paroxysmal Familial, 1|IVF
Finding|Gene or Genome|History of Present Illness|1123,1126|false|false|false|C1419864;C4321334|SCN5A gene;SCN5A wt Allele|IVF
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1123,1126|false|false|false|C0015915;C0872104|Assisted Reproductive Technologies;Fertilization in Vitro|IVF
Drug|Organic Chemical|History of Present Illness|1143,1151|false|false|false|C0039840;C3714802|Thiamine Drug Class;thiamine|thiamine
Drug|Pharmacologic Substance|History of Present Illness|1143,1151|false|false|false|C0039840;C3714802|Thiamine Drug Class;thiamine|thiamine
Drug|Vitamin|History of Present Illness|1143,1151|false|false|false|C0039840;C3714802|Thiamine Drug Class;thiamine|thiamine
Procedure|Laboratory Procedure|History of Present Illness|1143,1151|false|false|false|C0373727|Thiamine measurement|thiamine
Drug|Organic Chemical|Past Medical History|1188,1195|false|false|false|C0001962;C0001975|Alcohols;ethanol|Alcohol
Drug|Pharmacologic Substance|Past Medical History|1188,1195|false|false|false|C0001962;C0001975|Alcohols;ethanol|Alcohol
Finding|Intellectual Product|Past Medical History|1188,1195|false|false|false|C1547288|Alcohol - Recreational Drug Use Code|Alcohol
Disorder|Mental or Behavioral Dysfunction|Past Medical History|1188,1201|false|false|false|C0085762|Alcohol abuse|Alcohol abuse
Disorder|Mental or Behavioral Dysfunction|Past Medical History|1196,1201|false|false|false|C0013146|Drug abuse|abuse
Event|Event|Past Medical History|1196,1201|false|false|false|C1546935|Abuse|abuse
Finding|Finding|Past Medical History|1196,1201|false|false|false|C0562381|Victim of abuse (finding)|abuse
Finding|Intellectual Product|Past Medical History|1204,1211|false|false|false|C1547296|Chronic - Admission Level of Care Code|Chronic
Procedure|Health Care Activity|Past Medical History|1204,1211|false|false|false|C1555457|Provision of recurring care for chronic illness|Chronic
Finding|Sign or Symptom|Past Medical History|1204,1221|false|true|false|C0740418|Chronic back pain|Chronic back pain
Finding|Sign or Symptom|Past Medical History|1212,1221|false|true|false|C0004604|Back Pain|back pain
Attribute|Clinical Attribute|Past Medical History|1217,1221|false|false|false|C2598155||pain
Finding|Functional Concept|Past Medical History|1217,1221|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Past Medical History|1217,1221|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1260,1266|false|false|false|C0006141|Breast|Breast
Disorder|Neoplastic Process|Family Medical History|1260,1266|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|Breast
Finding|Finding|Family Medical History|1260,1266|false|false|false|C0567499|Breast problem|Breast
Procedure|Therapeutic or Preventive Procedure|Family Medical History|1260,1266|false|false|false|C0191838|Procedures on breast|Breast
Disorder|Neoplastic Process|Family Medical History|1260,1269|false|false|false|C0006142|Malignant neoplasm of breast|Breast Ca
Finding|Idea or Concept|Family Medical History|1273,1279|false|false|false|C1546508|Relationship - Mother|mother
Attribute|Clinical Attribute|Family Medical History|1280,1283|false|false|false|C1114365||age
Drug|Biologically Active Substance|Family Medical History|1280,1283|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|Family Medical History|1280,1283|false|false|false|C0162574|Glycation End Products, Advanced|age
Disorder|Disease or Syndrome|Family Medical History|1292,1295|true|false|false|C0021390;C0022104|Inflammatory Bowel Diseases;Irritable Bowel Syndrome|IBD
Drug|Organic Chemical|Family Medical History|1292,1295|true|false|false|C0123047|ibudilast|IBD
Drug|Pharmacologic Substance|Family Medical History|1292,1295|true|false|false|C0123047|ibudilast|IBD
Finding|Gene or Genome|Family Medical History|1292,1295|true|false|false|C5780974|ACAD8 wt Allele|IBD
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1297,1302|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|Family Medical History|1297,1302|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|Family Medical History|1297,1302|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|Family Medical History|1297,1302|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|Family Medical History|1297,1302|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|Family Medical History|1297,1302|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Finding|Finding|Family Medical History|1297,1302|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|Family Medical History|1297,1302|false|false|false|C0872387|Procedures on liver|liver
Disorder|Disease or Syndrome|Family Medical History|1297,1310|true|false|false|C0085605|Liver Failure|liver failure
Finding|Functional Concept|Family Medical History|1303,1310|true|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|Family Medical History|1303,1310|true|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|Family Medical History|1303,1310|true|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Disorder|Mental or Behavioral Dysfunction|Family Medical History|1338,1348|false|false|false|C0001973|Alcoholic Intoxication, Chronic|alcoholism
Finding|Classification|General Exam|1402,1405|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|GEN
Finding|Gene or Genome|General Exam|1402,1405|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|GEN
Finding|Mental Process|General Exam|1414,1422|false|false|false|C2987187|Pleasant|pleasant
Finding|Finding|General Exam|1437,1441|false|false|false|C5575035|Well (answer to question)|well
Anatomy|Body Location or Region|General Exam|1454,1459|false|false|false|C1512338|HEENT|HEENT
Disorder|Disease or Syndrome|General Exam|1464,1480|true|false|false|C1112303|Facial wasting|temporal wasting
Finding|Finding|General Exam|1464,1480|true|false|false|C2029785|Temporal wasting|temporal wasting
Disorder|Disease or Syndrome|General Exam|1473,1480|true|false|false|C0235394|Wasting|wasting
Finding|Sign or Symptom|General Exam|1473,1480|true|false|false|C0006625|Cachexia|wasting
Finding|Finding|General Exam|1482,1485|true|false|false|C0425687|Jugular venous engorgement|JVD
Anatomy|Body Location or Region|General Exam|1500,1504|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|General Exam|1500,1504|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|General Exam|1500,1504|true|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Anatomy|Body Part, Organ, or Organ Component|General Exam|1500,1510|false|false|false|C0226542;C4266538|Neck>Neck veins;Structure of vein of neck|neck veins
Anatomy|Body Part, Organ, or Organ Component|General Exam|1505,1510|false|false|false|C0042449|Veins|veins
Procedure|Therapeutic or Preventive Procedure|General Exam|1505,1510|false|false|false|C0398102|Procedure on vein|veins
Event|Activity|General Exam|1511,1515|false|false|false|C1708059|Fill|fill
Finding|Idea or Concept|General Exam|1522,1527|false|false|false|C1552828|Table Frame - above|above
Finding|Gene or Genome|General Exam|1543,1546|true|false|false|C1422304|MAS1L gene|MRG
Procedure|Health Care Activity|General Exam|1549,1553|false|false|false|C1315068|Pulmonary ventilator management|PULM
Drug|Organic Chemical|General Exam|1555,1559|false|false|false|C0951233|cetrimonium bromide|CTAB
Finding|Finding|General Exam|1564,1573|false|false|false|C0392756;C0442797|Decreasing;Reduced|decreased
Anatomy|Body Location or Region|General Exam|1582,1586|false|false|false|C2987514|Anatomical base|base
Drug|Biomedical or Dental Material|General Exam|1582,1586|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Chemical Viewed Functionally|General Exam|1582,1586|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|1582,1586|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Finding|Gene or Genome|General Exam|1582,1586|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Finding|Idea or Concept|General Exam|1582,1586|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Anatomy|Body Location or Region|General Exam|1590,1593|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|ABD
Disorder|Cell or Molecular Dysfunction|General Exam|1590,1593|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|ABD
Finding|Finding|General Exam|1595,1604|false|false|false|C0700124|Dilated|Distended
Procedure|Diagnostic Procedure|General Exam|1636,1645|false|false|false|C0030247|Palpation|palpation
Finding|Sign or Symptom|General Exam|1663,1673|false|false|false|C0016204|Flatulence|flatulence
Anatomy|Body Part, Organ, or Organ Component|General Exam|1677,1682|false|false|false|C0015385|Limb structure|LIMBS
Attribute|Clinical Attribute|General Exam|1687,1692|false|false|false|C1717255||edema
Finding|Pathologic Function|General Exam|1687,1692|false|false|false|C0013604|Edema|edema
Anatomy|Body Part, Organ, or Organ Component|General Exam|1700,1703|false|false|false|C0227192|Inferior esophageal sphincter structure|LEs
Finding|Classification|General Exam|1700,1703|false|false|false|C0023595|Lewis Blood-Group System|LEs
Anatomy|Body Location or Region|General Exam|1707,1711|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Anatomy|Body Part, Organ, or Organ Component|General Exam|1707,1711|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Anatomy|Body Space or Junction|General Exam|1707,1711|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Procedure|Diagnostic Procedure|General Exam|1707,1711|false|false|false|C0562271|Examination of knee joint|knee
Drug|Food|General Exam|1728,1734|false|false|false|C5890763||pulses
Finding|Physiologic Function|General Exam|1728,1734|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|General Exam|1728,1734|false|false|false|C0034107|Pulse taking|pulses
Finding|Sign or Symptom|General Exam|1763,1772|true|false|false|C0232766|Asterixis|asterixis
Finding|Finding|General Exam|1774,1783|true|false|false|C4036115|Very mild|very mild
Finding|Intellectual Product|General Exam|1779,1783|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Classification|General Exam|1784,1791|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|general
Procedure|Health Care Activity|General Exam|1784,1791|false|false|false|C3812897|General medical service|general
Finding|Sign or Symptom|General Exam|1792,1798|false|false|false|C0040822|Tremor|tremor
Disorder|Disease or Syndrome|General Exam|1836,1841|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|1836,1841|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|1842,1845|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|1852,1855|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|1852,1855|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|1852,1855|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|1862,1865|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|1862,1865|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|1862,1865|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|1862,1865|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|1871,1874|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|1871,1874|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|1881,1884|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|General Exam|1881,1884|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|1881,1884|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|1881,1884|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|1890,1893|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|1890,1893|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|General Exam|1890,1893|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|1890,1893|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|1890,1893|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|General Exam|1900,1904|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|1919,1922|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|1939,1944|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|1939,1944|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|1945,1948|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|1955,1958|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|1955,1958|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|1955,1958|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|1965,1968|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|1965,1968|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|1965,1968|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|1965,1968|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|1974,1977|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|1974,1977|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|1984,1987|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|General Exam|1984,1987|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|1984,1987|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|1984,1987|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|1993,1996|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|1993,1996|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|General Exam|1993,1996|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|1993,1996|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|1993,1996|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|General Exam|2003,2007|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|2022,2025|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|2042,2047|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|2042,2047|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|2048,2051|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|2058,2061|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|2058,2061|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|2058,2061|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|2068,2071|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|2068,2071|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|2068,2071|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|2068,2071|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|2077,2080|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|2077,2080|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|2087,2090|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|General Exam|2087,2090|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|2087,2090|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|2087,2090|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|2096,2099|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|2096,2099|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|General Exam|2096,2099|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|2096,2099|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|2096,2099|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|General Exam|2106,2110|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|2125,2128|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|2145,2150|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|2145,2150|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|2151,2154|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|2161,2164|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|2161,2164|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|2161,2164|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|2171,2174|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|2171,2174|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|2171,2174|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|2171,2174|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|2180,2183|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|2180,2183|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|2190,2193|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|General Exam|2190,2193|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|2190,2193|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|2190,2193|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|2199,2202|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|2199,2202|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|General Exam|2199,2202|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|2199,2202|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|2199,2202|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|General Exam|2209,2213|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|2228,2231|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|2248,2253|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|2248,2253|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|2254,2257|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|2264,2267|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|2264,2267|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|2264,2267|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|2274,2277|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|2274,2277|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|2274,2277|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|2274,2277|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|2284,2287|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|2284,2287|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|2295,2298|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|General Exam|2295,2298|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|2295,2298|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|2295,2298|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|2304,2307|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|2304,2307|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|General Exam|2304,2307|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|2304,2307|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|2304,2307|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|General Exam|2314,2318|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|2333,2336|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|2353,2358|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|2353,2358|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|2359,2362|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|2369,2372|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|2369,2372|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|2369,2372|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|2379,2382|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|2379,2382|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|2379,2382|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|2379,2382|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|2388,2391|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|2388,2391|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|2398,2401|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|General Exam|2398,2401|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|2398,2401|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|2398,2401|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|2407,2410|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|2407,2410|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|General Exam|2407,2410|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|2407,2410|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|2407,2410|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|General Exam|2417,2421|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|2436,2439|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|2456,2461|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|2456,2461|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Finding|Body Substance|General Exam|2474,2480|false|false|false|C0024202|Lymph|Lymphs
Drug|Antibiotic|General Exam|2487,2492|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|General Exam|2487,2492|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|General Exam|2487,2492|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|General Exam|2498,2501|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|Eos
Finding|Gene or Genome|General Exam|2498,2501|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|Eos
Disorder|Disease or Syndrome|General Exam|2527,2532|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|2527,2532|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|2533,2536|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|2553,2558|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|2553,2558|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|2563,2566|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Procedure|Laboratory Procedure|General Exam|2563,2566|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|General Exam|2585,2590|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|2585,2590|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|2591,2594|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|2611,2616|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|2611,2616|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|2621,2624|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Procedure|Laboratory Procedure|General Exam|2621,2624|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|General Exam|2647,2652|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|2647,2652|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|2653,2656|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|2673,2678|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|2673,2678|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|2683,2686|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Procedure|Laboratory Procedure|General Exam|2683,2686|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|General Exam|2708,2713|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|2708,2713|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|2714,2717|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|2734,2739|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|2734,2739|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|2744,2747|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Procedure|Laboratory Procedure|General Exam|2744,2747|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|General Exam|2769,2774|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|2769,2774|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|2775,2778|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|2795,2800|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|2795,2800|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|2805,2808|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Procedure|Laboratory Procedure|General Exam|2805,2808|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|General Exam|2830,2835|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|2830,2835|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|2836,2839|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|2856,2861|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|2856,2861|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|2856,2869|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|2856,2869|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|2856,2869|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|2862,2869|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|2862,2869|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|2862,2869|false|false|false|C0017725|glucose|Glucose
Lab|Laboratory or Test Result|General Exam|2862,2869|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|2862,2869|false|false|false|C0337438|Glucose measurement|Glucose
Disorder|Disease or Syndrome|General Exam|2946,2951|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|2946,2951|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|2946,2959|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|2946,2959|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|2946,2959|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|2952,2959|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|2952,2959|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|2952,2959|false|false|false|C0017725|glucose|Glucose
Lab|Laboratory or Test Result|General Exam|2952,2959|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|2952,2959|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|General Exam|3007,3011|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|3007,3011|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|General Exam|3007,3011|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|General Exam|3036,3041|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|3036,3041|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|3036,3049|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|3036,3049|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|3036,3049|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|3042,3049|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|3042,3049|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|3042,3049|false|false|false|C0017725|glucose|Glucose
Lab|Laboratory or Test Result|General Exam|3042,3049|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|3042,3049|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|General Exam|3094,3098|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|3094,3098|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|General Exam|3094,3098|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|General Exam|3123,3128|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|3123,3128|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|3123,3136|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|3123,3136|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|3123,3136|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|3129,3136|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|3129,3136|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|3129,3136|false|false|false|C0017725|glucose|Glucose
Lab|Laboratory or Test Result|General Exam|3129,3136|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|3129,3136|false|false|false|C0337438|Glucose measurement|Glucose
Disorder|Disease or Syndrome|General Exam|3212,3217|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|3212,3217|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|3212,3225|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|3212,3225|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|3212,3225|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|3218,3225|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|3218,3225|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|3218,3225|false|false|false|C0017725|glucose|Glucose
Lab|Laboratory or Test Result|General Exam|3218,3225|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|3218,3225|false|false|false|C0337438|Glucose measurement|Glucose
Disorder|Disease or Syndrome|General Exam|3299,3304|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|3299,3304|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|3299,3312|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|3299,3312|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|3299,3312|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|3305,3312|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|3305,3312|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|3305,3312|false|false|false|C0017725|glucose|Glucose
Lab|Laboratory or Test Result|General Exam|3305,3312|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|3305,3312|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|General Exam|3357,3361|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|3357,3361|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|General Exam|3357,3361|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|General Exam|3386,3391|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|3386,3391|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|3392,3395|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|General Exam|3392,3395|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|General Exam|3392,3395|false|false|false|C0001899|Alanine Transaminase|ALT
Finding|Gene or Genome|General Exam|3392,3395|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|General Exam|3392,3395|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|General Exam|3392,3395|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|General Exam|3392,3395|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|General Exam|3400,3403|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|General Exam|3400,3403|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|3400,3403|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|General Exam|3400,3403|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|General Exam|3400,3403|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Finding|Gene or Genome|General Exam|3400,3403|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|3409,3416|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|General Exam|3409,3416|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Disorder|Disease or Syndrome|General Exam|3448,3453|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|3448,3453|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|3454,3457|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|General Exam|3454,3457|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|General Exam|3454,3457|false|false|false|C0001899|Alanine Transaminase|ALT
Finding|Gene or Genome|General Exam|3454,3457|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|General Exam|3454,3457|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|General Exam|3454,3457|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|General Exam|3454,3457|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|General Exam|3462,3465|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|General Exam|3462,3465|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|3462,3465|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|General Exam|3462,3465|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|General Exam|3462,3465|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Finding|Gene or Genome|General Exam|3462,3465|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|3485,3492|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|General Exam|3485,3492|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Disorder|Disease or Syndrome|General Exam|3523,3528|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|3523,3528|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|3529,3532|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|General Exam|3529,3532|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|General Exam|3529,3532|false|false|false|C0001899|Alanine Transaminase|ALT
Finding|Gene or Genome|General Exam|3529,3532|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|General Exam|3529,3532|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|General Exam|3529,3532|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|General Exam|3529,3532|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|General Exam|3537,3540|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|General Exam|3537,3540|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|3537,3540|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|General Exam|3537,3540|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|General Exam|3537,3540|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Finding|Gene or Genome|General Exam|3537,3540|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|3546,3553|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|General Exam|3546,3553|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Disorder|Disease or Syndrome|General Exam|3585,3590|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|3585,3590|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|3591,3594|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|General Exam|3591,3594|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|General Exam|3591,3594|false|false|false|C0001899|Alanine Transaminase|ALT
Finding|Gene or Genome|General Exam|3591,3594|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|General Exam|3591,3594|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|General Exam|3591,3594|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|General Exam|3591,3594|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|General Exam|3599,3602|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|General Exam|3599,3602|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|3599,3602|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|General Exam|3599,3602|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|General Exam|3599,3602|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Finding|Gene or Genome|General Exam|3599,3602|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|3608,3615|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|General Exam|3608,3615|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Disorder|Disease or Syndrome|General Exam|3647,3652|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|3647,3652|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|3653,3656|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|General Exam|3653,3656|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|General Exam|3653,3656|false|false|false|C0001899|Alanine Transaminase|ALT
Finding|Gene or Genome|General Exam|3653,3656|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|General Exam|3653,3656|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|General Exam|3653,3656|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|General Exam|3653,3656|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|General Exam|3661,3664|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|General Exam|3661,3664|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|3661,3664|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|General Exam|3661,3664|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|General Exam|3661,3664|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Finding|Gene or Genome|General Exam|3661,3664|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|3673,3676|false|false|false|C0022917|Lactate Dehydrogenase|LDH
Drug|Enzyme|General Exam|3673,3676|false|false|false|C0022917|Lactate Dehydrogenase|LDH
Finding|Finding|General Exam|3673,3676|false|false|false|C0851148|Lifetime Drinking History|LDH
Procedure|Laboratory Procedure|General Exam|3673,3676|false|false|false|C0202113|Lactate dehydrogenase measurement|LDH
Drug|Amino Acid, Peptide, or Protein|General Exam|3684,3691|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|General Exam|3684,3691|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Disorder|Disease or Syndrome|General Exam|3722,3727|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|3722,3727|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|3728,3731|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|General Exam|3728,3731|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|General Exam|3728,3731|false|false|false|C0001899|Alanine Transaminase|ALT
Finding|Gene or Genome|General Exam|3728,3731|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|General Exam|3728,3731|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|General Exam|3728,3731|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|General Exam|3728,3731|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|General Exam|3736,3739|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|General Exam|3736,3739|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|3736,3739|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|General Exam|3736,3739|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|General Exam|3736,3739|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Finding|Gene or Genome|General Exam|3736,3739|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|3761,3764|false|false|false|C0010287|Creatine Kinase|CPK
Drug|Enzyme|General Exam|3761,3764|false|false|false|C0010287|Creatine Kinase|CPK
Finding|Gene or Genome|General Exam|3761,3764|false|false|false|C1418571|PIK3C2A gene|CPK
Procedure|Laboratory Procedure|General Exam|3761,3764|false|false|false|C0201973|Creatine kinase measurement|CPK
Drug|Amino Acid, Peptide, or Protein|General Exam|3770,3777|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|General Exam|3770,3777|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Disorder|Disease or Syndrome|General Exam|3807,3812|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|3807,3812|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|3813,3819|false|false|false|C0023764|lipase|Lipase
Drug|Enzyme|General Exam|3813,3819|false|false|false|C0023764|lipase|Lipase
Drug|Pharmacologic Substance|General Exam|3813,3819|false|false|false|C0023764|lipase|Lipase
Procedure|Laboratory Procedure|General Exam|3813,3819|false|false|false|C0373670|Lipase measurement|Lipase
Disorder|Disease or Syndrome|General Exam|3835,3840|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|3835,3840|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|3841,3847|false|false|false|C0023764|lipase|Lipase
Drug|Enzyme|General Exam|3841,3847|false|false|false|C0023764|lipase|Lipase
Drug|Pharmacologic Substance|General Exam|3841,3847|false|false|false|C0023764|lipase|Lipase
Procedure|Laboratory Procedure|General Exam|3841,3847|false|false|false|C0373670|Lipase measurement|Lipase
Drug|Amino Acid, Peptide, or Protein|General Exam|3851,3854|false|false|false|C0017040|Gamma-glutamyl transferase|GGT
Drug|Enzyme|General Exam|3851,3854|false|false|false|C0017040|Gamma-glutamyl transferase|GGT
Finding|Gene or Genome|General Exam|3851,3854|false|false|false|C1415053;C1415054|GGT1 gene;GGT2P gene|GGT
Procedure|Laboratory Procedure|General Exam|3851,3854|false|false|false|C0202035|Gamma glutamyl transferase measurement|GGT
Disorder|Disease or Syndrome|General Exam|3873,3878|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|3873,3878|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|3873,3886|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|General Exam|3879,3886|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|General Exam|3879,3886|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|General Exam|3879,3886|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|General Exam|3879,3886|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|General Exam|3879,3886|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Finding|Physiologic Function|General Exam|3879,3886|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|General Exam|3879,3886|false|false|false|C0201925|Calcium measurement|Calcium
Disorder|Disease or Syndrome|General Exam|3921,3926|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|3921,3926|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|3921,3934|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|General Exam|3927,3934|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|General Exam|3927,3934|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|General Exam|3927,3934|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|General Exam|3927,3934|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|General Exam|3927,3934|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Finding|Physiologic Function|General Exam|3927,3934|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|General Exam|3927,3934|false|false|false|C0201925|Calcium measurement|Calcium
Disorder|Disease or Syndrome|General Exam|3969,3974|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|3969,3974|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|3969,3982|false|false|false|C0853248|Blood albumin|BLOOD Albumin
Drug|Amino Acid, Peptide, or Protein|General Exam|3975,3982|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Biologically Active Substance|General Exam|3975,3982|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Pharmacologic Substance|General Exam|3975,3982|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Finding|Gene or Genome|General Exam|3975,3982|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Finding|Physiologic Function|General Exam|3975,3982|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Procedure|Laboratory Procedure|General Exam|3975,3982|false|false|false|C0201838|Albumin measurement|Albumin
Drug|Biologically Active Substance|General Exam|3988,3995|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|General Exam|3988,3995|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|General Exam|3988,3995|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|General Exam|3988,3995|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|General Exam|3988,3995|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Finding|Physiologic Function|General Exam|3988,3995|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|General Exam|3988,3995|false|false|false|C0201925|Calcium measurement|Calcium
Drug|Biologically Active Substance|General Exam|4019,4023|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Drug|Element, Ion, or Isotope|General Exam|4019,4023|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Drug|Pharmacologic Substance|General Exam|4019,4023|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Procedure|Laboratory Procedure|General Exam|4019,4023|false|false|false|C0337439|Iron measurement|Iron
Disorder|Disease or Syndrome|General Exam|4039,4044|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4039,4044|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|4039,4052|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|General Exam|4045,4052|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|General Exam|4045,4052|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|General Exam|4045,4052|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|General Exam|4045,4052|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|General Exam|4045,4052|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Finding|Physiologic Function|General Exam|4045,4052|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|General Exam|4045,4052|false|false|false|C0201925|Calcium measurement|Calcium
Disorder|Disease or Syndrome|General Exam|4087,4092|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4087,4092|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|4087,4100|false|false|false|C0853248|Blood albumin|BLOOD Albumin
Drug|Amino Acid, Peptide, or Protein|General Exam|4093,4100|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Biologically Active Substance|General Exam|4093,4100|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Pharmacologic Substance|General Exam|4093,4100|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Finding|Gene or Genome|General Exam|4093,4100|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Finding|Physiologic Function|General Exam|4093,4100|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Procedure|Laboratory Procedure|General Exam|4093,4100|false|false|false|C0201838|Albumin measurement|Albumin
Drug|Biologically Active Substance|General Exam|4106,4113|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|General Exam|4106,4113|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|General Exam|4106,4113|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|General Exam|4106,4113|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|General Exam|4106,4113|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Finding|Physiologic Function|General Exam|4106,4113|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|General Exam|4106,4113|false|false|false|C0201925|Calcium measurement|Calcium
Drug|Biologically Active Substance|General Exam|4137,4141|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Drug|Element, Ion, or Isotope|General Exam|4137,4141|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Drug|Pharmacologic Substance|General Exam|4137,4141|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Procedure|Laboratory Procedure|General Exam|4137,4141|false|false|false|C0337439|Iron measurement|Iron
Disorder|Disease or Syndrome|General Exam|4157,4162|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4157,4162|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|4157,4170|false|false|false|C0853248|Blood albumin|BLOOD Albumin
Drug|Amino Acid, Peptide, or Protein|General Exam|4163,4170|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Biologically Active Substance|General Exam|4163,4170|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Pharmacologic Substance|General Exam|4163,4170|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Finding|Gene or Genome|General Exam|4163,4170|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Finding|Physiologic Function|General Exam|4163,4170|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Procedure|Laboratory Procedure|General Exam|4163,4170|false|false|false|C0201838|Albumin measurement|Albumin
Disorder|Disease or Syndrome|General Exam|4188,4193|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4188,4193|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|4252,4255|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Drug|Biologically Active Substance|General Exam|4252,4255|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Drug|Hormone|General Exam|4252,4255|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Drug|Pharmacologic Substance|General Exam|4252,4255|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Finding|Gene or Genome|General Exam|4252,4255|false|false|false|C1334121;C1336604;C1705002|IL5 gene;TERF1 gene;TERF1 wt Allele|TRF
Disorder|Disease or Syndrome|General Exam|4273,4278|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4273,4278|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Attribute|Clinical Attribute|General Exam|4279,4282|false|false|false|C2708739||TSH
Drug|Amino Acid, Peptide, or Protein|General Exam|4279,4282|false|false|false|C0040160|thyrotropin|TSH
Drug|Hormone|General Exam|4279,4282|false|false|false|C0040160|thyrotropin|TSH
Drug|Pharmacologic Substance|General Exam|4279,4282|false|false|false|C0040160|thyrotropin|TSH
Procedure|Laboratory Procedure|General Exam|4279,4282|false|false|false|C0202230|Thyroid stimulating hormone measurement|TSH
Disorder|Disease or Syndrome|General Exam|4300,4305|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4300,4305|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Finding|Functional Concept|General Exam|4306,4310|false|false|false|C0332296|Free of (attribute)|Free
Procedure|Laboratory Procedure|General Exam|4306,4313|false|false|false|C0202225|T4 free measurement|Free T4
Disorder|Disease or Syndrome|General Exam|4330,4335|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4330,4335|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|4336,4341|false|false|false|C0019168;C0796320|Hepatitis B Antigen Vaccine;Hepatitis B Surface Antigens|HBsAg
Drug|Immunologic Factor|General Exam|4336,4341|false|false|false|C0019168;C0796320|Hepatitis B Antigen Vaccine;Hepatitis B Surface Antigens|HBsAg
Drug|Pharmacologic Substance|General Exam|4336,4341|false|false|false|C0019168;C0796320|Hepatitis B Antigen Vaccine;Hepatitis B Surface Antigens|HBsAg
Procedure|Laboratory Procedure|General Exam|4336,4341|false|false|false|C0201477|Hepatitis B surface antigen measurement|HBsAg
Finding|Classification|General Exam|4342,4350|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|NEGATIVE
Finding|Finding|General Exam|4342,4350|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|NEGATIVE
Lab|Laboratory or Test Result|General Exam|4342,4350|false|false|false|C5237010|Expression Negative|NEGATIVE
Drug|Amino Acid, Peptide, or Protein|General Exam|4351,4356|false|false|false|C0369334|Hepatitis B Virus Surface Antibody|HBsAb
Drug|Immunologic Factor|General Exam|4351,4356|false|false|false|C0369334|Hepatitis B Virus Surface Antibody|HBsAb
Disorder|Cell or Molecular Dysfunction|General Exam|4357,4365|false|false|false|C4727483|BRAF Gene Rearrangement|POSITIVE
Finding|Classification|General Exam|4357,4365|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|POSITIVE
Finding|Finding|General Exam|4357,4365|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|POSITIVE
Drug|Amino Acid, Peptide, or Protein|General Exam|4367,4372|false|false|false|C0312631|Antibody to hepatitis B core antigen|HBcAb
Drug|Immunologic Factor|General Exam|4367,4372|false|false|false|C0312631|Antibody to hepatitis B core antigen|HBcAb
Drug|Pharmacologic Substance|General Exam|4367,4372|false|false|false|C0312631|Antibody to hepatitis B core antigen|HBcAb
Finding|Classification|General Exam|4373,4381|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|NEGATIVE
Finding|Finding|General Exam|4373,4381|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|NEGATIVE
Lab|Laboratory or Test Result|General Exam|4373,4381|false|false|false|C5237010|Expression Negative|NEGATIVE
Disorder|Disease or Syndrome|General Exam|4382,4385|false|false|false|C0019159|Hepatitis A|HAV
Disorder|Cell or Molecular Dysfunction|General Exam|4389,4397|false|false|false|C4727483|BRAF Gene Rearrangement|POSITIVE
Finding|Classification|General Exam|4389,4397|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|POSITIVE
Finding|Finding|General Exam|4389,4397|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|POSITIVE
Drug|Amino Acid, Peptide, or Protein|General Exam|4398,4401|false|false|false|C0020861|Immunoglobulin M|IgM
Drug|Immunologic Factor|General Exam|4398,4401|false|false|false|C0020861|Immunoglobulin M|IgM
Finding|Gene or Genome|General Exam|4398,4401|false|false|false|C1706005|CD40LG wt Allele|IgM
Procedure|Laboratory Procedure|General Exam|4398,4401|false|false|false|C0202084|Immunoglobulin M measurement|IgM
Disorder|Disease or Syndrome|General Exam|4402,4405|false|false|false|C0019159|Hepatitis A|HAV
Finding|Classification|General Exam|4406,4414|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|NEGATIVE
Finding|Finding|General Exam|4406,4414|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|NEGATIVE
Lab|Laboratory or Test Result|General Exam|4406,4414|false|false|false|C5237010|Expression Negative|NEGATIVE
Disorder|Disease or Syndrome|General Exam|4427,4432|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4427,4432|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|General Exam|4433,4436|false|false|false|C5887323|HYPERTRICHOSIS, CONGENITAL GENERALIZED, 2|HCG
Drug|Amino Acid, Peptide, or Protein|General Exam|4433,4436|false|false|false|C1141639;C1527152|Recombinant Human Chorionic Gonadotropin;human chorionic gonadotropin|HCG
Drug|Hormone|General Exam|4433,4436|false|false|false|C1141639;C1527152|Recombinant Human Chorionic Gonadotropin;human chorionic gonadotropin|HCG
Drug|Pharmacologic Substance|General Exam|4433,4436|false|false|false|C1141639;C1527152|Recombinant Human Chorionic Gonadotropin;human chorionic gonadotropin|HCG
Finding|Gene or Genome|General Exam|4433,4436|false|false|false|C1413366;C1415796;C1424291;C4321295|CGA gene;CGA wt Allele;CGB5 gene;HTC2 gene|HCG
Disorder|Disease or Syndrome|General Exam|4452,4457|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4452,4457|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Finding|Finding|General Exam|4458,4461|false|false|false|C5891060|Against Medical Advice|AMA
Procedure|Therapeutic or Preventive Procedure|General Exam|4458,4461|false|false|false|C0279755|cytarabine/melphalan|AMA
Finding|Classification|General Exam|4462,4470|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|NEGATIVE
Finding|Finding|General Exam|4462,4470|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|NEGATIVE
Lab|Laboratory or Test Result|General Exam|4462,4470|false|false|false|C5237010|Expression Negative|NEGATIVE
Finding|Classification|General Exam|4478,4486|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|NEGATIVE
Finding|Finding|General Exam|4478,4486|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|NEGATIVE
Lab|Laboratory or Test Result|General Exam|4478,4486|false|false|false|C5237010|Expression Negative|NEGATIVE
Disorder|Disease or Syndrome|General Exam|4499,4504|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4499,4504|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|General Exam|4521,4526|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4521,4526|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|General Exam|4527,4530|false|false|false|C0019682;C0019693|HIV;HIV Infections|HIV
Disorder|Virus|General Exam|4527,4530|false|false|false|C0019682;C0019693|HIV;HIV Infections|HIV
Drug|Immunologic Factor|General Exam|4527,4530|false|false|false|C0086413|HIV Vaccine|HIV
Drug|Pharmacologic Substance|General Exam|4527,4530|false|false|false|C0086413|HIV Vaccine|HIV
Finding|Classification|General Exam|4534,4542|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|NEGATIVE
Finding|Finding|General Exam|4534,4542|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|NEGATIVE
Lab|Laboratory or Test Result|General Exam|4534,4542|false|false|false|C5237010|Expression Negative|NEGATIVE
Disorder|Disease or Syndrome|General Exam|4555,4560|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4555,4560|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|4561,4564|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Enzyme|General Exam|4561,4564|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Organic Chemical|General Exam|4561,4564|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Pharmacologic Substance|General Exam|4561,4564|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Finding|Gene or Genome|General Exam|4561,4564|false|false|false|C1412553|ARSA gene|ASA
Finding|Finding|General Exam|4565,4568|false|false|false|C5848551|Neg - answer|NEG
Finding|Finding|General Exam|4581,4584|false|false|false|C5848551|Neg - answer|NEG
Finding|Finding|General Exam|4594,4597|false|false|false|C5848551|Neg - answer|NEG
Finding|Finding|General Exam|4606,4609|false|false|false|C5848551|Neg - answer|NEG
Finding|Finding|General Exam|4618,4621|false|false|false|C5848551|Neg - answer|NEG
Disorder|Disease or Syndrome|General Exam|4634,4639|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4634,4639|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Event|Activity|General Exam|4648,4652|false|false|false|C1948035|Hold (action)|HOLD
Finding|Functional Concept|General Exam|4648,4652|false|false|false|C1553387;C3853841|Hold - dosing instruction fragment;hold - Data Operation|HOLD
Finding|Intellectual Product|General Exam|4648,4652|false|false|false|C1553387;C3853841|Hold - dosing instruction fragment;hold - Data Operation|HOLD
Disorder|Disease or Syndrome|General Exam|4665,4670|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4665,4670|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Event|Activity|General Exam|4679,4683|false|false|false|C1948035|Hold (action)|HOLD
Finding|Functional Concept|General Exam|4679,4683|false|false|false|C1553387;C3853841|Hold - dosing instruction fragment;hold - Data Operation|HOLD
Finding|Intellectual Product|General Exam|4679,4683|false|false|false|C1553387;C3853841|Hold - dosing instruction fragment;hold - Data Operation|HOLD
Disorder|Disease or Syndrome|General Exam|4696,4701|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4696,4701|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|General Exam|4702,4705|false|false|false|C0019196;C0220847|Hepatitis C;hepatitis C virus|HCV
Disorder|Virus|General Exam|4702,4705|false|false|false|C0019196;C0220847|Hepatitis C;hepatitis C virus|HCV
Finding|Classification|General Exam|4709,4717|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|NEGATIVE
Finding|Finding|General Exam|4709,4717|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|NEGATIVE
Lab|Laboratory or Test Result|General Exam|4709,4717|false|false|false|C5237010|Expression Negative|NEGATIVE
Disorder|Disease or Syndrome|General Exam|4730,4735|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4730,4735|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|4730,4743|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|4730,4743|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|4730,4743|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|4736,4743|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|4736,4743|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|4736,4743|false|false|false|C0017725|glucose|Glucose
Lab|Laboratory or Test Result|General Exam|4736,4743|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|4736,4743|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Organic Chemical|General Exam|4749,4756|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Drug|Pharmacologic Substance|General Exam|4749,4756|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Procedure|Laboratory Procedure|General Exam|4749,4756|false|false|false|C0202115|Lactic acid measurement|Lactate
Disorder|Disease or Syndrome|General Exam|4774,4779|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4774,4779|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|4780,4793|false|false|false|C0007841;C5441691|CP protein, human;Ceruloplasmin|CERULOPLASMIN
Drug|Enzyme|General Exam|4780,4793|false|false|false|C0007841;C5441691|CP protein, human;Ceruloplasmin|CERULOPLASMIN
Finding|Gene or Genome|General Exam|4780,4793|false|false|false|C1151847;C1439306|CP gene;ferroxidase activity|CERULOPLASMIN
Finding|Molecular Function|General Exam|4780,4793|false|false|false|C1151847;C1439306|CP gene;ferroxidase activity|CERULOPLASMIN
Procedure|Laboratory Procedure|General Exam|4780,4793|false|false|false|C0373573|Ceruloplasmin measurement|CERULOPLASMIN
Disorder|Disease or Syndrome|General Exam|4794,4797|false|false|false|C1956415|Paroxysmal nocturnal dyspnea|PND
Finding|Gene or Genome|General Exam|4794,4797|false|false|false|C1417807;C4552608|NPPA gene;NPPA wt Allele|PND
Disorder|Disease or Syndrome|General Exam|4810,4815|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4810,4815|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|4816,4821|false|false|false|C5400714|ALPHA (substance)|ALPHA
Drug|Pharmacologic Substance|General Exam|4816,4821|false|false|false|C5400714|ALPHA (substance)|ALPHA
Finding|Intellectual Product|General Exam|4816,4821|false|false|false|C0439095|Greek letter alpha (qualifier value)|ALPHA
Drug|Amino Acid, Peptide, or Protein|General Exam|4816,4823|false|false|false|C1979844|Alpha-1|ALPHA-1
Drug|Amino Acid, Peptide, or Protein|General Exam|4816,4835|false|false|false|C0002191;C1455316|SERPINA1 protein, human;alpha 1-antitrypsin|ALPHA-1-ANTITRYPSIN
Drug|Biologically Active Substance|General Exam|4816,4835|false|false|false|C0002191;C1455316|SERPINA1 protein, human;alpha 1-antitrypsin|ALPHA-1-ANTITRYPSIN
Drug|Pharmacologic Substance|General Exam|4816,4835|false|false|false|C0002191;C1455316|SERPINA1 protein, human;alpha 1-antitrypsin|ALPHA-1-ANTITRYPSIN
Finding|Gene or Genome|General Exam|4816,4835|false|false|false|C1418544|SERPINA1 gene|ALPHA-1-ANTITRYPSIN
Procedure|Laboratory Procedure|General Exam|4816,4835|false|false|false|C0201856|Alpha-1-antitrypsin measurement|ALPHA-1-ANTITRYPSIN
Drug|Amino Acid, Peptide, or Protein|General Exam|4824,4835|false|false|false|C2713669|SERPINA5 protein, human|ANTITRYPSIN
Drug|Biologically Active Substance|General Exam|4824,4835|false|false|false|C2713669|SERPINA5 protein, human|ANTITRYPSIN
Finding|Gene or Genome|General Exam|4824,4835|false|false|false|C1418544|SERPINA1 gene|ANTITRYPSIN
Disorder|Disease or Syndrome|General Exam|4836,4839|false|false|false|C1956415|Paroxysmal nocturnal dyspnea|PND
Finding|Gene or Genome|General Exam|4836,4839|false|false|false|C1417807;C4552608|NPPA gene;NPPA wt Allele|PND
Finding|Finding|General Exam|4841,4848|false|false|false|C0740845|Imaging problem|Imaging
Procedure|Diagnostic Procedure|General Exam|4841,4848|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|Imaging
Attribute|Clinical Attribute|General Exam|4853,4859|false|false|false|C0881797||US abd
Anatomy|Body Location or Region|General Exam|4856,4859|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|abd
Disorder|Cell or Molecular Dysfunction|General Exam|4856,4859|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|abd
Anatomy|Body Part, Organ, or Organ Component|General Exam|4860,4866|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Anatomy|Body Space or Junction|General Exam|4860,4866|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Disorder|Neoplastic Process|General Exam|4860,4866|false|false|false|C0153663|Malignant neoplasm of pelvis|pelvis
Finding|Finding|General Exam|4860,4866|false|false|false|C0812455|Pelvis problem|pelvis
Finding|Finding|Impression|4893,4902|false|false|false|C4697723|Echogenic|echogenic
Anatomy|Body Part, Organ, or Organ Component|Impression|4903,4908|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|Impression|4903,4908|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|Impression|4903,4908|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|Impression|4903,4908|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|Impression|4903,4908|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|Impression|4903,4908|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Finding|Finding|Impression|4903,4908|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|Impression|4903,4908|false|false|false|C0872387|Procedures on liver|liver
Finding|Functional Concept|Impression|4910,4920|false|false|false|C0332299|Suggestive of|suggestive
Finding|Functional Concept|Impression|4910,4923|false|false|false|C0332299|Suggestive of|suggestive of
Finding|Pathologic Function|Impression|4924,4942|false|false|false|C0333575|Fatty infiltration|fatty infiltration
Finding|Functional Concept|Impression|4930,4942|false|false|false|C0332448;C1523986;C3669041|Infiltration;Infiltration Route of Administration;Spread by direct extension|infiltration
Finding|Pathologic Function|Impression|4930,4942|false|false|false|C0332448;C1523986;C3669041|Infiltration;Infiltration Route of Administration;Spread by direct extension|infiltration
Procedure|Therapeutic or Preventive Procedure|Impression|4930,4942|false|false|false|C0702249|Infiltration (procedure)|infiltration
Anatomy|Body Part, Organ, or Organ Component|Impression|4960,4965|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|Impression|4960,4965|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|Impression|4960,4965|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|Impression|4960,4965|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|Impression|4960,4965|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|Impression|4960,4965|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Finding|Finding|Impression|4960,4965|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|Impression|4960,4965|false|false|false|C0872387|Procedures on liver|liver
Disorder|Disease or Syndrome|Impression|4960,4973|false|false|false|C0023895;C0267792|Hepatobiliary Disorder;Liver diseases|liver disease
Disorder|Disease or Syndrome|Impression|4966,4973|false|false|false|C0012634|Disease|disease
Anatomy|Body Part, Organ, or Organ Component|Impression|4992,4997|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|Impression|4992,4997|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|Impression|4992,4997|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|Impression|4992,4997|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|Impression|4992,4997|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|Impression|4992,4997|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Finding|Finding|Impression|4992,4997|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|Impression|4992,4997|false|false|false|C0872387|Procedures on liver|liver
Disorder|Disease or Syndrome|Impression|4992,5005|false|true|false|C0023895;C0267792|Hepatobiliary Disorder;Liver diseases|liver disease
Disorder|Disease or Syndrome|Impression|4998,5005|false|true|false|C0012634|Disease|disease
Finding|Pathologic Function|Impression|5017,5025|false|false|false|C0016059|Fibrosis|fibrosis
Disorder|Disease or Syndrome|Impression|5030,5039|false|false|false|C0023890;C1623038|Cirrhosis;Liver Cirrhosis|cirrhosis
Anatomy|Body Part, Organ, or Organ Component|Impression|5064,5072|false|false|false|C0934502|anatomical layer|Layering
Finding|Body Substance|Impression|5073,5079|false|false|false|C0750852|Physiological sludge|sludge
Phenomenon|Environmental Effect of Humans|Impression|5073,5079|false|false|false|C0282346|Environmental sludge|sludge
Anatomy|Body Part, Organ, or Organ Component|Impression|5091,5102|false|false|false|C0016976;C1524055;C4071903|Abdomen>Gallbladder;Gallbladder;Gallbladder (MMHCC)|gallbladder
Anatomy|Tissue|Impression|5091,5102|false|false|false|C0016976;C1524055;C4071903|Abdomen>Gallbladder;Gallbladder;Gallbladder (MMHCC)|gallbladder
Procedure|Health Care Activity|Impression|5091,5102|false|false|false|C2032932|examination of gallbladder|gallbladder
Finding|Intellectual Product|Impression|5109,5113|false|false|false|C1547225|Mild Severity of Illness Code|mild
Anatomy|Body Part, Organ, or Organ Component|Impression|5114,5125|false|false|false|C0016976;C1524055;C4071903|Abdomen>Gallbladder;Gallbladder;Gallbladder (MMHCC)|gallbladder
Anatomy|Tissue|Impression|5114,5125|false|false|false|C0016976;C1524055;C4071903|Abdomen>Gallbladder;Gallbladder;Gallbladder (MMHCC)|gallbladder
Procedure|Health Care Activity|Impression|5114,5125|false|false|false|C2032932|examination of gallbladder|gallbladder
Finding|Finding|Impression|5133,5143|false|false|false|C0205400|Thickened|thickening
Anatomy|Body Part, Organ, or Organ Component|Impression|5176,5181|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|Impression|5176,5181|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|Impression|5176,5181|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|Impression|5176,5181|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|Impression|5176,5181|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|Impression|5176,5181|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Finding|Finding|Impression|5176,5181|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|Impression|5176,5181|false|false|false|C0872387|Procedures on liver|liver
Disorder|Disease or Syndrome|Impression|5176,5189|false|false|false|C0023895;C0267792|Hepatobiliary Disorder;Liver diseases|liver disease
Disorder|Disease or Syndrome|Impression|5182,5189|false|false|false|C0012634|Disease|disease
Finding|Intellectual Product|Impression|5196,5202|false|false|false|C0030650|Legal patent|Patent
Anatomy|Body Location or Region|Impression|5203,5209|false|false|false|C0205054|Hepatic|portal
Anatomy|Body System|Impression|5203,5223|false|false|false|C0226727|Portal Venous System|portal venous system
Anatomy|Body Part, Organ, or Organ Component|Impression|5210,5216|false|false|false|C0042449|Veins|venous
Anatomy|Body System|Impression|5210,5223|false|false|false|C1267406|Venous system|venous system
Drug|Biomedical or Dental Material|Impression|5217,5223|false|false|false|C5671121|System (basic dose form)|system
Finding|Functional Concept|Impression|5217,5223|false|false|false|C0449913;C5441654|System;System, LOINC Axis 4|system
Finding|Finding|Impression|5229,5237|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Intellectual Product|Impression|5229,5237|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Disorder|Disease or Syndrome|Impression|5238,5245|false|false|false|C0003962|Ascites|ascites
Finding|Pathologic Function|Impression|5238,5245|false|false|false|C5441966|Peritoneal Effusion|ascites
Finding|Intellectual Product|Impression|5252,5257|false|false|false|C1705923|Study Object|study
Procedure|Research Activity|Impression|5252,5257|false|false|false|C0008972;C0947630;C2603343|Clinical Research;Scientific Study;Study|study
Attribute|Clinical Attribute|Impression|5266,5272|false|false|false|C4255046||report
Finding|Intellectual Product|Impression|5266,5272|false|false|false|C0684224|Report (document)|report
Procedure|Health Care Activity|Impression|5266,5272|false|false|false|C0700287|Reporting|report
Finding|Finding|Impression|5294,5299|false|false|false|C1551040|Encounter Special Courtesy - staff|staff
Finding|Intellectual Product|Impression|5300,5311|false|false|false|C1549438|Procedure Practitioner Identifier Code Type - Radiologist|radiologist
Attribute|Clinical Attribute|Impression|5316,5322|false|false|false|C1644645||CT abd
Anatomy|Body Location or Region|Impression|5319,5322|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|abd
Disorder|Cell or Molecular Dysfunction|Impression|5319,5322|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|abd
Anatomy|Body Part, Organ, or Organ Component|Impression|5323,5329|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Anatomy|Body Space or Junction|Impression|5323,5329|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Disorder|Neoplastic Process|Impression|5323,5329|false|false|false|C0153663|Malignant neoplasm of pelvis|pelvis
Finding|Finding|Impression|5323,5329|false|false|false|C0812455|Pelvis problem|pelvis
Finding|Gene or Genome|Impression|5350,5355|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|Large
Finding|Intellectual Product|Impression|5356,5362|false|false|false|C1705102|Volume (publication)|volume
Disorder|Disease or Syndrome|Impression|5363,5370|false|false|false|C0003962|Ascites|ascites
Finding|Pathologic Function|Impression|5363,5370|false|false|false|C5441966|Peritoneal Effusion|ascites
Procedure|Therapeutic or Preventive Procedure|Impression|5375,5383|false|false|false|C1293134|Enlargement procedure|enlarged
Finding|Pathologic Function|Impression|5384,5393|false|false|false|C0013604|Edema|edematous
Anatomy|Body Part, Organ, or Organ Component|Impression|5394,5399|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|Impression|5394,5399|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|Impression|5394,5399|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|Impression|5394,5399|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|Impression|5394,5399|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|Impression|5394,5399|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Finding|Finding|Impression|5394,5399|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|Impression|5394,5399|false|false|false|C0872387|Procedures on liver|liver
Finding|Functional Concept|Findings|5420,5430|false|false|false|C0332299|Suggestive of|suggestive
Finding|Functional Concept|Findings|5420,5433|false|false|false|C0332299|Suggestive of|suggestive of
Finding|Intellectual Product|Findings|5434,5439|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Disorder|Disease or Syndrome|Findings|5434,5449|false|false|false|C0267797|Acute hepatitis|acute hepatitis
Disorder|Disease or Syndrome|Findings|5440,5449|false|false|false|C0019158;C0019159|Hepatitis;Hepatitis A|hepatitis
Anatomy|Tissue|Findings|5472,5479|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|Findings|5472,5479|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Pathologic Function|Findings|5472,5489|false|false|false|C0032227|Pleural effusion (disorder)|pleural effusions
Finding|Pathologic Function|Findings|5480,5489|false|false|false|C0013687|effusion|effusions
Procedure|Health Care Activity|Findings|5492,5496|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Procedure|Therapeutic or Preventive Procedure|Findings|5492,5496|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Finding|Functional Concept|Findings|5506,5510|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Findings|5506,5517|false|false|false|C0225860|Left atrial structure|left atrium
Anatomy|Body Part, Organ, or Organ Component|Findings|5511,5517|false|false|false|C0018792|Heart Atrium|atrium
Finding|Functional Concept|Findings|5522,5527|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|Findings|5522,5534|false|false|false|C0225844|Right atrial structure|right atrium
Anatomy|Body Part, Organ, or Organ Component|Findings|5528,5534|false|false|false|C0018792|Heart Atrium|atrium
Anatomy|Body Space or Junction|Findings|5549,5555|false|false|false|C0333343|Body cavities|cavity
Disorder|Anatomical Abnormality|Findings|5549,5555|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Disorder|Disease or Syndrome|Findings|5549,5555|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Finding|Functional Concept|Findings|5562,5566|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|Findings|5568,5579|false|false|false|C0018827|Heart Ventricle|ventricular
Anatomy|Body Part, Organ, or Organ Component|Findings|5568,5584|false|false|false|C0507618|Wall of ventricle|ventricular wall
Finding|Finding|Findings|5568,5594|false|false|false|C2024242|cardiac evaluation of ventricular wall thickness|ventricular wall thickness
Anatomy|Body Space or Junction|Findings|5596,5602|false|false|false|C0333343|Body cavities|cavity
Disorder|Anatomical Abnormality|Findings|5596,5602|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Disorder|Disease or Syndrome|Findings|5596,5602|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Finding|Organ or Tissue Function|Findings|5629,5637|false|false|false|C0039155|Systole|systolic
Finding|Finding|Findings|5638,5646|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|Findings|5638,5646|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|Findings|5638,5646|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|Findings|5638,5646|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Attribute|Clinical Attribute|Findings|5659,5663|false|false|false|C0428772|Left ventricular ejection fraction|LVEF
Procedure|Diagnostic Procedure|Findings|5659,5663|false|false|false|C3837267|LVEF (procedure)|LVEF
Anatomy|Tissue|Findings|5687,5693|false|false|false|C0040300|Body tissue|tissue
Finding|Intellectual Product|Findings|5687,5693|false|false|false|C1547928|Tissue Specimen Code|tissue
Procedure|Diagnostic Procedure|Findings|5695,5702|false|false|false|C0554756|Doppler studies|Doppler
Finding|Finding|Findings|5703,5710|false|false|false|C0740845|Imaging problem|imaging
Procedure|Diagnostic Procedure|Findings|5703,5710|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|imaging
Attribute|Clinical Attribute|Findings|5727,5736|false|false|false|C0012000|Diastole|diastolic
Finding|Finding|Findings|5737,5745|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|Findings|5737,5745|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|Findings|5737,5745|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|Findings|5737,5745|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|Findings|5761,5765|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Findings|5766,5777|false|false|false|C0018827|Heart Ventricle|ventricular
Finding|Finding|Findings|5786,5794|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|Findings|5786,5794|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|Findings|5786,5794|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|Findings|5786,5794|false|false|false|C0033095||pressure
Attribute|Clinical Attribute|Findings|5796,5800|false|false|false|C0034094|Pulmonary Wedge Pressure|PCWP
Anatomy|Body Part, Organ, or Organ Component|Findings|5823,5834|false|false|false|C0018827|Heart Ventricle|ventricular
Disorder|Congenital Abnormality|Findings|5823,5848|false|false|false|C0018818|Ventricular Septal Defects|ventricular septal defect
Disorder|Anatomical Abnormality|Findings|5835,5848|false|false|false|C0018816;C5779791|Congenital septal defect of heart;Heart Septal Defects|septal defect
Disorder|Congenital Abnormality|Findings|5835,5848|false|false|false|C0018816;C5779791|Congenital septal defect of heart;Heart Septal Defects|septal defect
Disorder|Disease or Syndrome|Findings|5842,5848|false|false|false|C1861101|THYROID HORMONE PLASMA MEMBRANE TRANSPORT DEFECT|defect
Finding|Functional Concept|Findings|5842,5848|false|false|false|C1457869|Defect|defect
Finding|Functional Concept|Findings|5850,5855|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Anatomy|Body Part, Organ, or Organ Component|Findings|5856,5867|false|false|false|C0018827|Heart Ventricle|ventricular
Anatomy|Body Part, Organ, or Organ Component|Findings|5868,5875|false|false|false|C0935616|chamber [body part]|chamber
Finding|Functional Concept|Findings|5886,5890|false|false|false|C0332296|Free of (attribute)|free
Attribute|Clinical Attribute|Findings|5891,5902|false|false|false|C1980023|Wall motion|wall motion
Phenomenon|Natural Phenomenon or Process|Findings|5896,5902|false|false|false|C0026597|Motion|motion
Anatomy|Body Part, Organ, or Organ Component|Findings|5932,5937|false|false|false|C0003483;C4037978|Aorta;Chest+Abdomen>Aorta|aorta
Procedure|Health Care Activity|Findings|5932,5937|false|false|false|C0869784|Procedure on aorta|aorta
Anatomy|Body Space or Junction|Findings|5946,5951|false|false|false|C0030471;C1305231|Nasal sinus;Sinus - general anatomical term|sinus
Disorder|Anatomical Abnormality|Findings|5946,5951|false|false|false|C0016169|pathologic fistula|sinus
Drug|Organic Chemical|Findings|5946,5951|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Drug|Pharmacologic Substance|Findings|5946,5951|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Finding|Functional Concept|Findings|5953,5962|false|false|false|C1547175;C1962987|Ascend (action);Sequencing - Ascending|ascending
Anatomy|Body Location or Region|Findings|5967,5971|false|false|false|C0003741;C0230467;C0741204|ARCH;Arch of foot;Structure of nucleus infundibularis hypothalami|arch
Anatomy|Body Part, Organ, or Organ Component|Findings|5967,5971|false|false|false|C0003741;C0230467;C0741204|ARCH;Arch of foot;Structure of nucleus infundibularis hypothalami|arch
Anatomy|Body Space or Junction|Findings|5967,5971|false|false|false|C0003741;C0230467;C0741204|ARCH;Arch of foot;Structure of nucleus infundibularis hypothalami|arch
Finding|Finding|Findings|5967,5971|false|false|false|C1538146;C4722404|Age-Related Clonal Hematopoiesis;ZBTB8OS gene|arch
Finding|Gene or Genome|Findings|5967,5971|false|false|false|C1538146;C4722404|Age-Related Clonal Hematopoiesis;ZBTB8OS gene|arch
Anatomy|Body Part, Organ, or Organ Component|Findings|5995,6001|false|false|false|C0003483|Aorta|aortic
Anatomy|Body Part, Organ, or Organ Component|Findings|5995,6007|false|false|false|C0003501;C4533215|Aortic valve structure;Chest>Aortic valve|aortic valve
Anatomy|Body Part, Organ, or Organ Component|Findings|6002,6007|false|false|false|C1186983|Anatomical valve|valve
Finding|Idea or Concept|Findings|6054,6058|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Finding|Intellectual Product|Findings|6059,6066|false|false|false|C3273178|Leaflet|leaflet
Anatomy|Body Part, Organ, or Organ Component|Findings|6085,6091|false|false|false|C0003483|Aorta|aortic
Disorder|Disease or Syndrome|Findings|6085,6105|true|false|false|C0003504|Aortic Valve Insufficiency|aortic regurgitation
Finding|Finding|Findings|6092,6105|true|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|Findings|6092,6105|true|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|Findings|6092,6105|true|false|false|C0460152|Regurgitation - mechanism|regurgitation
Anatomy|Body Part, Organ, or Organ Component|Findings|6111,6123|false|false|false|C0026264|Mitral Valve|mitral valve
Anatomy|Body Part, Organ, or Organ Component|Findings|6118,6123|false|false|false|C1186983|Anatomical valve|valve
Disorder|Disease or Syndrome|Findings|6166,6186|false|false|false|C0026266|Mitral Valve Insufficiency|mitral regurgitation
Finding|Finding|Findings|6173,6186|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|Findings|6173,6186|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|Findings|6173,6186|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Anatomy|Body Part, Organ, or Organ Component|Findings|6201,6213|false|false|false|C0026264|Mitral Valve|mitral valve
Disorder|Disease or Syndrome|Findings|6201,6222|true|false|false|C0026267|Mitral Valve Prolapse Syndrome|mitral valve prolapse
Anatomy|Body Part, Organ, or Organ Component|Findings|6208,6213|false|false|false|C1186983|Anatomical valve|valve
Disorder|Disease or Syndrome|Findings|6214,6222|true|false|false|C0033377|Ptosis|prolapse
Anatomy|Body Location or Region|Findings|6236,6247|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Anatomy|Body Part, Organ, or Organ Component|Findings|6236,6247|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Disorder|Disease or Syndrome|Findings|6236,6256|true|false|false|C0031039|Pericardial effusion|pericardial effusion
Finding|Body Substance|Findings|6236,6256|true|false|false|C1253937|Pericardial effusion body substance|pericardial effusion
Finding|Body Substance|Findings|6248,6256|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|Findings|6248,6256|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|Findings|6248,6256|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|Findings|6260,6270|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|Findings|6260,6270|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Organ or Tissue Function|Findings|6313,6321|false|false|false|C0039155|Systole|systolic
Finding|Finding|Findings|6323,6331|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|Findings|6323,6331|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|Findings|6323,6331|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|Findings|6323,6331|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Attribute|Clinical Attribute|Findings|6336,6345|false|false|false|C0012000|Diastole|diastolic
Finding|Pathologic Function|Findings|6336,6357|true|false|false|C0520863|Diastolic dysfunction|diastolic dysfunction
Disorder|Disease or Syndrome|Findings|6346,6357|true|false|false|C3887505|DYSFUNCTION - SKIN DISORDERS|dysfunction
Finding|Conceptual Entity|Findings|6346,6357|true|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Functional Concept|Findings|6346,6357|true|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Pathologic Function|Findings|6346,6357|true|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Anatomy|Body Part, Organ, or Organ Component|Findings|6359,6368|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Findings|6359,6368|false|false|false|C2707265||pulmonary
Finding|Finding|Findings|6359,6368|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|Findings|6359,6381|true|false|false|C0020542|Pulmonary Hypertension|pulmonary hypertension
Disorder|Disease or Syndrome|Findings|6369,6381|true|false|false|C0020538|Hypertensive disease|hypertension
Finding|Functional Concept|Findings|6386,6396|false|false|false|C1521733|Pathologic|pathologic
Disorder|Disease or Syndrome|Findings|6397,6413|false|false|false|C3258293|Valvular disease|valvular disease
Disorder|Disease or Syndrome|Findings|6406,6413|false|false|false|C0012634|Disease|disease
Finding|Conceptual Entity|Hospital Course|6470,6477|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|6470,6477|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Hospital Course|6470,6477|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|6470,6480|false|false|false|C0262926|Medical History|history of
Drug|Organic Chemical|Hospital Course|6481,6485|false|false|false|C0001962|ethanol|EtOH
Drug|Pharmacologic Substance|Hospital Course|6481,6485|false|false|false|C0001962|ethanol|EtOH
Disorder|Disease or Syndrome|Hospital Course|6507,6512|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Finding|Hospital Course|6519,6522|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Hospital Course|6519,6522|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Finding|Hospital Course|6519,6528|false|false|false|C0746890|new onset|new onset
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6529,6534|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|Hospital Course|6529,6534|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|Hospital Course|6529,6534|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|Hospital Course|6529,6534|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|Hospital Course|6529,6534|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|Hospital Course|6529,6534|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Finding|Finding|Hospital Course|6529,6534|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|Hospital Course|6529,6534|false|false|false|C0872387|Procedures on liver|liver
Disorder|Disease or Syndrome|Hospital Course|6529,6542|false|false|false|C0085605|Liver Failure|liver failure
Finding|Functional Concept|Hospital Course|6535,6542|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|Hospital Course|6535,6542|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|Hospital Course|6535,6542|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Disorder|Disease or Syndrome|Hospital Course|6547,6554|false|false|false|C0003962|Ascites|ascites
Finding|Pathologic Function|Hospital Course|6547,6554|false|false|false|C5441966|Peritoneal Effusion|ascites
Disorder|Disease or Syndrome|Hospital Course|6564,6571|false|false|false|C0003962|Ascites|ASCITES
Finding|Pathologic Function|Hospital Course|6564,6571|false|false|false|C5441966|Peritoneal Effusion|ASCITES
Finding|Finding|Hospital Course|6579,6582|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|New
Finding|Idea or Concept|Hospital Course|6579,6582|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|New
Finding|Finding|Hospital Course|6579,6588|false|false|false|C0746890|new onset|New onset
Disorder|Disease or Syndrome|Hospital Course|6589,6596|false|false|false|C0003962|Ascites|ascites
Finding|Pathologic Function|Hospital Course|6589,6596|false|false|false|C5441966|Peritoneal Effusion|ascites
Lab|Laboratory or Test Result|Hospital Course|6602,6606|false|false|false|C4331276|Serum-Ascites Albumin Gradient|SAAG
Finding|Conceptual Entity|Hospital Course|6607,6617|false|false|false|C1521721|Supportive assistance|supportive
Anatomy|Body Location or Region|Hospital Course|6622,6628|false|false|false|C0205054|Hepatic|portal
Disorder|Disease or Syndrome|Hospital Course|6622,6641|false|false|false|C0020541|Portal Hypertension|portal hypertension
Disorder|Disease or Syndrome|Hospital Course|6629,6641|false|false|false|C0020538|Hypertensive disease|hypertension
Finding|Finding|Hospital Course|6644,6650|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Finding|Idea or Concept|Hospital Course|6644,6650|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Disorder|Disease or Syndrome|Hospital Course|6651,6670|false|true|false|C0019187|Hepatitis, Alcoholic|alcoholic hepatitis
Disorder|Disease or Syndrome|Hospital Course|6651,6683|false|true|false|C2887911|alcoholic hepatitis with ascites|alcoholic hepatitis with ascites
Disorder|Disease or Syndrome|Hospital Course|6661,6670|false|true|false|C0019158;C0019159|Hepatitis;Hepatitis A|hepatitis
Disorder|Disease or Syndrome|Hospital Course|6676,6683|false|false|false|C0003962|Ascites|ascites
Finding|Pathologic Function|Hospital Course|6676,6683|false|false|false|C5441966|Peritoneal Effusion|ascites
Disorder|Disease or Syndrome|Hospital Course|6704,6713|false|false|false|C0023890;C1623038|Cirrhosis;Liver Cirrhosis|cirrhosis
Drug|Organic Chemical|Hospital Course|6716,6724|false|false|false|C0038317|Steroids|Steroids
Drug|Pharmacologic Substance|Hospital Course|6716,6724|false|false|false|C0038317|Steroids|Steroids
Finding|Finding|Hospital Course|6769,6772|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|Hospital Course|6769,6772|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Conceptual Entity|Hospital Course|6786,6792|false|false|false|C1521761;C2827422;C5400797|Factor;Feelings about Genomic Testing Results;Mathematical Factor|factor
Finding|Functional Concept|Hospital Course|6786,6792|false|false|false|C1521761;C2827422;C5400797|Factor;Feelings about Genomic Testing Results;Mathematical Factor|factor
Finding|Intellectual Product|Hospital Course|6786,6792|false|false|false|C1521761;C2827422;C5400797|Factor;Feelings about Genomic Testing Results;Mathematical Factor|factor
Finding|Functional Concept|Hospital Course|6814,6824|false|false|false|C0015127|Etiology aspects|etiologies
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6828,6833|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|Hospital Course|6828,6833|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|Hospital Course|6828,6833|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|Hospital Course|6828,6833|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|Hospital Course|6828,6833|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|Hospital Course|6828,6833|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Finding|Finding|Hospital Course|6828,6833|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|Hospital Course|6828,6833|false|false|false|C0872387|Procedures on liver|liver
Disorder|Disease or Syndrome|Hospital Course|6828,6841|false|false|false|C0023895;C0267792|Hepatobiliary Disorder;Liver diseases|liver disease
Disorder|Disease or Syndrome|Hospital Course|6834,6841|false|false|false|C0012634|Disease|disease
Drug|Biologically Active Substance|Hospital Course|6843,6847|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Element, Ion, or Isotope|Hospital Course|6843,6847|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Pharmacologic Substance|Hospital Course|6843,6847|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Procedure|Laboratory Procedure|Hospital Course|6843,6847|false|false|false|C0337439|Iron measurement|iron
Attribute|Clinical Attribute|Hospital Course|6843,6853|false|false|false|C3870201||iron panel
Procedure|Laboratory Procedure|Hospital Course|6843,6853|false|false|false|C3484182|Iron panel|iron panel
Finding|Idea or Concept|Hospital Course|6848,6853|false|false|false|C0441833|Groups|panel
Finding|Idea or Concept|Hospital Course|6862,6872|true|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|Hospital Course|6862,6877|true|false|false|C0332290|Consistent with|consistent with
Disorder|Disease or Syndrome|Hospital Course|6879,6894|false|false|false|C0018995;C3469186|HEMOCHROMATOSIS, TYPE 1;Hemochromatosis|hemochromatosis
Finding|Gene or Genome|Hospital Course|6879,6894|false|false|false|C1384665|HFE gene|hemochromatosis
Finding|Finding|Hospital Course|6905,6908|false|false|false|C5891060|Against Medical Advice|AMA
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6905,6908|false|false|false|C0279755|cytarabine/melphalan|AMA
Finding|Classification|Hospital Course|6919,6927|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|6919,6927|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|6919,6927|false|false|false|C5237010|Expression Negative|negative
Finding|Functional Concept|Hospital Course|6937,6947|false|false|false|C0443146;C4551524|Autoimmune;Autoimmune reaction|autoimmune
Finding|Pathologic Function|Hospital Course|6937,6947|false|false|false|C0443146;C4551524|Autoimmune;Autoimmune reaction|autoimmune
Finding|Functional Concept|Hospital Course|6948,6954|false|false|false|C0015127;C1314792|Etiology;Etiology aspects|causes
Drug|Organic Chemical|Hospital Course|6966,6971|false|false|false|C5400714|ALPHA (substance)|Alpha
Drug|Pharmacologic Substance|Hospital Course|6966,6971|false|false|false|C5400714|ALPHA (substance)|Alpha
Finding|Intellectual Product|Hospital Course|6966,6971|false|false|false|C0439095|Greek letter alpha (qualifier value)|Alpha
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6966,6985|false|false|false|C0002191;C0795657|alpha 1-antitrypsin;alpha 1-proteinase inhibitor, human|Alpha 1 antitrypsin
Drug|Biologically Active Substance|Hospital Course|6966,6985|false|false|false|C0002191;C0795657|alpha 1-antitrypsin;alpha 1-proteinase inhibitor, human|Alpha 1 antitrypsin
Drug|Immunologic Factor|Hospital Course|6966,6985|false|false|false|C0002191;C0795657|alpha 1-antitrypsin;alpha 1-proteinase inhibitor, human|Alpha 1 antitrypsin
Drug|Pharmacologic Substance|Hospital Course|6966,6985|false|false|false|C0002191;C0795657|alpha 1-antitrypsin;alpha 1-proteinase inhibitor, human|Alpha 1 antitrypsin
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6974,6985|false|false|false|C2713669|SERPINA5 protein, human|antitrypsin
Drug|Biologically Active Substance|Hospital Course|6974,6985|false|false|false|C2713669|SERPINA5 protein, human|antitrypsin
Finding|Gene or Genome|Hospital Course|6974,6985|false|false|false|C1418544|SERPINA1 gene|antitrypsin
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6991,7004|false|false|false|C0007841;C5441691|CP protein, human;Ceruloplasmin|ceruloplasmin
Drug|Enzyme|Hospital Course|6991,7004|false|false|false|C0007841;C5441691|CP protein, human;Ceruloplasmin|ceruloplasmin
Finding|Gene or Genome|Hospital Course|6991,7004|false|false|false|C1151847;C1439306|CP gene;ferroxidase activity|ceruloplasmin
Finding|Molecular Function|Hospital Course|6991,7004|false|false|false|C1151847;C1439306|CP gene;ferroxidase activity|ceruloplasmin
Procedure|Laboratory Procedure|Hospital Course|6991,7004|false|false|false|C0373573|Ceruloplasmin measurement|ceruloplasmin
Finding|Functional Concept|Hospital Course|7019,7024|false|false|false|C0521026|Viral|Viral
Attribute|Clinical Attribute|Hospital Course|7019,7032|false|false|false|C4759974||Viral studies
Procedure|Laboratory Procedure|Hospital Course|7019,7032|false|false|false|C1273421|Viral studies (procedure)|Viral studies
Procedure|Research Activity|Hospital Course|7025,7032|false|false|false|C0947630|Scientific Study|studies
Finding|Organ or Tissue Function|Hospital Course|7038,7046|false|false|false|C0020964;C5234945|Immune response;Immune status|immunity
Finding|Physiologic Function|Hospital Course|7038,7046|false|false|false|C0020964;C5234945|Immune response;Immune status|immunity
Anatomy|Body Location or Region|Hospital Course|7050,7053|false|false|false|C0449198|HEP (body structure)|Hep
Disorder|Disease or Syndrome|Hospital Course|7050,7053|false|false|false|C0162569|Hepatoerythropoietic Porphyria|Hep
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7050,7053|false|false|false|C0540659|EPHB6 protein, human|Hep
Drug|Enzyme|Hospital Course|7050,7053|false|false|false|C0540659|EPHB6 protein, human|Hep
Finding|Gene or Genome|Hospital Course|7050,7053|false|false|false|C0540659;C1414432;C1705569;C2239359;C4723683|DNLZ gene;EPHB6 gene;EPHB6 protein, human;EPHB6 wt Allele, Human;HPSE wt Allele|Hep
Finding|Receptor|Hospital Course|7050,7053|false|false|false|C0540659;C1414432;C1705569;C2239359;C4723683|DNLZ gene;EPHB6 gene;EPHB6 protein, human;EPHB6 wt Allele, Human;HPSE wt Allele|Hep
Disorder|Disease or Syndrome|Hospital Course|7065,7068|false|false|false|C0019682;C0019693|HIV;HIV Infections|HIV
Disorder|Virus|Hospital Course|7065,7068|false|false|false|C0019682;C0019693|HIV;HIV Infections|HIV
Drug|Immunologic Factor|Hospital Course|7065,7068|false|false|false|C0086413|HIV Vaccine|HIV
Drug|Pharmacologic Substance|Hospital Course|7065,7068|false|false|false|C0086413|HIV Vaccine|HIV
Finding|Classification|Hospital Course|7073,7081|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|7073,7081|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|7073,7081|false|false|false|C5237010|Expression Negative|negative
Attribute|Clinical Attribute|Hospital Course|7092,7098|false|false|false|C1644645||CT abd
Anatomy|Body Location or Region|Hospital Course|7095,7098|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|abd
Disorder|Cell or Molecular Dysfunction|Hospital Course|7095,7098|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|abd
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7099,7105|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Anatomy|Body Space or Junction|Hospital Course|7099,7105|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Disorder|Neoplastic Process|Hospital Course|7099,7105|false|false|false|C0153663|Malignant neoplasm of pelvis|pelvis
Finding|Finding|Hospital Course|7099,7105|false|false|false|C0812455|Pelvis problem|pelvis
Finding|Functional Concept|Hospital Course|7116,7126|false|false|false|C0332299|Suggestive of|suggestive
Finding|Functional Concept|Hospital Course|7116,7129|false|false|false|C0332299|Suggestive of|suggestive of
Finding|Finding|Hospital Course|7130,7134|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|Hospital Course|7130,7134|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|Hospital Course|7130,7134|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Functional Concept|Hospital Course|7138,7149|false|false|false|C0549186|Obstructed|obstructive
Finding|Finding|Hospital Course|7150,7157|false|false|false|C0221198|Lesion|lesions
Finding|Body Substance|Hospital Course|7160,7167|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|7160,7167|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|7160,7167|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7185,7197|false|false|false|C0034115|Paracentesis|paracentesis
Finding|Idea or Concept|Hospital Course|7206,7209|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|7206,7209|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Body Substance|Hospital Course|7219,7228|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|7219,7228|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|7219,7228|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|7219,7228|false|false|false|C0030685|Patient Discharge|discharge
Finding|Finding|Hospital Course|7231,7234|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|Low
Finding|Intellectual Product|Hospital Course|7231,7234|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|Low
Procedure|Research Activity|Hospital Course|7231,7239|false|false|false|C1708745|Low-Dose Treatment|Low-dose
Drug|Organic Chemical|Hospital Course|7241,7255|false|false|false|C0037982|spironolactone|spironolactone
Drug|Pharmacologic Substance|Hospital Course|7241,7255|false|false|false|C0037982|spironolactone|spironolactone
Finding|Intellectual Product|Hospital Course|7312,7316|false|false|false|C1561540|Transaction counts and value totals - week|week
Disorder|Mental or Behavioral Dysfunction|Hospital Course|7324,7334|false|false|false|C0001973|Alcoholic Intoxication, Chronic|ALCOHOLISM
Procedure|Health Care Activity|Hospital Course|7340,7349|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Drug|Organic Chemical|Hospital Course|7351,7358|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Drug|Pharmacologic Substance|Hospital Course|7351,7358|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Finding|Intellectual Product|Hospital Course|7351,7358|false|false|false|C1547288|Alcohol - Recreational Drug Use Code|alcohol
Procedure|Laboratory Procedure|Hospital Course|7351,7364|false|false|false|C0202304|Ethanol measurement|alcohol level
Finding|Body Substance|Hospital Course|7381,7388|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|7381,7388|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|7381,7388|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Body Substance|Hospital Course|7412,7419|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|7412,7419|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|7412,7419|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|7439,7443|false|false|false|C0814193|clinical institute withdrawal assessment (CIWA) for alcohol|CIWA
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7445,7450|false|false|false|C0222045|Integumentary scale|scale
Event|Activity|Hospital Course|7445,7450|false|false|false|C1947916|Scaling|scale
Finding|Conceptual Entity|Hospital Course|7445,7450|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|scale
Finding|Intellectual Product|Hospital Course|7445,7450|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|scale
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7468,7471|false|false|false|C5417720|MVI Regimen|MVI
Drug|Organic Chemical|Hospital Course|7473,7481|false|false|false|C0039840;C3714802|Thiamine Drug Class;thiamine|thiamine
Drug|Pharmacologic Substance|Hospital Course|7473,7481|false|false|false|C0039840;C3714802|Thiamine Drug Class;thiamine|thiamine
Drug|Vitamin|Hospital Course|7473,7481|false|false|false|C0039840;C3714802|Thiamine Drug Class;thiamine|thiamine
Procedure|Laboratory Procedure|Hospital Course|7473,7481|false|false|false|C0373727|Thiamine measurement|thiamine
Drug|Organic Chemical|Hospital Course|7487,7493|false|false|false|C0178638|folate|folate
Drug|Pharmacologic Substance|Hospital Course|7487,7493|false|false|false|C0178638|folate|folate
Drug|Vitamin|Hospital Course|7487,7493|false|false|false|C0178638|folate|folate
Procedure|Laboratory Procedure|Hospital Course|7487,7493|false|false|false|C0523631|Folic acid measurement|folate
Finding|Functional Concept|Hospital Course|7513,7519|false|false|false|C0728831|Social|social
Event|Occupational Activity|Hospital Course|7520,7524|false|false|false|C0043227|Work|work
Event|Activity|Hospital Course|7539,7546|false|false|false|C3812666|Personal Contact|contact
Finding|Functional Concept|Hospital Course|7539,7546|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|contact
Finding|Idea or Concept|Hospital Course|7539,7546|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|contact
Finding|Intellectual Product|Hospital Course|7539,7546|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|contact
Phenomenon|Phenomenon or Process|Hospital Course|7539,7546|false|false|false|C0392367|Physical contact|contact
Finding|Conceptual Entity|Hospital Course|7539,7558|false|false|false|C1880174|Contact Information|contact information
Finding|Idea or Concept|Hospital Course|7547,7558|false|false|false|C0870705;C1533716;C1561527;C1561528|Acknowledgement Detail Type - Information;Error severity - Information;Information;control act - information|information
Finding|Intellectual Product|Hospital Course|7547,7558|false|false|false|C0870705;C1533716;C1561527;C1561528|Acknowledgement Detail Type - Information;Error severity - Information;Information;control act - information|information
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7563,7568|false|false|false|C0034991|Rehabilitation therapy|rehab
Finding|Body Substance|Hospital Course|7592,7599|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|7592,7599|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|7592,7599|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7629,7634|false|false|false|C0034991|Rehabilitation therapy|rehab
Finding|Classification|Hospital Course|7664,7674|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|7664,7674|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Procedure|Health Care Activity|Hospital Course|7664,7684|false|false|false|C0002423;C0086751|Ambulatory Care;Health Services, Outpatient|outpatient treatment
Finding|Conceptual Entity|Hospital Course|7675,7684|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|Hospital Course|7675,7684|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|Hospital Course|7675,7684|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7675,7684|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Disorder|Mental or Behavioral Dysfunction|Hospital Course|7694,7703|false|false|false|C0085281|Addictive Behavior|addiction
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7812,7817|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|Hospital Course|7812,7817|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|Hospital Course|7812,7817|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|Hospital Course|7812,7817|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|Hospital Course|7812,7817|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|Hospital Course|7812,7817|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Finding|Finding|Hospital Course|7812,7817|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|Hospital Course|7812,7817|false|false|false|C0872387|Procedures on liver|liver
Finding|Sign or Symptom|Hospital Course|7843,7852|false|false|false|C0004604|Back Pain|BACK PAIN
Attribute|Clinical Attribute|Hospital Course|7848,7852|false|false|false|C2598155||PAIN
Finding|Functional Concept|Hospital Course|7848,7852|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|PAIN
Finding|Sign or Symptom|Hospital Course|7848,7852|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|PAIN
Finding|Body Substance|Hospital Course|7855,7862|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|7855,7862|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|7855,7862|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Organic Chemical|Hospital Course|7880,7889|false|false|false|C0023660|lidocaine|lidocaine
Drug|Pharmacologic Substance|Hospital Course|7880,7889|false|false|false|C0023660|lidocaine|lidocaine
Procedure|Laboratory Procedure|Hospital Course|7880,7889|false|false|false|C0202404|Lidocaine measurement|lidocaine
Drug|Clinical Drug|Hospital Course|7880,7895|false|false|false|C1251704|Lidocaine Patch|lidocaine patch
Drug|Biomedical or Dental Material|Hospital Course|7890,7895|false|false|false|C0445403;C1533128;C1707974|Body tissue patch material;Human patch material;Patch - Extended Release Film|patch
Finding|Finding|Hospital Course|7890,7895|false|false|false|C0332461|Plaque (lesion)|patch
Drug|Organic Chemical|Hospital Course|7907,7916|false|false|false|C0030049|oxycodone|oxycodone
Drug|Pharmacologic Substance|Hospital Course|7907,7916|false|false|false|C0030049|oxycodone|oxycodone
Procedure|Laboratory Procedure|Hospital Course|7907,7916|false|false|false|C0524222|Oxycodone measurement|oxycodone
Finding|Sign or Symptom|Hospital Course|7921,7938|false|false|false|C1135120|Breakthrough Pain|breakthrough pain
Attribute|Clinical Attribute|Hospital Course|7934,7938|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|7934,7938|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|7934,7938|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Idea or Concept|Hospital Course|7952,7960|false|false|false|C1547192|Organization unit type - Hospital|hospital
Disorder|Disease or Syndrome|Hospital Course|7968,7980|false|false|false|C0023518|Leukocytosis|LEUKOCYTOSIS
Finding|Finding|Hospital Course|7968,7980|false|false|false|C0750426|Blood leukocyte number above reference range|LEUKOCYTOSIS
Finding|Finding|Hospital Course|7992,8003|false|true|false|C3811910|combination - answer to question|combination
Disorder|Disease or Syndrome|Hospital Course|8007,8026|false|false|false|C0019187|Hepatitis, Alcoholic|alcoholic hepatitis
Disorder|Disease or Syndrome|Hospital Course|8017,8026|false|false|false|C0019158;C0019159|Hepatitis;Hepatitis A|hepatitis
Disorder|Disease or Syndrome|Hospital Course|8032,8035|false|false|false|C0042029|Urinary tract infection|UTI
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8032,8035|false|false|false|C0077906|urinastatin|UTI
Drug|Pharmacologic Substance|Hospital Course|8032,8035|false|false|false|C0077906|urinastatin|UTI
Finding|Gene or Genome|Hospital Course|8032,8035|false|false|false|C1412376;C5780748|AMBP gene;AMBP wt Allele|UTI
Finding|Body Substance|Hospital Course|8037,8044|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|8037,8044|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|8037,8044|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Organic Chemical|Hospital Course|8060,8073|false|false|false|C0008809|ciprofloxacin|ciprofloxacin
Drug|Pharmacologic Substance|Hospital Course|8060,8073|false|false|false|C0008809|ciprofloxacin|ciprofloxacin
Disorder|Disease or Syndrome|Hospital Course|8082,8092|false|false|false|C0009450|Communicable Diseases|infectious
Event|Occupational Activity|Hospital Course|8094,8098|false|false|false|C0043227|Work|work
Procedure|Diagnostic Procedure|Hospital Course|8094,8101|false|false|false|C0750430|Work-up|work-up
Finding|Idea or Concept|Hospital Course|8123,8126|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|8123,8126|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Body Substance|Hospital Course|8136,8145|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|8136,8145|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|8136,8145|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|8136,8145|false|false|false|C0030685|Patient Discharge|discharge
Procedure|Health Care Activity|Hospital Course|8136,8154|false|false|false|C0030685|Patient Discharge|discharge, patient
Finding|Body Substance|Hospital Course|8147,8154|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|8147,8154|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|8147,8154|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Finding|Hospital Course|8165,8170|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|Hospital Course|8165,8170|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Anatomy|Cell Component|Hospital Course|8186,8189|false|false|false|C2244316|proteasome-activating nucleotidase complex|pan
Disorder|Disease or Syndrome|Hospital Course|8186,8189|false|false|false|C0031036|Polyarteritis Nodosa|pan
Finding|Gene or Genome|Hospital Course|8186,8189|false|false|false|C5401218|ADA2 wt Allele|pan
Procedure|Diagnostic Procedure|Hospital Course|8201,8204|false|false|false|C0039985|Plain chest X-ray|CXR
Finding|Body Substance|Hospital Course|8226,8231|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Functional Concept|Hospital Course|8226,8231|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Intellectual Product|Hospital Course|8226,8231|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Classification|Hospital Course|8236,8244|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|8236,8244|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|8236,8244|false|false|false|C5237010|Expression Negative|negative
Finding|Finding|Hospital Course|8236,8248|false|false|false|C0205160|Negative|negative for
Disorder|Disease or Syndrome|Hospital Course|8249,8258|false|false|false|C0009450|Communicable Diseases|infection
Finding|Pathologic Function|Hospital Course|8249,8258|false|false|false|C3714514|Infection|infection
Drug|Organic Chemical|Hospital Course|8269,8274|false|false|false|C0701042|Cipro|Cipro
Drug|Pharmacologic Substance|Hospital Course|8269,8274|false|false|false|C0701042|Cipro|Cipro
Drug|Antibiotic|Hospital Course|8304,8316|false|false|false|C0282386|levofloxacin|levofloxacin
Drug|Organic Chemical|Hospital Course|8304,8316|false|false|false|C0282386|levofloxacin|levofloxacin
Finding|Idea or Concept|Hospital Course|8325,8328|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|8325,8328|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Finding|Hospital Course|8343,8353|false|false|false|C0302845|Mean corpuscular volume above reference range|MACROCYTIC
Disorder|Disease or Syndrome|Hospital Course|8343,8360|false|false|false|C0002886|Anemia, Macrocytic|MACROCYTIC ANEMIA
Finding|Gene or Genome|Hospital Course|8343,8360|false|false|false|C1420653|TCN2 gene|MACROCYTIC ANEMIA
Disorder|Disease or Syndrome|Hospital Course|8354,8360|false|false|false|C0002871|Anemia|ANEMIA
Finding|Finding|Hospital Course|8363,8369|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Finding|Idea or Concept|Hospital Course|8363,8369|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Drug|Organic Chemical|Hospital Course|8375,8381|false|false|false|C0178638|folate|folate
Drug|Pharmacologic Substance|Hospital Course|8375,8381|false|false|false|C0178638|folate|folate
Drug|Vitamin|Hospital Course|8375,8381|false|false|false|C0178638|folate|folate
Procedure|Laboratory Procedure|Hospital Course|8375,8381|false|false|false|C0523631|Folic acid measurement|folate
Attribute|Clinical Attribute|Hospital Course|8386,8397|false|false|false|C2707262||nutritional
Disorder|Disease or Syndrome|Hospital Course|8399,8409|false|true|false|C0162429|Malnutrition|deficiency
Finding|Functional Concept|Hospital Course|8399,8409|false|true|false|C0011155|Deficiency|deficiency
Finding|Mental Process|Hospital Course|8413,8420|false|false|false|C0542559|contextual factors|setting
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8424,8434|false|false|false|C0001973|Alcoholic Intoxication, Chronic|alcoholism
Finding|Body Substance|Hospital Course|8437,8444|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|8437,8444|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|8437,8444|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Organic Chemical|Hospital Course|8465,8473|false|false|false|C0039840;C3714802|Thiamine Drug Class;thiamine|thiamine
Drug|Pharmacologic Substance|Hospital Course|8465,8473|false|false|false|C0039840;C3714802|Thiamine Drug Class;thiamine|thiamine
Drug|Vitamin|Hospital Course|8465,8473|false|false|false|C0039840;C3714802|Thiamine Drug Class;thiamine|thiamine
Procedure|Laboratory Procedure|Hospital Course|8465,8473|false|false|false|C0373727|Thiamine measurement|thiamine
Drug|Organic Chemical|Hospital Course|8479,8485|false|false|false|C0178638|folate|folate
Drug|Pharmacologic Substance|Hospital Course|8479,8485|false|false|false|C0178638|folate|folate
Drug|Vitamin|Hospital Course|8479,8485|false|false|false|C0178638|folate|folate
Procedure|Laboratory Procedure|Hospital Course|8479,8485|false|false|false|C0523631|Folic acid measurement|folate
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8479,8501|false|false|false|C4551652|Folate supplementation|folate supplementation
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8486,8501|false|false|false|C0242297|Dietary Supplementation|supplementation
Procedure|Laboratory Procedure|Hospital Course|8504,8507|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8504,8507|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Procedure|Health Care Activity|Hospital Course|8534,8543|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8549,8556|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|ANXIETY
Finding|Sign or Symptom|Hospital Course|8549,8556|false|false|false|C0860603|Anxiety symptoms|ANXIETY
Finding|Body Substance|Hospital Course|8559,8566|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|8559,8566|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|8559,8566|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8579,8586|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Finding|Sign or Symptom|Hospital Course|8579,8586|false|false|false|C0860603|Anxiety symptoms|anxiety
Finding|Finding|Hospital Course|8599,8605|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Hospital Course|8599,8605|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Classification|Hospital Course|8620,8630|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|8620,8630|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Finding|Hospital Course|8631,8638|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|Hospital Course|8631,8638|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8631,8638|false|false|false|C0087111|Therapeutic procedure|therapy
Drug|Pharmacologic Substance|Hospital Course|8646,8650|false|false|false|C0360105;C2911696|Selective Serotonin Reuptake Inhibitors;Serotonin Reuptake Inhibitor [EPC]|SSRI
Finding|Conceptual Entity|Hospital Course|8651,8660|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|Hospital Course|8651,8660|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|Hospital Course|8651,8660|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8651,8660|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Anatomy|Body Space or Junction|Hospital Course|8666,8671|false|false|false|C0030471;C1305231|Nasal sinus;Sinus - general anatomical term|SINUS
Disorder|Anatomical Abnormality|Hospital Course|8666,8671|false|false|false|C0016169|pathologic fistula|SINUS
Drug|Organic Chemical|Hospital Course|8666,8671|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|SINUS
Drug|Pharmacologic Substance|Hospital Course|8666,8671|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|SINUS
Disorder|Disease or Syndrome|Hospital Course|8666,8683|false|false|false|C0039239|Sinus Tachycardia|SINUS TACHYCARDIA
Finding|Finding|Hospital Course|8666,8683|false|false|false|C2108109;C5235163|Sinus Tachycardia by ECG Finding;continuous electrocardiogram sinus tachycardia|SINUS TACHYCARDIA
Finding|Finding|Hospital Course|8672,8683|false|false|false|C0039231;C3827868|Tachycardia;Tachycardia by ECG Finding|TACHYCARDIA
Finding|Finding|Hospital Course|8686,8692|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Finding|Idea or Concept|Hospital Course|8686,8692|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Finding|Idea or Concept|Hospital Course|8696,8703|false|true|false|C0449255;C0542559;C4281677|Application Context;Context;contextual factors|context
Finding|Intellectual Product|Hospital Course|8696,8703|false|true|false|C0449255;C0542559;C4281677|Application Context;Context;contextual factors|context
Finding|Mental Process|Hospital Course|8696,8703|false|true|false|C0449255;C0542559;C4281677|Application Context;Context;contextual factors|context
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8721,8726|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|Hospital Course|8721,8726|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|Hospital Course|8721,8726|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|Hospital Course|8721,8726|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|Hospital Course|8721,8726|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|Hospital Course|8721,8726|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Finding|Finding|Hospital Course|8721,8726|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|Hospital Course|8721,8726|false|false|false|C0872387|Procedures on liver|liver
Disorder|Disease or Syndrome|Hospital Course|8728,8735|false|false|false|C0012634|Disease|disease
Procedure|Health Care Activity|Hospital Course|8738,8742|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8738,8742|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Finding|Finding|Hospital Course|8747,8767|false|false|false|C0442816||within normal limits
Finding|Functional Concept|Hospital Course|8761,8767|false|false|false|C0439801|Limited (extensiveness)|limits
Finding|Body Substance|Hospital Course|8770,8777|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|8770,8777|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|8770,8777|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Procedure|Diagnostic Procedure|Hospital Course|8795,8804|false|false|false|C0039451|Telemetry|telemetry
Procedure|Health Care Activity|Hospital Course|8816,8831|false|false|false|C0019993|Hospitalization|hospitalization
Finding|Sign or Symptom|Hospital Course|8837,8849|false|false|false|C0009806|Constipation|CONSTIPATION
Finding|Body Substance|Hospital Course|8852,8859|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|8852,8859|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|8852,8859|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Organic Chemical|Hospital Course|8878,8883|false|false|false|C3489575|sennosides, USP|senna
Drug|Pharmacologic Substance|Hospital Course|8878,8883|false|false|false|C3489575|sennosides, USP|senna
Drug|Organic Chemical|Hospital Course|8888,8894|false|false|false|C0282139|Colace|colace
Drug|Pharmacologic Substance|Hospital Course|8888,8894|false|false|false|C0282139|Colace|colace
Attribute|Clinical Attribute|Hospital Course|8898,8909|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|8898,8909|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|Hospital Course|8898,8909|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|8898,8922|false|false|false|C1627937|Medications on admission|Medications on Admission
Procedure|Health Care Activity|Hospital Course|8913,8922|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Finding|Body Substance|Hospital Course|8932,8941|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|8932,8941|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|8932,8941|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|8932,8941|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|8932,8953|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|8942,8953|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|8942,8953|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|Hospital Course|8942,8953|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Hospital Course|8958,8970|false|false|false|C0301532|Multivitamin preparation|Multivitamin
Drug|Pharmacologic Substance|Hospital Course|8958,8970|false|false|false|C0301532|Multivitamin preparation|Multivitamin
Drug|Vitamin|Hospital Course|8958,8970|false|false|false|C0301532|Multivitamin preparation|Multivitamin
Drug|Pharmacologic Substance|Hospital Course|8958,8981|false|false|false|C0978787|Multivitamin tablet|Multivitamin     Tablet
Drug|Biomedical or Dental Material|Hospital Course|8975,8981|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|8995,9001|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|9029,9035|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|Hospital Course|9040,9047|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|9055,9065|false|false|false|C0016410|folic acid|Folic Acid
Drug|Pharmacologic Substance|Hospital Course|9055,9065|false|false|false|C0016410|folic acid|Folic Acid
Drug|Vitamin|Hospital Course|9055,9065|false|false|false|C0016410|folic acid|Folic Acid
Procedure|Laboratory Procedure|Hospital Course|9055,9065|false|false|false|C0523631|Folic acid measurement|Folic Acid
Drug|Biomedical or Dental Material|Hospital Course|9071,9077|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|9091,9097|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|9125,9131|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|Hospital Course|9136,9143|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|9151,9159|false|false|false|C0039840;C3714802|Thiamine Drug Class;thiamine|Thiamine
Drug|Pharmacologic Substance|Hospital Course|9151,9159|false|false|false|C0039840;C3714802|Thiamine Drug Class;thiamine|Thiamine
Drug|Vitamin|Hospital Course|9151,9159|false|false|false|C0039840;C3714802|Thiamine Drug Class;thiamine|Thiamine
Procedure|Laboratory Procedure|Hospital Course|9151,9159|false|false|false|C0373727|Thiamine measurement|Thiamine
Drug|Organic Chemical|Hospital Course|9151,9163|false|false|false|C0770309|thiamine hydrochloride|Thiamine HCl
Drug|Pharmacologic Substance|Hospital Course|9151,9163|false|false|false|C0770309|thiamine hydrochloride|Thiamine HCl
Drug|Vitamin|Hospital Course|9151,9163|false|false|false|C0770309|thiamine hydrochloride|Thiamine HCl
Disorder|Neoplastic Process|Hospital Course|9160,9163|false|false|false|C0023443|Hairy Cell Leukemia|HCl
Drug|Immunologic Factor|Hospital Course|9160,9163|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Inorganic Chemical|Hospital Course|9160,9163|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Pharmacologic Substance|Hospital Course|9160,9163|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Biomedical or Dental Material|Hospital Course|9171,9177|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|9191,9197|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|9226,9232|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|Hospital Course|9237,9244|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|9252,9261|false|false|false|C0023660|lidocaine|Lidocaine
Drug|Pharmacologic Substance|Hospital Course|9252,9261|false|false|false|C0023660|lidocaine|Lidocaine
Procedure|Laboratory Procedure|Hospital Course|9252,9261|false|false|false|C0202404|Lidocaine measurement|Lidocaine
Drug|Biomedical or Dental Material|Hospital Course|9273,9278|false|false|false|C0445403;C1533128;C1707974|Body tissue patch material;Human patch material;Patch - Extended Release Film|patch
Finding|Finding|Hospital Course|9273,9278|false|false|false|C0332461|Plaque (lesion)|patch
Drug|Biomedical or Dental Material|Hospital Course|9289,9294|false|false|false|C0445403;C1533128;C1707974|Body tissue patch material;Human patch material;Patch - Extended Release Film|Patch
Finding|Finding|Hospital Course|9289,9294|false|false|false|C0332461|Plaque (lesion)|Patch
Drug|Pharmacologic Substance|Hospital Course|9296,9305|false|false|false|C3812869|Medicated|Medicated
Finding|Finding|Hospital Course|9296,9305|false|false|false|C3812868|Medicated (finding)|Medicated
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9306,9309|false|false|false|C0262329|Short insular gyrus|Sig
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9306,9309|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Drug|Immunologic Factor|Hospital Course|9306,9309|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Finding|Receptor|Hospital Course|9306,9309|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Drug|Biomedical or Dental Material|Hospital Course|9329,9334|false|false|false|C0445403;C1533128;C1707974|Body tissue patch material;Human patch material;Patch - Extended Release Film|Patch
Finding|Finding|Hospital Course|9329,9334|false|false|false|C0332461|Plaque (lesion)|Patch
Drug|Pharmacologic Substance|Hospital Course|9336,9345|false|false|false|C3812869|Medicated|Medicated
Finding|Finding|Hospital Course|9336,9345|false|false|false|C3812868|Medicated (finding)|Medicated
Drug|Biomedical or Dental Material|Hospital Course|9346,9353|false|false|false|C1710439|Topical Dosage Form|Topical
Finding|Functional Concept|Hospital Course|9346,9353|false|false|false|C1522168|Topical Route of Administration|Topical
Finding|Functional Concept|Hospital Course|9369,9374|false|false|false|C1632850;C1879355;C4048755;C4521676|Apply;Apply (administration method);Apply (instruction)|Apply
Finding|Functional Concept|Hospital Course|9379,9387|false|false|false|C0392760;C1314939|Affecting;Involvement with|affected
Anatomy|Body Location or Region|Hospital Course|9379,9392|false|false|false|C4319771|Affected area of body|affected area
Finding|Finding|Hospital Course|9379,9392|false|false|false|C1879646|Affected Area|affected area
Event|Governmental or Regulatory Activity|Hospital Course|9388,9392|false|false|false|C1510751|Academic Research Enhancement Awards|area
Finding|Intellectual Product|Hospital Course|9393,9397|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Biomedical or Dental Material|Hospital Course|9435,9440|false|false|false|C0445403;C1533128;C1707974|Body tissue patch material;Human patch material;Patch - Extended Release Film|Patch
Finding|Finding|Hospital Course|9435,9440|false|false|false|C0332461|Plaque (lesion)|Patch
Drug|Pharmacologic Substance|Hospital Course|9442,9451|false|false|false|C3812869|Medicated|Medicated
Finding|Finding|Hospital Course|9442,9451|false|false|false|C3812868|Medicated (finding)|Medicated
Finding|Idea or Concept|Hospital Course|9456,9463|false|false|false|C0807726|refill|Refills
Drug|Hazardous or Poisonous Substance|Hospital Course|9471,9479|true|false|false|C0028040|nicotine|Nicotine
Drug|Organic Chemical|Hospital Course|9471,9479|true|false|false|C0028040|nicotine|Nicotine
Drug|Biomedical or Dental Material|Hospital Course|9492,9497|false|false|false|C0445403;C1533128;C1707974|Body tissue patch material;Human patch material;Patch - Extended Release Film|Patch
Finding|Finding|Hospital Course|9492,9497|false|false|false|C0332461|Plaque (lesion)|Patch
Drug|Biomedical or Dental Material|Hospital Course|9517,9522|false|false|false|C0445403;C1533128;C1707974|Body tissue patch material;Human patch material;Patch - Extended Release Film|Patch
Finding|Finding|Hospital Course|9517,9522|false|false|false|C0332461|Plaque (lesion)|Patch
Finding|Finding|Hospital Course|9530,9541|false|false|false|C0040652;C0694643;C4521342|Transdermal (intended site);Transdermal Route of Administration;transdermal|Transdermal
Finding|Functional Concept|Hospital Course|9530,9541|false|false|false|C0040652;C0694643;C4521342|Transdermal (intended site);Transdermal Route of Administration;transdermal|Transdermal
Finding|Intellectual Product|Hospital Course|9563,9567|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Biomedical or Dental Material|Hospital Course|9596,9601|false|false|false|C0445403;C1533128;C1707974|Body tissue patch material;Human patch material;Patch - Extended Release Film|Patch
Finding|Finding|Hospital Course|9596,9601|false|false|false|C0332461|Plaque (lesion)|Patch
Finding|Idea or Concept|Hospital Course|9612,9619|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|9627,9641|false|false|false|C0037982|spironolactone|Spironolactone
Drug|Pharmacologic Substance|Hospital Course|9627,9641|false|false|false|C0037982|spironolactone|Spironolactone
Drug|Biomedical or Dental Material|Hospital Course|9648,9654|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|9668,9674|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Intellectual Product|Hospital Course|9678,9682|false|false|false|C1720092|Once - dosing instruction fragment|once
Finding|Idea or Concept|Hospital Course|9686,9689|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|9686,9689|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Biomedical or Dental Material|Hospital Course|9700,9706|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|Hospital Course|9711,9718|false|false|false|C0807726|refill|Refills
Drug|Antibiotic|Hospital Course|9726,9738|false|false|false|C0282386|levofloxacin|Levofloxacin
Drug|Organic Chemical|Hospital Course|9726,9738|false|false|false|C0282386|levofloxacin|Levofloxacin
Drug|Biomedical or Dental Material|Hospital Course|9746,9752|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|9766,9772|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Intellectual Product|Hospital Course|9776,9780|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|Hospital Course|9776,9786|false|false|false|C3537736|Once A Day|once a day
Finding|Idea or Concept|Hospital Course|9783,9786|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|9783,9786|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Biomedical or Dental Material|Hospital Course|9808,9814|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|Hospital Course|9819,9826|false|false|false|C0807726|refill|Refills
Finding|Classification|Hospital Course|9834,9844|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|Outpatient
Finding|Idea or Concept|Hospital Course|9834,9844|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|Outpatient
Finding|Gene or Genome|Hospital Course|9845,9848|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|Lab
Finding|Intellectual Product|Hospital Course|9845,9848|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|Lab
Event|Occupational Activity|Hospital Course|9849,9853|false|false|false|C0043227|Work|Work
Disorder|Disease or Syndrome|Hospital Course|9866,9871|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|Hospital Course|9866,9871|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Body Substance|Hospital Course|9866,9879|false|false|false|C0178913|Blood specimen|blood samples
Anatomy|Cell Component|Hospital Course|9884,9887|false|false|false|C2263086|Nuclear cap binding complex location|CBC
Procedure|Laboratory Procedure|Hospital Course|9884,9887|false|false|false|C0009555|Complete Blood Count|CBC
Procedure|Laboratory Procedure|Hospital Course|9884,9905|false|false|false|C0545131|complete blood count with differential|CBC with differential
Finding|Idea or Concept|Hospital Course|9893,9905|false|false|false|C1549478|Amount type - Differential|differential
Anatomy|Body Space or Junction|Hospital Course|9907,9910|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|Hospital Course|9907,9910|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9907,9910|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|Hospital Course|9907,9910|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|Hospital Course|9907,9910|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Finding|Gene or Genome|Hospital Course|9907,9910|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Disorder|Neoplastic Process|Hospital Course|9911,9914|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9911,9914|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|Hospital Course|9911,9914|false|false|false|C0001899|Alanine Transaminase|ALT
Finding|Gene or Genome|Hospital Course|9911,9914|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|Hospital Course|9911,9914|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|Hospital Course|9911,9914|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9911,9914|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Drug|Biologically Active Substance|Hospital Course|9917,9932|false|false|false|C0005437|Bilirubin|total bilirubin
Drug|Organic Chemical|Hospital Course|9917,9932|false|false|false|C0005437|Bilirubin|total bilirubin
Finding|Physiologic Function|Hospital Course|9917,9932|false|false|false|C4553024|Total bilirubin metabolic function|total bilirubin
Lab|Laboratory or Test Result|Hospital Course|9917,9932|false|false|false|C0368753|Total bilirubin level|total bilirubin
Procedure|Laboratory Procedure|Hospital Course|9917,9932|false|false|false|C0201913|Bilirubin, total measurement|total bilirubin
Drug|Biologically Active Substance|Hospital Course|9923,9932|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|bilirubin
Drug|Organic Chemical|Hospital Course|9923,9932|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|bilirubin
Drug|Pharmacologic Substance|Hospital Course|9923,9932|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|bilirubin
Procedure|Laboratory Procedure|Hospital Course|9923,9932|false|false|false|C0201913;C0863174|Bilirubin, total measurement;blood bilirubin level test|bilirubin
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9934,9954|false|false|false|C0002059|Alkaline Phosphatase|alkaline phosphatase
Drug|Enzyme|Hospital Course|9934,9954|false|false|false|C0002059|Alkaline Phosphatase|alkaline phosphatase
Finding|Physiologic Function|Hospital Course|9934,9954|false|false|false|C4553029|Alkaline phosphatase metabolic function|alkaline phosphatase
Procedure|Laboratory Procedure|Hospital Course|9934,9954|false|false|false|C0201850|Alkaline phosphatase measurement|alkaline phosphatase
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9943,9954|false|false|false|C0031678|Phosphoric Monoester Hydrolases|phosphatase
Drug|Enzyme|Hospital Course|9943,9954|false|false|false|C0031678|Phosphoric Monoester Hydrolases|phosphatase
Finding|Molecular Function|Hospital Course|9943,9954|false|false|false|C1149880|phosphoric monoester hydrolase activity|phosphatase
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9956,9963|false|false|false|C0001924;C5966160|Albumin;Albumins|albumin
Drug|Biologically Active Substance|Hospital Course|9956,9963|false|false|false|C0001924;C5966160|Albumin;Albumins|albumin
Drug|Pharmacologic Substance|Hospital Course|9956,9963|false|false|false|C0001924;C5966160|Albumin;Albumins|albumin
Finding|Gene or Genome|Hospital Course|9956,9963|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|albumin
Finding|Physiologic Function|Hospital Course|9956,9963|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|albumin
Procedure|Laboratory Procedure|Hospital Course|9956,9963|false|false|false|C0201838|Albumin measurement|albumin
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9965,9968|false|false|false|C0022917|Lactate Dehydrogenase|LDH
Drug|Enzyme|Hospital Course|9965,9968|false|false|false|C0022917|Lactate Dehydrogenase|LDH
Finding|Finding|Hospital Course|9965,9968|false|false|false|C0851148|Lifetime Drinking History|LDH
Procedure|Laboratory Procedure|Hospital Course|9965,9968|false|false|false|C0202113|Lactate dehydrogenase measurement|LDH
Attribute|Clinical Attribute|Hospital Course|9970,9973|false|false|false|C0368980|Coagulation tissue factor induced.INR|INR
Procedure|Laboratory Procedure|Hospital Course|9970,9973|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9970,9973|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Disorder|Neoplastic Process|Hospital Course|9974,9977|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Procedure|Laboratory Procedure|Hospital Course|9974,9977|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Finding|Gene or Genome|Hospital Course|10014,10017|false|false|false|C1537987|MT-CO3 gene|CO3
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10019,10024|false|false|false|C0022646|Kidney|renal
Disorder|Disease or Syndrome|Hospital Course|10019,10024|false|false|false|C0042075|Urologic Diseases|renal
Finding|Organ or Tissue Function|Hospital Course|10019,10033|false|false|false|C0232804|Renal function|renal function
Procedure|Laboratory Procedure|Hospital Course|10019,10033|false|false|false|C0022662|Kidney Function Tests|renal function
Finding|Finding|Hospital Course|10025,10033|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|Hospital Course|10025,10033|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|Hospital Course|10025,10033|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|Hospital Course|10025,10033|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Drug|Biologically Active Substance|Hospital Course|10035,10042|false|false|false|C0017725|glucose|glucose
Drug|Organic Chemical|Hospital Course|10035,10042|false|false|false|C0017725|glucose|glucose
Drug|Pharmacologic Substance|Hospital Course|10035,10042|false|false|false|C0017725|glucose|glucose
Lab|Laboratory or Test Result|Hospital Course|10035,10042|false|false|false|C5781949|Glucose^1.5H post dose glucagon|glucose
Procedure|Laboratory Procedure|Hospital Course|10035,10042|false|false|false|C0337438|Glucose measurement|glucose
Finding|Body Substance|Hospital Course|10046,10055|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|10046,10055|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|10046,10055|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|10046,10055|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|10046,10067|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|10046,10067|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|10056,10067|false|false|false|C2926604||Disposition
Procedure|Health Care Activity|Hospital Course|10056,10067|false|false|false|C0184758|Patient disposition|Disposition
Finding|Idea or Concept|Hospital Course|10069,10073|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|10069,10073|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|10069,10073|false|false|false|C1553498|home health encounter|Home
Finding|Body Substance|Hospital Course|10076,10085|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|10076,10085|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|10076,10085|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|10076,10085|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|10076,10095|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|10086,10095|false|false|false|C0945731||Diagnosis
Finding|Classification|Hospital Course|10086,10095|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|10086,10095|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|10086,10095|false|false|false|C0011900|Diagnosis|Diagnosis
Drug|Organic Chemical|Principle Diagnosis|10118,10125|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Drug|Pharmacologic Substance|Principle Diagnosis|10118,10125|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Finding|Intellectual Product|Principle Diagnosis|10118,10125|false|false|false|C1547288|Alcohol - Recreational Drug Use Code|alcohol
Drug|Organic Chemical|Principle Diagnosis|10126,10133|false|false|false|C0163712|Relate - vinyl resin|related
Finding|Finding|Principle Diagnosis|10126,10133|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Finding|Functional Concept|Principle Diagnosis|10126,10133|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Disorder|Disease or Syndrome|Principle Diagnosis|10134,10143|false|false|false|C0019158;C0019159|Hepatitis;Hepatitis A|hepatitis
Disorder|Disease or Syndrome|Principle Diagnosis|10146,10153|false|false|false|C0003962|Ascites|ascites
Finding|Pathologic Function|Principle Diagnosis|10146,10153|false|false|false|C5441966|Peritoneal Effusion|ascites
Finding|Mental Process|Discharge Condition|10177,10183|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|10177,10190|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|10177,10190|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|10184,10190|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|10184,10190|false|false|false|C1546481|What subject filter - Status|Status
Finding|Idea or Concept|Discharge Condition|10192,10197|false|false|false|C1550016|Remote control command - Clear|Clear
Finding|Finding|Discharge Condition|10202,10210|false|false|false|C4068804|Coherent|coherent
Attribute|Clinical Attribute|Discharge Condition|10212,10234|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|10212,10234|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Finding|Finding|Discharge Condition|10221,10234|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|10221,10234|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|10236,10241|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|10236,10241|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|10236,10241|false|false|false|C0718338|Alert brand of caffeine|Alert
Finding|Finding|Discharge Condition|10236,10241|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|10236,10241|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|10236,10241|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|10246,10257|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|10259,10267|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|10259,10267|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|10259,10267|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|10268,10274|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|10268,10274|false|false|false|C1546481|What subject filter - Status|Status
Finding|Functional Concept|Discharge Condition|10276,10286|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|Discharge Condition|10276,10286|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|Discharge Condition|10276,10286|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|Discharge Condition|10276,10286|false|false|false|C1561560|ambulatory encounter|Ambulatory
Finding|Finding|Discharge Condition|10289,10300|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|Discharge Condition|10289,10300|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|Discharge Instructions|10353,10361|false|false|false|C1547192|Organization unit type - Hospital|hospital
Finding|Pathologic Function|Discharge Instructions|10366,10378|false|false|false|C0021368|Inflammation|inflammation
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|10386,10391|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|Discharge Instructions|10386,10391|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|Discharge Instructions|10386,10391|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|Discharge Instructions|10386,10391|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|Discharge Instructions|10386,10391|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|Discharge Instructions|10386,10391|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Finding|Finding|Discharge Instructions|10386,10391|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|Discharge Instructions|10386,10391|false|false|false|C0872387|Procedures on liver|liver
Finding|Finding|Discharge Instructions|10402,10408|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Discharge Instructions|10402,10408|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Drug|Organic Chemical|Discharge Instructions|10416,10423|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Drug|Pharmacologic Substance|Discharge Instructions|10416,10423|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Finding|Intellectual Product|Discharge Instructions|10416,10423|false|false|false|C1547288|Alcohol - Recreational Drug Use Code|alcohol
Finding|Finding|Discharge Instructions|10416,10435|false|false|false|C0001948;C2215684|Alcohol consumption;alcohol consumption (history)|alcohol consumption
Finding|Individual Behavior|Discharge Instructions|10416,10435|false|false|false|C0001948;C2215684|Alcohol consumption;alcohol consumption (history)|alcohol consumption
Disorder|Disease or Syndrome|Discharge Instructions|10424,10435|false|false|false|C0220811|Consumption-archaic term for TB|consumption
Event|Activity|Discharge Instructions|10424,10435|false|false|false|C0009830|Consumption of goods|consumption
Finding|Physiologic Function|Discharge Instructions|10424,10435|false|false|false|C1947907|biologic consumption|consumption
Finding|Finding|Discharge Instructions|10473,10482|false|false|false|C0392209;C0518896;C1442959|Nutrition (function);Nutrition outcomes;Nutritional status|nutrition
Finding|Intellectual Product|Discharge Instructions|10473,10482|false|false|false|C0392209;C0518896;C1442959|Nutrition (function);Nutrition outcomes;Nutritional status|nutrition
Finding|Organism Function|Discharge Instructions|10473,10482|false|false|false|C0392209;C0518896;C1442959|Nutrition (function);Nutrition outcomes;Nutritional status|nutrition
Procedure|Research Activity|Discharge Instructions|10473,10482|false|false|false|C0600072;C1521729|Feeding and dietary regimes;Nutritional Study|nutrition
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|10473,10482|false|false|false|C0600072;C1521729|Feeding and dietary regimes;Nutritional Study|nutrition
Drug|Pharmacologic Substance|Discharge Instructions|10505,10514|false|false|false|C0013227|Pharmaceutical Preparations|medicines
Drug|Organic Chemical|Discharge Instructions|10520,10527|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Drug|Pharmacologic Substance|Discharge Instructions|10520,10527|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Finding|Intellectual Product|Discharge Instructions|10520,10527|false|false|false|C1547288|Alcohol - Recreational Drug Use Code|alcohol
Disorder|Disease or Syndrome|Discharge Instructions|10520,10538|false|false|false|C0236663|Alcohol withdrawal syndrome|alcohol withdrawal
Disorder|Mental or Behavioral Dysfunction|Discharge Instructions|10528,10538|false|false|false|C2825032|Withdrawal (dysfunction)|withdrawal
Event|Activity|Discharge Instructions|10528,10538|false|false|false|C2349954|Withdraw (activity)|withdrawal
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|10528,10538|false|false|false|C3812880|Withdrawal - birth control|withdrawal
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|10558,10563|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|Discharge Instructions|10558,10563|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|Discharge Instructions|10558,10563|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|Discharge Instructions|10558,10563|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|Discharge Instructions|10558,10563|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|Discharge Instructions|10558,10563|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Finding|Finding|Discharge Instructions|10558,10563|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|Discharge Instructions|10558,10563|false|false|false|C0872387|Procedures on liver|liver
Finding|Organ or Tissue Function|Discharge Instructions|10558,10572|false|false|false|C0232741|Liver function|liver function
Finding|Finding|Discharge Instructions|10564,10572|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|Discharge Instructions|10564,10572|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|Discharge Instructions|10564,10572|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|Discharge Instructions|10564,10572|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Disorder|Disease or Syndrome|Discharge Instructions|10585,10590|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|Discharge Instructions|10585,10590|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Procedure|Laboratory Procedure|Discharge Instructions|10585,10596|false|false|false|C0018941|Hematologic Tests|blood tests
Finding|Intellectual Product|Discharge Instructions|10591,10596|false|false|false|C0392366|Tests (qualifier value)|tests
Procedure|Laboratory Procedure|Discharge Instructions|10591,10596|false|false|false|C0022885|Laboratory Procedures|tests
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|10616,10621|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|Discharge Instructions|10616,10621|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|Discharge Instructions|10616,10621|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|Discharge Instructions|10616,10621|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|Discharge Instructions|10616,10621|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|Discharge Instructions|10616,10621|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Finding|Finding|Discharge Instructions|10616,10621|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|Discharge Instructions|10616,10621|false|false|false|C0872387|Procedures on liver|liver
Finding|Organ or Tissue Function|Discharge Instructions|10616,10630|false|false|false|C0232741|Liver function|liver function
Finding|Finding|Discharge Instructions|10622,10630|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|Discharge Instructions|10622,10630|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|Discharge Instructions|10622,10630|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|Discharge Instructions|10622,10630|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Finding|Discharge Instructions|10649,10653|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Discharge Instructions|10649,10653|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Discharge Instructions|10649,10653|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Body Substance|Discharge Instructions|10657,10666|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Discharge Instructions|10657,10666|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Discharge Instructions|10657,10666|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Discharge Instructions|10657,10666|false|false|false|C0030685|Patient Discharge|discharge
Procedure|Health Care Activity|Discharge Instructions|10680,10689|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|10722,10729|false|false|false|C0042027|Urinary tract|urinary
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|10722,10735|false|false|false|C0042027;C1508753|Urinary system;Urinary tract|urinary tract
Anatomy|Body System|Discharge Instructions|10722,10735|false|false|false|C0042027;C1508753|Urinary system;Urinary tract|urinary tract
Disorder|Disease or Syndrome|Discharge Instructions|10722,10745|false|false|false|C0042029|Urinary tract infection|urinary tract infection
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|10730,10735|false|false|false|C1185740|Tract|tract
Disorder|Disease or Syndrome|Discharge Instructions|10736,10745|false|false|false|C0009450|Communicable Diseases|infection
Finding|Pathologic Function|Discharge Instructions|10736,10745|false|false|false|C3714514|Infection|infection
Disorder|Disease or Syndrome|Discharge Instructions|10752,10761|false|false|false|C0032285|Pneumonia|pneumonia
Drug|Organic Chemical|Discharge Instructions|10770,10778|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|Discharge Instructions|10770,10778|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|Discharge Instructions|10770,10778|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Finding|Functional Concept|Discharge Instructions|10770,10778|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|Discharge Instructions|10770,10778|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Antibiotic|Discharge Instructions|10798,10809|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Drug|Antibiotic|Discharge Instructions|10811,10823|false|false|false|C0282386|levofloxacin|levofloxacin
Drug|Organic Chemical|Discharge Instructions|10811,10823|false|false|false|C0282386|levofloxacin|levofloxacin
Disorder|Disease or Syndrome|Discharge Instructions|10841,10851|false|false|false|C0851162|Infection of musculoskeletal system|infections
Finding|Pathologic Function|Discharge Instructions|10841,10851|false|false|false|C3714514|Infection|infections
Finding|Finding|Discharge Instructions|10872,10875|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Discharge Instructions|10872,10875|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Drug|Pharmacologic Substance|Discharge Instructions|10876,10884|false|false|false|C0013227|Pharmaceutical Preparations|medicine
Drug|Substance|Discharge Instructions|10907,10912|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Discharge Instructions|10907,10912|false|false|false|C1546638|Fluid Specimen Code|fluid
Anatomy|Body Location or Region|Discharge Instructions|10923,10930|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|abdomen
Disorder|Neoplastic Process|Discharge Instructions|10923,10930|false|false|false|C0153662|Malignant neoplasm of abdomen|abdomen
Finding|Finding|Discharge Instructions|10923,10930|false|false|false|C0941288|Abdomen problem|abdomen
Anatomy|Body Location or Region|Discharge Instructions|10923,10934|false|false|false|C0000726|Abdomen|abdomen and
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|10935,10939|false|false|false|C1140621|Leg|legs
Attribute|Clinical Attribute|Discharge Instructions|10935,10939|false|false|false|C5781420||legs
Drug|Pharmacologic Substance|Discharge Instructions|10946,10954|false|false|false|C0013227|Pharmaceutical Preparations|medicine
Drug|Organic Chemical|Discharge Instructions|10965,10979|false|false|false|C0037982|spironolactone|spironolactone
Drug|Pharmacologic Substance|Discharge Instructions|10965,10979|false|false|false|C0037982|spironolactone|spironolactone
Drug|Pharmacologic Substance|Discharge Instructions|10993,11001|false|false|false|C0013227|Pharmaceutical Preparations|medicine
Drug|Biologically Active Substance|Discharge Instructions|11012,11021|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Element, Ion, or Isotope|Discharge Instructions|11012,11021|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Food|Discharge Instructions|11012,11021|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Inorganic Chemical|Discharge Instructions|11012,11021|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Pharmacologic Substance|Discharge Instructions|11012,11021|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Finding|Physiologic Function|Discharge Instructions|11012,11021|false|false|false|C4553027|Potassium metabolic function|potassium
Procedure|Laboratory Procedure|Discharge Instructions|11012,11021|false|false|false|C0202194|Potassium measurement|potassium
Disorder|Disease or Syndrome|Discharge Instructions|11036,11041|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|Discharge Instructions|11036,11041|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Disorder|Disease or Syndrome|Discharge Instructions|11075,11080|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|Discharge Instructions|11075,11080|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Event|Occupational Activity|Discharge Instructions|11081,11085|false|false|false|C0043227|Work|work
Finding|Idea or Concept|Discharge Instructions|11094,11098|false|false|false|C1552851|next - HtmlLinkType|next
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|11142,11148|false|false|false|C0018792|Heart Atrium|Atrium
Anatomy|Anatomical Structure|Discharge Instructions|11168,11173|false|false|false|C3714591|Floor (anatomic)|floor
Anatomy|Anatomical Structure|Discharge Instructions|11191,11196|false|false|false|C3714591|Floor (anatomic)|floor
Finding|Functional Concept|Discharge Instructions|11246,11253|false|false|false|C0392747|Changing|changes
Drug|Pharmacologic Substance|Discharge Instructions|11262,11271|false|false|false|C0013227|Pharmaceutical Preparations|medicines
Drug|Organic Chemical|Discharge Instructions|11284,11290|false|false|false|C0178638|folate|folate
Drug|Pharmacologic Substance|Discharge Instructions|11284,11290|false|false|false|C0178638|folate|folate
Drug|Vitamin|Discharge Instructions|11284,11290|false|false|false|C0178638|folate|folate
Procedure|Laboratory Procedure|Discharge Instructions|11284,11290|false|false|false|C0523631|Folic acid measurement|folate
Drug|Organic Chemical|Discharge Instructions|11292,11300|false|false|false|C0039840;C3714802|Thiamine Drug Class;thiamine|thiamine
Drug|Pharmacologic Substance|Discharge Instructions|11292,11300|false|false|false|C0039840;C3714802|Thiamine Drug Class;thiamine|thiamine
Drug|Vitamin|Discharge Instructions|11292,11300|false|false|false|C0039840;C3714802|Thiamine Drug Class;thiamine|thiamine
Procedure|Laboratory Procedure|Discharge Instructions|11292,11300|false|false|false|C0373727|Thiamine measurement|thiamine
Drug|Organic Chemical|Discharge Instructions|11306,11318|false|false|false|C0301532|Multivitamin preparation|multivitamin
Drug|Pharmacologic Substance|Discharge Instructions|11306,11318|false|false|false|C0301532|Multivitamin preparation|multivitamin
Drug|Vitamin|Discharge Instructions|11306,11318|false|false|false|C0301532|Multivitamin preparation|multivitamin
Finding|Classification|Discharge Instructions|11324,11331|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|general
Procedure|Health Care Activity|Discharge Instructions|11324,11331|false|false|false|C3812897|General medical service|general
Finding|Finding|Discharge Instructions|11333,11342|false|false|false|C0392209;C0518896;C1442959|Nutrition (function);Nutrition outcomes;Nutritional status|nutrition
Finding|Intellectual Product|Discharge Instructions|11333,11342|false|false|false|C0392209;C0518896;C1442959|Nutrition (function);Nutrition outcomes;Nutritional status|nutrition
Finding|Organism Function|Discharge Instructions|11333,11342|false|false|false|C0392209;C0518896;C1442959|Nutrition (function);Nutrition outcomes;Nutritional status|nutrition
Procedure|Research Activity|Discharge Instructions|11333,11342|false|false|false|C0600072;C1521729|Feeding and dietary regimes;Nutritional Study|nutrition
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|11333,11342|false|false|false|C0600072;C1521729|Feeding and dietary regimes;Nutritional Study|nutrition
Drug|Organic Chemical|Discharge Instructions|11355,11364|false|false|false|C0023660|lidocaine|lidocaine
Drug|Pharmacologic Substance|Discharge Instructions|11355,11364|false|false|false|C0023660|lidocaine|lidocaine
Procedure|Laboratory Procedure|Discharge Instructions|11355,11364|false|false|false|C0202404|Lidocaine measurement|lidocaine
Drug|Clinical Drug|Discharge Instructions|11355,11370|false|false|false|C1251704|Lidocaine Patch|lidocaine patch
Drug|Biomedical or Dental Material|Discharge Instructions|11365,11370|false|false|false|C0445403;C1533128;C1707974|Body tissue patch material;Human patch material;Patch - Extended Release Film|patch
Finding|Finding|Discharge Instructions|11365,11370|false|false|false|C0332461|Plaque (lesion)|patch
Attribute|Clinical Attribute|Discharge Instructions|11376,11380|false|false|false|C2598155||pain
Finding|Functional Concept|Discharge Instructions|11376,11380|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|11376,11380|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Hazardous or Poisonous Substance|Discharge Instructions|11393,11401|false|false|false|C0028040|nicotine|nicotine
Drug|Organic Chemical|Discharge Instructions|11393,11401|false|false|false|C0028040|nicotine|nicotine
Drug|Clinical Drug|Discharge Instructions|11393,11407|false|false|false|C0358855|Nicotine Transdermal Patch|nicotine patch
Drug|Biomedical or Dental Material|Discharge Instructions|11402,11407|false|false|false|C0445403;C1533128;C1707974|Body tissue patch material;Human patch material;Patch - Extended Release Film|patch
Finding|Finding|Discharge Instructions|11402,11407|false|false|false|C0332461|Plaque (lesion)|patch
Drug|Antibiotic|Discharge Instructions|11419,11431|false|false|false|C0282386|levofloxacin|levofloxacin
Drug|Organic Chemical|Discharge Instructions|11419,11431|false|false|false|C0282386|levofloxacin|levofloxacin
Drug|Antibiotic|Discharge Instructions|11433,11443|false|false|false|C0003232|Antibiotics|antibiotic
Disorder|Disease or Syndrome|Discharge Instructions|11448,11457|false|false|false|C0032285|Pneumonia|pneumonia
Drug|Organic Chemical|Discharge Instructions|11470,11484|false|false|false|C0037982|spironolactone|spironolactone
Drug|Pharmacologic Substance|Discharge Instructions|11470,11484|false|false|false|C0037982|spironolactone|spironolactone
Drug|Pharmacologic Substance|Discharge Instructions|11486,11494|false|false|false|C0012798;C5399719|Diuretic [APC];Diuretics|diuretic
Drug|Substance|Discharge Instructions|11506,11511|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Discharge Instructions|11506,11511|false|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Finding|Discharge Instructions|11513,11525|false|false|false|C4055506|Accumulation|accumulation
Finding|Functional Concept|Discharge Instructions|11547,11554|true|false|false|C0392747|Changing|changes
Drug|Pharmacologic Substance|Discharge Instructions|11563,11572|false|false|false|C0013227|Pharmaceutical Preparations|medicines
Event|Activity|Discharge Instructions|11590,11602|false|false|false|C0003629|Appointments|appointments
Procedure|Health Care Activity|Discharge Instructions|11644,11652|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|11653,11665|false|false|false|C3263700||Instructions
Finding|Intellectual Product|Discharge Instructions|11653,11665|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

