 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|43,52|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|43,52|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|43,57|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|77,86|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|77,86|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|77,91|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|133,136|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|144,151|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|144,151|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|153,161|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|SIMPLE_SEGMENT|164,173|false|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|164,173|false|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|164,173|false|false|false|C0020517|Hypersensitivity|Allergies
Attribute|Clinical Attribute|SIMPLE_SEGMENT|185,194|false|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|185,194|false|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|185,194|false|false|false|C0020517|Hypersensitivity|Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|197,219|true|false|false|C0041755|Adverse reaction to drug|Adverse Drug Reactions
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|205,209|false|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|Drug
Finding|Finding|SIMPLE_SEGMENT|205,209|false|false|false|C0740721|Drug problem|Drug
Finding|Pathologic Function|SIMPLE_SEGMENT|205,219|true|false|false|C0041755|Adverse reaction to drug|Drug Reactions
Event|Event|SIMPLE_SEGMENT|210,219|false|false|false|||Reactions
Event|Event|SIMPLE_SEGMENT|222,231|false|false|false|||Attending
Finding|Functional Concept|SIMPLE_SEGMENT|222,231|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|SIMPLE_SEGMENT|240,255|false|false|false|C0277786|Chief complaint (finding)|Chief Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|246,255|false|false|false|C3864418||Complaint
Event|Event|SIMPLE_SEGMENT|246,255|false|false|false|||Complaint
Finding|Finding|SIMPLE_SEGMENT|246,255|false|false|false|C5441521|Complaint (finding)|Complaint
Finding|Finding|SIMPLE_SEGMENT|257,265|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|Diarrhea
Finding|Sign or Symptom|SIMPLE_SEGMENT|257,265|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|Diarrhea
Event|Event|SIMPLE_SEGMENT|268,276|false|false|false|||Transfer
Finding|Functional Concept|SIMPLE_SEGMENT|268,276|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|Transfer
Finding|Idea or Concept|SIMPLE_SEGMENT|268,276|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|Transfer
Procedure|Health Care Activity|SIMPLE_SEGMENT|268,276|false|false|false|C4706767|Transfer (immobility management)|Transfer
Event|Event|SIMPLE_SEGMENT|280,284|false|false|false|||MICU
Event|Event|SIMPLE_SEGMENT|289,296|false|false|false|||Hypoxia
Finding|Finding|SIMPLE_SEGMENT|289,296|false|false|false|C0242184;C1963140|Hypoxia;Hypoxia, CTCAE|Hypoxia
Finding|Pathologic Function|SIMPLE_SEGMENT|289,296|false|false|false|C0242184;C1963140|Hypoxia;Hypoxia, CTCAE|Hypoxia
Finding|Classification|SIMPLE_SEGMENT|299,304|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|SIMPLE_SEGMENT|305,313|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|305,313|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|317,335|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|326,335|false|false|false|C0945766||Procedure
Event|Event|SIMPLE_SEGMENT|326,335|false|false|false|||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|326,335|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|326,335|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|326,335|false|false|false|C0184661|Interventional procedure|Procedure
Drug|Biologically Active Substance|SIMPLE_SEGMENT|341,345|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|341,345|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Substance|SIMPLE_SEGMENT|341,345|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Finding|Intellectual Product|SIMPLE_SEGMENT|341,345|false|false|false|C1546701|line source specimen code|line
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|341,355|false|false|false|C1519955|Vascular Access Device Placement|line placement
Event|Event|SIMPLE_SEGMENT|346,355|false|false|false|||placement
Procedure|Health Care Activity|SIMPLE_SEGMENT|346,355|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|346,355|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Finding|Functional Concept|SIMPLE_SEGMENT|356,361|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Anatomy|Tissue|SIMPLE_SEGMENT|370,377|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|370,377|false|false|false|C0032226|Pleural Diseases|pleural
Event|Event|SIMPLE_SEGMENT|378,386|false|false|false|||catheter
Finding|Intellectual Product|SIMPLE_SEGMENT|378,386|false|false|false|C1546572||catheter
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|378,396|false|false|false|C0883301|Catheter placement|catheter placement
Event|Event|SIMPLE_SEGMENT|387,396|false|false|false|||placement
Procedure|Health Care Activity|SIMPLE_SEGMENT|387,396|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|387,396|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Event|Event|SIMPLE_SEGMENT|399,406|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|399,406|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|399,406|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|399,406|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|399,409|false|false|false|C0262926|Medical History|History of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|399,425|false|false|false|C0488508||History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|399,425|false|false|false|C0262512|History of present illness (finding)|History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|410,417|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Idea or Concept|SIMPLE_SEGMENT|410,417|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Finding|SIMPLE_SEGMENT|410,425|false|false|false|C4264312|Present illness|Present Illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|418,425|false|false|false|C0221423|Illness (finding)|Illness
Finding|Idea or Concept|SIMPLE_SEGMENT|440,444|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|SIMPLE_SEGMENT|440,444|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Event|Event|SIMPLE_SEGMENT|445,448|false|false|false|||old
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|465,474|false|false|false|C1527336|Sjogren's Syndrome|Sjogren's
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|465,483|false|false|false|C1527336|Sjogren's Syndrome|Sjogren's syndrome
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|475,483|false|false|false|C0039082|Syndrome|syndrome
Event|Event|SIMPLE_SEGMENT|475,483|false|false|false|||syndrome
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|485,488|false|false|false|C0022104;C0432306|Ichthyosis Bullosa of Siemens;Irritable Bowel Syndrome|IBS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|485,488|false|false|false|C0022104;C0432306|Ichthyosis Bullosa of Siemens;Irritable Bowel Syndrome|IBS
Event|Event|SIMPLE_SEGMENT|485,488|false|false|false|||IBS
Event|Event|SIMPLE_SEGMENT|495,503|false|false|false|||presents
Event|Event|SIMPLE_SEGMENT|509,517|false|false|false|||diarrhea
Finding|Finding|SIMPLE_SEGMENT|509,517|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|SIMPLE_SEGMENT|509,517|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Event|Event|SIMPLE_SEGMENT|522,527|false|false|false|||fever
Finding|Finding|SIMPLE_SEGMENT|522,527|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|522,527|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Event|Event|SIMPLE_SEGMENT|537,545|false|false|false|||starting
Finding|Gene or Genome|SIMPLE_SEGMENT|608,611|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Event|Event|SIMPLE_SEGMENT|628,638|false|false|false|||persistent
Finding|Finding|SIMPLE_SEGMENT|650,654|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|650,654|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|650,654|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Finding|SIMPLE_SEGMENT|669,681|false|false|false|C3845714|Several days|several days
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|710,716|false|false|false|C0270814|Spastic syndrome|crampy
Event|Event|SIMPLE_SEGMENT|710,716|false|false|false|||crampy
Anatomy|Body Location or Region|SIMPLE_SEGMENT|721,726|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|721,726|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Location or Region|SIMPLE_SEGMENT|721,745|false|false|false|C0230184|Structure of lower abdominal quadrant|lower quadrant abdominal
Anatomy|Body Location or Region|SIMPLE_SEGMENT|736,745|false|false|false|C0000726|Abdomen|abdominal
Attribute|Clinical Attribute|SIMPLE_SEGMENT|747,751|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|747,751|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|747,751|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|747,751|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|756,766|false|false|false|||distension
Finding|Finding|SIMPLE_SEGMENT|756,766|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distension
Finding|Pathologic Function|SIMPLE_SEGMENT|756,766|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distension
Event|Event|SIMPLE_SEGMENT|778,787|false|false|false|||developed
Attribute|Clinical Attribute|SIMPLE_SEGMENT|788,798|false|false|false|C2979880||subjective
Finding|Finding|SIMPLE_SEGMENT|788,798|false|false|false|C2266644|subjective (symptom)|subjective
Finding|Sign or Symptom|SIMPLE_SEGMENT|788,804|false|false|false|C0743979|Subjective fever|subjective fever
Event|Event|SIMPLE_SEGMENT|799,804|false|false|false|||fever
Finding|Finding|SIMPLE_SEGMENT|799,804|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|799,804|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Event|Event|SIMPLE_SEGMENT|810,816|false|false|false|||rigors
Finding|Sign or Symptom|SIMPLE_SEGMENT|810,816|false|false|false|C0424790|Rigor - Temperature-associated observation|rigors
Finding|Finding|SIMPLE_SEGMENT|817,824|false|false|false|C4534363|At home|at home
Event|Event|SIMPLE_SEGMENT|820,824|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|820,824|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|820,824|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|820,824|false|false|false|C1553498|home health encounter|home
Event|Event|SIMPLE_SEGMENT|826,832|false|false|false|||Denies
Attribute|Clinical Attribute|SIMPLE_SEGMENT|833,839|false|false|false|C4255480||nausea
Event|Event|SIMPLE_SEGMENT|833,839|false|false|false|||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|833,839|false|false|false|C0027497|Nausea|nausea
Event|Event|SIMPLE_SEGMENT|841,849|false|false|false|||vomiting
Finding|Sign or Symptom|SIMPLE_SEGMENT|841,849|true|false|false|C0042963|Vomiting|vomiting
Event|Event|SIMPLE_SEGMENT|851,858|false|false|false|||dysuria
Finding|Sign or Symptom|SIMPLE_SEGMENT|851,858|false|false|false|C0013428|Dysuria|dysuria
Finding|Finding|SIMPLE_SEGMENT|860,869|false|false|false|C0392756;C0442797|Decreasing;Reduced|Decreased
Event|Event|SIMPLE_SEGMENT|871,879|false|false|false|||appetite
Finding|Organism Function|SIMPLE_SEGMENT|871,879|false|false|false|C0003618|Desire for food|appetite
Finding|Finding|SIMPLE_SEGMENT|890,894|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|890,894|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|890,894|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|SIMPLE_SEGMENT|895,901|false|false|false|||course
Finding|Idea or Concept|SIMPLE_SEGMENT|914,921|false|false|false|C1555582|Initial (abbreviation)|initial
Finding|Body Substance|SIMPLE_SEGMENT|956,963|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|956,963|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|956,963|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|965,970|false|false|false|||AAOx3
Event|Event|SIMPLE_SEGMENT|985,992|false|false|false|||febrile
Finding|Sign or Symptom|SIMPLE_SEGMENT|985,992|false|false|false|C0015967|Fever|febrile
Event|Event|SIMPLE_SEGMENT|1003,1007|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|1003,1007|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|1003,1007|false|false|false|C0582103|Medical Examination|Exam
Event|Event|SIMPLE_SEGMENT|1008,1018|false|false|false|||remarkable
Event|Event|SIMPLE_SEGMENT|1023,1027|false|false|false|||mild
Finding|Intellectual Product|SIMPLE_SEGMENT|1023,1027|false|false|false|C1547225|Mild Severity of Illness Code|mild
Event|Event|SIMPLE_SEGMENT|1029,1039|false|false|false|||discomfort
Finding|Sign or Symptom|SIMPLE_SEGMENT|1029,1039|false|false|false|C2364135|Discomfort|discomfort
Event|Event|SIMPLE_SEGMENT|1043,1052|false|false|false|||palpation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1043,1052|false|false|false|C0030247|Palpation|palpation
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1056,1059|false|false|false|C0230178|Structure of right lower quadrant of abdomen|RLQ
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1060,1063|false|false|false|C0230180|Structure of left lower quadrant of abdomen|LLQ
Event|Event|SIMPLE_SEGMENT|1065,1069|false|false|false|||Labs
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1065,1069|false|false|false|C0587081|Laboratory test finding|Labs
Event|Event|SIMPLE_SEGMENT|1070,1077|false|false|false|||notable
Anatomy|Cell|SIMPLE_SEGMENT|1082,1085|false|false|false|C0023516|Leukocytes|WBC
Event|Event|SIMPLE_SEGMENT|1103,1107|false|false|false|||PMNs
Drug|Organic Chemical|SIMPLE_SEGMENT|1128,1135|false|false|false|C0022924;C0376261|Lactates;lactate|lactate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1128,1135|false|false|false|C0022924;C0376261|Lactates;lactate|lactate
Event|Event|SIMPLE_SEGMENT|1128,1135|false|false|false|||lactate
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1128,1135|false|false|false|C0202115|Lactic acid measurement|lactate
Event|Event|SIMPLE_SEGMENT|1148,1152|false|false|false|||LFTs
Event|Event|SIMPLE_SEGMENT|1158,1164|false|false|false|||showed
Finding|Body Substance|SIMPLE_SEGMENT|1167,1174|false|false|false|C0020191|Hyalin Substance|hyaline
Finding|Body Substance|SIMPLE_SEGMENT|1167,1180|false|false|false|C0333121|Hyaline casts|hyaline casts
Event|Event|SIMPLE_SEGMENT|1175,1180|false|false|false|||casts
Finding|Body Substance|SIMPLE_SEGMENT|1175,1180|false|false|false|C0302143|cast body substance|casts
Event|Event|SIMPLE_SEGMENT|1185,1190|false|false|false|||mucus
Finding|Body Substance|SIMPLE_SEGMENT|1185,1190|true|false|false|C0026727;C1546714;C2753459|Mucus (substance);mucus layer|mucus
Finding|Intellectual Product|SIMPLE_SEGMENT|1185,1190|true|false|false|C0026727;C1546714;C2753459|Mucus (substance);mucus layer|mucus
Anatomy|Cell|SIMPLE_SEGMENT|1191,1194|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|1195,1198|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1195,1198|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1195,1198|false|false|false|C0014792|Erythrocytes|RBC
Finding|Idea or Concept|SIMPLE_SEGMENT|1199,1202|false|false|false|C1548556|Etc.|etc
Event|Event|SIMPLE_SEGMENT|1204,1207|false|false|false|||BCx
Event|Event|SIMPLE_SEGMENT|1216,1221|false|false|false|||drawn
Event|Event|SIMPLE_SEGMENT|1224,1226|false|false|false|||CT
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|1236,1244|false|false|false|C0009924|Contrast Media|contrast
Event|Event|SIMPLE_SEGMENT|1236,1244|false|false|false|||contrast
Event|Event|SIMPLE_SEGMENT|1245,1251|false|false|false|||showed
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1252,1262|false|false|false|C0868908|Pancolitis|pancolitis
Event|Event|SIMPLE_SEGMENT|1252,1262|false|false|false|||pancolitis
Event|Event|SIMPLE_SEGMENT|1272,1283|false|false|false|||perforation
Finding|Finding|SIMPLE_SEGMENT|1272,1283|false|false|false|C0549099|Perforation (morphologic abnormality)|perforation
Event|Event|SIMPLE_SEGMENT|1287,1298|false|false|false|||obstruction
Finding|Finding|SIMPLE_SEGMENT|1287,1298|false|false|false|C0028778|Obstruction|obstruction
Event|Event|SIMPLE_SEGMENT|1300,1312|false|false|false|||intrahepatic
Finding|Functional Concept|SIMPLE_SEGMENT|1300,1312|false|false|false|C1512952|Intrahepatic Route of Administration|intrahepatic
Finding|Functional Concept|SIMPLE_SEGMENT|1313,1320|false|false|false|C0521378|Biliary|biliary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1313,1325|false|false|false|C0005400|Bile duct structure|biliary duct
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1321,1325|false|false|false|C0687028;C1550227|Duct (organ) structure;canal [body parts]|duct
Event|Event|SIMPLE_SEGMENT|1326,1336|false|false|false|||dilatation
Finding|Finding|SIMPLE_SEGMENT|1326,1336|false|false|false|C0012359;C0700124|Dilated;Pathological Dilatation|dilatation
Finding|Pathologic Function|SIMPLE_SEGMENT|1326,1336|false|false|false|C0012359;C0700124|Dilated;Pathological Dilatation|dilatation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1326,1336|false|false|false|C1322279|Dilate procedure|dilatation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1352,1355|false|false|false|C3887938|Deuteranomaly|CBD
Drug|Organic Chemical|SIMPLE_SEGMENT|1352,1355|false|false|false|C0006863;C0006982|cannabidiol;carbidopa|CBD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1352,1355|false|false|false|C0006863;C0006982|cannabidiol;carbidopa|CBD
Event|Event|SIMPLE_SEGMENT|1352,1355|false|false|false|||CBD
Finding|Gene or Genome|SIMPLE_SEGMENT|1352,1355|false|false|false|C1415024|OPN1MW gene|CBD
Finding|Functional Concept|SIMPLE_SEGMENT|1357,1362|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1357,1367|false|false|false|C0225706|Right lung|right lung
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1357,1372|false|false|false|C0225708|Structure of base of right lung|right lung base
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1363,1367|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1363,1367|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1363,1367|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|SIMPLE_SEGMENT|1363,1367|false|false|false|C0740941|Lung Problem|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1363,1372|false|false|false|C0225704|Basal segment of lung|lung base
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1368,1372|false|false|false|C2987514|Anatomical base|base
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|1368,1372|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Chemical Viewed Functionally|SIMPLE_SEGMENT|1368,1372|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|1368,1372|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Finding|Gene or Genome|SIMPLE_SEGMENT|1368,1372|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Finding|Idea or Concept|SIMPLE_SEGMENT|1368,1372|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1373,1386|false|false|false|C0521530|Lung consolidation|consolidation
Event|Event|SIMPLE_SEGMENT|1373,1386|false|false|false|||consolidation
Event|Event|SIMPLE_SEGMENT|1388,1391|false|false|false|||CXR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1388,1391|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|SIMPLE_SEGMENT|1392,1398|false|false|false|||showed
Event|Event|SIMPLE_SEGMENT|1410,1419|false|false|false|||opacities
Finding|Finding|SIMPLE_SEGMENT|1410,1419|false|false|false|C0029053;C1265876|Abnormally opaque structure (morphologic abnormality);Decreased translucency|opacities
Finding|Pathologic Function|SIMPLE_SEGMENT|1410,1419|false|false|false|C0029053;C1265876|Abnormally opaque structure (morphologic abnormality);Decreased translucency|opacities
Procedure|Health Care Activity|SIMPLE_SEGMENT|1424,1428|false|false|false|C1315068|Pulmonary ventilator management|pulm
Finding|Pathologic Function|SIMPLE_SEGMENT|1424,1434|false|false|false|C0034063|Pulmonary Edema|pulm edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1429,1434|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|1429,1434|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|1429,1434|false|false|false|C0013604|Edema|edema
Finding|Finding|SIMPLE_SEGMENT|1448,1455|false|false|false|C0700124|Dilated|dilated
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1463,1468|false|false|false|C0021853|Intestines|bowel
Event|Event|SIMPLE_SEGMENT|1469,1474|false|false|false|||loops
Finding|Body Substance|SIMPLE_SEGMENT|1476,1483|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1476,1483|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1476,1483|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|1493,1495|false|false|false|||NS
Drug|Organic Chemical|SIMPLE_SEGMENT|1507,1512|false|false|false|C0701042|Cipro|Cipro
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1507,1512|false|false|false|C0701042|Cipro|Cipro
Event|Event|SIMPLE_SEGMENT|1507,1512|false|false|false|||Cipro
Drug|Organic Chemical|SIMPLE_SEGMENT|1517,1523|false|false|false|C0699678|Flagyl|Flagyl
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1517,1523|false|false|false|C0699678|Flagyl|Flagyl
Drug|Organic Chemical|SIMPLE_SEGMENT|1529,1536|false|false|false|C0699142|Tylenol|Tylenol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1529,1536|false|false|false|C0699142|Tylenol|Tylenol
Finding|Body Substance|SIMPLE_SEGMENT|1538,1545|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1538,1545|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1538,1545|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|1560,1568|false|false|false|||admitted
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1572,1580|false|false|false|C0013227|Pharmaceutical Preparations|medicine
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|1581,1586|false|false|false|C3714591|Floor (anatomic)|floor
Event|Event|SIMPLE_SEGMENT|1603,1610|false|false|false|||hypoxia
Finding|Finding|SIMPLE_SEGMENT|1603,1610|false|false|false|C0242184;C1963140|Hypoxia;Hypoxia, CTCAE|hypoxia
Finding|Pathologic Function|SIMPLE_SEGMENT|1603,1610|false|false|false|C0242184;C1963140|Hypoxia;Hypoxia, CTCAE|hypoxia
Finding|Finding|SIMPLE_SEGMENT|1631,1634|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|1631,1634|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Event|Event|SIMPLE_SEGMENT|1641,1652|false|false|false|||requirement
Finding|Functional Concept|SIMPLE_SEGMENT|1641,1652|false|false|false|C1514873|Requirement|requirement
Finding|Functional Concept|SIMPLE_SEGMENT|1665,1671|false|false|false|C0205341;C1705914|Repeat;Repeat Object|repeat
Event|Event|SIMPLE_SEGMENT|1672,1675|false|false|false|||CXR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1672,1675|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|SIMPLE_SEGMENT|1676,1683|false|false|false|||showing
Finding|Finding|SIMPLE_SEGMENT|1684,1692|false|false|false|C0332149|Possible|possible
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1693,1702|false|true|false|C0032285|Pneumonia|pneumonia
Event|Event|SIMPLE_SEGMENT|1693,1702|false|false|false|||pneumonia
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1707,1716|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1707,1716|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|1707,1716|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|SIMPLE_SEGMENT|1707,1722|false|false|false|C0034063|Pulmonary Edema|pulmonary edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1717,1722|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|1717,1722|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|1717,1722|false|false|false|C0013604|Edema|edema
Drug|Antibiotic|SIMPLE_SEGMENT|1738,1749|false|false|false|C0007561|ceftriaxone|ceftriaxone
Drug|Organic Chemical|SIMPLE_SEGMENT|1738,1749|false|false|false|C0007561|ceftriaxone|ceftriaxone
Event|Event|SIMPLE_SEGMENT|1738,1749|false|false|false|||ceftriaxone
Finding|Finding|SIMPLE_SEGMENT|1754,1762|false|false|false|C0332149|Possible|possible
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1763,1772|false|true|false|C0032285|Pneumonia|pneumonia
Event|Event|SIMPLE_SEGMENT|1763,1772|false|false|false|||pneumonia
Event|Event|SIMPLE_SEGMENT|1782,1793|false|false|false|||transferred
Event|Event|SIMPLE_SEGMENT|1797,1801|false|false|false|||MICU
Event|Activity|SIMPLE_SEGMENT|1808,1815|false|false|false|C1706079||arrival
Event|Event|SIMPLE_SEGMENT|1808,1815|false|false|false|||arrival
Finding|Functional Concept|SIMPLE_SEGMENT|1808,1815|false|false|false|C1555577|arrival - ActRelationshipType|arrival
Event|Event|SIMPLE_SEGMENT|1823,1827|false|false|false|||MICU
Finding|Body Substance|SIMPLE_SEGMENT|1829,1836|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1829,1836|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1829,1836|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Finding|SIMPLE_SEGMENT|1829,1858|false|false|false|C2051418|patient appears uncomfortable|patient appears uncomfortable
Event|Event|SIMPLE_SEGMENT|1845,1858|false|false|false|||uncomfortable
Event|Event|SIMPLE_SEGMENT|1867,1875|false|false|false|||rigoring
Finding|Sign or Symptom|SIMPLE_SEGMENT|1867,1875|false|false|false|C0424790|Rigor - Temperature-associated observation|rigoring
Event|Event|SIMPLE_SEGMENT|1881,1888|false|false|false|||reports
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1889,1895|false|false|false|C0270814|Spastic syndrome|crampy
Event|Event|SIMPLE_SEGMENT|1889,1895|false|false|false|||crampy
Finding|Sign or Symptom|SIMPLE_SEGMENT|1889,1910|false|false|false|C0000729;C3888418|Abdominal Cramps;Colicky Pain|crampy abdominal pain
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1896,1905|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|SIMPLE_SEGMENT|1896,1910|false|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1906,1910|false|true|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|1906,1910|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|1906,1910|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1906,1910|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1918,1923|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|1918,1923|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1925,1932|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|abdomen
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1925,1932|false|false|false|C0153662|Malignant neoplasm of abdomen|abdomen
Event|Event|SIMPLE_SEGMENT|1925,1932|false|false|false|||abdomen
Finding|Finding|SIMPLE_SEGMENT|1925,1932|false|false|false|C0941288|Abdomen problem|abdomen
Event|Event|SIMPLE_SEGMENT|1934,1940|false|false|false|||fevers
Finding|Sign or Symptom|SIMPLE_SEGMENT|1934,1940|false|false|false|C0015967|Fever|fevers
Event|Event|SIMPLE_SEGMENT|1946,1952|false|false|false|||rigors
Finding|Sign or Symptom|SIMPLE_SEGMENT|1946,1952|false|false|false|C0424790|Rigor - Temperature-associated observation|rigors
Event|Event|SIMPLE_SEGMENT|1958,1967|false|false|false|||continues
Finding|Intellectual Product|SIMPLE_SEGMENT|1971,1984|false|false|false|C3641756|Have Diarrhea|have diarrhea
Event|Event|SIMPLE_SEGMENT|1976,1984|false|false|false|||diarrhea
Finding|Finding|SIMPLE_SEGMENT|1976,1984|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|SIMPLE_SEGMENT|1976,1984|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1994,2000|true|false|false|C4255480||nausea
Event|Event|SIMPLE_SEGMENT|1994,2000|false|false|false|||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|1994,2000|true|false|false|C0027497|Nausea|nausea
Finding|Finding|SIMPLE_SEGMENT|1994,2012|true|false|false|C3843946|Nausea or vomiting|nausea or vomiting
Event|Event|SIMPLE_SEGMENT|2004,2012|false|false|false|||vomiting
Finding|Sign or Symptom|SIMPLE_SEGMENT|2004,2012|true|false|false|C0042963|Vomiting|vomiting
Finding|Intellectual Product|SIMPLE_SEGMENT|2014,2018|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Drug|Organic Chemical|SIMPLE_SEGMENT|2019,2024|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2019,2024|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|SIMPLE_SEGMENT|2019,2024|false|false|false|||cough
Finding|Sign or Symptom|SIMPLE_SEGMENT|2019,2024|false|false|false|C0010200|Coughing|cough
Finding|Finding|SIMPLE_SEGMENT|2019,2035|false|false|false|C0239134|Productive Cough|cough productive
Event|Event|SIMPLE_SEGMENT|2025,2035|false|false|false|||productive
Finding|Finding|SIMPLE_SEGMENT|2039,2051|false|false|false|C1997237|White sputum|white sputum
Event|Event|SIMPLE_SEGMENT|2045,2051|false|false|false|||sputum
Finding|Body Substance|SIMPLE_SEGMENT|2045,2051|false|false|false|C0038056;C1546789;C1576419|Specimen Type - Sputum;Sputum|sputum
Finding|Intellectual Product|SIMPLE_SEGMENT|2045,2051|false|false|false|C0038056;C1546789;C1576419|Specimen Type - Sputum;Sputum|sputum
Event|Event|SIMPLE_SEGMENT|2057,2061|false|false|false|||note
Finding|Body Substance|SIMPLE_SEGMENT|2063,2070|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|2063,2070|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|2063,2070|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Antibiotic|SIMPLE_SEGMENT|2085,2096|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|SIMPLE_SEGMENT|2085,2096|false|false|false|||antibiotics
Drug|Antibiotic|SIMPLE_SEGMENT|2106,2118|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Clinical Drug|SIMPLE_SEGMENT|2106,2118|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Organic Chemical|SIMPLE_SEGMENT|2106,2118|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Event|Event|SIMPLE_SEGMENT|2106,2118|false|false|false|||azithromycin
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|2123,2126|false|false|false|C1855179|CATARACT, ANTERIOR POLAR|CAP
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|2123,2126|false|false|false|C0006935|capsule (pharmacologic)|CAP
Event|Event|SIMPLE_SEGMENT|2123,2126|false|false|false|||CAP
Finding|Gene or Genome|SIMPLE_SEGMENT|2123,2126|false|false|false|C1416891;C1418551;C1419093;C1422073;C1422760;C2985259;C4522312|BRD4 gene;BRD4 wt Allele;CAP1 gene;HACD1 gene;LNPEP gene;SERPINB6 gene;SORBS1 gene|CAP
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2123,2126|false|false|false|C0278651;C0280547;C1879916|CAP Regimen;cisplatin/cyclophosphamide/doxorubicin protocol;cyclophosphamide/doxorubicin/prednisone protocol|CAP
Event|Event|SIMPLE_SEGMENT|2131,2137|false|false|false|||Review
Finding|Idea or Concept|SIMPLE_SEGMENT|2131,2137|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|Review
Finding|Intellectual Product|SIMPLE_SEGMENT|2131,2137|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|Review
Finding|Functional Concept|SIMPLE_SEGMENT|2131,2140|false|false|false|C0699752|Review of|Review of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2131,2148|false|false|false|C0488564;C0488565||Review of systems
Procedure|Health Care Activity|SIMPLE_SEGMENT|2131,2148|false|false|false|C0489633|Review of systems (procedure)|Review of systems
Event|Event|SIMPLE_SEGMENT|2141,2148|false|false|false|||systems
Finding|Functional Concept|SIMPLE_SEGMENT|2141,2148|false|false|false|C0449913|System|systems
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2158,2161|false|false|false|C0268529|Proline dehydrogenase deficiency|HPI
Event|Event|SIMPLE_SEGMENT|2158,2161|false|false|false|||HPI
Finding|Finding|SIMPLE_SEGMENT|2158,2161|false|false|false|C0262512;C1323983|History of present illness (finding);allene oxide synthase activity|HPI
Finding|Molecular Function|SIMPLE_SEGMENT|2158,2161|false|false|false|C0262512;C1323983|History of present illness (finding);allene oxide synthase activity|HPI
Event|Event|SIMPLE_SEGMENT|2166,2172|false|false|false|||Denies
Finding|Sign or Symptom|SIMPLE_SEGMENT|2173,2185|true|false|false|C0028081|Night sweats|night sweats
Event|Event|SIMPLE_SEGMENT|2179,2185|false|false|false|||sweats
Finding|Body Substance|SIMPLE_SEGMENT|2179,2185|true|false|false|C0038984;C0038990|Sweat;Sweating|sweats
Finding|Finding|SIMPLE_SEGMENT|2179,2185|true|false|false|C0038984;C0038990|Sweat;Sweating|sweats
Event|Event|SIMPLE_SEGMENT|2187,2193|false|false|false|||Denies
Event|Event|SIMPLE_SEGMENT|2194,2202|false|false|false|||headache
Finding|Sign or Symptom|SIMPLE_SEGMENT|2194,2202|true|false|false|C0018681|Headache|headache
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|2204,2209|false|false|false|C0030471;C1305231|Nasal sinus;Sinus - general anatomical term|sinus
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|2204,2209|false|false|false|C0016169|pathologic fistula|sinus
Drug|Organic Chemical|SIMPLE_SEGMENT|2204,2209|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2204,2209|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Event|Event|SIMPLE_SEGMENT|2210,2220|false|false|false|||tenderness
Finding|Mental Process|SIMPLE_SEGMENT|2210,2220|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|SIMPLE_SEGMENT|2210,2220|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Event|Event|SIMPLE_SEGMENT|2223,2233|false|false|false|||rhinorrhea
Finding|Sign or Symptom|SIMPLE_SEGMENT|2223,2233|false|false|false|C1260880|Rhinorrhea|rhinorrhea
Event|Event|SIMPLE_SEGMENT|2237,2247|false|false|false|||congestion
Finding|Pathologic Function|SIMPLE_SEGMENT|2237,2247|false|false|false|C0700148|Congestion|congestion
Event|Event|SIMPLE_SEGMENT|2249,2255|false|false|false|||Denies
Event|Event|SIMPLE_SEGMENT|2256,2265|false|false|false|||shortness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2256,2275|true|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|SIMPLE_SEGMENT|2256,2275|true|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|SIMPLE_SEGMENT|2269,2275|false|false|false|C0225386|Breath|breath
Event|Event|SIMPLE_SEGMENT|2281,2289|false|false|false|||wheezing
Finding|Sign or Symptom|SIMPLE_SEGMENT|2281,2289|false|false|false|C0043144|Wheezing|wheezing
Event|Event|SIMPLE_SEGMENT|2291,2297|false|false|false|||Denies
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2298,2303|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|2298,2303|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2298,2308|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|2298,2308|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2304,2308|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|2304,2308|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|2304,2308|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|2304,2308|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|2304,2315|false|false|false|C0008031|Chest Pain|pain, chest
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2310,2315|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|2310,2315|false|false|false|C0741025|Chest problem|chest
Finding|Sign or Symptom|SIMPLE_SEGMENT|2310,2324|false|false|false|C0438716|Chest pressure|chest pressure
Event|Event|SIMPLE_SEGMENT|2316,2324|false|false|false|||pressure
Finding|Finding|SIMPLE_SEGMENT|2316,2324|true|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|SIMPLE_SEGMENT|2316,2324|true|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|2316,2324|true|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|2316,2324|true|false|false|C0033095||pressure
Event|Event|SIMPLE_SEGMENT|2326,2338|false|false|false|||palpitations
Finding|Finding|SIMPLE_SEGMENT|2326,2338|false|false|false|C0030252|Palpitations|palpitations
Event|Event|SIMPLE_SEGMENT|2344,2352|false|false|false|||weakness
Finding|Sign or Symptom|SIMPLE_SEGMENT|2344,2352|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Event|Event|SIMPLE_SEGMENT|2354,2360|false|false|false|||Denies
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2361,2367|false|false|false|C4255480||nausea
Event|Event|SIMPLE_SEGMENT|2361,2367|false|false|false|||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|2361,2367|false|false|false|C0027497|Nausea|nausea
Event|Event|SIMPLE_SEGMENT|2369,2377|false|false|false|||vomiting
Finding|Sign or Symptom|SIMPLE_SEGMENT|2369,2377|true|false|false|C0042963|Vomiting|vomiting
Event|Event|SIMPLE_SEGMENT|2379,2385|false|false|false|||Denies
Event|Event|SIMPLE_SEGMENT|2386,2393|false|false|false|||dysuria
Finding|Sign or Symptom|SIMPLE_SEGMENT|2386,2393|false|false|false|C0013428|Dysuria|dysuria
Event|Event|SIMPLE_SEGMENT|2395,2404|false|false|false|||frequency
Finding|Intellectual Product|SIMPLE_SEGMENT|2395,2404|true|false|false|C3898838;C4321352|Frequency;How Often|frequency
Event|Event|SIMPLE_SEGMENT|2410,2417|false|false|false|||urgency
Event|Event|SIMPLE_SEGMENT|2419,2425|false|false|false|||Denies
Event|Event|SIMPLE_SEGMENT|2426,2437|false|false|false|||arthralgias
Finding|Sign or Symptom|SIMPLE_SEGMENT|2426,2437|true|false|false|C0003862|Arthralgia|arthralgias
Event|Event|SIMPLE_SEGMENT|2441,2449|false|false|false|||myalgias
Finding|Sign or Symptom|SIMPLE_SEGMENT|2441,2449|true|false|false|C0231528|Myalgia|myalgias
Event|Event|SIMPLE_SEGMENT|2451,2457|false|false|false|||Denies
Event|Event|SIMPLE_SEGMENT|2458,2464|false|false|false|||rashes
Finding|Sign or Symptom|SIMPLE_SEGMENT|2458,2464|true|false|false|C0015230;C5779628|Exanthema;Skin rash|rashes
Anatomy|Body System|SIMPLE_SEGMENT|2468,2472|false|false|false|C1123023;C4520765|Skin;Skin, Human|skin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2468,2472|true|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2468,2472|true|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Event|Event|SIMPLE_SEGMENT|2468,2472|false|false|false|||skin
Finding|Body Substance|SIMPLE_SEGMENT|2468,2472|true|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Finding|Intellectual Product|SIMPLE_SEGMENT|2468,2472|true|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Event|Event|SIMPLE_SEGMENT|2474,2481|false|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|2474,2481|false|false|false|C0392747|Changing|changes
Finding|Finding|SIMPLE_SEGMENT|2484,2504|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Event|Event|SIMPLE_SEGMENT|2489,2496|false|false|false|||Medical
Finding|Functional Concept|SIMPLE_SEGMENT|2489,2496|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|2489,2496|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|2489,2496|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|2489,2496|false|false|false|C0199168|Medical service|Medical
Finding|Finding|SIMPLE_SEGMENT|2489,2504|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2497,2504|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2497,2504|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2497,2504|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2506,2512|false|false|false|C0002871|Anemia|Anemia
Event|Event|SIMPLE_SEGMENT|2506,2512|false|false|false|||Anemia
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2513,2535|false|false|false|C0694540|borderline cholesterol|Borderline cholesterol
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2524,2535|false|false|false|C0008377|cholesterol|cholesterol
Drug|Organic Chemical|SIMPLE_SEGMENT|2524,2535|false|false|false|C0008377|cholesterol|cholesterol
Event|Event|SIMPLE_SEGMENT|2524,2535|false|false|false|||cholesterol
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2524,2535|false|false|false|C0201950|Cholesterol measurement|cholesterol
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2544,2549|false|false|false|C0018787;C4037974|Chest>Heart;Heart|Heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2544,2549|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|Heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|2544,2549|false|false|false|C0795691|HEART PROBLEM|Heart
Finding|Finding|SIMPLE_SEGMENT|2544,2556|false|false|false|C0018808|Heart murmur|Heart Murmur
Event|Event|SIMPLE_SEGMENT|2550,2556|false|false|false|||Murmur
Finding|Finding|SIMPLE_SEGMENT|2550,2556|false|false|false|C0018808|Heart murmur|Murmur
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2557,2569|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|SIMPLE_SEGMENT|2557,2569|false|false|false|||Hypertension
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2570,2584|false|false|false|C0020676|Hypothyroidism|Hypothyroidism
Event|Event|SIMPLE_SEGMENT|2570,2584|false|false|false|||Hypothyroidism
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2585,2605|false|false|false|C0026266|Mitral Valve Insufficiency|Mitral Regurgitation
Event|Event|SIMPLE_SEGMENT|2592,2605|false|false|false|||Regurgitation
Finding|Finding|SIMPLE_SEGMENT|2592,2605|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|Regurgitation
Finding|Sign or Symptom|SIMPLE_SEGMENT|2592,2605|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|Regurgitation
Phenomenon|Biologic Function|SIMPLE_SEGMENT|2592,2605|false|false|false|C0460152|Regurgitation - mechanism|Regurgitation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2606,2618|false|false|false|C0029456|Osteoporosis|Osteoporosis
Event|Event|SIMPLE_SEGMENT|2606,2618|false|false|false|||Osteoporosis
Finding|Finding|SIMPLE_SEGMENT|2606,2618|false|false|false|C2911643|Encounter due to family history of osteoporosis|Osteoporosis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2619,2628|false|false|false|C0032285|Pneumonia|Pneumonia
Event|Event|SIMPLE_SEGMENT|2619,2628|false|false|false|||Pneumonia
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2629,2638|false|false|false|C0037199|Sinusitis|Sinusitis
Event|Event|SIMPLE_SEGMENT|2629,2638|false|false|false|||Sinusitis
Finding|Functional Concept|SIMPLE_SEGMENT|2646,2652|false|false|false|C0728831|Social|Social
Finding|Finding|SIMPLE_SEGMENT|2646,2660|false|false|false|C0424945;C3714536|Social History;Social and personal history|Social History
Event|Event|SIMPLE_SEGMENT|2653,2660|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2653,2660|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2653,2660|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2653,2660|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Classification|SIMPLE_SEGMENT|2666,2672|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|SIMPLE_SEGMENT|2666,2672|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|SIMPLE_SEGMENT|2666,2672|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|SIMPLE_SEGMENT|2666,2672|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Finding|SIMPLE_SEGMENT|2666,2680|false|false|false|C0241889|Family Medical History|Family History
Event|Event|SIMPLE_SEGMENT|2673,2680|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2673,2680|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2673,2680|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2673,2680|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Event|Event|SIMPLE_SEGMENT|2687,2694|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|2687,2694|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|2687,2694|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|2687,2694|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|2687,2697|false|false|false|C0262926|Medical History|history of
Finding|Finding|SIMPLE_SEGMENT|2687,2710|false|false|false|C0455527||history of hypertension
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2698,2710|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|SIMPLE_SEGMENT|2698,2710|false|false|false|||hypertension
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2714,2724|false|false|false|C3812393|ErbB Receptors|her family
Drug|Enzyme|SIMPLE_SEGMENT|2714,2724|false|false|false|C3812393|ErbB Receptors|her family
Finding|Receptor|SIMPLE_SEGMENT|2714,2724|false|false|false|C3812393|ErbB Receptors|her family
Event|Event|SIMPLE_SEGMENT|2718,2724|false|false|false|||family
Finding|Classification|SIMPLE_SEGMENT|2718,2724|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|2718,2724|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|2718,2724|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|2718,2724|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2736,2742|false|false|false|C4255046||report
Event|Event|SIMPLE_SEGMENT|2736,2742|false|false|false|||report
Finding|Intellectual Product|SIMPLE_SEGMENT|2736,2742|false|false|false|C0684224|Report (document)|report
Procedure|Health Care Activity|SIMPLE_SEGMENT|2736,2742|false|false|false|C0700287|Reporting|report
Event|Event|SIMPLE_SEGMENT|2753,2759|false|false|false|||father
Finding|Conceptual Entity|SIMPLE_SEGMENT|2753,2759|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|father
Finding|Idea or Concept|SIMPLE_SEGMENT|2753,2759|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|father
Finding|Classification|SIMPLE_SEGMENT|2762,2768|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|2762,2768|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|2762,2768|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|2762,2768|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Event|Event|SIMPLE_SEGMENT|2775,2782|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|2775,2782|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|2775,2782|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|2775,2782|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|2775,2785|false|false|false|C0262926|Medical History|history of
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2795,2802|false|false|false|C0006826|Malignant Neoplasms|cancers
Event|Event|SIMPLE_SEGMENT|2795,2802|false|false|false|||cancers
Event|Event|SIMPLE_SEGMENT|2816,2827|false|false|false|||grandfather
Event|Event|SIMPLE_SEGMENT|2835,2842|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|2835,2842|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|2835,2842|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|2835,2842|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|2835,2845|false|false|false|C0262926|Medical History|history of
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2846,2853|false|false|false|C0038351;C3714551;C4266636|Abdomen>Stomach;Stomach;Stomach structure|stomach
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2846,2853|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2846,2853|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Event|Event|SIMPLE_SEGMENT|2846,2853|false|false|false|||stomach
Finding|Finding|SIMPLE_SEGMENT|2846,2853|false|false|false|C0577027|Stomach problem|stomach
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2846,2853|false|false|false|C0872393|Procedure on stomach|stomach
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2846,2860|false|false|false|C0024623;C0699791|Malignant neoplasm of stomach;Stomach Carcinoma|stomach cancer
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2854,2860|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|SIMPLE_SEGMENT|2854,2860|false|false|false|||cancer
Event|Event|SIMPLE_SEGMENT|2882,2889|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|2882,2889|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|2882,2889|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|2882,2889|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|2882,2892|false|false|false|C0262926|Medical History|history of
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2893,2899|false|false|false|C0031354;C0230069;C3665375|Anterior portion of neck;Pharyngeal structure;Throat|throat
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2893,2899|false|false|false|C0031354;C0230069;C3665375|Anterior portion of neck;Pharyngeal structure;Throat|throat
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2893,2899|false|false|false|C1950455|Throat Homeopathic Medication|throat
Finding|Body Substance|SIMPLE_SEGMENT|2893,2899|false|false|false|C1547926;C1550663|Specimen Type - Throat|throat
Finding|Intellectual Product|SIMPLE_SEGMENT|2893,2899|false|false|false|C1547926;C1550663|Specimen Type - Throat|throat
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2893,2906|false|false|false|C0740339|Throat cancer|throat cancer
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2900,2906|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|SIMPLE_SEGMENT|2900,2906|false|false|false|||cancer
Event|Event|SIMPLE_SEGMENT|2913,2919|false|false|false|||denies
Event|Event|SIMPLE_SEGMENT|2924,2931|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|2924,2931|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|2924,2931|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|2924,2931|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|2924,2934|true|false|false|C0262926|Medical History|history of
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2936,2941|false|false|false|C0009368;C4071907|Abdomen+Pelvis>Colon;Colon structure (body structure)|colon
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2936,2941|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2936,2941|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Finding|Finding|SIMPLE_SEGMENT|2936,2941|false|false|false|C0750873|COLON PROBLEM|colon
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2936,2949|false|false|false|C0007102|Malignant tumor of colon|colon cancers
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2942,2949|false|false|false|C0006826|Malignant Neoplasms|cancers
Event|Event|SIMPLE_SEGMENT|2942,2949|false|false|false|||cancers
Finding|Conceptual Entity|SIMPLE_SEGMENT|2951,2957|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Idea or Concept|SIMPLE_SEGMENT|2951,2957|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2962,2968|false|false|false|C0038454|Cerebrovascular accident|stroke
Event|Event|SIMPLE_SEGMENT|2962,2968|false|false|false|||stroke
Finding|Finding|SIMPLE_SEGMENT|2962,2968|false|false|false|C5977286|Stroke (heart beat)|stroke
Finding|Classification|SIMPLE_SEGMENT|2973,2979|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|2973,2979|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|2973,2979|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|2973,2979|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|2988,2994|false|false|false|C1546508|Relationship - Mother|Mother
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3002,3007|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3002,3007|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|3002,3007|false|false|false|C0795691|HEART PROBLEM|heart
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3002,3013|false|false|false|C0018826;C1305961|Heart Valves|heart valve
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3008,3013|false|false|false|C1186983|Anatomical valve|valve
Event|Event|SIMPLE_SEGMENT|3014,3022|false|false|false|||replaced
Event|Event|SIMPLE_SEGMENT|3031,3035|false|false|false|||sure
Finding|Intellectual Product|SIMPLE_SEGMENT|3031,3035|true|false|false|C4724437|SURE Test|sure
Event|Event|SIMPLE_SEGMENT|3051,3059|false|false|false|||Physical
Finding|Finding|SIMPLE_SEGMENT|3051,3059|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|3051,3059|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|3051,3059|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|3051,3064|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|3051,3064|false|false|false|C0031809|Physical Examination|Physical Exam
Event|Event|SIMPLE_SEGMENT|3060,3064|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|3060,3064|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|3060,3064|false|false|false|C0582103|Medical Examination|Exam
Event|Event|SIMPLE_SEGMENT|3066,3075|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|3066,3075|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Event|Event|SIMPLE_SEGMENT|3076,3080|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|3076,3080|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|3076,3080|false|false|false|C0582103|Medical Examination|Exam
Event|Event|SIMPLE_SEGMENT|3082,3089|false|false|false|||General
Finding|Classification|SIMPLE_SEGMENT|3082,3089|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|SIMPLE_SEGMENT|3082,3089|false|false|false|C3812897|General medical service|General
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3091,3096|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|3091,3096|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3091,3096|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|SIMPLE_SEGMENT|3091,3096|false|false|false|||Alert
Finding|Finding|SIMPLE_SEGMENT|3091,3096|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|3091,3096|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|3091,3096|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|SIMPLE_SEGMENT|3098,3106|false|false|false|||oriented
Event|Event|SIMPLE_SEGMENT|3108,3116|false|false|false|||rigoring
Finding|Sign or Symptom|SIMPLE_SEGMENT|3108,3116|false|false|false|C0424790|Rigor - Temperature-associated observation|rigoring
Event|Event|SIMPLE_SEGMENT|3126,3139|false|false|false|||uncomfortable
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3140,3145|false|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3147,3153|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3147,3153|false|false|false|C0036412|Scleral Diseases|Sclera
Procedure|Health Care Activity|SIMPLE_SEGMENT|3147,3153|false|false|false|C2228481|examination of sclera|Sclera
Event|Event|SIMPLE_SEGMENT|3154,3163|false|false|false|||anicteric
Finding|Finding|SIMPLE_SEGMENT|3154,3163|false|false|false|C0205180|Anicteric|anicteric
Finding|Body Substance|SIMPLE_SEGMENT|3169,3174|false|false|false|C0026727;C1546714;C2753459|Mucus (substance);mucus layer|mucus
Finding|Intellectual Product|SIMPLE_SEGMENT|3169,3174|false|false|false|C0026727;C1546714;C2753459|Mucus (substance);mucus layer|mucus
Anatomy|Tissue|SIMPLE_SEGMENT|3175,3184|false|false|false|C0025255|Membrane Tissue|membranes
Event|Event|SIMPLE_SEGMENT|3186,3190|false|false|false|||EOMI
Event|Event|SIMPLE_SEGMENT|3192,3197|false|false|false|||PERRL
Finding|Finding|SIMPLE_SEGMENT|3192,3197|false|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3198,3202|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Anatomy|Cell Component|SIMPLE_SEGMENT|3198,3202|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Finding|Finding|SIMPLE_SEGMENT|3198,3202|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|Neck
Event|Event|SIMPLE_SEGMENT|3204,3210|false|false|false|||supple
Finding|Functional Concept|SIMPLE_SEGMENT|3204,3210|false|false|false|C0332254|Supple|supple
Event|Event|SIMPLE_SEGMENT|3212,3215|false|false|false|||JVP
Finding|Finding|SIMPLE_SEGMENT|3212,3215|false|false|false|C0428897|Jugular venous pressure|JVP
Event|Event|SIMPLE_SEGMENT|3220,3228|false|false|false|||elevated
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3233,3236|true|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3233,3236|true|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|SIMPLE_SEGMENT|3233,3236|false|false|false|||LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|3233,3236|true|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Finding|Finding|SIMPLE_SEGMENT|3262,3281|false|false|false|C0232258|Pansystolic murmur|holosystolic murmur
Event|Event|SIMPLE_SEGMENT|3275,3281|false|false|false|||murmur
Finding|Finding|SIMPLE_SEGMENT|3275,3281|false|false|false|C0018808|Heart murmur|murmur
Anatomy|Cell Component|SIMPLE_SEGMENT|3285,3289|false|false|false|C3890171|dinoflagellate apex|apex
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3285,3289|false|false|false|C0140145|APEX1 protein, human|apex
Drug|Enzyme|SIMPLE_SEGMENT|3285,3289|false|false|false|C0140145|APEX1 protein, human|apex
Finding|Gene or Genome|SIMPLE_SEGMENT|3285,3289|false|false|false|C1332102|APEX1 gene|apex
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3290,3295|false|false|false|C0024109|Lung|Lungs
Event|Event|SIMPLE_SEGMENT|3305,3312|false|false|false|||rhonchi
Finding|Finding|SIMPLE_SEGMENT|3305,3312|false|false|false|C0035508|Rhonchi|rhonchi
Event|Event|SIMPLE_SEGMENT|3317,3324|false|false|false|||wheezes
Finding|Sign or Symptom|SIMPLE_SEGMENT|3317,3324|true|false|false|C0043144|Wheezing|wheezes
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3325,3332|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3325,3332|false|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Event|Event|SIMPLE_SEGMENT|3325,3332|false|false|false|||Abdomen
Finding|Finding|SIMPLE_SEGMENT|3325,3332|false|false|false|C0941288|Abdomen problem|Abdomen
Event|Event|SIMPLE_SEGMENT|3345,3354|false|false|false|||distended
Finding|Finding|SIMPLE_SEGMENT|3345,3354|false|false|false|C0700124|Dilated|distended
Event|Event|SIMPLE_SEGMENT|3356,3362|false|false|false|||tender
Event|Event|SIMPLE_SEGMENT|3366,3375|false|false|false|||palpation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3366,3375|false|false|false|C0030247|Palpation|palpation
Finding|Functional Concept|SIMPLE_SEGMENT|3379,3384|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Finding|Functional Concept|SIMPLE_SEGMENT|3390,3394|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3390,3409|false|false|false|C0230180|Structure of left lower quadrant of abdomen|left lower quadrant
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3395,3400|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|3395,3400|false|false|false|C2003888|Lower (action)|lower
Event|Event|SIMPLE_SEGMENT|3414,3421|false|false|false|||rebound
Event|Event|SIMPLE_SEGMENT|3422,3430|false|false|false|||guarding
Finding|Finding|SIMPLE_SEGMENT|3422,3430|true|false|false|C0427198|Protective muscle spasm|guarding
Event|Event|SIMPLE_SEGMENT|3435,3440|false|false|false|||foley
Event|Activity|SIMPLE_SEGMENT|3444,3449|false|false|false|C1882509|put - instruction imperative|place
Event|Event|SIMPLE_SEGMENT|3444,3449|false|false|false|||place
Finding|Functional Concept|SIMPLE_SEGMENT|3444,3449|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|SIMPLE_SEGMENT|3444,3449|false|false|false|C1533810||place
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|3450,3453|false|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Event|Event|SIMPLE_SEGMENT|3450,3453|false|false|false|||Ext
Finding|Gene or Genome|SIMPLE_SEGMENT|3450,3453|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Event|Event|SIMPLE_SEGMENT|3455,3459|false|false|false|||warm
Finding|Finding|SIMPLE_SEGMENT|3455,3459|false|false|false|C0582051|Feels warm|warm
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3455,3459|false|false|false|C0687712|warming process|warm
Finding|Finding|SIMPLE_SEGMENT|3461,3465|false|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|3466,3474|false|false|false|||perfused
Drug|Food|SIMPLE_SEGMENT|3479,3485|false|false|false|C5890763||pulses
Event|Event|SIMPLE_SEGMENT|3479,3485|false|false|false|||pulses
Finding|Physiologic Function|SIMPLE_SEGMENT|3479,3485|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|SIMPLE_SEGMENT|3479,3485|false|false|false|C0034107|Pulse taking|pulses
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|3490,3498|true|false|false|C0149651|Clubbing|clubbing
Event|Event|SIMPLE_SEGMENT|3490,3498|false|false|false|||clubbing
Event|Event|SIMPLE_SEGMENT|3500,3508|false|false|false|||cyanosis
Finding|Sign or Symptom|SIMPLE_SEGMENT|3500,3508|true|false|false|C0010520|Cyanosis|cyanosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3513,3518|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|3513,3518|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|3513,3518|false|false|false|C0013604|Edema|edema
Event|Event|SIMPLE_SEGMENT|3535,3541|false|false|false|||intact
Finding|Finding|SIMPLE_SEGMENT|3535,3541|false|false|false|C1554187|Gender Status - Intact|intact
Event|Event|SIMPLE_SEGMENT|3543,3549|false|false|false|||moving
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3550,3565|false|false|false|C0278454|All extremities|all extremities
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3554,3565|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Event|Event|SIMPLE_SEGMENT|3568,3577|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|3568,3577|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|3568,3577|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|3568,3577|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|3568,3577|false|false|false|C0030685|Patient Discharge|Discharge
Event|Event|SIMPLE_SEGMENT|3578,3582|false|false|false|||exam
Finding|Functional Concept|SIMPLE_SEGMENT|3578,3582|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|3578,3582|false|false|false|C0582103|Medical Examination|exam
Event|Event|SIMPLE_SEGMENT|3585,3594|false|false|false|||unchanged
Finding|Finding|SIMPLE_SEGMENT|3585,3594|false|false|false|C0442739||unchanged
Finding|Idea or Concept|SIMPLE_SEGMENT|3600,3605|false|false|false|C1552828|Table Frame - above|above
Event|Event|SIMPLE_SEGMENT|3624,3631|false|false|false|||General
Finding|Classification|SIMPLE_SEGMENT|3624,3631|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|SIMPLE_SEGMENT|3624,3631|false|false|false|C3812897|General medical service|General
Event|Event|SIMPLE_SEGMENT|3633,3638|false|false|false|||tired
Finding|Finding|SIMPLE_SEGMENT|3633,3638|false|false|false|C0015672;C0849970;C3539029|Fatigue;Feel Tired question;Feeling tired|tired
Finding|Intellectual Product|SIMPLE_SEGMENT|3633,3638|false|false|false|C0015672;C0849970;C3539029|Fatigue;Feel Tired question;Feeling tired|tired
Finding|Sign or Symptom|SIMPLE_SEGMENT|3633,3638|false|false|false|C0015672;C0849970;C3539029|Fatigue;Feel Tired question;Feeling tired|tired
Event|Event|SIMPLE_SEGMENT|3643,3652|false|false|false|||arousable
Event|Event|SIMPLE_SEGMENT|3656,3661|false|false|false|||voice
Finding|Idea or Concept|SIMPLE_SEGMENT|3656,3661|false|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Finding|Intellectual Product|SIMPLE_SEGMENT|3656,3661|false|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Finding|Organism Function|SIMPLE_SEGMENT|3656,3661|false|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Event|Event|SIMPLE_SEGMENT|3663,3674|false|false|false|||appropriate
Event|Event|SIMPLE_SEGMENT|3679,3682|false|false|false|||RRR
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|3688,3696|false|false|false|C0039155|Systole|systolic
Finding|Finding|SIMPLE_SEGMENT|3688,3703|false|false|false|C0232257|Systolic Murmurs|systolic murmur
Event|Event|SIMPLE_SEGMENT|3697,3703|false|false|false|||murmur
Finding|Finding|SIMPLE_SEGMENT|3697,3703|false|false|false|C0018808|Heart murmur|murmur
Anatomy|Cell Component|SIMPLE_SEGMENT|3711,3715|false|false|false|C3890171|dinoflagellate apex|apex
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3711,3715|false|false|false|C0140145|APEX1 protein, human|apex
Drug|Enzyme|SIMPLE_SEGMENT|3711,3715|false|false|false|C0140145|APEX1 protein, human|apex
Finding|Gene or Genome|SIMPLE_SEGMENT|3711,3715|false|false|false|C1332102|APEX1 gene|apex
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3716,3721|false|false|false|C0024109|Lung|Lungs
Event|Event|SIMPLE_SEGMENT|3732,3741|false|false|false|||decreased
Finding|Finding|SIMPLE_SEGMENT|3732,3755|false|false|false|C0238844|Decreased breath sounds|decreased breath sounds
Finding|Body Substance|SIMPLE_SEGMENT|3742,3748|false|false|false|C0225386|Breath|breath
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3742,3755|false|false|false|C0035234;C3484186|Respiratory Sounds|breath sounds
Event|Event|SIMPLE_SEGMENT|3749,3755|false|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3749,3755|false|false|false|C0037709||sounds
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3763,3767|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3763,3767|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3763,3767|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|SIMPLE_SEGMENT|3763,3767|false|false|false|C0740941|Lung Problem|lung
Drug|Chemical Viewed Functionally|SIMPLE_SEGMENT|3768,3773|false|false|false|C0178499|Base|bases
Event|Event|SIMPLE_SEGMENT|3768,3773|false|false|false|||bases
Event|Event|SIMPLE_SEGMENT|3775,3780|false|false|false|||right
Finding|Functional Concept|SIMPLE_SEGMENT|3775,3780|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Event|Event|SIMPLE_SEGMENT|3790,3798|false|false|false|||catheter
Finding|Intellectual Product|SIMPLE_SEGMENT|3790,3798|false|false|false|C1546572||catheter
Event|Activity|SIMPLE_SEGMENT|3802,3807|false|false|false|C1882509|put - instruction imperative|place
Event|Event|SIMPLE_SEGMENT|3802,3807|false|false|false|||place
Finding|Functional Concept|SIMPLE_SEGMENT|3802,3807|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|SIMPLE_SEGMENT|3802,3807|false|false|false|C1533810||place
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3808,3811|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|Abd
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|3808,3811|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|Abd
Finding|Finding|SIMPLE_SEGMENT|3813,3823|false|false|false|C0086439|Hypokinesia|Hypoactive
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3828,3832|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|SIMPLE_SEGMENT|3828,3832|false|false|false|||soft
Event|Event|SIMPLE_SEGMENT|3853,3862|false|false|false|||distended
Finding|Finding|SIMPLE_SEGMENT|3853,3862|false|false|false|C0700124|Dilated|distended
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3872,3877|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|3872,3877|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|3872,3877|false|false|false|C0013604|Edema|edema
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3885,3890|false|false|false|C0039866;C4299091|Lower extremity>Thigh;Thigh structure|thigh
Procedure|Health Care Activity|SIMPLE_SEGMENT|3924,3933|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Event|Event|SIMPLE_SEGMENT|3934,3938|false|false|false|||Labs
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3934,3938|false|false|false|C0587081|Laboratory test finding|Labs
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3952,3957|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3952,3957|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3952,3957|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|3958,3961|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|3969,3972|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3969,3972|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3969,3972|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3979,3982|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3979,3982|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|3979,3982|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3979,3982|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3989,3992|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3989,3992|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|3999,4002|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|3999,4002|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3999,4002|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3999,4002|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3999,4002|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|4006,4009|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4006,4009|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|4006,4009|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|4006,4009|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|4006,4009|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4006,4009|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|SIMPLE_SEGMENT|4015,4019|false|false|false|||MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4015,4019|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4034,4037|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4054,4059|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4054,4059|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4054,4059|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4072,4078|false|false|false|C0024202|Lymph|Lymphs
Drug|Antibiotic|SIMPLE_SEGMENT|4084,4089|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4084,4089|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|SIMPLE_SEGMENT|4084,4089|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4094,4097|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|Eos
Event|Event|SIMPLE_SEGMENT|4094,4097|false|false|false|||Eos
Finding|Gene or Genome|SIMPLE_SEGMENT|4094,4097|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|Eos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4124,4129|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4124,4129|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4124,4129|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4134,4137|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|SIMPLE_SEGMENT|4134,4137|false|false|false|||PTT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4134,4137|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4159,4164|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4159,4164|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4159,4164|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|4159,4172|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4159,4172|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4159,4172|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4165,4172|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|4165,4172|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4165,4172|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|4165,4172|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4165,4172|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4165,4172|false|false|false|C0337438|Glucose measurement|Glucose
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4248,4253|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4248,4253|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4248,4253|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4254,4257|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4254,4257|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|SIMPLE_SEGMENT|4254,4257|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|SIMPLE_SEGMENT|4254,4257|false|false|false|||ALT
Finding|Gene or Genome|SIMPLE_SEGMENT|4254,4257|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|SIMPLE_SEGMENT|4254,4257|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|SIMPLE_SEGMENT|4254,4257|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4254,4257|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4261,4264|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4261,4264|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4261,4264|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4261,4264|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|SIMPLE_SEGMENT|4261,4264|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|SIMPLE_SEGMENT|4261,4264|false|false|false|||AST
Finding|Gene or Genome|SIMPLE_SEGMENT|4261,4264|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4268,4275|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|SIMPLE_SEGMENT|4268,4275|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4303,4308|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4303,4308|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4303,4308|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4309,4315|false|false|false|C0023764|lipase|Lipase
Drug|Enzyme|SIMPLE_SEGMENT|4309,4315|false|false|false|C0023764|lipase|Lipase
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4309,4315|false|false|false|C0023764|lipase|Lipase
Event|Event|SIMPLE_SEGMENT|4309,4315|false|false|false|||Lipase
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4309,4315|false|false|false|C0373670|Lipase measurement|Lipase
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4331,4336|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4331,4336|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4331,4336|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4331,4344|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4337,4344|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4337,4344|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4337,4344|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4337,4344|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|4337,4344|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|SIMPLE_SEGMENT|4337,4344|false|false|false|||Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|4337,4344|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4337,4344|false|false|false|C0201925|Calcium measurement|Calcium
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4380,4385|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4380,4385|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4380,4385|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4380,4393|false|false|false|C0853248|Blood albumin|BLOOD Albumin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4386,4393|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4386,4393|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4386,4393|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Event|Event|SIMPLE_SEGMENT|4386,4393|false|false|false|||Albumin
Finding|Gene or Genome|SIMPLE_SEGMENT|4386,4393|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Finding|Physiologic Function|SIMPLE_SEGMENT|4386,4393|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4386,4393|false|false|false|C0201838|Albumin measurement|Albumin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4410,4415|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4410,4415|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4410,4415|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4410,4423|false|false|false|C3824990|lactate in blood (lab test)|BLOOD Lactate
Drug|Organic Chemical|SIMPLE_SEGMENT|4416,4423|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4416,4423|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4416,4423|false|false|false|C0202115|Lactic acid measurement|Lactate
Event|Event|SIMPLE_SEGMENT|4430,4439|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|4430,4439|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|4430,4439|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|4430,4439|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|4430,4439|false|false|false|C0030685|Patient Discharge|Discharge
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4440,4444|false|false|false|C0587081|Laboratory test finding|Labs
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4458,4463|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4458,4463|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4458,4463|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|4464,4467|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|4472,4475|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4472,4475|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4472,4475|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4482,4485|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4482,4485|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|4482,4485|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4482,4485|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4491,4494|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4491,4494|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|4502,4505|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|4502,4505|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4502,4505|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4502,4505|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4502,4505|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|4509,4512|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4509,4512|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|4509,4512|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|4509,4512|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|4509,4512|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4509,4512|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|SIMPLE_SEGMENT|4518,4522|false|false|false|||MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4518,4522|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4538,4541|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4558,4563|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4558,4563|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4558,4563|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|4558,4571|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4558,4571|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4558,4571|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4564,4571|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|4564,4571|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4564,4571|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|4564,4571|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4564,4571|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4564,4571|false|false|false|C0337438|Glucose measurement|Glucose
Event|Event|SIMPLE_SEGMENT|4637,4642|false|false|false|||Micro
Finding|Conceptual Entity|SIMPLE_SEGMENT|4637,4642|false|false|false|C3811161;C4049106|Micro (prefix);Microbiology - Laboratory Class|Micro
Finding|Intellectual Product|SIMPLE_SEGMENT|4637,4642|false|false|false|C3811161;C4049106|Micro (prefix);Microbiology - Laboratory Class|Micro
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4637,4642|false|false|false|C0085672|Microbiology procedure|Micro
Finding|Body Substance|SIMPLE_SEGMENT|4644,4649|false|false|false|C0015733|Feces|Stool
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4644,4657|false|false|false|C0430414|Stool culture|Stool Culture
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4650,4657|false|false|false|C1706355|Culture Dose Form|Culture
Event|Event|SIMPLE_SEGMENT|4650,4657|false|false|false|||Culture
Finding|Functional Concept|SIMPLE_SEGMENT|4650,4657|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|Culture
Finding|Idea or Concept|SIMPLE_SEGMENT|4650,4657|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|Culture
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4650,4657|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|Culture
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4681,4684|false|false|false|C0012854|DNA|DNA
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|4681,4684|false|false|false|C0012854|DNA|DNA
Finding|Genetic Function|SIMPLE_SEGMENT|4681,4698|false|false|false|C0683230|dna amplification|DNA amplification
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|4685,4698|false|false|false|C1705759|Gene Amplification Abnormality|amplification
Event|Event|SIMPLE_SEGMENT|4685,4698|false|false|false|||amplification
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|4685,4698|false|false|false|C1521871|Amplification|amplification
Procedure|Molecular Biology Research Technique|SIMPLE_SEGMENT|4685,4698|false|false|false|C1517480|Gene Amplification Technique|amplification
Event|Event|SIMPLE_SEGMENT|4699,4704|false|false|false|||assay
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4699,4704|false|false|false|C0005507;C1510438|Assay;Biological Assay|assay
Finding|Idea or Concept|SIMPLE_SEGMENT|4706,4711|false|false|false|C1546485|Diagnosis Type - Final|Final
Event|Event|SIMPLE_SEGMENT|4724,4732|false|false|false|||Reported
Event|Event|SIMPLE_SEGMENT|4740,4744|false|false|false|||read
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|4820,4828|false|false|false|C4727483|BRAF Gene Rearrangement|Positive
Event|Event|SIMPLE_SEGMENT|4820,4828|false|false|false|||Positive
Finding|Classification|SIMPLE_SEGMENT|4820,4828|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|Positive
Finding|Finding|SIMPLE_SEGMENT|4820,4828|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|Positive
Finding|Finding|SIMPLE_SEGMENT|4820,4832|false|false|false|C1446409|Positive|Positive for
Finding|Intellectual Product|SIMPLE_SEGMENT|4833,4842|false|false|false|C0445332|Toxigenic|toxigenic
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4875,4878|false|false|false|C0012854|DNA|DNA
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|4875,4878|false|false|false|C0012854|DNA|DNA
Event|Event|SIMPLE_SEGMENT|4875,4878|false|false|false|||DNA
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|4888,4901|false|false|false|C1705759|Gene Amplification Abnormality|amplification
Event|Event|SIMPLE_SEGMENT|4888,4901|false|false|false|||amplification
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|4888,4901|false|false|false|C1521871|Amplification|amplification
Procedure|Molecular Biology Research Technique|SIMPLE_SEGMENT|4888,4901|false|false|false|C1517480|Gene Amplification Technique|amplification
Finding|Conceptual Entity|SIMPLE_SEGMENT|4915,4924|false|false|false|C1514811;C1561577;C1706462;C3244318;C4266518|Bibliographic Reference;Reference - HL7UpdateMode;Reference - MdfHmdMetSourceType;Reference Object;Reference source|Reference
Finding|Idea or Concept|SIMPLE_SEGMENT|4915,4924|false|false|false|C1514811;C1561577;C1706462;C3244318;C4266518|Bibliographic Reference;Reference - HL7UpdateMode;Reference - MdfHmdMetSourceType;Reference Object;Reference source|Reference
Finding|Intellectual Product|SIMPLE_SEGMENT|4915,4924|false|false|false|C1514811;C1561577;C1706462;C3244318;C4266518|Bibliographic Reference;Reference - HL7UpdateMode;Reference - MdfHmdMetSourceType;Reference Object;Reference source|Reference
Finding|Intellectual Product|SIMPLE_SEGMENT|4925,4930|false|false|false|C3542016|Concept model range (foundation metadata concept)|Range
Event|Event|SIMPLE_SEGMENT|4931,4939|false|false|false|||Negative
Finding|Classification|SIMPLE_SEGMENT|4931,4939|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|Negative
Finding|Finding|SIMPLE_SEGMENT|4931,4939|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|Negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4931,4939|false|false|false|C5237010|Expression Negative|Negative
Finding|Body Substance|SIMPLE_SEGMENT|4947,4952|false|false|false|C0015733|Feces|FECAL
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4947,4960|false|false|false|C0430414|Stool culture|FECAL CULTURE
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4953,4960|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|SIMPLE_SEGMENT|4953,4960|false|false|false|||CULTURE
Finding|Functional Concept|SIMPLE_SEGMENT|4953,4960|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|SIMPLE_SEGMENT|4953,4960|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4953,4960|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Event|Event|SIMPLE_SEGMENT|4962,4967|false|false|false|||Final
Finding|Idea or Concept|SIMPLE_SEGMENT|4962,4967|false|false|false|C1546485|Diagnosis Type - Final|Final
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4979,4989|true|false|false|C0036117|Salmonella infections|SALMONELLA
Event|Event|SIMPLE_SEGMENT|4979,4989|false|false|false|||SALMONELLA
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4993,5001|true|false|false|C0013371|Shigella Infections|SHIGELLA
Event|Event|SIMPLE_SEGMENT|4993,5001|false|false|false|||SHIGELLA
Event|Event|SIMPLE_SEGMENT|5003,5008|false|false|false|||FOUND
Finding|Finding|SIMPLE_SEGMENT|5003,5008|false|false|false|C0150312|Present|FOUND
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5015,5036|false|false|false|C1294214|Campylobacter culture|CAMPYLOBACTER CULTURE
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5029,5036|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|SIMPLE_SEGMENT|5029,5036|false|false|false|||CULTURE
Finding|Functional Concept|SIMPLE_SEGMENT|5029,5036|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|SIMPLE_SEGMENT|5029,5036|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5029,5036|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Finding|Idea or Concept|SIMPLE_SEGMENT|5038,5043|false|false|false|C1546485|Diagnosis Type - Final|Final
Event|Event|SIMPLE_SEGMENT|5070,5075|false|false|false|||FOUND
Finding|Finding|SIMPLE_SEGMENT|5070,5075|false|false|false|C0150312|Present|FOUND
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5091,5099|false|false|false|C3161394|Mini-bronchoalveolar lavage|Mini-BAL
Finding|Idea or Concept|SIMPLE_SEGMENT|5131,5136|false|false|false|C1546485|Diagnosis Type - Final|FINAL
Finding|Intellectual Product|SIMPLE_SEGMENT|5131,5143|false|false|false|C0460114|Final report|FINAL REPORT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5137,5143|false|false|false|C4255046||REPORT
Event|Event|SIMPLE_SEGMENT|5137,5143|false|false|false|||REPORT
Finding|Intellectual Product|SIMPLE_SEGMENT|5137,5143|false|false|false|C0684224|Report (document)|REPORT
Procedure|Health Care Activity|SIMPLE_SEGMENT|5137,5143|false|false|false|C0700287|Reporting|REPORT
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|5152,5162|false|false|false|C0061856|Gram's stain|GRAM STAIN
Drug|Organic Chemical|SIMPLE_SEGMENT|5152,5162|false|false|false|C0061856|Gram's stain|GRAM STAIN
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5152,5162|false|false|false|C0200966|Bacterial stain, routine|GRAM STAIN
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|5157,5162|false|false|false|C0038128|Stains|STAIN
Event|Event|SIMPLE_SEGMENT|5157,5162|false|false|false|||STAIN
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5157,5162|false|false|false|C0487602|Staining method|STAIN
Finding|Idea or Concept|SIMPLE_SEGMENT|5164,5169|false|false|false|C1546485|Diagnosis Type - Final|Final
Event|Event|SIMPLE_SEGMENT|5202,5207|false|false|false|||FIELD
Finding|Conceptual Entity|SIMPLE_SEGMENT|5202,5207|false|false|false|C1521738;C2346620;C2349184|Field;Force Field;Knowledge Field|FIELD
Procedure|Health Care Activity|SIMPLE_SEGMENT|5202,5207|false|false|false|C1553496|field - patient encounter|FIELD
Event|Event|SIMPLE_SEGMENT|5212,5229|false|false|false|||POLYMORPHONUCLEAR
Anatomy|Cell|SIMPLE_SEGMENT|5231,5241|false|false|false|C0023516|Leukocytes|LEUKOCYTES
Event|Event|SIMPLE_SEGMENT|5231,5241|false|false|false|||LEUKOCYTES
Finding|Body Substance|SIMPLE_SEGMENT|5231,5241|false|false|false|C1547962;C1550647|Specimen Type - Leukocytes|LEUKOCYTES
Finding|Intellectual Product|SIMPLE_SEGMENT|5231,5241|false|false|false|C1547962;C1550647|Specimen Type - Leukocytes|LEUKOCYTES
Finding|Finding|SIMPLE_SEGMENT|5253,5272|false|false|false|C2924473|Microorganisms seen|MICROORGANISMS SEEN
Event|Event|SIMPLE_SEGMENT|5268,5272|false|false|false|||SEEN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5279,5290|false|false|false|C0231832|Respiratory rate|RESPIRATORY
Finding|Body Substance|SIMPLE_SEGMENT|5279,5290|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|RESPIRATORY
Finding|Functional Concept|SIMPLE_SEGMENT|5279,5290|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|RESPIRATORY
Finding|Intellectual Product|SIMPLE_SEGMENT|5279,5290|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|RESPIRATORY
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5279,5298|false|false|false|C4282127|Respiratory culture|RESPIRATORY CULTURE
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5291,5298|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|SIMPLE_SEGMENT|5291,5298|false|false|false|||CULTURE
Finding|Functional Concept|SIMPLE_SEGMENT|5291,5298|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|SIMPLE_SEGMENT|5291,5298|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5291,5298|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Finding|Idea or Concept|SIMPLE_SEGMENT|5300,5305|false|false|false|C1546485|Diagnosis Type - Final|Final
Event|Event|SIMPLE_SEGMENT|5317,5323|false|false|false|||GROWTH
Finding|Finding|SIMPLE_SEGMENT|5317,5323|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|5317,5323|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organism Function|SIMPLE_SEGMENT|5317,5323|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Physiologic Function|SIMPLE_SEGMENT|5317,5323|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|5317,5323|true|false|false|C2911660|Growth action|GROWTH
Event|Event|SIMPLE_SEGMENT|5332,5335|false|false|false|||CFU
Anatomy|Tissue|SIMPLE_SEGMENT|5355,5362|false|false|false|C0032225|Pleura|PLEURAL
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5355,5362|false|false|false|C0032226|Pleural Diseases|PLEURAL
Finding|Body Substance|SIMPLE_SEGMENT|5355,5368|false|false|false|C0225778|Pleural fluid|PLEURAL FLUID
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5355,5368|false|false|false|C2242629|Pleural fluid analysis|PLEURAL FLUID
Drug|Substance|SIMPLE_SEGMENT|5363,5368|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|FLUID
Event|Event|SIMPLE_SEGMENT|5363,5368|false|false|false|||FLUID
Finding|Intellectual Product|SIMPLE_SEGMENT|5363,5368|false|false|false|C1546638|Fluid Specimen Code|FLUID
Finding|Body Substance|SIMPLE_SEGMENT|5363,5381|false|false|false|C0225778|Pleural fluid|FLUID      PLEURAL
Anatomy|Tissue|SIMPLE_SEGMENT|5374,5381|false|false|false|C0032225|Pleura|PLEURAL
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5374,5381|false|false|false|C0032226|Pleural Diseases|PLEURAL
Finding|Body Substance|SIMPLE_SEGMENT|5374,5387|false|false|false|C0225778|Pleural fluid|PLEURAL FLUID
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5374,5387|false|false|false|C2242629|Pleural fluid analysis|PLEURAL FLUID
Drug|Substance|SIMPLE_SEGMENT|5382,5387|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|FLUID
Event|Event|SIMPLE_SEGMENT|5382,5387|false|false|false|||FLUID
Finding|Intellectual Product|SIMPLE_SEGMENT|5382,5387|false|false|false|C1546638|Fluid Specimen Code|FLUID
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|5394,5404|false|false|false|C0061856|Gram's stain|GRAM STAIN
Drug|Organic Chemical|SIMPLE_SEGMENT|5394,5404|false|false|false|C0061856|Gram's stain|GRAM STAIN
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5394,5404|false|false|false|C0200966|Bacterial stain, routine|GRAM STAIN
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|5399,5404|false|false|false|C0038128|Stains|STAIN
Event|Event|SIMPLE_SEGMENT|5399,5404|false|false|false|||STAIN
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5399,5404|false|false|false|C0487602|Staining method|STAIN
Finding|Idea or Concept|SIMPLE_SEGMENT|5406,5411|false|false|false|C1546485|Diagnosis Type - Final|Final
Event|Event|SIMPLE_SEGMENT|5443,5448|false|false|false|||FIELD
Finding|Conceptual Entity|SIMPLE_SEGMENT|5443,5448|false|false|false|C1521738;C2346620;C2349184|Field;Force Field;Knowledge Field|FIELD
Procedure|Health Care Activity|SIMPLE_SEGMENT|5443,5448|false|false|false|C1553496|field - patient encounter|FIELD
Event|Event|SIMPLE_SEGMENT|5453,5470|false|false|false|||POLYMORPHONUCLEAR
Anatomy|Cell|SIMPLE_SEGMENT|5472,5482|false|false|false|C0023516|Leukocytes|LEUKOCYTES
Event|Event|SIMPLE_SEGMENT|5472,5482|false|false|false|||LEUKOCYTES
Finding|Body Substance|SIMPLE_SEGMENT|5472,5482|false|false|false|C1547962;C1550647|Specimen Type - Leukocytes|LEUKOCYTES
Finding|Intellectual Product|SIMPLE_SEGMENT|5472,5482|false|false|false|C1547962;C1550647|Specimen Type - Leukocytes|LEUKOCYTES
Finding|Finding|SIMPLE_SEGMENT|5494,5513|false|false|false|C2924473|Microorganisms seen|MICROORGANISMS SEEN
Event|Event|SIMPLE_SEGMENT|5509,5513|false|false|false|||SEEN
Event|Activity|SIMPLE_SEGMENT|5545,5550|false|false|false|C1947932|Smear - instruction imperative|smear
Event|Event|SIMPLE_SEGMENT|5545,5550|false|false|false|||smear
Finding|Functional Concept|SIMPLE_SEGMENT|5545,5550|false|false|false|C3872789|Smearing technique|smear
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5545,5550|false|false|false|C0444186|Smear test|smear
Event|Event|SIMPLE_SEGMENT|5568,5574|false|false|false|||method
Finding|Functional Concept|SIMPLE_SEGMENT|5568,5574|false|false|false|C0025663;C0449851;C2828387|Method, LOINC Axis 6;Methods;Techniques|method
Finding|Intellectual Product|SIMPLE_SEGMENT|5568,5574|false|false|false|C0025663;C0449851;C2828387|Method, LOINC Axis 6;Methods;Techniques|method
Event|Event|SIMPLE_SEGMENT|5599,5609|false|false|false|||hematology
Finding|Intellectual Product|SIMPLE_SEGMENT|5599,5609|false|false|false|C1547985|Diagnostic Service Section ID - Hematology|hematology
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5599,5609|false|false|false|C0018941;C0200627;C2183233|Hematologic Tests;Hematology procedure;diagnostic service sources hematology (procedure)|hematology
Anatomy|Cell|SIMPLE_SEGMENT|5629,5645|false|false|false|C0023516|Leukocytes|white blood cell
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5629,5651|false|false|false|C0427512||white blood cell count
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5629,5651|false|false|false|C0023508|White Blood Cell Count procedure|white blood cell count
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5635,5640|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|SIMPLE_SEGMENT|5635,5640|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Anatomy|Cell|SIMPLE_SEGMENT|5635,5645|false|false|false|C0005773|Blood Cells|blood cell
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5635,5651|false|false|false|C0005771;C0009555|Blood Cell Count;Complete Blood Count|blood cell count
Anatomy|Cell|SIMPLE_SEGMENT|5641,5645|false|false|false|C0007634|Cells|cell
Finding|Gene or Genome|SIMPLE_SEGMENT|5641,5645|false|false|false|C1413336;C1413337|CEL gene;CELP gene|cell
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5641,5651|false|false|false|C0007584|Cell Count|cell count
Event|Event|SIMPLE_SEGMENT|5646,5651|false|false|false|||count
Drug|Substance|SIMPLE_SEGMENT|5659,5664|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|FLUID
Event|Event|SIMPLE_SEGMENT|5659,5664|false|false|false|||FLUID
Finding|Intellectual Product|SIMPLE_SEGMENT|5659,5664|false|false|false|C1546638|Fluid Specimen Code|FLUID
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5665,5672|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|SIMPLE_SEGMENT|5665,5672|false|false|false|||CULTURE
Finding|Functional Concept|SIMPLE_SEGMENT|5665,5672|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|SIMPLE_SEGMENT|5665,5672|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5665,5672|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Event|Event|SIMPLE_SEGMENT|5674,5679|false|false|false|||Final
Finding|Idea or Concept|SIMPLE_SEGMENT|5674,5679|false|false|false|C1546485|Diagnosis Type - Final|Final
Event|Event|SIMPLE_SEGMENT|5691,5697|false|false|false|||GROWTH
Finding|Finding|SIMPLE_SEGMENT|5691,5697|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|5691,5697|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organism Function|SIMPLE_SEGMENT|5691,5697|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Physiologic Function|SIMPLE_SEGMENT|5691,5697|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|5691,5697|true|false|false|C2911660|Growth action|GROWTH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5704,5721|false|false|false|C1273935|Anaerobic microbial culture|ANAEROBIC CULTURE
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5714,5721|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|SIMPLE_SEGMENT|5714,5721|false|false|false|||CULTURE
Finding|Functional Concept|SIMPLE_SEGMENT|5714,5721|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|SIMPLE_SEGMENT|5714,5721|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5714,5721|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Event|Event|SIMPLE_SEGMENT|5743,5749|false|false|false|||GROWTH
Finding|Finding|SIMPLE_SEGMENT|5743,5749|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|5743,5749|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organism Function|SIMPLE_SEGMENT|5743,5749|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Physiologic Function|SIMPLE_SEGMENT|5743,5749|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|5743,5749|true|false|false|C2911660|Growth action|GROWTH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5753,5779|false|false|false|C2721555|Legionella urinary antigen|Legionella Urinary Antigen
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5764,5771|false|false|false|C0042027|Urinary tract|Urinary
Drug|Immunologic Factor|SIMPLE_SEGMENT|5772,5779|false|false|false|C0003320|Antigens|Antigen
Event|Event|SIMPLE_SEGMENT|5772,5779|false|false|false|||Antigen
Event|Event|SIMPLE_SEGMENT|5787,5790|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|5787,5790|false|false|false|C5848551|Neg - answer|NEG
Event|Event|SIMPLE_SEGMENT|5795,5805|false|false|false|||LEGIONELLA
Finding|Intellectual Product|SIMPLE_SEGMENT|5807,5816|false|false|false|C0449543|Serogroup|SEROGROUP
Finding|Body Substance|SIMPLE_SEGMENT|5826,5831|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Finding|Functional Concept|SIMPLE_SEGMENT|5826,5831|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Finding|Intellectual Product|SIMPLE_SEGMENT|5826,5831|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5826,5839|false|false|false|C0430404|Urine culture|Urine Culture
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5832,5839|false|false|false|C1706355|Culture Dose Form|Culture
Event|Event|SIMPLE_SEGMENT|5832,5839|false|false|false|||Culture
Finding|Functional Concept|SIMPLE_SEGMENT|5832,5839|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|Culture
Finding|Idea or Concept|SIMPLE_SEGMENT|5832,5839|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|Culture
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5832,5839|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|Culture
Event|Event|SIMPLE_SEGMENT|5841,5849|false|false|false|||negative
Finding|Classification|SIMPLE_SEGMENT|5841,5849|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|5841,5849|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5841,5849|false|false|false|C5237010|Expression Negative|negative
Drug|Food|SIMPLE_SEGMENT|5853,5858|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|yeast
Drug|Immunologic Factor|SIMPLE_SEGMENT|5853,5858|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|yeast
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|5853,5858|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|yeast
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5853,5858|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|yeast
Event|Event|SIMPLE_SEGMENT|5853,5858|false|false|false|||yeast
Event|Event|SIMPLE_SEGMENT|5871,5879|false|false|false|||cultures
Finding|Idea or Concept|SIMPLE_SEGMENT|5871,5879|true|true|false|C0010453|Culture (Anthropological)|cultures
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5881,5886|false|false|false|C0851353|Blood and lymphatic system disorders|Blood
Event|Event|SIMPLE_SEGMENT|5881,5886|false|false|false|||Blood
Finding|Body Substance|SIMPLE_SEGMENT|5881,5886|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5881,5895|false|true|false|C0200949|Blood culture|Blood Cultures
Event|Event|SIMPLE_SEGMENT|5887,5895|false|false|false|||Cultures
Finding|Idea or Concept|SIMPLE_SEGMENT|5887,5895|false|false|false|C0010453|Culture (Anthropological)|Cultures
Event|Event|SIMPLE_SEGMENT|5897,5901|false|false|false|||NGTD
Event|Event|SIMPLE_SEGMENT|5905,5913|false|false|false|||negative
Finding|Classification|SIMPLE_SEGMENT|5905,5913|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|5905,5913|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5905,5913|false|false|false|C5237010|Expression Negative|negative
Event|Event|SIMPLE_SEGMENT|5926,5934|false|false|false|||cultures
Finding|Idea or Concept|SIMPLE_SEGMENT|5926,5934|true|true|false|C0010453|Culture (Anthropological)|cultures
Event|Event|SIMPLE_SEGMENT|5936,5943|false|false|false|||Imaging
Finding|Finding|SIMPLE_SEGMENT|5936,5943|false|false|false|C0740845|Imaging problem|Imaging
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5936,5943|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|Imaging
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5945,5951|false|false|false|C1644645||CT Abd
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5948,5951|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|Abd
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|5948,5951|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|Abd
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|5964,5972|false|false|false|C0009924|Contrast Media|Contrast
Event|Event|SIMPLE_SEGMENT|5964,5972|false|false|false|||Contrast
Event|Event|SIMPLE_SEGMENT|5980,5990|false|false|false|||IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|5980,5990|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|5980,5990|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6004,6011|false|false|false|C0009368|Colon structure (body structure)|colonic
Anatomy|Tissue|SIMPLE_SEGMENT|6012,6019|false|false|false|C0026724|Mucous Membrane|mucosal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6041,6046|false|false|false|C0021853|Intestines|bowel
Event|Event|SIMPLE_SEGMENT|6053,6063|false|false|false|||thickening
Finding|Finding|SIMPLE_SEGMENT|6053,6063|false|false|false|C0205400|Thickened|thickening
Event|Event|SIMPLE_SEGMENT|6067,6077|false|false|false|||consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|6067,6077|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|6067,6082|false|false|false|C0332290|Consistent with|consistent with
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6083,6093|false|false|false|C0868908|Pancolitis|pancolitis
Event|Event|SIMPLE_SEGMENT|6083,6093|false|false|false|||pancolitis
Finding|Finding|SIMPLE_SEGMENT|6099,6121|false|false|false|C5539411|Ground glass opacity|Ground-glass opacities
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6106,6111|false|false|false|C2676739|Chromosome 2q32-Q33 Deletion Syndrome|glass
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|6106,6111|false|false|false|C0025611|methamphetamine|glass
Drug|Organic Chemical|SIMPLE_SEGMENT|6106,6111|false|false|false|C0025611|methamphetamine|glass
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6106,6111|false|false|false|C0025611|methamphetamine|glass
Event|Event|SIMPLE_SEGMENT|6112,6121|false|false|false|||opacities
Finding|Finding|SIMPLE_SEGMENT|6112,6121|false|false|false|C0029053;C1265876|Abnormally opaque structure (morphologic abnormality);Decreased translucency|opacities
Finding|Pathologic Function|SIMPLE_SEGMENT|6112,6121|false|false|false|C0029053;C1265876|Abnormally opaque structure (morphologic abnormality);Decreased translucency|opacities
Finding|Functional Concept|SIMPLE_SEGMENT|6133,6138|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Finding|Intellectual Product|SIMPLE_SEGMENT|6139,6145|false|false|false|C1552826|Table Cell Vertical Align - middle|middle
Finding|Functional Concept|SIMPLE_SEGMENT|6150,6155|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6157,6162|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|6157,6162|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6163,6168|false|false|false|C0796494|lobe|lobes
Event|Event|SIMPLE_SEGMENT|6169,6179|false|false|false|||compatible
Finding|Idea or Concept|SIMPLE_SEGMENT|6169,6179|false|false|false|C0332290|Consistent with|compatible
Finding|Idea or Concept|SIMPLE_SEGMENT|6169,6184|false|false|false|C0332290|Consistent with|compatible with
Finding|Intellectual Product|SIMPLE_SEGMENT|6185,6190|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6185,6200|false|false|false|C0275518|Acute infectious disease|acute infection
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6191,6200|false|true|false|C0009450|Communicable Diseases|infection
Event|Event|SIMPLE_SEGMENT|6191,6200|false|false|false|||infection
Finding|Pathologic Function|SIMPLE_SEGMENT|6191,6200|false|true|false|C3714514|Infection|infection
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|6208,6218|false|false|false|C1720922|Respiratory Aspiration|aspiration
Event|Event|SIMPLE_SEGMENT|6208,6218|false|false|false|||aspiration
Finding|Finding|SIMPLE_SEGMENT|6208,6218|false|false|false|C0220787;C0700198;C2712334|Aspiration into respiratory tract;Endotracheal aspiration;Pulmonary aspiration|aspiration
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|6208,6218|false|false|false|C0220787;C0700198;C2712334|Aspiration into respiratory tract;Endotracheal aspiration;Pulmonary aspiration|aspiration
Finding|Pathologic Function|SIMPLE_SEGMENT|6208,6218|false|false|false|C0220787;C0700198;C2712334|Aspiration into respiratory tract;Endotracheal aspiration;Pulmonary aspiration|aspiration
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6208,6218|false|false|false|C0349707||aspiration
Finding|Finding|SIMPLE_SEGMENT|6221,6229|false|false|false|C0332149|Possible|Possible
Finding|Intellectual Product|SIMPLE_SEGMENT|6231,6235|false|false|false|C1547225|Mild Severity of Illness Code|mild
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6236,6245|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6236,6245|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|6236,6245|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6246,6251|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|6246,6251|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|6246,6251|false|false|false|C0013604|Edema|edema
Finding|Functional Concept|SIMPLE_SEGMENT|6257,6269|false|false|false|C1512952|Intrahepatic Route of Administration|Intrahepatic
Finding|Functional Concept|SIMPLE_SEGMENT|6270,6277|false|false|false|C0521378|Biliary|biliary
Event|Event|SIMPLE_SEGMENT|6285,6295|false|false|false|||dilatation
Finding|Finding|SIMPLE_SEGMENT|6285,6295|false|false|false|C0012359;C0700124|Dilated;Pathological Dilatation|dilatation
Finding|Pathologic Function|SIMPLE_SEGMENT|6285,6295|false|false|false|C0012359;C0700124|Dilated;Pathological Dilatation|dilatation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6285,6295|false|false|false|C1322279|Dilate procedure|dilatation
Event|Event|SIMPLE_SEGMENT|6300,6310|false|false|false|||prominence
Finding|Functional Concept|SIMPLE_SEGMENT|6319,6325|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Finding|Intellectual Product|SIMPLE_SEGMENT|6319,6325|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Event|Event|SIMPLE_SEGMENT|6326,6330|false|false|false|||bile
Finding|Body Substance|SIMPLE_SEGMENT|6326,6330|false|false|false|C0005388|Bile fluid|bile
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6335,6345|false|false|false|C0030274|Pancreas|pancreatic
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6335,6345|false|false|false|C0030292|Pancreatic Hormones|pancreatic
Drug|Hormone|SIMPLE_SEGMENT|6335,6345|false|false|false|C0030292|Pancreatic Hormones|pancreatic
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6335,6345|false|false|false|C0030292|Pancreatic Hormones|pancreatic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6335,6351|false|false|false|C0030288|Pancreatic duct|pancreatic ducts
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6346,6351|false|false|false|C0687028|Duct (organ) structure|ducts
Finding|Idea or Concept|SIMPLE_SEGMENT|6361,6367|false|true|false|C1550462|Observation Interpretation - better|better
Event|Activity|SIMPLE_SEGMENT|6368,6381|false|true|false|C1880022|Characterization|characterized
Event|Event|SIMPLE_SEGMENT|6368,6381|false|false|false|||characterized
Event|Event|SIMPLE_SEGMENT|6401,6405|false|false|false|||MRCP
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6401,6405|false|false|false|C0994163|Cholangiopancreatography, Magnetic Resonance|MRCP
Event|Event|SIMPLE_SEGMENT|6408,6411|false|false|false|||CXR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6408,6411|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|SIMPLE_SEGMENT|6419,6429|false|false|false|||IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|6419,6429|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|6419,6429|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Event|Event|SIMPLE_SEGMENT|6445,6454|false|false|false|||opacities
Finding|Finding|SIMPLE_SEGMENT|6445,6454|false|false|false|C0029053;C1265876|Abnormally opaque structure (morphologic abnormality);Decreased translucency|opacities
Finding|Pathologic Function|SIMPLE_SEGMENT|6445,6454|false|false|false|C0029053;C1265876|Abnormally opaque structure (morphologic abnormality);Decreased translucency|opacities
Event|Event|SIMPLE_SEGMENT|6464,6474|false|false|false|||consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|6464,6474|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|6464,6479|false|false|false|C0332290|Consistent with|consistent with
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6480,6489|false|true|false|C0032285|Pneumonia|pneumonia
Event|Event|SIMPLE_SEGMENT|6480,6489|false|false|false|||pneumonia
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|6498,6508|false|false|false|C1720922|Respiratory Aspiration|aspiration
Event|Event|SIMPLE_SEGMENT|6498,6508|false|false|false|||aspiration
Finding|Finding|SIMPLE_SEGMENT|6498,6508|false|false|false|C0220787;C0700198;C2712334|Aspiration into respiratory tract;Endotracheal aspiration;Pulmonary aspiration|aspiration
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|6498,6508|false|false|false|C0220787;C0700198;C2712334|Aspiration into respiratory tract;Endotracheal aspiration;Pulmonary aspiration|aspiration
Finding|Pathologic Function|SIMPLE_SEGMENT|6498,6508|false|false|false|C0220787;C0700198;C2712334|Aspiration into respiratory tract;Endotracheal aspiration;Pulmonary aspiration|aspiration
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6498,6508|false|false|false|C0349707||aspiration
Finding|Functional Concept|SIMPLE_SEGMENT|6516,6521|false|true|false|C1552823|Table Cell Horizontal Align - right|right
Finding|Intellectual Product|SIMPLE_SEGMENT|6522,6530|false|false|false|C1315013|Clinical NEC (not elsewhere classified in LNC)|clinical
Event|Event|SIMPLE_SEGMENT|6531,6538|false|false|false|||setting
Finding|Mental Process|SIMPLE_SEGMENT|6531,6538|false|false|false|C0542559|contextual factors|setting
Finding|Finding|SIMPLE_SEGMENT|6541,6547|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Finding|Idea or Concept|SIMPLE_SEGMENT|6541,6547|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6554,6563|false|false|false|C1179435|Protein Component|component
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6554,6563|false|false|false|C1179435|Protein Component|component
Event|Event|SIMPLE_SEGMENT|6554,6563|false|false|false|||component
Finding|Conceptual Entity|SIMPLE_SEGMENT|6554,6563|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Finding|Idea or Concept|SIMPLE_SEGMENT|6554,6563|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Finding|Intellectual Product|SIMPLE_SEGMENT|6554,6563|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6567,6576|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6567,6576|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|6567,6576|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|SIMPLE_SEGMENT|6567,6582|false|false|false|C0034063|Pulmonary Edema|pulmonary edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6577,6582|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|6577,6582|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|6577,6582|false|false|false|C0013604|Edema|edema
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6593,6605|false|false|false|C0596790|interstitial|interstitial
Finding|Functional Concept|SIMPLE_SEGMENT|6593,6605|false|false|false|C1522203|Interstitial Route of Administration|interstitial
Finding|Finding|SIMPLE_SEGMENT|6593,6616|false|false|false|C2750120|Interstitial thickening|interstitial thickening
Event|Event|SIMPLE_SEGMENT|6606,6616|false|false|false|||thickening
Finding|Finding|SIMPLE_SEGMENT|6606,6616|false|false|false|C0205400|Thickened|thickening
Finding|Finding|SIMPLE_SEGMENT|6631,6638|false|false|false|C0700124|Dilated|dilated
Finding|Finding|SIMPLE_SEGMENT|6631,6644|false|false|false|C4697734|Dilated loops|dilated loops
Event|Event|SIMPLE_SEGMENT|6639,6644|false|false|false|||loops
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6648,6659|false|false|false|C0021852;C4319010|Abdomen>Small bowel;Intestines, Small|small bowel
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6648,6659|false|false|false|C0021852;C4319010|Abdomen>Small bowel;Intestines, Small|small bowel
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6654,6659|false|false|false|C0021853|Intestines|bowel
Event|Event|SIMPLE_SEGMENT|6664,6673|false|false|false|||represent
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6674,6679|false|false|false|C1258215;C4019039|Ileus;Intestinal obstruction co-occurrent and due to decreased peristalsis|ileus
Event|Event|SIMPLE_SEGMENT|6674,6679|false|false|false|||ileus
Event|Event|SIMPLE_SEGMENT|6684,6695|false|false|false|||obstruction
Finding|Finding|SIMPLE_SEGMENT|6684,6695|false|false|false|C0028778|Obstruction|obstruction
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6707,6716|false|false|false|C0000726|Abdomen|abdominal
Event|Event|SIMPLE_SEGMENT|6717,6727|false|false|false|||radiograph
Finding|Intellectual Product|SIMPLE_SEGMENT|6717,6727|false|false|false|C1548003|Diagnostic Service Section ID - Radiograph|radiograph
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6717,6727|false|false|false|C1306645|Plain x-ray|radiograph
Finding|Idea or Concept|SIMPLE_SEGMENT|6750,6756|false|false|false|C1550462|Observation Interpretation - better|better
Event|Activity|SIMPLE_SEGMENT|6757,6773|false|false|false|C1880022|Characterization|characterization
Event|Event|SIMPLE_SEGMENT|6757,6773|false|false|false|||characterization
Event|Event|SIMPLE_SEGMENT|6776,6780|false|false|false|||ECHO
Procedure|Health Care Activity|SIMPLE_SEGMENT|6776,6780|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6776,6780|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Finding|Functional Concept|SIMPLE_SEGMENT|6788,6792|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6788,6809|false|false|false|C0504053|Wall of left ventricle|Left ventricular wall
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6793,6804|false|false|false|C0018827|Heart Ventricle|ventricular
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6793,6809|false|false|false|C0507618|Wall of ventricle|ventricular wall
Event|Event|SIMPLE_SEGMENT|6810,6821|false|false|false|||thicknesses
Event|Event|SIMPLE_SEGMENT|6826,6832|false|false|false|||normal
Finding|Functional Concept|SIMPLE_SEGMENT|6834,6838|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6839,6850|false|false|false|C0018827|Heart Ventricle|ventricular
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|6852,6860|false|false|false|C0039155|Systole|systolic
Event|Event|SIMPLE_SEGMENT|6861,6869|false|false|false|||function
Finding|Finding|SIMPLE_SEGMENT|6861,6869|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|SIMPLE_SEGMENT|6861,6869|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|SIMPLE_SEGMENT|6861,6869|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|SIMPLE_SEGMENT|6861,6869|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Event|Event|SIMPLE_SEGMENT|6873,6885|false|false|false|||hyperdynamic
Finding|Intellectual Product|SIMPLE_SEGMENT|6907,6911|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Functional Concept|SIMPLE_SEGMENT|6921,6925|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6921,6945|false|false|false|C0225912|Outflow tract of left ventricle|left ventricular outflow
Finding|Finding|SIMPLE_SEGMENT|6921,6945|false|false|false|C0455821|Left ventricular outflow|left ventricular outflow
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6921,6951|false|false|false|C1305766;C4284103|Left Ventricular Outflow Tract|left ventricular outflow tract
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6921,6951|false|false|false|C5212772|Blood flow velocity.max.left ventricular outflow tract|left ventricular outflow tract
Finding|Finding|SIMPLE_SEGMENT|6921,6951|false|false|false|C4288824|Left Ventricular Outflow Tract Velocity Time Integral|left ventricular outflow tract
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6921,6963|false|false|false|C0023213|Ventricular Outflow Obstruction, Left|left ventricular outflow tract obstruction
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6926,6937|false|false|false|C0018827|Heart Ventricle|ventricular
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|6926,6951|false|false|false|C0507070|Outflow part of ventricle|ventricular outflow tract
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6946,6951|false|false|false|C1185740|Tract|tract
Event|Event|SIMPLE_SEGMENT|6952,6963|false|false|false|||obstruction
Finding|Finding|SIMPLE_SEGMENT|6952,6963|false|false|false|C0028778|Obstruction|obstruction
Finding|Functional Concept|SIMPLE_SEGMENT|6965,6970|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6972,6983|false|false|false|C0018827|Heart Ventricle|ventricular
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6984,6991|false|false|false|C0935616|chamber [body part]|chamber
Event|Event|SIMPLE_SEGMENT|6992,6996|false|false|false|||size
Event|Event|SIMPLE_SEGMENT|7001,7005|false|false|false|||free
Finding|Functional Concept|SIMPLE_SEGMENT|7001,7005|false|false|false|C0332296|Free of (attribute)|free
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7006,7017|false|false|false|C1980023|Wall motion|wall motion
Event|Event|SIMPLE_SEGMENT|7011,7017|false|false|false|||motion
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|7011,7017|false|false|false|C0026597|Motion|motion
Event|Event|SIMPLE_SEGMENT|7022,7028|false|false|false|||normal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7035,7041|false|false|false|C0003483|Aorta|aortic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7035,7047|false|false|false|C0003501;C4533215|Aortic valve structure;Chest>Aortic valve|aortic valve
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7042,7047|false|false|false|C1186983|Anatomical valve|valve
Event|Event|SIMPLE_SEGMENT|7048,7056|false|false|false|||leaflets
Event|Event|SIMPLE_SEGMENT|7072,7081|false|false|false|||thickened
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7087,7099|false|false|false|C0026264|Mitral Valve|mitral valve
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7094,7099|false|false|false|C1186983|Anatomical valve|valve
Event|Event|SIMPLE_SEGMENT|7101,7109|false|false|false|||leaflets
Event|Event|SIMPLE_SEGMENT|7121,7130|false|false|false|||thickened
Finding|Finding|SIMPLE_SEGMENT|7141,7147|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|SIMPLE_SEGMENT|7141,7147|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Event|Event|SIMPLE_SEGMENT|7164,7177|false|false|false|||calcification
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|7164,7177|false|false|false|C0006660;C0006663;C1533591|Calcification;Calcinosis;Physiologic calcification|calcification
Finding|Pathologic Function|SIMPLE_SEGMENT|7164,7177|false|false|false|C0006660;C0006663;C1533591|Calcification;Calcinosis;Physiologic calcification|calcification
Finding|Finding|SIMPLE_SEGMENT|7188,7196|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|SIMPLE_SEGMENT|7188,7196|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Conceptual Entity|SIMPLE_SEGMENT|7197,7207|false|false|false|C0205245;C0542341;C2700217|Function (attribute);Functional;Functional Relationship|functional
Finding|Functional Concept|SIMPLE_SEGMENT|7197,7207|false|false|false|C0205245;C0542341;C2700217|Function (attribute);Functional;Functional Relationship|functional
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7208,7223|false|false|false|C0026269;C0264766|Mitral Valve Stenosis;Rheumatic mitral stenosis|mitral stenosis
Event|Event|SIMPLE_SEGMENT|7215,7223|false|false|false|||stenosis
Finding|Pathologic Function|SIMPLE_SEGMENT|7215,7223|false|false|false|C1261287|Stenosis|stenosis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7255,7283|false|false|false|C0428811|Mitral valve annular calcification|mitral annular calcification
Finding|Finding|SIMPLE_SEGMENT|7255,7283|false|false|false|C1835130|Premature calcification of mitral annulus|mitral annular calcification
Event|Event|SIMPLE_SEGMENT|7270,7283|false|false|false|||calcification
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|7270,7283|false|false|false|C0006660;C0006663;C1533591|Calcification;Calcinosis;Physiologic calcification|calcification
Finding|Pathologic Function|SIMPLE_SEGMENT|7270,7283|false|false|false|C0006660;C0006663;C1533591|Calcification;Calcinosis;Physiologic calcification|calcification
Finding|Intellectual Product|SIMPLE_SEGMENT|7285,7289|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Finding|Finding|SIMPLE_SEGMENT|7294,7302|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|SIMPLE_SEGMENT|7294,7302|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7309,7329|false|false|false|C0026266|Mitral Valve Insufficiency|mitral regurgitation
Event|Event|SIMPLE_SEGMENT|7316,7329|false|false|false|||regurgitation
Finding|Finding|SIMPLE_SEGMENT|7316,7329|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|SIMPLE_SEGMENT|7316,7329|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|SIMPLE_SEGMENT|7316,7329|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Event|Event|SIMPLE_SEGMENT|7333,7337|false|false|false|||seen
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|7348,7356|false|false|false|C0001166|Acoustics|acoustic
Finding|Finding|SIMPLE_SEGMENT|7348,7366|false|false|false|C1719833|Acoustic shadowing|acoustic shadowing
Event|Event|SIMPLE_SEGMENT|7357,7366|false|false|false|||shadowing
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7357,7366|false|false|false|C0085195;C0600111|Shadowing (Histology);Shadowing (regime/therapy)|shadowing
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7357,7366|false|false|false|C0085195;C0600111|Shadowing (Histology);Shadowing (regime/therapy)|shadowing
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7384,7404|false|false|false|C0026266|Mitral Valve Insufficiency|mitral regurgitation
Event|Event|SIMPLE_SEGMENT|7391,7404|false|false|false|||regurgitation
Finding|Finding|SIMPLE_SEGMENT|7391,7404|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|SIMPLE_SEGMENT|7391,7404|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|SIMPLE_SEGMENT|7391,7404|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Event|Event|SIMPLE_SEGMENT|7427,7441|false|false|false|||UNDERestimated
Finding|Functional Concept|SIMPLE_SEGMENT|7448,7452|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7453,7464|false|false|false|C0018827|Heart Ventricle|ventricular
Event|Event|SIMPLE_SEGMENT|7465,7471|false|false|false|||inflow
Event|Event|SIMPLE_SEGMENT|7473,7480|false|false|false|||pattern
Event|Event|SIMPLE_SEGMENT|7481,7489|false|false|false|||suggests
Event|Event|SIMPLE_SEGMENT|7490,7498|false|false|false|||impaired
Event|Activity|SIMPLE_SEGMENT|7499,7509|false|false|false|C0035028|Relaxation|relaxation
Event|Event|SIMPLE_SEGMENT|7499,7509|false|false|false|||relaxation
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7515,7530|false|false|false|C0040960|Tricuspid valve structure|tricuspid valve
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7525,7530|false|false|false|C1186983|Anatomical valve|valve
Event|Event|SIMPLE_SEGMENT|7532,7540|false|false|false|||leaflets
Event|Event|SIMPLE_SEGMENT|7552,7561|false|false|false|||thickened
Finding|Finding|SIMPLE_SEGMENT|7563,7571|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Intellectual Product|SIMPLE_SEGMENT|7563,7571|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Event|Event|SIMPLE_SEGMENT|7588,7601|false|false|false|||regurgitation
Finding|Finding|SIMPLE_SEGMENT|7588,7601|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|SIMPLE_SEGMENT|7588,7601|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|SIMPLE_SEGMENT|7588,7601|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Event|Event|SIMPLE_SEGMENT|7605,7609|false|false|false|||seen
Finding|Intellectual Product|SIMPLE_SEGMENT|7620,7624|false|false|false|C1547225|Mild Severity of Illness Code|mild
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7625,7634|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7625,7634|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|7625,7634|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7625,7641|false|false|false|C0034052|Pulmonary artery structure|pulmonary artery
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7635,7641|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|SIMPLE_SEGMENT|7635,7641|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Event|Event|SIMPLE_SEGMENT|7642,7650|false|false|false|||systolic
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|7642,7650|false|false|false|C0039155|Systole|systolic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7652,7664|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|SIMPLE_SEGMENT|7652,7664|false|false|false|||hypertension
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7678,7689|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7678,7689|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7678,7698|true|false|false|C0031039|Pericardial effusion|pericardial effusion
Finding|Body Substance|SIMPLE_SEGMENT|7678,7698|true|false|false|C1253937|Pericardial effusion body substance|pericardial effusion
Event|Event|SIMPLE_SEGMENT|7690,7698|false|false|false|||effusion
Finding|Body Substance|SIMPLE_SEGMENT|7690,7698|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|SIMPLE_SEGMENT|7690,7698|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|7690,7698|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Event|Event|SIMPLE_SEGMENT|7725,7730|false|false|false|||study
Finding|Intellectual Product|SIMPLE_SEGMENT|7725,7730|false|false|false|C1705923|Study Object|study
Procedure|Research Activity|SIMPLE_SEGMENT|7725,7730|false|false|false|C0008972;C0947630;C2603343|Clinical Research;Scientific Study;Study|study
Event|Event|SIMPLE_SEGMENT|7739,7747|false|false|false|||reviewed
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7758,7778|false|false|false|C0026266|Mitral Valve Insufficiency|mitral regurgitation
Event|Event|SIMPLE_SEGMENT|7765,7778|false|false|false|||regurgitation
Finding|Finding|SIMPLE_SEGMENT|7765,7778|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|SIMPLE_SEGMENT|7765,7778|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|SIMPLE_SEGMENT|7765,7778|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Event|Event|SIMPLE_SEGMENT|7791,7800|false|false|false|||prominent
Event|Event|SIMPLE_SEGMENT|7821,7829|false|false|false|||gradient
Event|Event|SIMPLE_SEGMENT|7833,7840|false|false|false|||similar
Event|Event|SIMPLE_SEGMENT|7855,7863|false|false|false|||reported
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7881,7887|false|false|false|C4255046||report
Event|Event|SIMPLE_SEGMENT|7881,7887|false|false|false|||report
Finding|Intellectual Product|SIMPLE_SEGMENT|7881,7887|false|false|false|C0684224|Report (document)|report
Procedure|Health Care Activity|SIMPLE_SEGMENT|7881,7887|false|false|false|C0700287|Reporting|report
Event|Event|SIMPLE_SEGMENT|7892,7895|false|false|false|||AXR
Finding|Finding|SIMPLE_SEGMENT|7915,7940|true|false|false|C0749093|SUBDIAPHRAGMATIC FREE AIR|subdiaphragmatic free air
Finding|Functional Concept|SIMPLE_SEGMENT|7932,7936|false|false|false|C0332296|Free of (attribute)|free
Drug|Inorganic Chemical|SIMPLE_SEGMENT|7937,7940|true|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7937,7940|true|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|SIMPLE_SEGMENT|7937,7940|true|false|false|C0001861;C3536832|Air (substance);air|air
Event|Event|SIMPLE_SEGMENT|7937,7940|false|false|false|||air
Finding|Finding|SIMPLE_SEGMENT|7937,7940|true|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|SIMPLE_SEGMENT|7937,7940|true|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|SIMPLE_SEGMENT|7937,7940|true|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Finding|SIMPLE_SEGMENT|7963,7972|false|false|false|C0700124|Dilated|distended
Event|Event|SIMPLE_SEGMENT|7973,7978|false|false|false|||loops
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7982,7987|false|false|false|C0021853|Intestines|bowel
Finding|Idea or Concept|SIMPLE_SEGMENT|7989,8000|false|false|false|C0750501|most likely|most likely
Finding|Finding|SIMPLE_SEGMENT|7994,8000|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|7994,8000|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|SIMPLE_SEGMENT|8001,8013|false|false|false|||representing
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8019,8024|false|false|false|C0009368;C4071907|Abdomen+Pelvis>Colon;Colon structure (body structure)|colon
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8019,8024|false|true|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Disorder|Neoplastic Process|SIMPLE_SEGMENT|8019,8024|false|true|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Event|Event|SIMPLE_SEGMENT|8019,8024|false|false|false|||colon
Finding|Finding|SIMPLE_SEGMENT|8019,8024|false|true|false|C0750873|COLON PROBLEM|colon
Anatomy|Body Location or Region|SIMPLE_SEGMENT|8030,8041|false|false|false|C0021852;C4319010|Abdomen>Small bowel;Intestines, Small|small bowel
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8030,8041|false|false|false|C0021852;C4319010|Abdomen>Small bowel;Intestines, Small|small bowel
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8036,8041|false|false|false|C0021853|Intestines|bowel
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8044,8052|false|false|false|C2926606||Findings
Event|Event|SIMPLE_SEGMENT|8044,8052|false|false|false|||Findings
Finding|Functional Concept|SIMPLE_SEGMENT|8044,8052|false|false|false|C2607943|findings aspects|Findings
Event|Event|SIMPLE_SEGMENT|8062,8072|false|false|false|||consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|8062,8072|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|8062,8077|false|false|false|C0332290|Consistent with|consistent with
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8081,8086|false|false|false|C1258215;C4019039|Ileus;Intestinal obstruction co-occurrent and due to decreased peristalsis|ileus
Event|Event|SIMPLE_SEGMENT|8081,8086|false|false|false|||ileus
Drug|Inorganic Chemical|SIMPLE_SEGMENT|8090,8093|true|false|false|C0001861;C3536832|Air (substance);air|Air
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8090,8093|true|false|false|C0001861;C3536832|Air (substance);air|Air
Drug|Substance|SIMPLE_SEGMENT|8090,8093|true|false|false|C0001861;C3536832|Air (substance);air|Air
Event|Event|SIMPLE_SEGMENT|8090,8093|false|false|false|||Air
Finding|Finding|SIMPLE_SEGMENT|8090,8093|true|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|Air
Finding|Gene or Genome|SIMPLE_SEGMENT|8090,8093|true|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|Air
Finding|Intellectual Product|SIMPLE_SEGMENT|8090,8093|true|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|Air
Drug|Substance|SIMPLE_SEGMENT|8094,8099|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|8094,8099|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|8100,8106|false|false|false|||levels
Event|Event|SIMPLE_SEGMENT|8111,8115|false|false|false|||seen
Finding|Functional Concept|SIMPLE_SEGMENT|8123,8127|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8136,8145|false|false|false|C4554531|Pressure injury|decubitus
Event|Event|SIMPLE_SEGMENT|8152,8162|false|false|false|||IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|8152,8162|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|8152,8162|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Finding|SIMPLE_SEGMENT|8165,8172|false|false|false|C0700124|Dilated|Dilated
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8173,8178|false|false|false|C0009368;C4071907|Abdomen+Pelvis>Colon;Colon structure (body structure)|colon
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8173,8178|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Disorder|Neoplastic Process|SIMPLE_SEGMENT|8173,8178|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Event|Event|SIMPLE_SEGMENT|8173,8178|false|false|false|||colon
Finding|Finding|SIMPLE_SEGMENT|8173,8178|false|false|false|C0750873|COLON PROBLEM|colon
Anatomy|Body Location or Region|SIMPLE_SEGMENT|8183,8194|false|false|false|C0021852;C4319010|Abdomen>Small bowel;Intestines, Small|small bowel
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8183,8194|false|false|false|C0021852;C4319010|Abdomen>Small bowel;Intestines, Small|small bowel
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8189,8194|false|false|false|C0021853|Intestines|bowel
Event|Event|SIMPLE_SEGMENT|8195,8205|false|false|false|||consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|8195,8205|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|8195,8210|false|false|false|C0332290|Consistent with|consistent with
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8212,8217|false|false|false|C1258215;C4019039|Ileus;Intestinal obstruction co-occurrent and due to decreased peristalsis|ileus
Event|Event|SIMPLE_SEGMENT|8212,8217|false|false|false|||ileus
Anatomy|Body Location or Region|SIMPLE_SEGMENT|8220,8224|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|Head
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8220,8224|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|Head
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8220,8224|false|false|false|C0362076|Problems with head|Head
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8220,8224|false|false|false|C0876917|Procedure on head|Head
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8220,8227|false|false|false|C0202691|CAT scan of head|Head CT
Event|Event|SIMPLE_SEGMENT|8225,8227|false|false|false|||CT
Event|Event|SIMPLE_SEGMENT|8235,8245|false|false|false|||IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|8235,8245|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|8235,8245|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|8251,8256|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Anatomy|Body Location or Region|SIMPLE_SEGMENT|8257,8269|false|false|false|C0524466|Intracranial|intracranial
Finding|Functional Concept|SIMPLE_SEGMENT|8257,8269|false|false|false|C1522213|Intracranial Route of Administration|intracranial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8270,8277|false|false|false|C1184743|bony process|process
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8270,8277|true|false|false|C1951340|Process Pharmacologic Substance|process
Event|Event|SIMPLE_SEGMENT|8270,8277|false|false|false|||process
Finding|Functional Concept|SIMPLE_SEGMENT|8270,8277|true|false|false|C4521054|Process (qualifier value)|process
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|8270,8277|true|false|false|C1522240|Process|process
Event|Event|SIMPLE_SEGMENT|8280,8284|false|false|false|||ECHO
Procedure|Health Care Activity|SIMPLE_SEGMENT|8280,8284|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8280,8284|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Finding|Functional Concept|SIMPLE_SEGMENT|8296,8300|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8296,8307|false|false|false|C0225860|Left atrial structure|left atrium
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8301,8307|false|false|false|C0018792|Heart Atrium|atrium
Event|Event|SIMPLE_SEGMENT|8311,8317|false|false|false|||normal
Finding|Intellectual Product|SIMPLE_SEGMENT|8336,8340|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Conceptual Entity|SIMPLE_SEGMENT|8341,8350|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Finding|SIMPLE_SEGMENT|8341,8350|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Functional Concept|SIMPLE_SEGMENT|8351,8355|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8357,8368|false|false|false|C0018827|Heart Ventricle|ventricular
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8357,8380|false|false|false|C0340279|Ventricular hypertrophy|ventricular hypertrophy
Event|Event|SIMPLE_SEGMENT|8369,8380|false|false|false|||hypertrophy
Finding|Pathologic Function|SIMPLE_SEGMENT|8369,8380|false|false|false|C0020564|Hypertrophy|hypertrophy
Finding|Functional Concept|SIMPLE_SEGMENT|8386,8390|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|8386,8409|false|false|false|C0503990|Cavity of left ventricle|left ventricular cavity
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8391,8402|false|false|false|C0018827|Heart Ventricle|ventricular
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|8391,8409|false|false|false|C0507083|Cavity of ventricle|ventricular cavity
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|8403,8409|false|false|false|C0333343|Body cavities|cavity
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|8403,8409|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8403,8409|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Event|Event|SIMPLE_SEGMENT|8424,8429|false|false|false|||small
Finding|Functional Concept|SIMPLE_SEGMENT|8431,8435|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8436,8447|false|false|false|C0018827|Heart Ventricle|ventricular
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|8448,8456|false|false|false|C0039155|Systole|systolic
Event|Event|SIMPLE_SEGMENT|8457,8465|false|false|false|||function
Finding|Finding|SIMPLE_SEGMENT|8457,8465|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|SIMPLE_SEGMENT|8457,8465|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|SIMPLE_SEGMENT|8457,8465|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|SIMPLE_SEGMENT|8457,8465|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Event|Event|SIMPLE_SEGMENT|8470,8482|false|false|false|||hyperdynamic
Finding|Functional Concept|SIMPLE_SEGMENT|8493,8498|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8499,8510|false|false|false|C0018827|Heart Ventricle|ventricular
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8511,8518|false|false|false|C0935616|chamber [body part]|chamber
Event|Event|SIMPLE_SEGMENT|8528,8532|false|false|false|||free
Finding|Functional Concept|SIMPLE_SEGMENT|8528,8532|false|false|false|C0332296|Free of (attribute)|free
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8534,8545|false|false|false|C1980023|Wall motion|wall motion
Event|Event|SIMPLE_SEGMENT|8539,8545|false|false|false|||motion
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|8539,8545|false|false|false|C0026597|Motion|motion
Event|Event|SIMPLE_SEGMENT|8550,8556|false|false|false|||normal
Finding|Intellectual Product|SIMPLE_SEGMENT|8567,8571|false|false|false|C1547225|Mild Severity of Illness Code|mild
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8567,8593|false|false|false|C3276923|Mild aortic valve stenosis|mild aortic valve stenosis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8572,8578|false|false|false|C0003483|Aorta|aortic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8572,8584|false|false|false|C0003501;C4533215|Aortic valve structure;Chest>Aortic valve|aortic valve
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|8572,8593|false|false|false|C5193127;C5700069|AORTIC VALVE DISEASE 3;Stenosis of aorta|aortic valve stenosis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8572,8593|false|false|false|C5193127;C5700069|AORTIC VALVE DISEASE 3;Stenosis of aorta|aortic valve stenosis
Finding|Pathologic Function|SIMPLE_SEGMENT|8572,8593|false|false|false|C0003507|Aortic Valve Stenosis|aortic valve stenosis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8579,8584|false|false|false|C1186983|Anatomical valve|valve
Event|Event|SIMPLE_SEGMENT|8585,8593|false|false|false|||stenosis
Finding|Pathologic Function|SIMPLE_SEGMENT|8585,8593|false|false|false|C1261287|Stenosis|stenosis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8596,8601|false|false|false|C1186983|Anatomical valve|valve
Finding|Finding|SIMPLE_SEGMENT|8596,8606|false|false|false|C4687749|Valve Area|valve area
Event|Governmental or Regulatory Activity|SIMPLE_SEGMENT|8602,8606|false|false|false|C1510751|Academic Research Enhancement Awards|area
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|8611,8614|false|false|false|C0555206|Chiari malformation type II|cm2
Event|Event|SIMPLE_SEGMENT|8651,8657|false|false|false|||nature
Finding|Functional Concept|SIMPLE_SEGMENT|8651,8657|false|false|false|C0349590;C1262865|Nature;Natures|nature
Finding|Idea or Concept|SIMPLE_SEGMENT|8651,8657|false|false|false|C0349590;C1262865|Nature;Natures|nature
Event|Event|SIMPLE_SEGMENT|8667,8672|false|false|false|||study
Finding|Intellectual Product|SIMPLE_SEGMENT|8667,8672|false|false|false|C1705923|Study Object|study
Procedure|Research Activity|SIMPLE_SEGMENT|8667,8672|false|false|false|C0008972;C0947630;C2603343|Clinical Research;Scientific Study;Study|study
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8674,8690|false|false|false|C0023213|Ventricular Outflow Obstruction, Left|LVOT obstruction
Event|Event|SIMPLE_SEGMENT|8679,8690|false|false|false|||obstruction
Finding|Finding|SIMPLE_SEGMENT|8679,8690|false|true|false|C0028778|Obstruction|obstruction
Event|Event|SIMPLE_SEGMENT|8701,8709|false|false|false|||excluded
Event|Event|SIMPLE_SEGMENT|8716,8725|false|false|false|||certainty
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8731,8743|false|false|false|C0026264|Mitral Valve|mitral valve
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8738,8743|false|false|false|C1186983|Anatomical valve|valve
Event|Event|SIMPLE_SEGMENT|8744,8752|false|false|false|||leaflets
Event|Event|SIMPLE_SEGMENT|8764,8773|false|false|false|||thickened
Finding|Finding|SIMPLE_SEGMENT|8785,8791|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|SIMPLE_SEGMENT|8785,8791|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8792,8820|false|false|false|C0428811|Mitral valve annular calcification|mitral annular calcification
Finding|Finding|SIMPLE_SEGMENT|8792,8820|false|false|false|C1835130|Premature calcification of mitral annulus|mitral annular calcification
Event|Event|SIMPLE_SEGMENT|8807,8820|false|false|false|||calcification
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|8807,8820|false|false|false|C0006660;C0006663;C1533591|Calcification;Calcinosis;Physiologic calcification|calcification
Finding|Pathologic Function|SIMPLE_SEGMENT|8807,8820|false|false|false|C0006660;C0006663;C1533591|Calcification;Calcinosis;Physiologic calcification|calcification
Event|Event|SIMPLE_SEGMENT|8829,8836|false|false|false|||exclude
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8837,8846|false|true|false|C0751438|Posterior pituitary disease|posterior
Event|Event|SIMPLE_SEGMENT|8837,8846|false|false|false|||posterior
Finding|Intellectual Product|SIMPLE_SEGMENT|8848,8855|false|false|false|C3273178|Leaflet|leaflet
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8856,8859|false|false|false|C0026267|Mitral Valve Prolapse Syndrome|MVP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8856,8859|false|false|false|C1097902|MVP protein, human|MVP
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8856,8859|false|false|false|C1097902|MVP protein, human|MVP
Event|Event|SIMPLE_SEGMENT|8856,8859|false|false|false|||MVP
Finding|Finding|SIMPLE_SEGMENT|8856,8859|false|false|false|C1417509;C1513287|MVP gene;Microvascular Proliferation|MVP
Finding|Gene or Genome|SIMPLE_SEGMENT|8856,8859|false|false|false|C1417509;C1513287|MVP gene;Microvascular Proliferation|MVP
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8856,8859|false|false|false|C0084989;C0280017;C0280018;C0280540;C0280541;C1880093|Cisplatin-Mitomycin-Vinblastine Regimen;cisplatin, etoposide, and methotrexate chemotherapy protocol;cisplatin/mitomycin/vinblastine protocol;cisplatin/mitomycin/vindesine protocol;medroxyprogesterone/mitomycin/vinblastine;procarbazine/semustine/vincristine protocol|MVP
Finding|Finding|SIMPLE_SEGMENT|8862,8870|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Intellectual Product|SIMPLE_SEGMENT|8862,8870|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8876,8896|false|false|false|C0026266|Mitral Valve Insufficiency|mitral regurgitation
Event|Event|SIMPLE_SEGMENT|8883,8896|false|false|false|||regurgitation
Finding|Finding|SIMPLE_SEGMENT|8883,8896|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|SIMPLE_SEGMENT|8883,8896|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|SIMPLE_SEGMENT|8883,8896|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Event|Event|SIMPLE_SEGMENT|8900,8904|false|false|false|||seen
Finding|Functional Concept|SIMPLE_SEGMENT|8907,8910|false|false|false|C0678226;C3146286|Due;Due to|Due
Finding|Idea or Concept|SIMPLE_SEGMENT|8907,8910|false|false|false|C0678226;C3146286|Due;Due to|Due
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|8915,8923|false|false|false|C0001166|Acoustics|acoustic
Finding|Finding|SIMPLE_SEGMENT|8915,8933|false|false|false|C1719833|Acoustic shadowing|acoustic shadowing
Event|Event|SIMPLE_SEGMENT|8924,8933|false|false|false|||shadowing
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8924,8933|false|false|false|C0085195;C0600111|Shadowing (Histology);Shadowing (regime/therapy)|shadowing
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8924,8933|false|false|false|C0085195;C0600111|Shadowing (Histology);Shadowing (regime/therapy)|shadowing
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8951,8971|false|false|false|C0026266|Mitral Valve Insufficiency|mitral regurgitation
Finding|Finding|SIMPLE_SEGMENT|8958,8971|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|SIMPLE_SEGMENT|8958,8971|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|SIMPLE_SEGMENT|8958,8971|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Event|Event|SIMPLE_SEGMENT|8994,9008|false|false|false|||UNDERestimated
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9023,9034|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9023,9034|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Event|Event|SIMPLE_SEGMENT|9036,9044|false|false|false|||effusion
Finding|Body Substance|SIMPLE_SEGMENT|9036,9044|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|SIMPLE_SEGMENT|9036,9044|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|9036,9044|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9055,9061|false|false|false|C1644645||CT Abd
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9058,9061|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|Abd
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|9058,9061|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|Abd
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9062,9068|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|Pelvis
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|9062,9068|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|Pelvis
Disorder|Neoplastic Process|SIMPLE_SEGMENT|9062,9068|false|false|false|C0153663|Malignant neoplasm of pelvis|Pelvis
Finding|Finding|SIMPLE_SEGMENT|9062,9068|false|false|false|C0812455|Pelvis problem|Pelvis
Event|Event|SIMPLE_SEGMENT|9076,9086|false|false|false|||IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|9076,9086|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|9076,9086|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|9089,9097|false|false|false|C1552654|Parameterized Data Type - Interval|Interval
Event|Event|SIMPLE_SEGMENT|9098,9106|false|false|false|||increase
Finding|Functional Concept|SIMPLE_SEGMENT|9098,9106|false|false|false|C0442805|Increase|increase
Anatomy|Tissue|SIMPLE_SEGMENT|9120,9127|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9120,9127|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Pathologic Function|SIMPLE_SEGMENT|9120,9137|false|false|false|C0032227|Pleural effusion (disorder)|pleural effusions
Event|Event|SIMPLE_SEGMENT|9128,9137|false|false|false|||effusions
Finding|Pathologic Function|SIMPLE_SEGMENT|9128,9137|false|false|false|C0013687|effusion|effusions
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9148,9157|false|false|false|C0000726|Abdomen|abdominal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9148,9165|false|false|false|C0003962|Ascites|abdominal ascites
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9158,9165|false|false|false|C0003962|Ascites|ascites
Event|Event|SIMPLE_SEGMENT|9158,9165|false|false|false|||ascites
Finding|Pathologic Function|SIMPLE_SEGMENT|9158,9165|false|false|false|C5441966|Peritoneal Effusion|ascites
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9172,9177|false|false|false|C0009368;C4071907|Abdomen+Pelvis>Colon;Colon structure (body structure)|colon
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9172,9177|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Disorder|Neoplastic Process|SIMPLE_SEGMENT|9172,9177|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Event|Event|SIMPLE_SEGMENT|9172,9177|false|false|false|||colon
Finding|Finding|SIMPLE_SEGMENT|9172,9177|false|false|false|C0750873|COLON PROBLEM|colon
Event|Event|SIMPLE_SEGMENT|9186,9193|false|false|false|||dilated
Finding|Finding|SIMPLE_SEGMENT|9186,9193|false|false|false|C0700124|Dilated|dilated
Event|Event|SIMPLE_SEGMENT|9198,9207|false|false|false|||ahaustral
Event|Event|SIMPLE_SEGMENT|9213,9220|false|false|false|||keeping
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9239,9246|false|false|false|C0009319|Colitis|colitis
Event|Event|SIMPLE_SEGMENT|9239,9246|false|false|false|||colitis
Event|Event|SIMPLE_SEGMENT|9250,9253|false|false|false|||CXR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|9250,9253|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|SIMPLE_SEGMENT|9281,9285|false|false|false|||tube
Finding|Functional Concept|SIMPLE_SEGMENT|9281,9285|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|tube
Finding|Gene or Genome|SIMPLE_SEGMENT|9281,9285|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|tube
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9292,9298|false|false|false|C4522154|Distal Resection Margin|distal
Event|Event|SIMPLE_SEGMENT|9299,9302|false|false|false|||tip
Finding|Gene or Genome|SIMPLE_SEGMENT|9299,9302|false|false|false|C1705504;C1823282;C1825626;C1825978|ITFG1 gene;KAT5 wt Allele;METTL8 gene;TIPRL gene|tip
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9299,9302|false|false|false|C0673828|TIP regimen|tip
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|9313,9317|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9313,9317|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Finding|Intellectual Product|SIMPLE_SEGMENT|9313,9317|false|false|false|C1551342|Document Body|body
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9326,9333|false|false|false|C0038351;C3714551;C4266636|Abdomen>Stomach;Stomach;Stomach structure|stomach
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9326,9333|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Disorder|Neoplastic Process|SIMPLE_SEGMENT|9326,9333|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Event|Event|SIMPLE_SEGMENT|9326,9333|false|false|false|||stomach
Finding|Finding|SIMPLE_SEGMENT|9326,9333|false|false|false|C0577027|Stomach problem|stomach
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9326,9333|false|false|false|C0872393|Procedure on stomach|stomach
Anatomy|Tissue|SIMPLE_SEGMENT|9357,9364|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9357,9364|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Pathologic Function|SIMPLE_SEGMENT|9357,9374|false|false|false|C0032227|Pleural effusion (disorder)|pleural effusions
Event|Event|SIMPLE_SEGMENT|9365,9374|false|false|false|||effusions
Finding|Pathologic Function|SIMPLE_SEGMENT|9365,9374|false|false|false|C0013687|effusion|effusions
Finding|Functional Concept|SIMPLE_SEGMENT|9388,9393|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Tissue|SIMPLE_SEGMENT|9401,9408|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9401,9408|false|false|false|C0032226|Pleural Diseases|pleural
Event|Event|SIMPLE_SEGMENT|9415,9423|false|false|false|||catheter
Finding|Intellectual Product|SIMPLE_SEGMENT|9415,9423|false|false|false|C1546572||catheter
Event|Event|SIMPLE_SEGMENT|9438,9452|false|false|false|||pneumothoraces
Event|Event|SIMPLE_SEGMENT|9456,9461|false|false|false|||signs
Finding|Finding|SIMPLE_SEGMENT|9456,9461|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|SIMPLE_SEGMENT|9456,9461|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9473,9482|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9473,9482|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|9473,9482|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|SIMPLE_SEGMENT|9473,9488|false|false|false|C0034063|Pulmonary Edema|pulmonary edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9483,9488|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|9483,9488|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|9483,9488|false|false|false|C0013604|Edema|edema
Finding|Intellectual Product|SIMPLE_SEGMENT|9491,9498|false|false|false|C0282416|Overall Publication Type|Overall
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9506,9514|false|false|false|C2926606||findings
Event|Event|SIMPLE_SEGMENT|9506,9514|false|false|false|||findings
Finding|Functional Concept|SIMPLE_SEGMENT|9506,9514|false|false|false|C2607943|findings aspects|findings
Event|Event|SIMPLE_SEGMENT|9519,9525|false|false|false|||stable
Finding|Intellectual Product|SIMPLE_SEGMENT|9519,9525|false|false|false|C1547311|Patient Condition Code - Stable|stable
Event|Event|SIMPLE_SEGMENT|9539,9544|false|false|false|||study
Finding|Intellectual Product|SIMPLE_SEGMENT|9539,9544|false|false|false|C1705923|Study Object|study
Procedure|Research Activity|SIMPLE_SEGMENT|9539,9544|false|false|false|C0008972;C0947630;C2603343|Clinical Research;Scientific Study;Study|study
Finding|Intellectual Product|SIMPLE_SEGMENT|9559,9564|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|Brief
Finding|Idea or Concept|SIMPLE_SEGMENT|9565,9573|false|false|false|C1547192|Organization unit type - Hospital|Hospital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9565,9580|false|false|false|C0488549||Hospital Course
Finding|Finding|SIMPLE_SEGMENT|9565,9580|false|false|false|C0489547|Hospital course|Hospital Course
Finding|Idea or Concept|SIMPLE_SEGMENT|9595,9599|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|SIMPLE_SEGMENT|9595,9599|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Event|Event|SIMPLE_SEGMENT|9600,9603|false|false|false|||old
Event|Event|SIMPLE_SEGMENT|9615,9622|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|9615,9622|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|9615,9622|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|9615,9622|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|9615,9625|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9626,9635|false|false|false|C1527336|Sjogren's Syndrome|Sjogren's
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9626,9644|false|false|false|C1527336|Sjogren's Syndrome|Sjogren's syndrome
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9636,9644|false|false|false|C0039082|Syndrome|syndrome
Event|Event|SIMPLE_SEGMENT|9636,9644|false|false|false|||syndrome
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|9650,9653|false|false|false|C0022104;C0432306|Ichthyosis Bullosa of Siemens;Irritable Bowel Syndrome|IBS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9650,9653|false|false|false|C0022104;C0432306|Ichthyosis Bullosa of Siemens;Irritable Bowel Syndrome|IBS
Event|Event|SIMPLE_SEGMENT|9650,9653|false|false|false|||IBS
Event|Event|SIMPLE_SEGMENT|9654,9664|false|false|false|||presenting
Event|Event|SIMPLE_SEGMENT|9670,9676|false|false|false|||fevers
Finding|Sign or Symptom|SIMPLE_SEGMENT|9670,9676|false|false|false|C0015967|Fever|fevers
Event|Event|SIMPLE_SEGMENT|9678,9686|false|false|false|||diarrhea
Finding|Finding|SIMPLE_SEGMENT|9678,9686|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|SIMPLE_SEGMENT|9678,9686|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Event|Event|SIMPLE_SEGMENT|9688,9699|false|false|false|||tachycardia
Finding|Finding|SIMPLE_SEGMENT|9688,9699|false|false|false|C0039231;C3827868|Tachycardia;Tachycardia by ECG Finding|tachycardia
Event|Event|SIMPLE_SEGMENT|9702,9713|false|false|false|||hypotension
Finding|Finding|SIMPLE_SEGMENT|9702,9713|false|false|false|C0020649|Hypotension|hypotension
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9715,9727|false|false|false|C0023518|Leukocytosis|leukocytosis
Event|Event|SIMPLE_SEGMENT|9715,9727|false|false|false|||leukocytosis
Finding|Finding|SIMPLE_SEGMENT|9715,9727|false|false|false|C0750426|Blood leukocyte number above reference range|leukocytosis
Event|Event|SIMPLE_SEGMENT|9729,9736|false|false|false|||hypoxia
Finding|Finding|SIMPLE_SEGMENT|9729,9736|false|false|false|C0242184;C1963140|Hypoxia;Hypoxia, CTCAE|hypoxia
Finding|Pathologic Function|SIMPLE_SEGMENT|9729,9736|false|false|false|C0242184;C1963140|Hypoxia;Hypoxia, CTCAE|hypoxia
Event|Event|SIMPLE_SEGMENT|9738,9743|false|false|false|||found
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9752,9762|false|false|false|C0868908|Pancolitis|pancolitis
Event|Event|SIMPLE_SEGMENT|9752,9762|false|false|false|||pancolitis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9768,9777|false|false|false|C0032285|Pneumonia|pneumonia
Event|Event|SIMPLE_SEGMENT|9768,9777|false|false|false|||pneumonia
Finding|Functional Concept|SIMPLE_SEGMENT|9782,9788|false|false|false|C0333534|septic|Septic
Finding|Pathologic Function|SIMPLE_SEGMENT|9782,9794|false|false|false|C0036983|Septic Shock|Septic Shock
Event|Event|SIMPLE_SEGMENT|9789,9794|false|false|false|||Shock
Finding|Pathologic Function|SIMPLE_SEGMENT|9789,9794|false|false|false|C0036974|Shock|Shock
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9808,9815|false|false|false|C0009319|Colitis|Colitis
Event|Event|SIMPLE_SEGMENT|9808,9815|false|false|false|||Colitis
Event|Event|SIMPLE_SEGMENT|9820,9829|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|9820,9829|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|9830,9834|false|false|false|C1550543|Fulfill|meet
Event|Event|SIMPLE_SEGMENT|9835,9843|false|false|false|||criteria
Finding|Idea or Concept|SIMPLE_SEGMENT|9835,9843|false|false|false|C0243161|criteria|criteria
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9849,9855|false|false|false|C0036690;C0243026|Sepsis;Septicemia|sepsis
Event|Event|SIMPLE_SEGMENT|9862,9867|false|false|false|||fever
Finding|Finding|SIMPLE_SEGMENT|9862,9867|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|9862,9867|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Event|Event|SIMPLE_SEGMENT|9869,9880|false|false|false|||tachycardia
Finding|Finding|SIMPLE_SEGMENT|9869,9880|false|false|false|C0039231;C3827868|Tachycardia;Tachycardia by ECG Finding|tachycardia
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9882,9894|false|false|false|C0023518|Leukocytosis|leukocytosis
Event|Event|SIMPLE_SEGMENT|9882,9894|false|false|false|||leukocytosis
Finding|Finding|SIMPLE_SEGMENT|9882,9894|false|false|false|C0750426|Blood leukocyte number above reference range|leukocytosis
Finding|Finding|SIMPLE_SEGMENT|9899,9905|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|9899,9905|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|SIMPLE_SEGMENT|9907,9913|false|false|false|||source
Finding|Finding|SIMPLE_SEGMENT|9907,9913|false|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Finding|Functional Concept|SIMPLE_SEGMENT|9907,9913|false|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Finding|Intellectual Product|SIMPLE_SEGMENT|9907,9913|false|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9920,9927|false|false|false|C0009319|Colitis|colitis
Event|Event|SIMPLE_SEGMENT|9920,9927|false|false|false|||colitis
Event|Event|SIMPLE_SEGMENT|9929,9931|false|false|false|||BP
Event|Event|SIMPLE_SEGMENT|9932,9940|false|false|false|||remained
Event|Event|SIMPLE_SEGMENT|9941,9944|false|false|false|||low
Finding|Finding|SIMPLE_SEGMENT|9941,9944|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|SIMPLE_SEGMENT|9941,9944|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Body Substance|SIMPLE_SEGMENT|9949,9956|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|9949,9956|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|9949,9956|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|9957,9965|false|false|false|||remained
Event|Event|SIMPLE_SEGMENT|9974,9985|false|false|false|||tachycardic
Finding|Idea or Concept|SIMPLE_SEGMENT|9990,9994|false|false|false|C1552851|next - HtmlLinkType|next
Event|Event|SIMPLE_SEGMENT|9999,10008|false|false|false|||requiring
Finding|Individual Behavior|SIMPLE_SEGMENT|10009,10019|false|false|false|C0001807;C1547300;C1548760|Aggressive behavior;Precaution Code - Aggressive;Risk Codes - Aggressive|aggressive
Finding|Intellectual Product|SIMPLE_SEGMENT|10009,10019|false|false|false|C0001807;C1547300;C1548760|Aggressive behavior;Precaution Code - Aggressive;Risk Codes - Aggressive|aggressive
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|10020,10023|false|false|false|C0016520|Structure of interventricular foramen|IVF
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10020,10023|false|false|false|C2751898|Ventricular Fibrillation, Paroxysmal Familial, 1|IVF
Event|Event|SIMPLE_SEGMENT|10020,10023|false|false|false|||IVF
Finding|Gene or Genome|SIMPLE_SEGMENT|10020,10023|false|false|false|C1419864;C4321334|SCN5A gene;SCN5A wt Allele|IVF
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10020,10023|false|false|false|C0015915;C0872104|Assisted Reproductive Technologies;Fertilization in Vitro|IVF
Event|Event|SIMPLE_SEGMENT|10065,10072|false|false|false|||started
Finding|Finding|SIMPLE_SEGMENT|10073,10078|false|false|false|C3714655|On IV|on IV
Drug|Organic Chemical|SIMPLE_SEGMENT|10079,10085|false|false|false|C0699678|Flagyl|flagyl
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10079,10085|false|false|false|C0699678|Flagyl|flagyl
Event|Event|SIMPLE_SEGMENT|10079,10085|false|false|false|||flagyl
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10090,10095|false|false|false|C0042313|vancomycin|vanco
Drug|Antibiotic|SIMPLE_SEGMENT|10090,10095|false|false|false|C0042313|vancomycin|vanco
Finding|Finding|SIMPLE_SEGMENT|10112,10120|false|false|false|C0332149|Possible|possible
Event|Event|SIMPLE_SEGMENT|10121,10126|false|false|false|||Cdiff
Finding|Finding|SIMPLE_SEGMENT|10130,10134|false|false|false|C5575035|Well (answer to question)|well
Drug|Antibiotic|SIMPLE_SEGMENT|10138,10150|false|false|false|C0282386|levofloxacin|levofloxacin
Drug|Organic Chemical|SIMPLE_SEGMENT|10138,10150|false|false|false|C0282386|levofloxacin|levofloxacin
Event|Event|SIMPLE_SEGMENT|10138,10150|false|false|false|||levofloxacin
Event|Event|SIMPLE_SEGMENT|10157,10164|false|false|false|||concern
Finding|Idea or Concept|SIMPLE_SEGMENT|10157,10164|false|false|false|C2699424|Concern|concern
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|10169,10172|false|false|false|C0600500|Peptide Nucleic Acids|PNA
Event|Event|SIMPLE_SEGMENT|10169,10172|false|false|false|||PNA
Event|Event|SIMPLE_SEGMENT|10196,10201|false|false|false|||Stool
Finding|Body Substance|SIMPLE_SEGMENT|10196,10201|false|false|false|C0015733|Feces|Stool
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|10224,10232|false|false|false|C4727483|BRAF Gene Rearrangement|positive
Event|Event|SIMPLE_SEGMENT|10224,10232|false|false|false|||positive
Finding|Classification|SIMPLE_SEGMENT|10224,10232|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|SIMPLE_SEGMENT|10224,10232|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Drug|Antibiotic|SIMPLE_SEGMENT|10237,10249|false|false|false|C0282386|levofloxacin|levofloxacin
Drug|Organic Chemical|SIMPLE_SEGMENT|10237,10249|false|false|false|C0282386|levofloxacin|levofloxacin
Event|Event|SIMPLE_SEGMENT|10237,10249|false|false|false|||levofloxacin
Event|Event|SIMPLE_SEGMENT|10250,10257|false|false|false|||changed
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10261,10264|false|false|false|C0238052|Xanthomatosis, Cerebrotendinous|CTX
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10261,10264|false|false|false|C0010377;C0010583;C5574748|C-Terminal Telopeptide Type 1 Collagen, human;Crotoxin;cyclophosphamide|CTX
Drug|Biologically Active Substance|SIMPLE_SEGMENT|10261,10264|false|false|false|C0010377;C0010583;C5574748|C-Terminal Telopeptide Type 1 Collagen, human;Crotoxin;cyclophosphamide|CTX
Drug|Enzyme|SIMPLE_SEGMENT|10261,10264|false|false|false|C0010377;C0010583;C5574748|C-Terminal Telopeptide Type 1 Collagen, human;Crotoxin;cyclophosphamide|CTX
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|10261,10264|false|false|false|C0010377;C0010583;C5574748|C-Terminal Telopeptide Type 1 Collagen, human;Crotoxin;cyclophosphamide|CTX
Drug|Organic Chemical|SIMPLE_SEGMENT|10261,10264|false|false|false|C0010377;C0010583;C5574748|C-Terminal Telopeptide Type 1 Collagen, human;Crotoxin;cyclophosphamide|CTX
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10261,10264|false|false|false|C0010377;C0010583;C5574748|C-Terminal Telopeptide Type 1 Collagen, human;Crotoxin;cyclophosphamide|CTX
Event|Event|SIMPLE_SEGMENT|10261,10264|false|false|false|||CTX
Finding|Gene or Genome|SIMPLE_SEGMENT|10261,10264|false|false|false|C1413864;C3539598|CYP27A1 gene;CYP27A1 wt Allele|CTX
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10274,10277|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|10274,10277|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|10274,10277|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10274,10277|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|SIMPLE_SEGMENT|10274,10277|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|10274,10277|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|SIMPLE_SEGMENT|10274,10277|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10274,10277|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|SIMPLE_SEGMENT|10274,10277|false|false|false|||PCP
Finding|Gene or Genome|SIMPLE_SEGMENT|10274,10277|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|SIMPLE_SEGMENT|10274,10277|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Event|SIMPLE_SEGMENT|10288,10295|false|false|false|||visited
Event|Event|SIMPLE_SEGMENT|10300,10304|false|false|false|||said
Finding|Finding|SIMPLE_SEGMENT|10313,10319|false|false|false|C1549493;C3812891|All of the Time;Always - AcknowledgementCondition|always
Finding|Idea or Concept|SIMPLE_SEGMENT|10313,10319|false|false|false|C1549493;C3812891|All of the Time;Always - AcknowledgementCondition|always
Event|Event|SIMPLE_SEGMENT|10324,10327|false|false|false|||CXR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10324,10327|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|SIMPLE_SEGMENT|10328,10338|false|false|false|||infiltrate
Finding|Functional Concept|SIMPLE_SEGMENT|10328,10338|false|false|false|C0332448;C1546677;C1549537|Administration Method - Infiltrate;Infiltration|infiltrate
Finding|Intellectual Product|SIMPLE_SEGMENT|10328,10338|false|false|false|C0332448;C1546677;C1549537|Administration Method - Infiltrate;Infiltration|infiltrate
Finding|Pathologic Function|SIMPLE_SEGMENT|10328,10338|false|false|false|C0332448;C1546677;C1549537|Administration Method - Infiltrate;Infiltration|infiltrate
Event|Event|SIMPLE_SEGMENT|10343,10346|false|false|false|||abx
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10351,10354|false|false|false|C0238052|Xanthomatosis, Cerebrotendinous|CTX
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10351,10354|false|false|false|C0010377;C0010583;C5574748|C-Terminal Telopeptide Type 1 Collagen, human;Crotoxin;cyclophosphamide|CTX
Drug|Biologically Active Substance|SIMPLE_SEGMENT|10351,10354|false|false|false|C0010377;C0010583;C5574748|C-Terminal Telopeptide Type 1 Collagen, human;Crotoxin;cyclophosphamide|CTX
Drug|Enzyme|SIMPLE_SEGMENT|10351,10354|false|false|false|C0010377;C0010583;C5574748|C-Terminal Telopeptide Type 1 Collagen, human;Crotoxin;cyclophosphamide|CTX
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|10351,10354|false|false|false|C0010377;C0010583;C5574748|C-Terminal Telopeptide Type 1 Collagen, human;Crotoxin;cyclophosphamide|CTX
Drug|Organic Chemical|SIMPLE_SEGMENT|10351,10354|false|false|false|C0010377;C0010583;C5574748|C-Terminal Telopeptide Type 1 Collagen, human;Crotoxin;cyclophosphamide|CTX
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10351,10354|false|false|false|C0010377;C0010583;C5574748|C-Terminal Telopeptide Type 1 Collagen, human;Crotoxin;cyclophosphamide|CTX
Event|Event|SIMPLE_SEGMENT|10351,10354|false|false|false|||CTX
Finding|Gene or Genome|SIMPLE_SEGMENT|10351,10354|false|false|false|C1413864;C3539598|CYP27A1 gene;CYP27A1 wt Allele|CTX
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10367,10376|false|false|false|C0032285|Pneumonia|pneumonia
Event|Event|SIMPLE_SEGMENT|10367,10376|false|false|false|||pneumonia
Event|Event|SIMPLE_SEGMENT|10377,10384|false|false|false|||stopped
Event|Event|SIMPLE_SEGMENT|10428,10437|false|false|false|||treatment
Finding|Conceptual Entity|SIMPLE_SEGMENT|10428,10437|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|SIMPLE_SEGMENT|10428,10437|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|SIMPLE_SEGMENT|10428,10437|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10428,10437|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Drug|Organic Chemical|SIMPLE_SEGMENT|10439,10446|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10439,10446|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Event|Event|SIMPLE_SEGMENT|10439,10446|false|false|false|||Lactate
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10439,10446|false|false|false|C0202115|Lactic acid measurement|Lactate
Anatomy|Cell|SIMPLE_SEGMENT|10451,10454|false|false|false|C0023516|Leukocytes|WBC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10451,10460|false|false|false|C0023508|White Blood Cell Count procedure|WBC count
Event|Event|SIMPLE_SEGMENT|10455,10460|false|false|false|||count
Event|Event|SIMPLE_SEGMENT|10462,10469|false|false|false|||trended
Finding|Body Substance|SIMPLE_SEGMENT|10492,10499|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|10492,10499|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|10492,10499|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|10500,10509|false|false|false|||developed
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10510,10515|false|false|false|C1258215;C4019039|Ileus;Intestinal obstruction co-occurrent and due to decreased peristalsis|ileus
Event|Event|SIMPLE_SEGMENT|10510,10515|false|false|false|||ileus
Anatomy|Body Location or Region|SIMPLE_SEGMENT|10520,10529|false|false|false|C0000726|Abdomen|abdominal
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10520,10537|false|false|false|C4481095|abdominal imaging|abdominal imaging
Event|Event|SIMPLE_SEGMENT|10530,10537|false|false|false|||imaging
Finding|Finding|SIMPLE_SEGMENT|10530,10537|false|false|false|C0740845|Imaging problem|imaging
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10530,10537|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|imaging
Event|Event|SIMPLE_SEGMENT|10543,10552|false|false|false|||worsening
Finding|Idea or Concept|SIMPLE_SEGMENT|10543,10552|false|false|false|C1546960|Patient Outcome - Worsening|worsening
Event|Event|SIMPLE_SEGMENT|10553,10563|false|false|false|||distension
Finding|Finding|SIMPLE_SEGMENT|10553,10563|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distension
Finding|Pathologic Function|SIMPLE_SEGMENT|10553,10563|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distension
Finding|Classification|SIMPLE_SEGMENT|10572,10575|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Finding|Gene or Genome|SIMPLE_SEGMENT|10572,10575|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Event|Event|SIMPLE_SEGMENT|10576,10580|false|false|false|||Surg
Finding|Functional Concept|SIMPLE_SEGMENT|10576,10580|false|false|false|C0038895|Surgical aspects|Surg
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10576,10580|false|false|false|C0543467;C1948041|Operative Surgical Procedures;Surgical and medical procedures|Surg
Event|Event|SIMPLE_SEGMENT|10603,10606|false|false|false|||NPO
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10603,10606|false|false|false|C0419179|NPO - Nothing by mouth|NPO
Event|Event|SIMPLE_SEGMENT|10633,10640|false|false|false|||illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|10633,10640|false|false|false|C0221423|Illness (finding)|illness
Event|Event|SIMPLE_SEGMENT|10642,10648|false|false|false|||turned
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|10674,10677|false|false|false|C0016520|Structure of interventricular foramen|IVF
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10674,10677|false|false|false|C2751898|Ventricular Fibrillation, Paroxysmal Familial, 1|IVF
Event|Event|SIMPLE_SEGMENT|10674,10677|false|false|false|||IVF
Finding|Gene or Genome|SIMPLE_SEGMENT|10674,10677|false|false|false|C1419864;C4321334|SCN5A gene;SCN5A wt Allele|IVF
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10674,10677|false|false|false|C0015915;C0872104|Assisted Reproductive Technologies;Fertilization in Vitro|IVF
Finding|Finding|SIMPLE_SEGMENT|10682,10686|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|10682,10686|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|10682,10686|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|10690,10693|false|false|false|C0228479|Structure of intraculminate fissure|ICU
Finding|Intellectual Product|SIMPLE_SEGMENT|10690,10693|false|false|false|C4554035|Inventory of Callous-Unemotional Traits|ICU
Event|Event|SIMPLE_SEGMENT|10694,10698|false|false|false|||call
Finding|Functional Concept|SIMPLE_SEGMENT|10694,10698|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|call
Finding|Gene or Genome|SIMPLE_SEGMENT|10694,10698|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|call
Finding|Intellectual Product|SIMPLE_SEGMENT|10694,10698|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|call
Finding|Mental Process|SIMPLE_SEGMENT|10694,10698|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|call
Event|Event|SIMPLE_SEGMENT|10712,10722|false|false|false|||stabilized
Finding|Finding|SIMPLE_SEGMENT|10712,10722|false|false|false|C0184512|Stabilized (qualifier value)|stabilized
Drug|Substance|SIMPLE_SEGMENT|10741,10747|false|false|false|C0302908|Liquid substance|fluids
Event|Event|SIMPLE_SEGMENT|10741,10747|false|false|false|||fluids
Finding|Body Substance|SIMPLE_SEGMENT|10741,10747|false|false|false|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10741,10747|false|false|false|C0016286|Fluid Therapy|fluids
Anatomy|Body Location or Region|SIMPLE_SEGMENT|10752,10761|false|false|false|C0000726|Abdomen|abdominal
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10752,10766|false|false|false|C0562238|Examination of abdomen|abdominal exam
Event|Event|SIMPLE_SEGMENT|10762,10766|false|false|false|||exam
Finding|Functional Concept|SIMPLE_SEGMENT|10762,10766|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|10762,10766|false|false|false|C0582103|Medical Examination|exam
Event|Event|SIMPLE_SEGMENT|10772,10781|false|false|false|||improving
Event|Event|SIMPLE_SEGMENT|10787,10799|false|false|false|||downtrending
Anatomy|Cell|SIMPLE_SEGMENT|10800,10803|false|false|false|C0023516|Leukocytes|WBC
Event|Event|SIMPLE_SEGMENT|10805,10809|false|false|false|||Came
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|10818,10821|false|false|false|C0228479|Structure of intraculminate fissure|ICU
Finding|Intellectual Product|SIMPLE_SEGMENT|10818,10821|false|false|false|C4554035|Inventory of Callous-Unemotional Traits|ICU
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10837,10848|false|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|SIMPLE_SEGMENT|10837,10848|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|SIMPLE_SEGMENT|10837,10848|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|SIMPLE_SEGMENT|10837,10848|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Sign or Symptom|SIMPLE_SEGMENT|10837,10857|false|false|false|C0476273|Respiratory distress|respiratory distress
Event|Event|SIMPLE_SEGMENT|10849,10857|false|false|false|||distress
Finding|Finding|SIMPLE_SEGMENT|10849,10857|false|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|SIMPLE_SEGMENT|10849,10857|false|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Event|Event|SIMPLE_SEGMENT|10862,10869|false|false|false|||hypoxia
Finding|Finding|SIMPLE_SEGMENT|10862,10869|false|false|false|C0242184;C1963140|Hypoxia;Hypoxia, CTCAE|hypoxia
Finding|Pathologic Function|SIMPLE_SEGMENT|10862,10869|false|false|false|C0242184;C1963140|Hypoxia;Hypoxia, CTCAE|hypoxia
Event|Event|SIMPLE_SEGMENT|10886,10893|false|false|false|||started
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10903,10911|false|false|false|C0237795|Pressors|pressors
Event|Event|SIMPLE_SEGMENT|10903,10911|false|false|false|||pressors
Drug|Organic Chemical|SIMPLE_SEGMENT|10923,10936|false|false|false|C0031469|phenylephrine|phenylephrine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10923,10936|false|false|false|C0031469|phenylephrine|phenylephrine
Event|Event|SIMPLE_SEGMENT|10923,10936|false|false|false|||phenylephrine
Finding|Intellectual Product|SIMPLE_SEGMENT|10941,10945|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|SIMPLE_SEGMENT|10955,10962|false|false|false|||stopped
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10967,10978|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10984,10988|false|false|false|C0009443;C0024117|Chronic Obstructive Airway Disease;Common Cold|cold
Drug|Organic Chemical|SIMPLE_SEGMENT|10984,10988|false|false|false|C0719425|Cold brand of chlorpheniramine-phenylpropanolamine|cold
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10984,10988|false|false|false|C0719425|Cold brand of chlorpheniramine-phenylpropanolamine|cold
Event|Event|SIMPLE_SEGMENT|10984,10988|false|false|false|||cold
Finding|Organism Function|SIMPLE_SEGMENT|10984,10988|false|false|false|C0234192|Cold Sensation|cold
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|10984,10988|false|false|false|C0009264|Cold Temperature|cold
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10984,10988|false|false|false|C0010412|Cold Therapy|cold
Event|Event|SIMPLE_SEGMENT|10993,11000|false|false|false|||mottled
Finding|Finding|SIMPLE_SEGMENT|10993,11000|false|false|false|C0302133|Mottling|mottled
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11002,11010|false|false|false|C0237795|Pressors|Pressors
Event|Event|SIMPLE_SEGMENT|11002,11010|false|false|false|||Pressors
Event|Event|SIMPLE_SEGMENT|11011,11018|false|false|false|||changed
Event|Event|SIMPLE_SEGMENT|11023,11037|false|false|false|||Norepinephrine
Event|Event|SIMPLE_SEGMENT|11042,11050|false|false|false|||mottling
Finding|Finding|SIMPLE_SEGMENT|11042,11050|false|false|false|C0302133|Mottling|mottling
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|11054,11057|false|false|false|C0015306|Hereditary Multiple Exostoses|ext
Event|Event|SIMPLE_SEGMENT|11054,11057|false|false|false|||ext
Finding|Gene or Genome|SIMPLE_SEGMENT|11054,11057|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|ext
Event|Event|SIMPLE_SEGMENT|11066,11074|false|false|false|||resolved
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|11076,11080|false|false|false|C0428176|Venous oxygen saturation measurement|SVO2
Event|Event|SIMPLE_SEGMENT|11086,11090|false|false|false|||ECHO
Procedure|Health Care Activity|SIMPLE_SEGMENT|11086,11090|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11086,11090|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Event|Event|SIMPLE_SEGMENT|11095,11105|false|false|false|||consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|11095,11105|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|11095,11110|false|false|false|C0332290|Consistent with|consistent with
Finding|Pathologic Function|SIMPLE_SEGMENT|11111,11128|false|true|false|C0036980|Shock, Cardiogenic|cardiogenic shock
Event|Event|SIMPLE_SEGMENT|11123,11128|false|false|false|||shock
Finding|Pathologic Function|SIMPLE_SEGMENT|11123,11128|false|true|false|C0036974|Shock|shock
Event|Event|SIMPLE_SEGMENT|11133,11136|false|false|false|||EKG
Finding|Intellectual Product|SIMPLE_SEGMENT|11133,11136|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|11133,11136|false|false|false|C1623258|Electrocardiography|EKG
Event|Event|SIMPLE_SEGMENT|11149,11157|false|false|false|||negative
Finding|Classification|SIMPLE_SEGMENT|11149,11157|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|11149,11157|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|11149,11157|false|false|false|C5237010|Expression Negative|negative
Event|Event|SIMPLE_SEGMENT|11162,11165|false|false|false|||saw
Event|Event|SIMPLE_SEGMENT|11169,11176|false|false|false|||consult
Procedure|Health Care Activity|SIMPLE_SEGMENT|11169,11176|false|false|false|C0009818|Consultation|consult
Event|Event|SIMPLE_SEGMENT|11181,11192|false|false|false|||recommended
Finding|Idea or Concept|SIMPLE_SEGMENT|11181,11192|false|false|false|C0034866|Recommendation|recommended
Drug|Antibiotic|SIMPLE_SEGMENT|11202,11213|false|false|false|C1260298|tigecycline|Tigecycline
Drug|Organic Chemical|SIMPLE_SEGMENT|11202,11213|false|false|false|C1260298|tigecycline|Tigecycline
Event|Event|SIMPLE_SEGMENT|11202,11213|false|false|false|||Tigecycline
Event|Event|SIMPLE_SEGMENT|11218,11222|false|false|false|||help
Event|Event|SIMPLE_SEGMENT|11223,11228|false|false|false|||cover
Event|Event|SIMPLE_SEGMENT|11245,11254|false|false|false|||completed
Finding|Idea or Concept|SIMPLE_SEGMENT|11260,11263|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|11260,11263|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|11264,11270|false|false|false|||course
Anatomy|Body Location or Region|SIMPLE_SEGMENT|11276,11285|false|false|false|C0000726|Abdomen|Abdominal
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|11276,11290|false|false|false|C0562238|Examination of abdomen|Abdominal exam
Event|Event|SIMPLE_SEGMENT|11286,11290|false|false|false|||exam
Finding|Functional Concept|SIMPLE_SEGMENT|11286,11290|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|11286,11290|false|false|false|C0582103|Medical Examination|exam
Event|Event|SIMPLE_SEGMENT|11291,11299|false|false|false|||improved
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11304,11309|false|false|false|C1258215;C4019039|Ileus;Intestinal obstruction co-occurrent and due to decreased peristalsis|ileus
Event|Event|SIMPLE_SEGMENT|11304,11309|false|false|false|||ileus
Event|Event|SIMPLE_SEGMENT|11310,11318|false|false|false|||resolved
Event|Event|SIMPLE_SEGMENT|11320,11326|false|false|false|||Doboff
Event|Event|SIMPLE_SEGMENT|11331,11337|false|false|false|||placed
Finding|Functional Concept|SIMPLE_SEGMENT|11350,11354|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|tube
Finding|Gene or Genome|SIMPLE_SEGMENT|11350,11354|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|tube
Event|Event|SIMPLE_SEGMENT|11355,11360|false|false|false|||feeds
Finding|Functional Concept|SIMPLE_SEGMENT|11355,11360|false|false|false|C1510670|Feeds|feeds
Event|Event|SIMPLE_SEGMENT|11366,11373|false|false|false|||started
Finding|Intellectual Product|SIMPLE_SEGMENT|11378,11382|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|poor
Event|Event|SIMPLE_SEGMENT|11383,11390|false|false|false|||ability
Finding|Functional Concept|SIMPLE_SEGMENT|11383,11390|false|false|false|C5891046|Oral Intake Ability|ability
Finding|Intellectual Product|SIMPLE_SEGMENT|11383,11393|false|false|false|C5420000|Ability Question|ability to
Event|Event|SIMPLE_SEGMENT|11394,11398|false|false|false|||keep
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11410,11421|false|false|false|C2707262||nutritional
Event|Event|SIMPLE_SEGMENT|11422,11434|false|false|false|||requirements
Drug|Organic Chemical|SIMPLE_SEGMENT|11436,11449|false|false|false|C0025872|metronidazole|Metronidazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11436,11449|false|false|false|C0025872|metronidazole|Metronidazole
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11464,11468|false|false|false|C0270724|Infantile Neuroaxonal Dystrophy|Plan
Event|Event|SIMPLE_SEGMENT|11464,11468|false|false|false|||Plan
Finding|Functional Concept|SIMPLE_SEGMENT|11464,11468|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|Plan
Finding|Intellectual Product|SIMPLE_SEGMENT|11464,11468|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|Plan
Finding|Mental Process|SIMPLE_SEGMENT|11464,11468|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|Plan
Event|Event|SIMPLE_SEGMENT|11473,11481|false|false|false|||continue
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|11482,11492|false|false|false|C0042313|vancomycin|Vancomycin
Drug|Antibiotic|SIMPLE_SEGMENT|11482,11492|false|false|false|C0042313|vancomycin|Vancomycin
Event|Event|SIMPLE_SEGMENT|11482,11492|false|false|false|||Vancomycin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|11482,11492|false|false|false|C0489941|Vancomycin measurement|Vancomycin
Event|Event|SIMPLE_SEGMENT|11493,11498|false|false|false|||500mg
Event|Event|SIMPLE_SEGMENT|11502,11504|false|false|false|||Q6
Finding|Finding|SIMPLE_SEGMENT|11535,11544|false|false|false|C5425799|All other|all other
Drug|Antibiotic|SIMPLE_SEGMENT|11545,11556|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|SIMPLE_SEGMENT|11545,11556|false|false|false|||antibiotics
Event|Event|SIMPLE_SEGMENT|11562,11569|false|false|false|||stopped
Finding|Idea or Concept|SIMPLE_SEGMENT|11576,11579|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|11576,11579|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Finding|SIMPLE_SEGMENT|11588,11595|false|false|false|C0242184;C1963140|Hypoxia;Hypoxia, CTCAE|Hypoxia
Finding|Pathologic Function|SIMPLE_SEGMENT|11588,11595|false|false|false|C0242184;C1963140|Hypoxia;Hypoxia, CTCAE|Hypoxia
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11600,11609|true|false|false|C5885990||breathing
Finding|Finding|SIMPLE_SEGMENT|11600,11609|true|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|SIMPLE_SEGMENT|11600,11609|true|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|SIMPLE_SEGMENT|11600,11609|true|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|SIMPLE_SEGMENT|11600,11609|true|false|false|C1160636|respiratory system process|breathing
Event|Event|SIMPLE_SEGMENT|11610,11616|false|false|false|||issues
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|11620,11628|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|SIMPLE_SEGMENT|11620,11628|false|false|false|||baseline
Finding|Idea or Concept|SIMPLE_SEGMENT|11620,11628|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Event|Event|SIMPLE_SEGMENT|11633,11642|false|false|false|||developed
Event|Event|SIMPLE_SEGMENT|11643,11650|false|false|false|||hypoxia
Finding|Finding|SIMPLE_SEGMENT|11643,11650|false|false|false|C0242184;C1963140|Hypoxia;Hypoxia, CTCAE|hypoxia
Finding|Pathologic Function|SIMPLE_SEGMENT|11643,11650|false|false|false|C0242184;C1963140|Hypoxia;Hypoxia, CTCAE|hypoxia
Event|Event|SIMPLE_SEGMENT|11652,11661|false|false|false|||requiring
Event|Event|SIMPLE_SEGMENT|11665,11667|false|false|false|||NC
Event|Event|SIMPLE_SEGMENT|11687,11695|false|false|false|||admitted
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|11703,11706|false|false|false|C0228479|Structure of intraculminate fissure|ICU
Finding|Intellectual Product|SIMPLE_SEGMENT|11703,11706|false|false|false|C4554035|Inventory of Callous-Unemotional Traits|ICU
Finding|Idea or Concept|SIMPLE_SEGMENT|11708,11715|false|false|false|C1555582|Initial (abbreviation)|Initial
Event|Event|SIMPLE_SEGMENT|11717,11724|false|false|false|||concern
Finding|Idea or Concept|SIMPLE_SEGMENT|11717,11724|false|false|false|C2699424|Concern|concern
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11729,11732|false|false|false|C1261075|Structure of right lower lobe of lung|RLL
Finding|Finding|SIMPLE_SEGMENT|11729,11732|false|false|false|C5703311|Radiolucent Lines|RLL
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|11733,11736|false|false|false|C0600500|Peptide Nucleic Acids|PNA
Event|Event|SIMPLE_SEGMENT|11733,11736|false|false|false|||PNA
Event|Event|SIMPLE_SEGMENT|11740,11743|false|false|false|||CXR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|11740,11743|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|SIMPLE_SEGMENT|11774,11779|false|false|false|||noted
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11793,11796|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|11793,11796|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|11793,11796|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|11793,11796|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|SIMPLE_SEGMENT|11793,11796|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|11793,11796|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|SIMPLE_SEGMENT|11793,11796|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11793,11796|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|SIMPLE_SEGMENT|11793,11796|false|false|false|||PCP
Finding|Gene or Genome|SIMPLE_SEGMENT|11793,11796|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|SIMPLE_SEGMENT|11793,11796|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Event|SIMPLE_SEGMENT|11797,11805|false|false|false|||informed
Event|Event|SIMPLE_SEGMENT|11811,11815|false|false|false|||team
Event|Event|SIMPLE_SEGMENT|11821,11831|false|false|false|||infiltrate
Finding|Functional Concept|SIMPLE_SEGMENT|11821,11831|false|false|false|C0332448;C1546677;C1549537|Administration Method - Infiltrate;Infiltration|infiltrate
Finding|Intellectual Product|SIMPLE_SEGMENT|11821,11831|false|false|false|C0332448;C1546677;C1549537|Administration Method - Infiltrate;Infiltration|infiltrate
Finding|Pathologic Function|SIMPLE_SEGMENT|11821,11831|false|false|false|C0332448;C1546677;C1549537|Administration Method - Infiltrate;Infiltration|infiltrate
Event|Event|SIMPLE_SEGMENT|11842,11849|false|false|false|||present
Finding|Finding|SIMPLE_SEGMENT|11842,11849|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|SIMPLE_SEGMENT|11842,11849|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Finding|SIMPLE_SEGMENT|11859,11863|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|11859,11863|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|11859,11863|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|SIMPLE_SEGMENT|11865,11872|false|false|false|||Thought
Event|Event|SIMPLE_SEGMENT|11878,11885|false|false|false|||hypoxia
Finding|Finding|SIMPLE_SEGMENT|11878,11885|false|false|false|C0242184;C1963140|Hypoxia;Hypoxia, CTCAE|hypoxia
Finding|Pathologic Function|SIMPLE_SEGMENT|11878,11885|false|false|false|C0242184;C1963140|Hypoxia;Hypoxia, CTCAE|hypoxia
Event|Event|SIMPLE_SEGMENT|11886,11895|false|false|false|||developed
Finding|Mental Process|SIMPLE_SEGMENT|11899,11906|false|false|false|C0542559|contextual factors|setting
Finding|Individual Behavior|SIMPLE_SEGMENT|11911,11921|false|false|false|C0001807;C1547300;C1548760|Aggressive behavior;Precaution Code - Aggressive;Risk Codes - Aggressive|aggressive
Finding|Intellectual Product|SIMPLE_SEGMENT|11911,11921|false|false|false|C0001807;C1547300;C1548760|Aggressive behavior;Precaution Code - Aggressive;Risk Codes - Aggressive|aggressive
Drug|Substance|SIMPLE_SEGMENT|11922,11928|false|false|false|C0302908|Liquid substance|fluids
Event|Event|SIMPLE_SEGMENT|11922,11928|false|false|false|||fluids
Finding|Body Substance|SIMPLE_SEGMENT|11922,11928|false|false|false|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11922,11928|false|false|false|C0016286|Fluid Therapy|fluids
Finding|Body Substance|SIMPLE_SEGMENT|11932,11939|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|11932,11939|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|11932,11939|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|11945,11956|false|false|false|C0750502|Significant|significant
Event|Event|SIMPLE_SEGMENT|11964,11970|false|false|false|||regurg
Finding|Intellectual Product|SIMPLE_SEGMENT|11990,11994|false|false|false|C1720594|Then - dosing instruction fragment|then
Finding|Individual Behavior|SIMPLE_SEGMENT|11995,12005|false|false|false|C0001807;C1547300;C1548760|Aggressive behavior;Precaution Code - Aggressive;Risk Codes - Aggressive|aggressive
Finding|Intellectual Product|SIMPLE_SEGMENT|11995,12005|false|false|false|C0001807;C1547300;C1548760|Aggressive behavior;Precaution Code - Aggressive;Risk Codes - Aggressive|aggressive
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|12006,12009|false|false|false|C0016520|Structure of interventricular foramen|IVF
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12006,12009|false|false|false|C2751898|Ventricular Fibrillation, Paroxysmal Familial, 1|IVF
Event|Event|SIMPLE_SEGMENT|12006,12009|false|false|false|||IVF
Finding|Gene or Genome|SIMPLE_SEGMENT|12006,12009|false|false|false|C1419864;C4321334|SCN5A gene;SCN5A wt Allele|IVF
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|12006,12009|false|false|false|C0015915;C0872104|Assisted Reproductive Technologies;Fertilization in Vitro|IVF
Event|Event|SIMPLE_SEGMENT|12035,12046|false|false|false|||development
Finding|Functional Concept|SIMPLE_SEGMENT|12035,12046|false|false|false|C0018271;C0243107;C0678723;C1527148|Development;Growth and Development function;biological development;development aspects|development
Finding|Organism Function|SIMPLE_SEGMENT|12035,12046|false|false|false|C0018271;C0243107;C0678723;C1527148|Development;Growth and Development function;biological development;development aspects|development
Anatomy|Tissue|SIMPLE_SEGMENT|12050,12057|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12050,12057|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Pathologic Function|SIMPLE_SEGMENT|12050,12067|false|false|false|C0032227|Pleural effusion (disorder)|pleural effusions
Event|Event|SIMPLE_SEGMENT|12058,12067|false|false|false|||effusions
Finding|Pathologic Function|SIMPLE_SEGMENT|12058,12067|false|false|false|C0013687|effusion|effusions
Event|Event|SIMPLE_SEGMENT|12073,12080|false|false|false|||started
Event|Event|SIMPLE_SEGMENT|12081,12089|false|false|false|||diuresis
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|12081,12089|false|false|false|C0012797|Diuresis|diuresis
Event|Event|SIMPLE_SEGMENT|12093,12097|false|false|false|||MICU
Event|Event|SIMPLE_SEGMENT|12099,12106|false|false|false|||callout
Finding|Intellectual Product|SIMPLE_SEGMENT|12118,12122|false|false|false|C1720594|Then - dosing instruction fragment|then
Finding|Functional Concept|SIMPLE_SEGMENT|12129,12135|false|false|false|C1948027|Couple (action)|couple
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|12144,12149|false|false|false|C3714591|Floor (anatomic)|floor
Event|Event|SIMPLE_SEGMENT|12151,12160|false|false|false|||triggered
Event|Event|SIMPLE_SEGMENT|12166,12173|false|false|false|||hypoxia
Finding|Finding|SIMPLE_SEGMENT|12166,12173|false|false|false|C0242184;C1963140|Hypoxia;Hypoxia, CTCAE|hypoxia
Finding|Pathologic Function|SIMPLE_SEGMENT|12166,12173|false|false|false|C0242184;C1963140|Hypoxia;Hypoxia, CTCAE|hypoxia
Finding|Finding|SIMPLE_SEGMENT|12178,12187|false|false|false|C0442805;C5236002|Increase;Increased (finding)|increased
Finding|Functional Concept|SIMPLE_SEGMENT|12178,12187|false|false|false|C0442805;C5236002|Increase;Increased (finding)|increased
Event|Event|SIMPLE_SEGMENT|12188,12192|false|false|false|||work
Event|Occupational Activity|SIMPLE_SEGMENT|12188,12192|false|false|false|C0043227|Work|work
Event|Event|SIMPLE_SEGMENT|12196,12205|false|false|false|||breathing
Finding|Finding|SIMPLE_SEGMENT|12214,12219|false|false|false|C0150312|Present|Found
Finding|Idea or Concept|SIMPLE_SEGMENT|12229,12240|false|false|false|C0750502|Significant|significant
Event|Event|SIMPLE_SEGMENT|12241,12250|false|false|false|||worsening
Finding|Idea or Concept|SIMPLE_SEGMENT|12241,12250|false|false|false|C1546960|Patient Outcome - Worsening|worsening
Anatomy|Tissue|SIMPLE_SEGMENT|12256,12263|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12256,12263|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Body Substance|SIMPLE_SEGMENT|12256,12272|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Finding|Finding|SIMPLE_SEGMENT|12256,12272|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|12256,12272|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Event|Event|SIMPLE_SEGMENT|12264,12272|false|false|false|||effusion
Finding|Body Substance|SIMPLE_SEGMENT|12264,12272|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|SIMPLE_SEGMENT|12264,12272|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|12264,12272|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Event|Event|SIMPLE_SEGMENT|12277,12288|false|false|false|||development
Finding|Functional Concept|SIMPLE_SEGMENT|12277,12288|false|false|false|C0018271;C0243107;C0678723;C1527148|Development;Growth and Development function;biological development;development aspects|development
Finding|Organism Function|SIMPLE_SEGMENT|12277,12288|false|false|false|C0018271;C0243107;C0678723;C1527148|Development;Growth and Development function;biological development;development aspects|development
Anatomy|Tissue|SIMPLE_SEGMENT|12295,12302|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12295,12302|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Body Substance|SIMPLE_SEGMENT|12295,12311|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Finding|Finding|SIMPLE_SEGMENT|12295,12311|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|12295,12311|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Event|Event|SIMPLE_SEGMENT|12303,12311|false|false|false|||effusion
Finding|Body Substance|SIMPLE_SEGMENT|12303,12311|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|SIMPLE_SEGMENT|12303,12311|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|12303,12311|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Finding|SIMPLE_SEGMENT|12313,12332|false|false|false|C5555338|Intubation Required|Required intubation
Event|Event|SIMPLE_SEGMENT|12322,12332|false|false|false|||intubation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|12322,12332|false|false|false|C0021925|Intubation (procedure)|intubation
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12337,12348|false|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|SIMPLE_SEGMENT|12337,12348|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|SIMPLE_SEGMENT|12337,12348|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|SIMPLE_SEGMENT|12337,12348|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Event|Event|SIMPLE_SEGMENT|12349,12354|false|false|false|||state
Finding|Functional Concept|SIMPLE_SEGMENT|12349,12354|false|false|false|C1442792|State|state
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|12364,12371|false|false|false|C0018787|Heart|Cardiac
Event|Event|SIMPLE_SEGMENT|12364,12371|false|false|false|||Cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|12364,12371|false|false|false|C1314974|Cardiac attachment|Cardiac
Event|Event|SIMPLE_SEGMENT|12376,12382|false|false|false|||showed
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|12398,12407|true|false|false|C1179435|Protein Component|component
Drug|Biologically Active Substance|SIMPLE_SEGMENT|12398,12407|true|false|false|C1179435|Protein Component|component
Event|Event|SIMPLE_SEGMENT|12398,12407|false|false|false|||component
Finding|Conceptual Entity|SIMPLE_SEGMENT|12398,12407|true|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Finding|Idea or Concept|SIMPLE_SEGMENT|12398,12407|true|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Finding|Intellectual Product|SIMPLE_SEGMENT|12398,12407|true|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Event|Event|SIMPLE_SEGMENT|12425,12430|false|false|false|||fever
Finding|Finding|SIMPLE_SEGMENT|12425,12430|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|12425,12430|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Event|Event|SIMPLE_SEGMENT|12438,12445|false|false|false|||started
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|12457,12461|false|false|false|C0535219|SMC3 protein, human|HCAP
Drug|Biologically Active Substance|SIMPLE_SEGMENT|12457,12461|false|false|false|C0535219|SMC3 protein, human|HCAP
Event|Event|SIMPLE_SEGMENT|12457,12461|false|false|false|||HCAP
Finding|Gene or Genome|SIMPLE_SEGMENT|12457,12461|false|false|false|C1419431;C1422826;C1704469;C1822780|DCD gene;RNGTT gene;SMC3 gene;SMC3 wt Allele|HCAP
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|12457,12461|false|false|false|C0056451|Cyclophosphamide/Altretamine/Doxorubicin/Cisplatin Regimen|HCAP
Event|Event|SIMPLE_SEGMENT|12462,12470|false|false|false|||coverage
Finding|Functional Concept|SIMPLE_SEGMENT|12462,12470|false|false|false|C1551362;C1999244;C3854012|coverage - HL7PublishingDomain;coverage - financial contract|coverage
Finding|Idea or Concept|SIMPLE_SEGMENT|12462,12470|false|false|false|C1551362;C1999244;C3854012|coverage - HL7PublishingDomain;coverage - financial contract|coverage
Finding|Intellectual Product|SIMPLE_SEGMENT|12462,12470|false|false|false|C1551362;C1999244;C3854012|coverage - HL7PublishingDomain;coverage - financial contract|coverage
Event|Event|SIMPLE_SEGMENT|12478,12486|false|false|false|||mini-BAL
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|12478,12486|false|false|false|C3161394|Mini-bronchoalveolar lavage|mini-BAL
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|12502,12516|false|false|false|C0184661;C2183254|Interventional procedure;interventional (invasive) radiology|Interventional
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|12502,12516|false|false|false|C0184661;C2183254|Interventional procedure;interventional (invasive) radiology|Interventional
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|12517,12526|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12517,12526|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|12517,12526|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Event|Event|SIMPLE_SEGMENT|12532,12541|false|false|false|||consulted
Finding|Functional Concept|SIMPLE_SEGMENT|12564,12569|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Event|Event|SIMPLE_SEGMENT|12576,12589|false|false|false|||thoracentesis
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|12576,12589|false|false|false|C0189477|Thoracentesis|thoracentesis
Event|Event|SIMPLE_SEGMENT|12604,12613|false|false|false|||placement
Procedure|Health Care Activity|SIMPLE_SEGMENT|12604,12613|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|12604,12613|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Event|Event|SIMPLE_SEGMENT|12618,12621|false|false|false|||saw
Drug|Inorganic Chemical|SIMPLE_SEGMENT|12645,12653|false|false|false|C0723457|Stop brand of fluoride|stopping
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12645,12653|false|false|false|C0723457|Stop brand of fluoride|stopping
Event|Event|SIMPLE_SEGMENT|12645,12653|false|false|false|||stopping
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|12655,12660|false|false|false|C0042313|vancomycin|Vanco
Drug|Antibiotic|SIMPLE_SEGMENT|12655,12660|false|false|false|C0042313|vancomycin|Vanco
Event|Event|SIMPLE_SEGMENT|12655,12660|false|false|false|||Vanco
Drug|Antibiotic|SIMPLE_SEGMENT|12661,12669|false|false|false|C0055003|cefepime|cefepime
Drug|Organic Chemical|SIMPLE_SEGMENT|12661,12669|false|false|false|C0055003|cefepime|cefepime
Event|Event|SIMPLE_SEGMENT|12661,12669|false|false|false|||cefepime
Event|Event|SIMPLE_SEGMENT|12673,12680|false|false|false|||unclear
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12691,12700|false|false|false|C0032285|Pneumonia|pneumonia
Event|Event|SIMPLE_SEGMENT|12691,12700|false|false|false|||pneumonia
Event|Event|SIMPLE_SEGMENT|12705,12713|false|false|false|||starting
Drug|Antibiotic|SIMPLE_SEGMENT|12715,12726|false|false|false|C1260298|tigecycline|Tigecycline
Drug|Organic Chemical|SIMPLE_SEGMENT|12715,12726|false|false|false|C1260298|tigecycline|Tigecycline
Event|Event|SIMPLE_SEGMENT|12715,12726|false|false|false|||Tigecycline
Finding|Functional Concept|SIMPLE_SEGMENT|12736,12741|false|false|false|C1999244||cover
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|12747,12751|false|false|false|C0535219|SMC3 protein, human|HCAP
Drug|Biologically Active Substance|SIMPLE_SEGMENT|12747,12751|false|false|false|C0535219|SMC3 protein, human|HCAP
Event|Event|SIMPLE_SEGMENT|12747,12751|false|false|false|||HCAP
Finding|Gene or Genome|SIMPLE_SEGMENT|12747,12751|false|false|false|C1419431;C1422826;C1704469;C1822780|DCD gene;RNGTT gene;SMC3 gene;SMC3 wt Allele|HCAP
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|12747,12751|false|false|false|C0056451|Cyclophosphamide/Altretamine/Doxorubicin/Cisplatin Regimen|HCAP
Event|Event|SIMPLE_SEGMENT|12752,12761|false|false|false|||organisms
Event|Event|SIMPLE_SEGMENT|12771,12776|false|false|false|||treat
Event|Event|SIMPLE_SEGMENT|12785,12793|false|false|false|||Mini-BAL
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|12785,12793|false|false|false|C3161394|Mini-bronchoalveolar lavage|Mini-BAL
Anatomy|Tissue|SIMPLE_SEGMENT|12798,12805|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12798,12805|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Body Substance|SIMPLE_SEGMENT|12798,12811|false|false|false|C0225778|Pleural fluid|pleural fluid
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|12798,12811|false|false|false|C2242629|Pleural fluid analysis|pleural fluid
Drug|Substance|SIMPLE_SEGMENT|12806,12811|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|12806,12811|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|12806,12811|false|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Classification|SIMPLE_SEGMENT|12817,12825|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|12817,12825|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|12817,12825|false|false|false|C5237010|Expression Negative|negative
Event|Event|SIMPLE_SEGMENT|12826,12834|false|false|false|||cultures
Finding|Idea or Concept|SIMPLE_SEGMENT|12826,12834|false|true|false|C0010453|Culture (Anthropological)|cultures
Event|Event|SIMPLE_SEGMENT|12845,12853|false|false|false|||diuresis
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|12845,12853|false|false|false|C0012797|Diuresis|diuresis
Event|Event|SIMPLE_SEGMENT|12878,12884|false|false|false|||weaned
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12889,12897|false|false|false|C0237795|Pressors|pressors
Event|Event|SIMPLE_SEGMENT|12889,12897|false|false|false|||pressors
Event|Event|SIMPLE_SEGMENT|12903,12912|false|false|false|||extubated
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|12903,12912|false|false|false|C0553891|Tracheal Extubation|extubated
Event|Event|SIMPLE_SEGMENT|12922,12928|false|false|false|||weaned
Drug|Biologically Active Substance|SIMPLE_SEGMENT|12937,12943|false|false|false|C0030054|oxygen|oxygen
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|12937,12943|false|false|false|C0030054|oxygen|oxygen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12937,12943|false|false|false|C0030054|oxygen|oxygen
Event|Event|SIMPLE_SEGMENT|12937,12943|false|false|false|||oxygen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|12937,12943|false|false|false|C0184633|Oxygen Therapy Care|oxygen
Finding|Finding|SIMPLE_SEGMENT|12951,12955|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|12951,12955|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|12951,12955|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|SIMPLE_SEGMENT|12960,12969|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|12960,12969|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|12960,12969|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|12960,12969|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|12960,12969|false|false|false|C0030685|Patient Discharge|discharge
Finding|Functional Concept|SIMPLE_SEGMENT|12974,12979|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12988,12993|false|false|false|C1410088|Still|still
Event|Event|SIMPLE_SEGMENT|12994,13002|false|false|false|||draining
Finding|Idea or Concept|SIMPLE_SEGMENT|13017,13020|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|13017,13020|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|13028,13034|false|false|false|||follow
Event|Event|SIMPLE_SEGMENT|13052,13061|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|13052,13061|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|13052,13061|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|13052,13061|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|13052,13061|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|SIMPLE_SEGMENT|13073,13080|false|false|false|||require
Finding|Idea or Concept|SIMPLE_SEGMENT|13082,13089|false|false|false|C0549178|Continuous|ongoing
Event|Event|SIMPLE_SEGMENT|13090,13098|false|false|false|||diuresis
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|13090,13098|false|false|false|C0012797|Diuresis|diuresis
Finding|Idea or Concept|SIMPLE_SEGMENT|13109,13120|false|false|false|C0750502|Significant|significant
Finding|Intellectual Product|SIMPLE_SEGMENT|13121,13127|false|false|false|C1705102|Volume (publication)|volume
Finding|Pathologic Function|SIMPLE_SEGMENT|13121,13136|false|false|false|C0546817|Hypervolemia (finding)|volume overload
Event|Event|SIMPLE_SEGMENT|13128,13136|false|false|false|||overload
Event|Event|SIMPLE_SEGMENT|13143,13151|false|false|false|||responds
Finding|Finding|SIMPLE_SEGMENT|13152,13156|false|false|false|C5575035|Well (answer to question)|well
Drug|Organic Chemical|SIMPLE_SEGMENT|13167,13172|false|false|false|C0699992|Lasix|Lasix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13167,13172|false|false|false|C0699992|Lasix|Lasix
Event|Event|SIMPLE_SEGMENT|13190,13198|false|false|false|||negative
Finding|Classification|SIMPLE_SEGMENT|13190,13198|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|13190,13198|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|13190,13198|false|false|false|C5237010|Expression Negative|negative
Event|Event|SIMPLE_SEGMENT|13212,13219|false|false|false|||leading
Event|Event|SIMPLE_SEGMENT|13226,13235|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|13226,13235|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|13226,13235|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|13226,13235|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|13226,13235|false|false|false|C0030685|Patient Discharge|discharge
Finding|Mental Process|SIMPLE_SEGMENT|13248,13254|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13248,13261|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|SIMPLE_SEGMENT|13248,13261|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13255,13261|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|13255,13261|false|false|false|C1546481|What subject filter - Status|Status
Finding|Mental Process|SIMPLE_SEGMENT|13267,13274|false|false|false|C0542559|contextual factors|setting
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13278,13285|false|false|false|C0032930|Precipitating Factors|trigger
Event|Event|SIMPLE_SEGMENT|13278,13285|false|false|false|||trigger
Event|Event|SIMPLE_SEGMENT|13290,13297|false|false|false|||hypoxia
Finding|Finding|SIMPLE_SEGMENT|13290,13297|false|false|false|C0242184;C1963140|Hypoxia;Hypoxia, CTCAE|hypoxia
Finding|Pathologic Function|SIMPLE_SEGMENT|13290,13297|false|false|false|C0242184;C1963140|Hypoxia;Hypoxia, CTCAE|hypoxia
Event|Event|SIMPLE_SEGMENT|13307,13315|false|false|false|||transfer
Finding|Functional Concept|SIMPLE_SEGMENT|13307,13315|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|SIMPLE_SEGMENT|13307,13315|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|SIMPLE_SEGMENT|13307,13315|false|false|false|C4706767|Transfer (immobility management)|transfer
Event|Event|SIMPLE_SEGMENT|13335,13342|false|false|false|||concern
Finding|Idea or Concept|SIMPLE_SEGMENT|13335,13342|false|false|false|C2699424|Concern|concern
Event|Event|SIMPLE_SEGMENT|13361,13371|false|false|false|||responsive
Finding|Functional Concept|SIMPLE_SEGMENT|13361,13371|false|false|false|C0205342|Responsive|responsive
Event|Event|SIMPLE_SEGMENT|13377,13384|false|false|false|||concern
Finding|Idea or Concept|SIMPLE_SEGMENT|13377,13384|false|false|false|C2699424|Concern|concern
Event|Event|SIMPLE_SEGMENT|13396,13404|false|false|false|||defecits
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|13406,13410|false|false|false|C1366753|STAT protein|Stat
Drug|Biologically Active Substance|SIMPLE_SEGMENT|13406,13410|false|false|false|C1366753|STAT protein|Stat
Finding|Gene or Genome|SIMPLE_SEGMENT|13406,13410|false|false|false|C1335960;C1420304;C1547583;C1548425;C1561443|Extended Priority Codes - Stat;Referral priority - STAT;Report priority - Stat;SOAT1 gene;STAT family gene|Stat
Finding|Idea or Concept|SIMPLE_SEGMENT|13406,13410|false|false|false|C1335960;C1420304;C1547583;C1548425;C1561443|Extended Priority Codes - Stat;Referral priority - STAT;Report priority - Stat;SOAT1 gene;STAT family gene|Stat
Finding|Intellectual Product|SIMPLE_SEGMENT|13406,13410|false|false|false|C1335960;C1420304;C1547583;C1548425;C1561443|Extended Priority Codes - Stat;Referral priority - STAT;Report priority - Stat;SOAT1 gene;STAT family gene|Stat
Anatomy|Body Location or Region|SIMPLE_SEGMENT|13411,13415|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|13411,13415|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13411,13415|false|false|false|C0362076|Problems with head|head
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|13411,13415|false|false|false|C0876917|Procedure on head|head
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|13411,13418|false|false|false|C0202691|CAT scan of head|head CT
Event|Event|SIMPLE_SEGMENT|13416,13418|false|false|false|||CT
Event|Event|SIMPLE_SEGMENT|13427,13435|false|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|13427,13435|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|13427,13438|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13439,13445|true|false|false|C0038454|Cerebrovascular accident|stroke
Event|Event|SIMPLE_SEGMENT|13439,13445|false|false|false|||stroke
Finding|Finding|SIMPLE_SEGMENT|13439,13445|true|false|false|C5977286|Stroke (heart beat)|stroke
Event|Event|SIMPLE_SEGMENT|13450,13455|false|false|false|||bleed
Finding|Pathologic Function|SIMPLE_SEGMENT|13450,13455|false|false|false|C0019080|Hemorrhage|bleed
Event|Event|SIMPLE_SEGMENT|13467,13476|false|false|false|||consulted
Event|Event|SIMPLE_SEGMENT|13481,13485|false|false|false|||said
Event|Event|SIMPLE_SEGMENT|13486,13493|false|false|false|||nothing
Event|Event|SIMPLE_SEGMENT|13504,13512|false|false|false|||deficits
Event|Event|SIMPLE_SEGMENT|13514,13522|false|false|false|||resolved
Finding|Idea or Concept|SIMPLE_SEGMENT|13528,13532|false|false|false|C1552851|next - HtmlLinkType|next
Event|Event|SIMPLE_SEGMENT|13538,13541|false|false|false|||EEG
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|13538,13541|false|false|false|C0013819|Electroencephalography|EEG
Event|Event|SIMPLE_SEGMENT|13552,13559|false|false|false|||ordered
Finding|Intellectual Product|SIMPLE_SEGMENT|13564,13568|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|SIMPLE_SEGMENT|13570,13578|false|false|false|||canceled
Event|Event|SIMPLE_SEGMENT|13585,13595|false|false|false|||discussion
Finding|Social Behavior|SIMPLE_SEGMENT|13585,13595|false|false|false|C2584313|Discussion (communication)|discussion
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|13585,13595|false|false|false|C0557061|Discussion (procedure)|discussion
Event|Event|SIMPLE_SEGMENT|13601,13606|false|false|false|||neuro
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|13608,13612|false|false|false|C1742913|REST protein, human|Rest
Drug|Biologically Active Substance|SIMPLE_SEGMENT|13608,13612|false|false|false|C1742913|REST protein, human|Rest
Event|Event|SIMPLE_SEGMENT|13608,13612|false|false|false|||Rest
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|13608,13612|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|Rest
Finding|Gene or Genome|SIMPLE_SEGMENT|13608,13612|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|Rest
Finding|Molecular Function|SIMPLE_SEGMENT|13608,13612|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|Rest
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|13616,13619|false|false|false|C0228479|Structure of intraculminate fissure|ICU
Finding|Intellectual Product|SIMPLE_SEGMENT|13616,13619|false|false|false|C4554035|Inventory of Callous-Unemotional Traits|ICU
Event|Event|SIMPLE_SEGMENT|13643,13651|false|false|false|||delerium
Event|Event|SIMPLE_SEGMENT|13668,13677|false|false|false|||requiring
Event|Event|SIMPLE_SEGMENT|13683,13688|false|false|false|||doses
Drug|Organic Chemical|SIMPLE_SEGMENT|13693,13703|false|false|false|C0171023|olanzapine|Olanzapine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13693,13703|false|false|false|C0171023|olanzapine|Olanzapine
Event|Event|SIMPLE_SEGMENT|13693,13703|false|false|false|||Olanzapine
Event|Event|SIMPLE_SEGMENT|13718,13726|false|false|false|||improved
Finding|Finding|SIMPLE_SEGMENT|13730,13734|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|13730,13734|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|13730,13734|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|13738,13741|false|false|false|C0228479|Structure of intraculminate fissure|ICU
Finding|Intellectual Product|SIMPLE_SEGMENT|13738,13741|false|false|false|C4554035|Inventory of Callous-Unemotional Traits|ICU
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13755,13760|false|false|false|C1410088|Still|still
Event|Event|SIMPLE_SEGMENT|13755,13760|false|false|false|||still
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|13771,13781|false|false|false|C1142436|Sundowning|sundowning
Event|Event|SIMPLE_SEGMENT|13771,13781|false|false|false|||sundowning
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13786,13798|false|false|false|C0020625|Hyponatremia|Hyponatremia
Event|Event|SIMPLE_SEGMENT|13786,13798|false|false|false|||Hyponatremia
Finding|Body Substance|SIMPLE_SEGMENT|13800,13807|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|13800,13807|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|13800,13807|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Finding|SIMPLE_SEGMENT|13830,13836|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Finding|Idea or Concept|SIMPLE_SEGMENT|13830,13836|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|13837,13848|false|true|false|C0752266|Hypovolemic|hypovolemic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13850,13862|false|true|false|C0020625|Hyponatremia|hyponatremia
Event|Event|SIMPLE_SEGMENT|13850,13862|false|false|false|||hyponatremia
Event|Event|SIMPLE_SEGMENT|13866,13873|false|false|false|||setting
Finding|Mental Process|SIMPLE_SEGMENT|13866,13873|false|false|false|C0542559|contextual factors|setting
Event|Event|SIMPLE_SEGMENT|13877,13885|false|false|false|||diarrhea
Finding|Finding|SIMPLE_SEGMENT|13877,13885|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|SIMPLE_SEGMENT|13877,13885|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Intellectual Product|SIMPLE_SEGMENT|13886,13890|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|poor
Event|Event|SIMPLE_SEGMENT|13894,13900|false|false|false|||intake
Finding|Functional Concept|SIMPLE_SEGMENT|13894,13900|false|false|false|C1512806|Intake|intake
Procedure|Health Care Activity|SIMPLE_SEGMENT|13894,13900|false|false|false|C3251814;C4521161|Intake (treatment);Measurement of fluid intake|intake
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13917,13922|false|false|false|C0021141|Inappropriate ADH Syndrome|SIADH
Event|Event|SIMPLE_SEGMENT|13917,13922|false|false|false|||SIADH
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13929,13938|false|true|false|C0032285|Pneumonia|pneumonia
Event|Event|SIMPLE_SEGMENT|13929,13938|false|false|false|||pneumonia
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13940,13944|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|13940,13944|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|13940,13944|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|13940,13944|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|13951,13957|false|false|false|||review
Finding|Idea or Concept|SIMPLE_SEGMENT|13951,13957|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Finding|Intellectual Product|SIMPLE_SEGMENT|13951,13957|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Finding|Functional Concept|SIMPLE_SEGMENT|13951,13960|false|false|false|C0699752|Review of|review of
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|13965,13969|false|false|false|C0587081|Laboratory test finding|labs
Finding|Body Substance|SIMPLE_SEGMENT|13971,13978|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|13971,13978|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|13971,13978|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|13980,13985|false|false|false|C4050225|Often - answer to question|often
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13986,13998|false|false|false|C0857122|Hyponatraemic|hyponatremic
Event|Event|SIMPLE_SEGMENT|13986,13998|false|false|false|||hyponatremic
Event|Event|SIMPLE_SEGMENT|14002,14012|false|false|false|||outpatient
Finding|Classification|SIMPLE_SEGMENT|14002,14012|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|14002,14012|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Finding|SIMPLE_SEGMENT|14016,14020|false|false|false|C5575035|Well (answer to question)|well
Finding|Body Substance|SIMPLE_SEGMENT|14022,14027|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Finding|Functional Concept|SIMPLE_SEGMENT|14022,14027|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Finding|Intellectual Product|SIMPLE_SEGMENT|14022,14027|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Event|Event|SIMPLE_SEGMENT|14034,14043|false|false|false|||confusing
Finding|Mental Process|SIMPLE_SEGMENT|14048,14055|false|false|false|C0542559|contextual factors|setting
Finding|Pathologic Function|SIMPLE_SEGMENT|14059,14064|false|false|false|C0036974|Shock|shock
Finding|Body Substance|SIMPLE_SEGMENT|14068,14073|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Functional Concept|SIMPLE_SEGMENT|14068,14073|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Intellectual Product|SIMPLE_SEGMENT|14068,14073|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Event|Event|SIMPLE_SEGMENT|14101,14109|false|false|false|||question
Finding|Intellectual Product|SIMPLE_SEGMENT|14101,14109|false|false|false|C1522634|Question (inquiry)|question
Drug|Biologically Active Substance|SIMPLE_SEGMENT|14114,14120|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|14114,14120|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14114,14120|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Event|Event|SIMPLE_SEGMENT|14114,14120|false|false|false|||sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|14114,14120|false|false|false|C4553025|Sodium metabolic function|sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|14114,14120|false|false|false|C0337443|Sodium measurement|sodium
Event|Event|SIMPLE_SEGMENT|14121,14128|false|false|false|||wasting
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|14129,14134|false|false|false|C0022646|Kidney|renal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14129,14134|false|false|false|C0042075|Urologic Diseases|renal
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|14129,14141|false|false|false|C0160420|Injury of kidney|renal injury
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|14135,14141|false|false|false|C3263722;C3263723|Traumatic AND/OR non-traumatic injury;Traumatic injury|injury
Event|Event|SIMPLE_SEGMENT|14135,14141|false|false|false|||injury
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14143,14155|false|false|false|C0020625|Hyponatremia|Hyponatremia
Event|Event|SIMPLE_SEGMENT|14143,14155|false|false|false|||Hyponatremia
Event|Event|SIMPLE_SEGMENT|14156,14163|false|false|false|||started
Event|Event|SIMPLE_SEGMENT|14167,14174|false|false|false|||resolve
Finding|Conceptual Entity|SIMPLE_SEGMENT|14167,14174|false|false|false|C2699488|Resolution|resolve
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|14167,14174|false|false|false|C5401470|RESOLVE Multishot Diffusion Weighted Echoplanar Imaging|resolve
Finding|Intellectual Product|SIMPLE_SEGMENT|14179,14186|false|false|false|C0282416|Overall Publication Type|overall
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14187,14196|false|false|false|C3864998||condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14187,14196|false|false|false|C0012634|Disease|condition
Event|Event|SIMPLE_SEGMENT|14187,14196|false|false|false|||condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|14187,14196|false|false|false|C1705253|Logical Condition|condition
Event|Event|SIMPLE_SEGMENT|14197,14205|false|false|false|||improved
Event|Event|SIMPLE_SEGMENT|14218,14228|false|false|false|||re-develop
Event|Event|SIMPLE_SEGMENT|14238,14245|false|false|false|||setting
Finding|Mental Process|SIMPLE_SEGMENT|14238,14245|false|false|false|C0542559|contextual factors|setting
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|14253,14256|false|false|false|C0228479|Structure of intraculminate fissure|ICU
Finding|Intellectual Product|SIMPLE_SEGMENT|14253,14256|false|false|false|C4554035|Inventory of Callous-Unemotional Traits|ICU
Event|Event|SIMPLE_SEGMENT|14257,14268|false|false|false|||readmission
Procedure|Health Care Activity|SIMPLE_SEGMENT|14257,14268|false|false|false|C4489276|Readmission|readmission
Event|Event|SIMPLE_SEGMENT|14273,14280|false|false|false|||hypoxia
Finding|Finding|SIMPLE_SEGMENT|14273,14280|false|false|false|C0242184;C1963140|Hypoxia;Hypoxia, CTCAE|hypoxia
Finding|Pathologic Function|SIMPLE_SEGMENT|14273,14280|false|false|false|C0242184;C1963140|Hypoxia;Hypoxia, CTCAE|hypoxia
Finding|Body Substance|SIMPLE_SEGMENT|14290,14297|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|14290,14297|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|14290,14297|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Biologically Active Substance|SIMPLE_SEGMENT|14303,14313|false|false|false|C0010294|creatinine|creatinine
Drug|Organic Chemical|SIMPLE_SEGMENT|14303,14313|false|false|false|C0010294|creatinine|creatinine
Event|Event|SIMPLE_SEGMENT|14303,14313|false|false|false|||creatinine
Finding|Physiologic Function|SIMPLE_SEGMENT|14303,14313|false|false|false|C4551889|Creatinine metabolic function|creatinine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|14303,14313|false|false|false|C0201975|Creatinine measurement|creatinine
Finding|Finding|SIMPLE_SEGMENT|14321,14333|false|false|false|C4533677|at admission|at admission
Event|Event|SIMPLE_SEGMENT|14324,14333|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|14324,14333|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|14350,14358|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|SIMPLE_SEGMENT|14350,14358|false|false|false|||baseline
Finding|Idea or Concept|SIMPLE_SEGMENT|14350,14358|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Finding|Finding|SIMPLE_SEGMENT|14373,14379|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Finding|Idea or Concept|SIMPLE_SEGMENT|14373,14379|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Finding|Conceptual Entity|SIMPLE_SEGMENT|14390,14398|false|true|false|C0015127;C1314792;C1524003|Etiology;Etiology aspects;Science of Etiology|etiology
Finding|Functional Concept|SIMPLE_SEGMENT|14390,14398|false|true|false|C0015127;C1314792;C1524003|Etiology;Etiology aspects;Science of Etiology|etiology
Event|Event|SIMPLE_SEGMENT|14403,14410|false|false|false|||setting
Finding|Mental Process|SIMPLE_SEGMENT|14403,14410|false|false|false|C0542559|contextual factors|setting
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14414,14423|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|SIMPLE_SEGMENT|14414,14423|false|false|false|||infection
Finding|Pathologic Function|SIMPLE_SEGMENT|14414,14423|false|false|false|C3714514|Infection|infection
Event|Event|SIMPLE_SEGMENT|14425,14433|false|false|false|||diarrhea
Finding|Finding|SIMPLE_SEGMENT|14425,14433|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|SIMPLE_SEGMENT|14425,14433|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Intellectual Product|SIMPLE_SEGMENT|14435,14439|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|poor
Event|Event|SIMPLE_SEGMENT|14443,14449|false|false|false|||intake
Finding|Functional Concept|SIMPLE_SEGMENT|14443,14449|false|false|false|C1512806|Intake|intake
Procedure|Health Care Activity|SIMPLE_SEGMENT|14443,14449|false|false|false|C3251814;C4521161|Intake (treatment);Measurement of fluid intake|intake
Finding|Finding|SIMPLE_SEGMENT|14496,14502|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|14496,14502|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Intellectual Product|SIMPLE_SEGMENT|14508,14512|false|true|false|C1547225|Mild Severity of Illness Code|mild
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14513,14516|false|true|false|C4551504|Oculocutaneous albinism type 1A|ATN
Event|Event|SIMPLE_SEGMENT|14513,14516|false|false|false|||ATN
Finding|Gene or Genome|SIMPLE_SEGMENT|14513,14516|false|true|false|C1710338|TYR wt Allele|ATN
Finding|Mental Process|SIMPLE_SEGMENT|14520,14527|false|false|false|C0542559|contextual factors|setting
Event|Event|SIMPLE_SEGMENT|14555,14566|false|false|false|||hypotension
Finding|Finding|SIMPLE_SEGMENT|14555,14566|false|false|false|C0020649|Hypotension|hypotension
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|14568,14578|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14568,14578|false|false|false|C0065374|lisinopril|Lisinopril
Event|Event|SIMPLE_SEGMENT|14568,14578|false|false|false|||Lisinopril
Event|Event|SIMPLE_SEGMENT|14583,14587|false|false|false|||held
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|14598,14601|false|false|false|C0228479|Structure of intraculminate fissure|ICU
Finding|Intellectual Product|SIMPLE_SEGMENT|14598,14601|false|false|false|C4554035|Inventory of Callous-Unemotional Traits|ICU
Event|Event|SIMPLE_SEGMENT|14615,14626|false|false|false|||hypotension
Finding|Finding|SIMPLE_SEGMENT|14615,14626|false|false|false|C0020649|Hypotension|hypotension
Event|Event|SIMPLE_SEGMENT|14631,14638|false|false|false|||trended
Event|Event|SIMPLE_SEGMENT|14639,14643|false|false|false|||back
Event|Event|SIMPLE_SEGMENT|14669,14675|false|false|false|||stayed
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|14686,14690|false|false|false|C1742913|REST protein, human|rest
Drug|Biologically Active Substance|SIMPLE_SEGMENT|14686,14690|false|false|false|C1742913|REST protein, human|rest
Event|Event|SIMPLE_SEGMENT|14686,14690|false|false|false|||rest
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|14686,14690|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Gene or Genome|SIMPLE_SEGMENT|14686,14690|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Molecular Function|SIMPLE_SEGMENT|14686,14690|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Event|Event|SIMPLE_SEGMENT|14694,14709|false|false|false|||hospitalization
Procedure|Health Care Activity|SIMPLE_SEGMENT|14694,14709|false|true|false|C0019993|Hospitalization|hospitalization
Finding|Mental Process|SIMPLE_SEGMENT|14718,14725|false|false|false|C0542559|contextual factors|setting
Finding|Functional Concept|SIMPLE_SEGMENT|14730,14736|false|false|false|C1522484;C1561503;C1705190|Precision - second;Second Suffix;metastatic qualifier|second
Finding|Idea or Concept|SIMPLE_SEGMENT|14730,14736|false|false|false|C1522484;C1561503;C1705190|Precision - second;Second Suffix;metastatic qualifier|second
Finding|Intellectual Product|SIMPLE_SEGMENT|14730,14736|false|false|false|C1522484;C1561503;C1705190|Precision - second;Second Suffix;metastatic qualifier|second
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|14737,14740|false|false|false|C0228479|Structure of intraculminate fissure|ICU
Finding|Intellectual Product|SIMPLE_SEGMENT|14737,14740|false|false|false|C4554035|Inventory of Callous-Unemotional Traits|ICU
Event|Event|SIMPLE_SEGMENT|14741,14752|false|false|false|||readmission
Procedure|Health Care Activity|SIMPLE_SEGMENT|14741,14752|false|false|false|C4489276|Readmission|readmission
Finding|Finding|SIMPLE_SEGMENT|14757,14765|false|false|false|C1547420;C1608263;C1608264;C3244313;C3834263;C3890554|Certificate Status - Inactive;Edit Status - Inactive;Immunization Registry Status - Inactive;Inactive - answer to question;Inactive Healthcare Coverage;Physical Inactivity|Inactive
Finding|Idea or Concept|SIMPLE_SEGMENT|14757,14765|false|false|false|C1547420;C1608263;C1608264;C3244313;C3834263;C3890554|Certificate Status - Inactive;Edit Status - Inactive;Immunization Registry Status - Inactive;Inactive - answer to question;Inactive Healthcare Coverage;Physical Inactivity|Inactive
Event|Event|SIMPLE_SEGMENT|14766,14772|false|false|false|||issues
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14778,14792|false|false|false|C0020676|Hypothyroidism|Hypothyroidism
Event|Event|SIMPLE_SEGMENT|14778,14792|false|false|false|||Hypothyroidism
Event|Event|SIMPLE_SEGMENT|14794,14803|false|false|false|||Continued
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|14804,14817|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Hormone|SIMPLE_SEGMENT|14804,14817|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Organic Chemical|SIMPLE_SEGMENT|14804,14817|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14804,14817|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Event|Event|SIMPLE_SEGMENT|14804,14817|false|false|false|||levothyroxine
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14834,14846|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|SIMPLE_SEGMENT|14834,14846|false|false|false|||Hypertension
Event|Event|SIMPLE_SEGMENT|14855,14866|false|false|false|||hypotension
Finding|Finding|SIMPLE_SEGMENT|14855,14866|false|false|false|C0020649|Hypotension|hypotension
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14872,14878|false|false|false|C0036690;C0243026|Sepsis;Septicemia|sepsis
Event|Event|SIMPLE_SEGMENT|14872,14878|false|false|false|||sepsis
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|14880,14890|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14880,14890|false|false|false|C0065374|lisinopril|lisinopril
Event|Event|SIMPLE_SEGMENT|14880,14890|false|false|false|||lisinopril
Event|Event|SIMPLE_SEGMENT|14896,14900|false|false|false|||held
Event|Event|SIMPLE_SEGMENT|14906,14914|false|false|false|||remained
Finding|Finding|SIMPLE_SEGMENT|14915,14919|false|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|14920,14930|false|false|false|||controlled
Event|Event|SIMPLE_SEGMENT|14945,14953|false|false|false|||continue
Event|Event|SIMPLE_SEGMENT|14961,14965|false|false|false|||held
Event|Event|SIMPLE_SEGMENT|14969,14978|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|14969,14978|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|14969,14978|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|14969,14978|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|14969,14978|false|false|false|C0030685|Patient Discharge|discharge
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14983,14987|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Event|Event|SIMPLE_SEGMENT|14983,14987|false|false|false|||GERD
Drug|Organic Chemical|SIMPLE_SEGMENT|14989,14999|false|false|false|C0028978|omeprazole|Omeprazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14989,14999|false|false|false|C0028978|omeprazole|Omeprazole
Event|Event|SIMPLE_SEGMENT|15000,15007|false|false|false|||stopped
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|15029,15037|false|false|false|C4727483|BRAF Gene Rearrangement|positive
Event|Event|SIMPLE_SEGMENT|15029,15037|false|false|false|||positive
Finding|Classification|SIMPLE_SEGMENT|15029,15037|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|SIMPLE_SEGMENT|15029,15037|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|SIMPLE_SEGMENT|15044,15048|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|15044,15048|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|15044,15048|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|SIMPLE_SEGMENT|15053,15056|false|false|false|||put
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|15060,15070|false|false|false|C0019593|Histamine H2 Antagonists|H2 blocker
Event|Event|SIMPLE_SEGMENT|15063,15070|false|false|false|||blocker
Event|Event|SIMPLE_SEGMENT|15078,15089|false|false|false|||prophylaxis
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|15078,15089|false|false|false|C0199176|Prophylactic treatment|prophylaxis
Event|Event|SIMPLE_SEGMENT|15099,15106|false|false|false|||stopped
Event|Event|SIMPLE_SEGMENT|15133,15140|false|false|false|||started
Event|Event|SIMPLE_SEGMENT|15141,15149|false|false|false|||feeeding
Event|Event|SIMPLE_SEGMENT|15154,15158|false|false|false|||Code
Event|Occupational Activity|SIMPLE_SEGMENT|15154,15158|false|false|false|C0009219|Coding|Code
Finding|Intellectual Product|SIMPLE_SEGMENT|15154,15158|false|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|Code
Event|Event|SIMPLE_SEGMENT|15166,15175|false|false|false|||confirmed
Finding|Body Substance|SIMPLE_SEGMENT|15181,15188|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|15181,15188|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|15181,15188|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Gene or Genome|SIMPLE_SEGMENT|15190,15193|false|false|false|C1420310|SON gene|son
Finding|Intellectual Product|SIMPLE_SEGMENT|15197,15200|false|false|false|C1947938|Law (document)|law
Finding|Idea or Concept|SIMPLE_SEGMENT|15205,15217|false|false|false|C1548597|Marketing basis - Transitional|Transitional
Event|Event|SIMPLE_SEGMENT|15218,15224|false|false|false|||issues
Finding|Functional Concept|SIMPLE_SEGMENT|15226,15231|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Anatomy|Tissue|SIMPLE_SEGMENT|15240,15247|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15240,15247|false|false|false|C0032226|Pleural Diseases|pleural
Event|Event|SIMPLE_SEGMENT|15248,15256|false|false|false|||catheter
Finding|Intellectual Product|SIMPLE_SEGMENT|15248,15256|false|false|false|C1546572||catheter
Event|Activity|SIMPLE_SEGMENT|15260,15265|false|false|false|C1882509|put - instruction imperative|place
Event|Event|SIMPLE_SEGMENT|15260,15265|false|false|false|||place
Finding|Functional Concept|SIMPLE_SEGMENT|15260,15265|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|SIMPLE_SEGMENT|15260,15265|false|false|false|C1533810||place
Event|Event|SIMPLE_SEGMENT|15269,15278|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|15269,15278|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|15269,15278|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|15269,15278|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|15269,15278|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|SIMPLE_SEGMENT|15290,15296|false|false|false|||follow
Event|Event|SIMPLE_SEGMENT|15305,15319|false|false|false|||interventional
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|15305,15319|false|false|false|C0184661;C2183254|Interventional procedure;interventional (invasive) radiology|interventional
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|15305,15319|false|false|false|C0184661;C2183254|Interventional procedure;interventional (invasive) radiology|interventional
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|15320,15329|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|15320,15329|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|15320,15329|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Event|Event|SIMPLE_SEGMENT|15336,15345|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|15336,15345|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|15336,15345|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|15336,15345|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|15336,15345|false|false|false|C0030685|Patient Discharge|discharge
Finding|Functional Concept|SIMPLE_SEGMENT|15347,15351|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|Tube
Finding|Gene or Genome|SIMPLE_SEGMENT|15347,15351|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|Tube
Event|Event|SIMPLE_SEGMENT|15360,15367|false|false|false|||removed
Event|Event|SIMPLE_SEGMENT|15373,15379|false|false|false|||output
Finding|Conceptual Entity|SIMPLE_SEGMENT|15373,15379|false|false|false|C1709366|system output|output
Procedure|Health Care Activity|SIMPLE_SEGMENT|15373,15379|false|false|false|C3251815|Measurement of fluid output|output
Finding|Idea or Concept|SIMPLE_SEGMENT|15394,15397|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|15394,15397|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|15405,15409|false|false|false|||need
Finding|Idea or Concept|SIMPLE_SEGMENT|15410,15417|false|false|false|C0549178|Continuous|ongoing
Event|Event|SIMPLE_SEGMENT|15418,15426|false|false|false|||diuresis
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|15418,15426|false|false|false|C0012797|Diuresis|diuresis
Finding|Gene or Genome|SIMPLE_SEGMENT|15433,15438|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Event|Event|SIMPLE_SEGMENT|15439,15445|false|false|false|||volume
Finding|Intellectual Product|SIMPLE_SEGMENT|15439,15445|false|false|false|C1705102|Volume (publication)|volume
Drug|Substance|SIMPLE_SEGMENT|15449,15455|false|false|false|C0302908|Liquid substance|fluids
Event|Event|SIMPLE_SEGMENT|15449,15455|false|false|false|||fluids
Finding|Body Substance|SIMPLE_SEGMENT|15449,15455|false|false|false|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|15449,15455|false|false|false|C0016286|Fluid Therapy|fluids
Event|Event|SIMPLE_SEGMENT|15461,15469|false|false|false|||received
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|15477,15480|false|false|false|C0228479|Structure of intraculminate fissure|ICU
Finding|Intellectual Product|SIMPLE_SEGMENT|15477,15480|false|false|false|C4554035|Inventory of Callous-Unemotional Traits|ICU
Event|Event|SIMPLE_SEGMENT|15486,15495|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|15486,15495|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|SIMPLE_SEGMENT|15501,15509|false|false|false|||responds
Event|Event|SIMPLE_SEGMENT|15510,15514|false|false|false|||well
Finding|Finding|SIMPLE_SEGMENT|15510,15514|false|false|false|C5575035|Well (answer to question)|well
Drug|Organic Chemical|SIMPLE_SEGMENT|15518,15523|false|false|false|C0699992|Lasix|Lasix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|15518,15523|false|false|false|C0699992|Lasix|Lasix
Event|Event|SIMPLE_SEGMENT|15518,15523|false|false|false|||Lasix
Finding|Idea or Concept|SIMPLE_SEGMENT|15534,15538|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|Goal
Finding|Intellectual Product|SIMPLE_SEGMENT|15534,15538|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|Goal
Event|Event|SIMPLE_SEGMENT|15543,15551|false|false|false|||negative
Finding|Classification|SIMPLE_SEGMENT|15543,15551|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|15543,15551|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|15543,15551|false|false|false|C5237010|Expression Negative|negative
Event|Event|SIMPLE_SEGMENT|15558,15567|false|false|false|||tolerates
Event|Event|SIMPLE_SEGMENT|15575,15583|false|false|false|||continue
Finding|Finding|SIMPLE_SEGMENT|15587,15591|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|SIMPLE_SEGMENT|15587,15591|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|SIMPLE_SEGMENT|15587,15591|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Event|Event|SIMPLE_SEGMENT|15592,15596|false|false|false|||dose
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|15600,15610|false|false|false|C0042313|vancomycin|vancomycin
Drug|Antibiotic|SIMPLE_SEGMENT|15600,15610|false|false|false|C0042313|vancomycin|vancomycin
Event|Event|SIMPLE_SEGMENT|15600,15610|false|false|false|||vancomycin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|15600,15610|false|false|false|C0489941|Vancomycin measurement|vancomycin
Event|Event|SIMPLE_SEGMENT|15642,15649|false|false|false|||stopped
Event|Event|SIMPLE_SEGMENT|15663,15671|false|false|false|||continue
Event|Event|SIMPLE_SEGMENT|15672,15676|false|false|false|||tube
Finding|Functional Concept|SIMPLE_SEGMENT|15672,15676|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|tube
Finding|Gene or Genome|SIMPLE_SEGMENT|15672,15676|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|tube
Event|Event|SIMPLE_SEGMENT|15716,15723|false|false|false|||benefit
Finding|Idea or Concept|SIMPLE_SEGMENT|15729,15736|false|false|false|C0549178|Continuous|ongoing
Finding|Finding|SIMPLE_SEGMENT|15737,15746|false|false|false|C0392209;C0518896;C1442959|Nutrition (function);Nutrition outcomes;Nutritional status|nutrition
Finding|Intellectual Product|SIMPLE_SEGMENT|15737,15746|false|false|false|C0392209;C0518896;C1442959|Nutrition (function);Nutrition outcomes;Nutritional status|nutrition
Finding|Organism Function|SIMPLE_SEGMENT|15737,15746|false|false|false|C0392209;C0518896;C1442959|Nutrition (function);Nutrition outcomes;Nutritional status|nutrition
Procedure|Research Activity|SIMPLE_SEGMENT|15737,15746|false|false|false|C0600072;C1521729|Feeding and dietary regimes;Nutritional Study|nutrition
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|15737,15746|false|false|false|C0600072;C1521729|Feeding and dietary regimes;Nutritional Study|nutrition
Event|Event|SIMPLE_SEGMENT|15747,15757|false|false|false|||evaluation
Finding|Idea or Concept|SIMPLE_SEGMENT|15747,15757|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|SIMPLE_SEGMENT|15747,15757|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Attribute|Clinical Attribute|SIMPLE_SEGMENT|15760,15771|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|15760,15771|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|15760,15771|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|15760,15771|false|false|false|C4284232|Medications|Medications
Finding|Finding|SIMPLE_SEGMENT|15760,15784|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|SIMPLE_SEGMENT|15775,15784|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|15775,15784|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Organic Chemical|SIMPLE_SEGMENT|15786,15797|false|false|false|C0082607|fluticasone|fluticasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|15786,15797|false|false|false|C0082607|fluticasone|fluticasone
Event|Event|SIMPLE_SEGMENT|15786,15797|false|false|false|||fluticasone
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|15811,15816|false|false|false|C0028429||nasal
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|15811,15816|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Organic Chemical|SIMPLE_SEGMENT|15811,15816|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|15811,15816|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Finding|Finding|SIMPLE_SEGMENT|15811,15816|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Functional Concept|SIMPLE_SEGMENT|15811,15816|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|15817,15823|false|false|false|C0233601|Spraying behavior|sprays
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|15817,15823|false|false|false|C1154182|Spray Dosage Form|sprays
Event|Event|SIMPLE_SEGMENT|15817,15823|false|false|false|||sprays
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|15824,15827|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|15824,15827|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|15824,15827|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|15824,15827|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|15824,15827|false|false|false|C1332410|BID gene|BID
Finding|Gene or Genome|SIMPLE_SEGMENT|15828,15831|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|15832,15841|false|false|false|C1717415||allergies
Event|Event|SIMPLE_SEGMENT|15832,15841|false|false|false|||allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|15832,15841|false|false|false|C0020517|Hypersensitivity|allergies
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|15842,15855|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Hormone|SIMPLE_SEGMENT|15842,15855|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Organic Chemical|SIMPLE_SEGMENT|15842,15855|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|15842,15855|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Event|Event|SIMPLE_SEGMENT|15842,15855|false|false|false|||levothyroxine
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|15869,15879|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|15869,15879|false|false|false|C0065374|lisinopril|lisinopril
Event|Event|SIMPLE_SEGMENT|15869,15879|false|false|false|||lisinopril
Drug|Inorganic Chemical|SIMPLE_SEGMENT|15902,15909|false|false|false|C0006222|Bromides|bromide
Event|Event|SIMPLE_SEGMENT|15902,15909|false|false|false|||bromide
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|15902,15909|false|false|false|C0202341|Bromides measurement|bromide
Drug|Biologically Active Substance|SIMPLE_SEGMENT|15923,15930|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|15923,15930|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|15923,15930|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|15923,15930|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|15923,15930|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|SIMPLE_SEGMENT|15923,15930|false|false|false|||Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|15923,15930|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|15923,15930|false|false|false|C0201925|Calcium measurement|Calcium
Drug|Organic Chemical|SIMPLE_SEGMENT|15931,15943|false|false|false|C0301532|Multivitamin preparation|multivitamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|15931,15943|false|false|false|C0301532|Multivitamin preparation|multivitamin
Drug|Vitamin|SIMPLE_SEGMENT|15931,15943|false|false|false|C0301532|Multivitamin preparation|multivitamin
Event|Event|SIMPLE_SEGMENT|15931,15943|false|false|false|||multivitamin
Drug|Organic Chemical|SIMPLE_SEGMENT|15944,15954|false|false|false|C0028978|omeprazole|omeprazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|15944,15954|false|false|false|C0028978|omeprazole|omeprazole
Event|Event|SIMPLE_SEGMENT|15944,15954|false|false|false|||omeprazole
Drug|Organic Chemical|SIMPLE_SEGMENT|15967,15980|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|15967,15980|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Event|Event|SIMPLE_SEGMENT|15967,15980|false|false|false|||acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|15967,15980|false|false|false|C0373527|Acetaminophen measurement|acetaminophen
Finding|Gene or Genome|SIMPLE_SEGMENT|15981,15984|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|15985,15989|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|15985,15989|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|15985,15989|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|15985,15989|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|15993,16002|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|15993,16002|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|15993,16002|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|15993,16002|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|15993,16002|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|15993,16014|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|16003,16014|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|16003,16014|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|16003,16014|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|16003,16014|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|SIMPLE_SEGMENT|16019,16030|false|false|false|C0082607|fluticasone|fluticasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|16019,16030|false|false|false|C0082607|fluticasone|fluticasone
Event|Event|SIMPLE_SEGMENT|16019,16030|false|false|false|||fluticasone
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|16048,16053|false|false|false|C1154182|Spray Dosage Form|Spray
Event|Activity|SIMPLE_SEGMENT|16048,16053|false|false|false|C2003858|Spray (action)|Spray
Event|Event|SIMPLE_SEGMENT|16048,16053|false|false|false|||Spray
Finding|Functional Concept|SIMPLE_SEGMENT|16048,16053|false|false|false|C4521772|Spray (administration method)|Spray
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|16048,16065|false|false|false|C1710170|SPRAY, SUSPENSION|Spray, Suspension
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|16055,16065|false|false|false|C0038960;C1382107|Suspension substance;Suspensions|Suspension
Drug|Substance|SIMPLE_SEGMENT|16055,16065|false|false|false|C0038960;C1382107|Suspension substance;Suspensions|Suspension
Event|Event|SIMPLE_SEGMENT|16055,16065|false|false|false|||Suspension
Finding|Functional Concept|SIMPLE_SEGMENT|16055,16065|false|false|false|C1705537|Suspension (action)|Suspension
Event|Event|SIMPLE_SEGMENT|16075,16080|false|false|false|||puffs
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|16082,16087|false|false|false|C0028429||Nasal
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|16082,16087|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Organic Chemical|SIMPLE_SEGMENT|16082,16087|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|16082,16087|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Finding|Finding|SIMPLE_SEGMENT|16082,16087|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Finding|Functional Concept|SIMPLE_SEGMENT|16082,16087|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Finding|Idea or Concept|SIMPLE_SEGMENT|16096,16099|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|16096,16099|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|16103,16109|false|false|false|||needed
Attribute|Clinical Attribute|SIMPLE_SEGMENT|16114,16123|false|false|false|C1717415||allergies
Event|Event|SIMPLE_SEGMENT|16114,16123|false|false|false|||allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|16114,16123|false|false|false|C0020517|Hypersensitivity|allergies
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|16130,16143|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Hormone|SIMPLE_SEGMENT|16130,16143|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Organic Chemical|SIMPLE_SEGMENT|16130,16143|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|16130,16143|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Event|Event|SIMPLE_SEGMENT|16130,16143|false|false|false|||levothyroxine
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|16151,16157|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|16151,16157|false|false|false|||Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|16171,16177|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|16171,16177|false|false|false|||Tablet
Drug|Organic Chemical|SIMPLE_SEGMENT|16202,16215|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|16202,16215|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Event|Event|SIMPLE_SEGMENT|16202,16215|false|false|false|||acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|16202,16215|false|false|false|C0373527|Acetaminophen measurement|acetaminophen
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|16223,16229|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|16239,16246|false|false|false|C0039225|Tablet Dosage Form|Tablets
Event|Event|SIMPLE_SEGMENT|16239,16246|false|false|false|||Tablets
Event|Event|SIMPLE_SEGMENT|16275,16281|false|false|false|||needed
Attribute|Clinical Attribute|SIMPLE_SEGMENT|16286,16290|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|16286,16290|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|16286,16290|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|16286,16290|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|16297,16306|false|false|false|C0032629|Polyvinyls|polyvinyl
Drug|Organic Chemical|SIMPLE_SEGMENT|16297,16306|false|false|false|C0032629|Polyvinyls|polyvinyl
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|16297,16314|false|false|false|C0032623|polyvinyl alcohol|polyvinyl alcohol
Drug|Organic Chemical|SIMPLE_SEGMENT|16307,16314|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|16307,16314|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Event|Event|SIMPLE_SEGMENT|16307,16314|false|false|false|||alcohol
Finding|Intellectual Product|SIMPLE_SEGMENT|16307,16314|false|false|false|C1547288|Alcohol - Recreational Drug Use Code|alcohol
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|16321,16326|false|false|false|C0991568|Drops - Drug Form|Drops
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|16340,16344|false|false|false|C0991568|Drops - Drug Form|drop
Event|Activity|SIMPLE_SEGMENT|16340,16344|false|false|false|C1705648|Dropping|drop
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|16345,16355|false|false|false|C0015392|Eye|Ophthalmic
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|16345,16355|false|false|false|C2347396|Ophthalmic Dosage Form|Ophthalmic
Event|Event|SIMPLE_SEGMENT|16345,16355|false|false|false|||Ophthalmic
Finding|Functional Concept|SIMPLE_SEGMENT|16345,16355|false|false|false|C1522230|Ophthalmic Route of Administration|Ophthalmic
Event|Event|SIMPLE_SEGMENT|16381,16387|false|false|false|||needed
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|16392,16400|false|false|false|C0013238;C0022575|Dry Eye Syndromes;Keratoconjunctivitis Sicca|dry eyes
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|16392,16400|false|false|false|C0720056|Dry Eyes brand of ocular lubricant|dry eyes
Finding|Sign or Symptom|SIMPLE_SEGMENT|16392,16400|false|false|false|C0314719|Dryness of eye|dry eyes
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|16396,16400|false|false|false|C0015392|Eye|eyes
Attribute|Clinical Attribute|SIMPLE_SEGMENT|16396,16400|false|false|false|C5848506||eyes
Event|Event|SIMPLE_SEGMENT|16396,16400|false|false|false|||eyes
Drug|Biologically Active Substance|SIMPLE_SEGMENT|16407,16414|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Organic Chemical|SIMPLE_SEGMENT|16407,16414|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|16407,16414|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Event|Event|SIMPLE_SEGMENT|16407,16414|false|false|false|||heparin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|16407,16423|false|false|false|C0770546|heparin, porcine|heparin, porcine
Drug|Organic Chemical|SIMPLE_SEGMENT|16407,16423|false|false|false|C0770546|heparin, porcine|heparin, porcine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|16407,16423|false|false|false|C0770546|heparin, porcine|heparin, porcine
Event|Event|SIMPLE_SEGMENT|16416,16423|false|false|false|||porcine
Finding|Finding|SIMPLE_SEGMENT|16416,16423|false|false|false|C4554819|Porcine prosthetic valve|porcine
Event|Event|SIMPLE_SEGMENT|16448,16451|false|false|false|||Sig
Finding|Functional Concept|SIMPLE_SEGMENT|16465,16476|false|false|false|C1522726|Intravenous Route of Administration|Intravenous
Event|Event|SIMPLE_SEGMENT|16477,16480|false|false|false|||PRN
Finding|Gene or Genome|SIMPLE_SEGMENT|16477,16480|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|SIMPLE_SEGMENT|16485,16491|false|false|false|||needed
Event|Event|SIMPLE_SEGMENT|16496,16502|false|false|false|||needed
Drug|Biologically Active Substance|SIMPLE_SEGMENT|16507,16511|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|16507,16511|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Substance|SIMPLE_SEGMENT|16507,16511|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Finding|Intellectual Product|SIMPLE_SEGMENT|16507,16511|false|false|false|C1546701|line source specimen code|line
Attribute|Clinical Attribute|SIMPLE_SEGMENT|16507,16517|false|false|false|C4036660||line flush
Event|Event|SIMPLE_SEGMENT|16512,16517|false|false|false|||flush
Finding|Functional Concept|SIMPLE_SEGMENT|16512,16517|false|false|false|C0016382;C1696091|Flush - RouteOfAdministration;Flushing|flush
Finding|Sign or Symptom|SIMPLE_SEGMENT|16512,16517|false|false|false|C0016382;C1696091|Flush - RouteOfAdministration;Flushing|flush
Drug|Biologically Active Substance|SIMPLE_SEGMENT|16524,16531|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Organic Chemical|SIMPLE_SEGMENT|16524,16531|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|16524,16531|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Event|Event|SIMPLE_SEGMENT|16524,16531|false|false|false|||heparin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|16524,16541|false|false|false|C0770546|heparin, porcine|heparin (porcine)
Drug|Organic Chemical|SIMPLE_SEGMENT|16524,16541|false|false|false|C0770546|heparin, porcine|heparin (porcine)
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|16524,16541|false|false|false|C0770546|heparin, porcine|heparin (porcine)
Event|Event|SIMPLE_SEGMENT|16533,16540|false|false|false|||porcine
Finding|Finding|SIMPLE_SEGMENT|16533,16540|false|false|false|C4554819|Porcine prosthetic valve|porcine
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|16556,16564|false|false|false|C0037633;C0525069;C1382100|Pharmaceutical Solutions;Solution Dosage Form;Solutions|Solution
Drug|Substance|SIMPLE_SEGMENT|16556,16564|false|false|false|C0037633;C0525069;C1382100|Pharmaceutical Solutions;Solution Dosage Form;Solutions|Solution
Event|Event|SIMPLE_SEGMENT|16556,16564|false|false|false|||Solution
Finding|Conceptual Entity|SIMPLE_SEGMENT|16556,16564|false|false|false|C2699488|Resolution|Solution
Event|Event|SIMPLE_SEGMENT|16565,16568|false|false|false|||Sig
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|16589,16598|false|false|false|C1272883|Injection|Injection
Event|Event|SIMPLE_SEGMENT|16589,16598|false|false|false|||Injection
Finding|Functional Concept|SIMPLE_SEGMENT|16589,16598|false|false|false|C1828121|Injection Route of Administration|Injection
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|16589,16598|false|false|false|C0021485;C1533685|Injection of therapeutic agent;Injection procedure|Injection
Finding|Idea or Concept|SIMPLE_SEGMENT|16607,16610|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|16607,16610|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|16617,16624|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|SIMPLE_SEGMENT|16617,16624|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|16617,16624|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|SIMPLE_SEGMENT|16617,16624|false|false|false|||insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|16617,16624|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|16617,16624|false|false|false|C0202098|Insulin measurement|insulin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|16617,16631|false|false|false|C0293359|insulin lispro|insulin lispro
Drug|Hormone|SIMPLE_SEGMENT|16617,16631|false|false|false|C0293359|insulin lispro|insulin lispro
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|16617,16631|false|false|false|C0293359|insulin lispro|insulin lispro
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|16625,16631|false|false|false|C0293359|insulin lispro|lispro
Drug|Hormone|SIMPLE_SEGMENT|16625,16631|false|false|false|C0293359|insulin lispro|lispro
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|16625,16631|false|false|false|C0293359|insulin lispro|lispro
Event|Event|SIMPLE_SEGMENT|16625,16631|false|false|false|||lispro
Event|Event|SIMPLE_SEGMENT|16636,16640|false|false|false|||unit
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|16644,16652|false|false|false|C0037633;C0525069;C1382100|Pharmaceutical Solutions;Solution Dosage Form;Solutions|Solution
Drug|Substance|SIMPLE_SEGMENT|16644,16652|false|false|false|C0037633;C0525069;C1382100|Pharmaceutical Solutions;Solution Dosage Form;Solutions|Solution
Event|Event|SIMPLE_SEGMENT|16644,16652|false|false|false|||Solution
Finding|Conceptual Entity|SIMPLE_SEGMENT|16644,16652|false|false|false|C2699488|Resolution|Solution
Event|Event|SIMPLE_SEGMENT|16658,16665|false|false|false|||sliding
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|16666,16671|false|false|false|C0222045|Integumentary scale|scale
Event|Activity|SIMPLE_SEGMENT|16666,16671|false|false|false|C1947916|Scaling|scale
Finding|Conceptual Entity|SIMPLE_SEGMENT|16666,16671|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|scale
Finding|Intellectual Product|SIMPLE_SEGMENT|16666,16671|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|scale
Event|Event|SIMPLE_SEGMENT|16672,16677|false|false|false|||units
Finding|Functional Concept|SIMPLE_SEGMENT|16679,16691|false|false|false|C1522438|Subcutaneous Route of Administration|Subcutaneous
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|16698,16703|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|SIMPLE_SEGMENT|16706,16709|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|16706,16709|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Functional Concept|SIMPLE_SEGMENT|16711,16718|false|false|false|C0332246|Sliding|Sliding
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|16711,16724|false|false|false|C2937251|sliding scale|Sliding scale
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|16719,16724|false|false|false|C0222045|Integumentary scale|scale
Event|Activity|SIMPLE_SEGMENT|16719,16724|false|false|false|C1947916|Scaling|scale
Finding|Conceptual Entity|SIMPLE_SEGMENT|16719,16724|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|scale
Finding|Intellectual Product|SIMPLE_SEGMENT|16719,16724|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|scale
Event|Event|SIMPLE_SEGMENT|16847,16851|false|false|false|||call
Finding|Functional Concept|SIMPLE_SEGMENT|16847,16851|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|call
Finding|Gene or Genome|SIMPLE_SEGMENT|16847,16851|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|call
Finding|Intellectual Product|SIMPLE_SEGMENT|16847,16851|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|call
Finding|Mental Process|SIMPLE_SEGMENT|16847,16851|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|call
Drug|Organic Chemical|SIMPLE_SEGMENT|16861,16871|false|false|false|C0025942|miconazole|miconazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|16861,16871|false|false|false|C0025942|miconazole|miconazole
Event|Event|SIMPLE_SEGMENT|16861,16871|false|false|false|||miconazole
Drug|Organic Chemical|SIMPLE_SEGMENT|16861,16879|false|false|false|C0086620|miconazole nitrate|miconazole nitrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|16861,16879|false|false|false|C0086620|miconazole nitrate|miconazole nitrate
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|16872,16879|false|false|false|C0028125;C0699857;C3848573|Nitrate;Nitrates;nitrate ion|nitrate
Drug|Inorganic Chemical|SIMPLE_SEGMENT|16872,16879|false|false|false|C0028125;C0699857;C3848573|Nitrate;Nitrates;nitrate ion|nitrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|16872,16879|false|false|false|C0028125;C0699857;C3848573|Nitrate;Nitrates;nitrate ion|nitrate
Event|Event|SIMPLE_SEGMENT|16872,16879|false|false|false|||nitrate
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|16884,16890|false|false|false|C0032861;C1382110|Powder dose form;powder physical state|Powder
Drug|Substance|SIMPLE_SEGMENT|16884,16890|false|false|false|C0032861;C1382110|Powder dose form;powder physical state|Powder
Finding|Gene or Genome|SIMPLE_SEGMENT|16904,16908|false|false|false|C1858559|APPL1 gene|Appl
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|16909,16916|false|false|false|C1710439|Topical Dosage Form|Topical
Finding|Functional Concept|SIMPLE_SEGMENT|16909,16916|false|false|false|C1522168|Topical Route of Administration|Topical
Event|Event|SIMPLE_SEGMENT|16917,16920|false|false|false|||TID
Finding|Finding|SIMPLE_SEGMENT|16923,16930|false|false|false|C4035626|3 times|3 times
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|16925,16930|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Event|Event|SIMPLE_SEGMENT|16925,16930|false|false|false|||times
Finding|Idea or Concept|SIMPLE_SEGMENT|16933,16936|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|16933,16936|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|16941,16947|false|false|false|||needed
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|16952,16956|false|false|false|C5779629|Eruption of skin (disorder)|rash
Event|Event|SIMPLE_SEGMENT|16952,16956|false|false|false|||rash
Finding|Pathologic Function|SIMPLE_SEGMENT|16952,16956|false|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Sign or Symptom|SIMPLE_SEGMENT|16952,16956|false|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Drug|Organic Chemical|SIMPLE_SEGMENT|16963,16974|false|false|false|C0061851|ondansetron|ondansetron
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|16963,16974|false|false|false|C0061851|ondansetron|ondansetron
Event|Event|SIMPLE_SEGMENT|16963,16974|false|false|false|||ondansetron
Drug|Organic Chemical|SIMPLE_SEGMENT|16963,16978|false|false|false|C0700478|ondansetron hydrochloride|ondansetron HCl
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|16963,16978|false|false|false|C0700478|ondansetron hydrochloride|ondansetron HCl
Disorder|Neoplastic Process|SIMPLE_SEGMENT|16975,16978|false|false|false|C0023443|Hairy Cell Leukemia|HCl
Drug|Immunologic Factor|SIMPLE_SEGMENT|16975,16978|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Inorganic Chemical|SIMPLE_SEGMENT|16975,16978|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|16975,16978|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Event|Event|SIMPLE_SEGMENT|16975,16978|false|false|false|||HCl
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|16987,16995|false|false|false|C0037633;C0525069;C1382100|Pharmaceutical Solutions;Solution Dosage Form;Solutions|Solution
Drug|Substance|SIMPLE_SEGMENT|16987,16995|false|false|false|C0037633;C0525069;C1382100|Pharmaceutical Solutions;Solution Dosage Form;Solutions|Solution
Event|Event|SIMPLE_SEGMENT|16987,16995|false|false|false|||Solution
Finding|Conceptual Entity|SIMPLE_SEGMENT|16987,16995|false|false|false|C2699488|Resolution|Solution
Event|Event|SIMPLE_SEGMENT|17013,17024|false|false|false|||Intravenous
Finding|Functional Concept|SIMPLE_SEGMENT|17013,17024|false|false|false|C1522726|Intravenous Route of Administration|Intravenous
Event|Event|SIMPLE_SEGMENT|17051,17057|false|false|false|||needed
Attribute|Clinical Attribute|SIMPLE_SEGMENT|17062,17068|false|false|false|C4255480||nausea
Event|Event|SIMPLE_SEGMENT|17062,17068|false|false|false|||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|17062,17068|false|false|false|C0027497|Nausea|nausea
Drug|Organic Chemical|SIMPLE_SEGMENT|17076,17086|false|false|false|C0171023|olanzapine|olanzapine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|17076,17086|false|false|false|C0171023|olanzapine|olanzapine
Event|Event|SIMPLE_SEGMENT|17076,17086|false|false|false|||olanzapine
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|17094,17100|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|17114,17120|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|17114,17120|false|false|false|||Tablet
Event|Event|SIMPLE_SEGMENT|17144,17150|false|false|false|||needed
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|17155,17162|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Event|Event|SIMPLE_SEGMENT|17155,17162|false|false|false|||anxiety
Finding|Sign or Symptom|SIMPLE_SEGMENT|17155,17162|false|false|false|C0860603|Anxiety symptoms|anxiety
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|17163,17171|false|false|false|C1950154|Insomnia homeopathic medication|insomnia
Event|Event|SIMPLE_SEGMENT|17163,17171|false|false|false|||insomnia
Finding|Sign or Symptom|SIMPLE_SEGMENT|17163,17171|false|false|false|C0917801|Sleeplessness|insomnia
Drug|Organic Chemical|SIMPLE_SEGMENT|17179,17189|false|false|false|C0171023|olanzapine|olanzapine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|17179,17189|false|false|false|C0171023|olanzapine|olanzapine
Event|Event|SIMPLE_SEGMENT|17179,17189|false|false|false|||olanzapine
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|17197,17203|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|17217,17223|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|17217,17223|false|false|false|||Tablet
Event|Event|SIMPLE_SEGMENT|17245,17251|false|false|false|||needed
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|17256,17263|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Event|Event|SIMPLE_SEGMENT|17256,17263|false|false|false|||anxiety
Finding|Sign or Symptom|SIMPLE_SEGMENT|17256,17263|false|false|false|C0860603|Anxiety symptoms|anxiety
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|17271,17281|false|false|false|C0042313|vancomycin|vancomycin
Drug|Antibiotic|SIMPLE_SEGMENT|17271,17281|false|false|false|C0042313|vancomycin|vancomycin
Event|Event|SIMPLE_SEGMENT|17271,17281|false|false|false|||vancomycin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|17271,17281|false|false|false|C0489941|Vancomycin measurement|vancomycin
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|17289,17296|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|SIMPLE_SEGMENT|17289,17296|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|17289,17296|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|17310,17317|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|SIMPLE_SEGMENT|17310,17317|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|17310,17317|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Finding|Intellectual Product|SIMPLE_SEGMENT|17326,17331|false|false|false|C1720374|Every - dosing instruction fragment|every
Event|Event|SIMPLE_SEGMENT|17355,17363|false|false|false|||Continue
Event|Event|SIMPLE_SEGMENT|17382,17391|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|17382,17391|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|17382,17391|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|17382,17391|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|17382,17391|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|17382,17403|false|false|false|C4019243||Discharge Disposition
Finding|Finding|SIMPLE_SEGMENT|17382,17403|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|17392,17403|false|false|false|C2926604||Disposition
Event|Event|SIMPLE_SEGMENT|17392,17403|false|false|false|||Disposition
Procedure|Health Care Activity|SIMPLE_SEGMENT|17392,17403|false|false|false|C0184758|Patient disposition|Disposition
Finding|Finding|SIMPLE_SEGMENT|17405,17413|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|SIMPLE_SEGMENT|17405,17413|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Procedure|Health Care Activity|SIMPLE_SEGMENT|17405,17418|false|false|false|C0023977|long-term care|Extended Care
Event|Activity|SIMPLE_SEGMENT|17414,17418|false|false|false|C1947933|care activity|Care
Event|Event|SIMPLE_SEGMENT|17414,17418|false|false|false|||Care
Finding|Finding|SIMPLE_SEGMENT|17414,17418|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|SIMPLE_SEGMENT|17414,17418|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Event|Event|SIMPLE_SEGMENT|17421,17429|false|false|false|||Facility
Finding|Intellectual Product|SIMPLE_SEGMENT|17421,17429|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|SIMPLE_SEGMENT|17437,17446|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|17437,17446|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|17437,17446|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|17437,17446|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|17437,17446|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|17437,17456|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|17447,17456|false|false|false|C0945731||Diagnosis
Event|Event|SIMPLE_SEGMENT|17447,17456|false|false|false|||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|17447,17456|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|17447,17456|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|17447,17456|false|false|false|C0011900|Diagnosis|Diagnosis
Event|Event|SIMPLE_SEGMENT|17466,17475|false|false|false|||diagnoses
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|17466,17475|false|false|false|C0011900|Diagnosis|diagnoses
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|17477,17506|false|false|false|C0238106|Clostridium difficile colitis|Clostridium difficile colitis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|17499,17506|false|false|false|C0009319|Colitis|colitis
Event|Event|SIMPLE_SEGMENT|17499,17506|false|false|false|||colitis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|17511,17517|false|false|false|C0036690;C0243026|Sepsis;Septicemia|sepsis
Event|Event|SIMPLE_SEGMENT|17511,17517|false|false|false|||sepsis
Anatomy|Tissue|SIMPLE_SEGMENT|17518,17525|false|false|false|C0032225|Pleura|Pleural
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|17518,17525|false|false|false|C0032226|Pleural Diseases|Pleural
Finding|Body Substance|SIMPLE_SEGMENT|17518,17534|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|Pleural effusion
Finding|Finding|SIMPLE_SEGMENT|17518,17534|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|Pleural effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|17518,17534|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|Pleural effusion
Event|Event|SIMPLE_SEGMENT|17526,17534|false|false|false|||effusion
Finding|Body Substance|SIMPLE_SEGMENT|17526,17534|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|SIMPLE_SEGMENT|17526,17534|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|17526,17534|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Event|Event|SIMPLE_SEGMENT|17548,17556|false|false|false|||catheter
Finding|Intellectual Product|SIMPLE_SEGMENT|17548,17556|false|false|false|C1546572||catheter
Event|Event|SIMPLE_SEGMENT|17557,17563|false|false|false|||placed
Event|Event|SIMPLE_SEGMENT|17567,17576|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|17567,17576|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|17567,17576|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|17567,17576|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|17567,17576|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|17577,17586|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|17577,17586|false|false|false|C0012634|Disease|Condition
Event|Event|SIMPLE_SEGMENT|17577,17586|false|false|false|||Condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|17577,17586|false|false|false|C1705253|Logical Condition|Condition
Finding|Mental Process|SIMPLE_SEGMENT|17588,17594|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|17588,17601|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|SIMPLE_SEGMENT|17588,17601|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|17595,17601|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|17595,17601|false|false|false|C1546481|What subject filter - Status|Status
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|17603,17611|false|false|false|C0009676|Confusion|Confused
Event|Event|SIMPLE_SEGMENT|17603,17611|false|false|false|||Confused
Finding|Finding|SIMPLE_SEGMENT|17603,17611|false|false|false|C0683369;C1547301|Clouded consciousness;Precaution Code - Confused|Confused
Finding|Intellectual Product|SIMPLE_SEGMENT|17603,17611|false|false|false|C0683369;C1547301|Clouded consciousness;Precaution Code - Confused|Confused
Event|Event|SIMPLE_SEGMENT|17625,17630|false|false|false|||Level
Attribute|Clinical Attribute|SIMPLE_SEGMENT|17625,17647|false|false|false|C4050479||Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|17625,17647|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|SIMPLE_SEGMENT|17634,17647|false|false|false|||Consciousness
Finding|Finding|SIMPLE_SEGMENT|17634,17647|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|SIMPLE_SEGMENT|17634,17647|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Event|Event|SIMPLE_SEGMENT|17649,17658|false|false|false|||Lethargic
Finding|Sign or Symptom|SIMPLE_SEGMENT|17649,17658|false|false|false|C0023380|Lethargy|Lethargic
Event|Event|SIMPLE_SEGMENT|17663,17672|false|false|false|||arousable
Event|Activity|SIMPLE_SEGMENT|17674,17682|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|17674,17682|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|SIMPLE_SEGMENT|17674,17682|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|SIMPLE_SEGMENT|17683,17689|false|false|false|C5889824||Status
Event|Event|SIMPLE_SEGMENT|17683,17689|false|false|false|||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|17683,17689|false|false|false|C1546481|What subject filter - Status|Status
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|17698,17701|false|false|false|C3159311|BORNHOLM EYE DISEASE|Bed
Event|Event|SIMPLE_SEGMENT|17698,17701|false|false|false|||Bed
Finding|Intellectual Product|SIMPLE_SEGMENT|17698,17701|false|false|false|C2346952|Bachelor of Education|Bed
Event|Event|SIMPLE_SEGMENT|17707,17717|false|false|false|||assistance
Finding|Social Behavior|SIMPLE_SEGMENT|17707,17717|false|false|false|C0018896|Helping Behavior|assistance
Event|Event|SIMPLE_SEGMENT|17731,17741|false|false|false|||wheelchair
Finding|Finding|SIMPLE_SEGMENT|17731,17741|false|false|false|C2135586;C4321408|Wheelchair Usually Used;has wheelchair at home (history)|wheelchair
Event|Event|SIMPLE_SEGMENT|17746,17755|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|17746,17755|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|17746,17755|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|17746,17755|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|17746,17755|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|17746,17768|false|false|false|C3669312||Discharge Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|17746,17768|false|false|false|C4282220|Discharge instructions|Discharge Instructions
Procedure|Health Care Activity|SIMPLE_SEGMENT|17746,17768|false|false|false|C2266673|hospital discharge instructions (treatment)|Discharge Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|17756,17768|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|17756,17768|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|17756,17768|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Finding|Gene or Genome|SIMPLE_SEGMENT|17770,17774|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Event|Event|SIMPLE_SEGMENT|17794,17802|false|false|false|||pleasure
Finding|Intellectual Product|SIMPLE_SEGMENT|17794,17802|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|SIMPLE_SEGMENT|17794,17802|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|SIMPLE_SEGMENT|17810,17814|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|17810,17814|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|17810,17814|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|17810,17814|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|17810,17817|false|false|false|C1555558|care of - AddressPartType|care of
Event|Event|SIMPLE_SEGMENT|17834,17843|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|17834,17843|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Anatomy|Body Location or Region|SIMPLE_SEGMENT|17856,17865|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|SIMPLE_SEGMENT|17856,17870|false|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|17866,17870|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|17866,17870|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|17866,17870|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|17866,17870|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|17882,17887|false|false|false|||found
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|17899,17908|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|SIMPLE_SEGMENT|17899,17908|false|false|false|||infection
Finding|Pathologic Function|SIMPLE_SEGMENT|17899,17908|false|false|false|C3714514|Infection|infection
Event|Event|SIMPLE_SEGMENT|17910,17916|false|false|false|||called
Event|Event|SIMPLE_SEGMENT|17936,17943|false|false|false|||treated
Drug|Antibiotic|SIMPLE_SEGMENT|17949,17960|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|SIMPLE_SEGMENT|17949,17960|false|false|false|||antibiotics
Event|Event|SIMPLE_SEGMENT|17977,17985|false|false|false|||continue
Event|Event|SIMPLE_SEGMENT|17992,18001|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|17992,18001|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|17992,18001|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|17992,18001|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|17992,18001|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|SIMPLE_SEGMENT|18017,18026|false|false|false|||shortness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|18017,18036|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|SIMPLE_SEGMENT|18017,18036|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|SIMPLE_SEGMENT|18030,18036|false|false|false|C0225386|Breath|breath
Event|Event|SIMPLE_SEGMENT|18047,18052|false|false|false|||found
Finding|Gene or Genome|SIMPLE_SEGMENT|18063,18068|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Event|Event|SIMPLE_SEGMENT|18069,18079|false|false|false|||collection
Finding|Conceptual Entity|SIMPLE_SEGMENT|18069,18079|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|SIMPLE_SEGMENT|18069,18079|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|SIMPLE_SEGMENT|18069,18079|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|SIMPLE_SEGMENT|18069,18079|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Drug|Substance|SIMPLE_SEGMENT|18083,18088|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|18083,18088|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|18083,18088|false|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Functional Concept|SIMPLE_SEGMENT|18102,18107|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|18102,18112|false|false|false|C0225706|Right lung|right lung
Anatomy|Body Location or Region|SIMPLE_SEGMENT|18108,18112|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|18108,18112|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|18108,18112|false|false|false|C0024115|Lung diseases|lung
Event|Event|SIMPLE_SEGMENT|18108,18112|false|false|false|||lung
Finding|Finding|SIMPLE_SEGMENT|18108,18112|false|false|false|C0740941|Lung Problem|lung
Event|Event|SIMPLE_SEGMENT|18119,18127|false|false|false|||catheter
Finding|Intellectual Product|SIMPLE_SEGMENT|18119,18127|false|false|false|C1546572||catheter
Event|Event|SIMPLE_SEGMENT|18132,18138|false|false|false|||placed
Event|Event|SIMPLE_SEGMENT|18142,18147|false|false|false|||drain
Drug|Substance|SIMPLE_SEGMENT|18153,18158|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|18153,18158|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|18153,18158|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|18167,18175|false|false|false|||catheter
Finding|Intellectual Product|SIMPLE_SEGMENT|18167,18175|false|false|false|C1546572||catheter
Event|Event|SIMPLE_SEGMENT|18181,18187|false|false|false|||remain
Event|Activity|SIMPLE_SEGMENT|18191,18196|false|false|false|C1882509|put - instruction imperative|place
Event|Event|SIMPLE_SEGMENT|18191,18196|false|false|false|||place
Finding|Functional Concept|SIMPLE_SEGMENT|18191,18196|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|SIMPLE_SEGMENT|18191,18196|false|false|false|C1533810||place
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|18212,18217|false|false|false|C0034991|Rehabilitation therapy|rehab
Event|Event|SIMPLE_SEGMENT|18232,18238|false|false|false|||follow
Anatomy|Body Location or Region|SIMPLE_SEGMENT|18251,18255|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|18251,18255|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|18251,18255|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|SIMPLE_SEGMENT|18251,18255|false|false|false|C0740941|Lung Problem|lung
Event|Event|SIMPLE_SEGMENT|18256,18263|false|false|false|||doctors
Event|Event|SIMPLE_SEGMENT|18290,18297|false|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|18290,18297|false|false|false|C0392747|Changing|changes
Event|Event|SIMPLE_SEGMENT|18308,18312|false|false|false|||made
Attribute|Clinical Attribute|SIMPLE_SEGMENT|18321,18332|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|18321,18332|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|18321,18332|false|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|18321,18332|false|false|false|C4284232|Medications|medications
Drug|Inorganic Chemical|SIMPLE_SEGMENT|18334,18338|false|false|false|C0723457|Stop brand of fluoride|STOP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|18334,18338|false|false|false|C0723457|Stop brand of fluoride|STOP
Event|Activity|SIMPLE_SEGMENT|18334,18338|false|false|false|C1947925|Stop (Instruction Imperative)|STOP
Event|Event|SIMPLE_SEGMENT|18334,18338|false|false|false|||STOP
Finding|Gene or Genome|SIMPLE_SEGMENT|18334,18338|false|false|false|C1417022|MAP6 gene|STOP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|18339,18349|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|18339,18349|false|false|false|C0065374|lisinopril|lisinopril
Event|Event|SIMPLE_SEGMENT|18339,18349|false|false|false|||lisinopril
Drug|Inorganic Chemical|SIMPLE_SEGMENT|18350,18354|false|false|false|C0723457|Stop brand of fluoride|STOP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|18350,18354|false|false|false|C0723457|Stop brand of fluoride|STOP
Event|Activity|SIMPLE_SEGMENT|18350,18354|false|false|false|C1947925|Stop (Instruction Imperative)|STOP
Event|Event|SIMPLE_SEGMENT|18350,18354|false|false|false|||STOP
Finding|Gene or Genome|SIMPLE_SEGMENT|18350,18354|false|false|false|C1417022|MAP6 gene|STOP
Drug|Organic Chemical|SIMPLE_SEGMENT|18355,18365|false|false|false|C0028978|omeprazole|omeprazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|18355,18365|false|false|false|C0028978|omeprazole|omeprazole
Event|Event|SIMPLE_SEGMENT|18355,18365|false|false|false|||omeprazole
Drug|Inorganic Chemical|SIMPLE_SEGMENT|18366,18370|false|false|false|C0723457|Stop brand of fluoride|STOP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|18366,18370|false|false|false|C0723457|Stop brand of fluoride|STOP
Event|Activity|SIMPLE_SEGMENT|18366,18370|false|false|false|C1947925|Stop (Instruction Imperative)|STOP
Event|Event|SIMPLE_SEGMENT|18366,18370|false|false|false|||STOP
Finding|Gene or Genome|SIMPLE_SEGMENT|18366,18370|false|false|false|C1417022|MAP6 gene|STOP
Drug|Organic Chemical|SIMPLE_SEGMENT|18371,18381|false|false|false|C0213771|tiotropium|tiotropium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|18371,18381|false|false|false|C0213771|tiotropium|tiotropium
Event|Event|SIMPLE_SEGMENT|18371,18381|false|false|false|||tiotropium
Drug|Food|SIMPLE_SEGMENT|18382,18387|false|false|false|C0452588|Start brand of breakfast cereal|START
Event|Event|SIMPLE_SEGMENT|18382,18387|false|false|false|||START
Finding|Intellectual Product|SIMPLE_SEGMENT|18382,18387|false|false|false|C1552850|start - HtmlLinkType|START
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|18382,18387|false|false|false|C5447432|Collagen Tile Brachytherapy|START
Drug|Organic Chemical|SIMPLE_SEGMENT|18388,18394|false|false|false|C0206046|Zofran|Zofran
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|18388,18394|false|false|false|C0206046|Zofran|Zofran
Drug|Food|SIMPLE_SEGMENT|18403,18408|false|false|false|C0452588|Start brand of breakfast cereal|START
Event|Event|SIMPLE_SEGMENT|18403,18408|false|false|false|||START
Finding|Intellectual Product|SIMPLE_SEGMENT|18403,18408|false|false|false|C1552850|start - HtmlLinkType|START
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|18403,18408|false|false|false|C5447432|Collagen Tile Brachytherapy|START
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|18409,18419|false|false|false|C0042313|vancomycin|vancomycin
Drug|Antibiotic|SIMPLE_SEGMENT|18409,18419|false|false|false|C0042313|vancomycin|vancomycin
Event|Event|SIMPLE_SEGMENT|18409,18419|false|false|false|||vancomycin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|18409,18419|false|false|false|C0489941|Vancomycin measurement|vancomycin
Event|Event|SIMPLE_SEGMENT|18420,18425|false|false|false|||500mg
Finding|Functional Concept|SIMPLE_SEGMENT|18426,18434|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|18429,18434|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|18429,18434|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Food|SIMPLE_SEGMENT|18461,18466|false|false|false|C0452588|Start brand of breakfast cereal|START
Event|Event|SIMPLE_SEGMENT|18461,18466|false|false|false|||START
Finding|Intellectual Product|SIMPLE_SEGMENT|18461,18466|false|false|false|C1552850|start - HtmlLinkType|START
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|18461,18466|false|false|false|C5447432|Collagen Tile Brachytherapy|START
Drug|Organic Chemical|SIMPLE_SEGMENT|18467,18477|false|false|false|C0171023|olanzapine|olanzapine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|18467,18477|false|false|false|C0171023|olanzapine|olanzapine
Event|Event|SIMPLE_SEGMENT|18467,18477|false|false|false|||olanzapine
Event|Event|SIMPLE_SEGMENT|18499,18505|false|false|false|||needed
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|18510,18517|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Event|Event|SIMPLE_SEGMENT|18510,18517|false|false|false|||anxiety
Finding|Sign or Symptom|SIMPLE_SEGMENT|18510,18517|false|false|false|C0860603|Anxiety symptoms|anxiety
Procedure|Health Care Activity|SIMPLE_SEGMENT|18520,18528|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|18529,18541|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|18529,18541|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|18529,18541|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

