 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|26,30
No|31,33
:|33,34
_|37,38
_|38,39
_|39,40
<EOL>|40,41
<EOL>|42,43
Admission|43,52
Date|53,57
:|57,58
_|60,61
_|61,62
_|62,63
Discharge|77,86
Date|87,91
:|91,92
_|95,96
_|96,97
_|97,98
<EOL>|98,99
<EOL>|100,101
Date|101,105
of|106,108
Birth|109,114
:|114,115
_|117,118
_|118,119
_|119,120
Sex|133,136
:|136,137
F|140,141
<EOL>|141,142
<EOL>|143,144
Service|144,151
:|151,152
MEDICINE|153,161
<EOL>|161,162
<EOL>|163,164
No|176,178
Known|179,184
Allergies|185,194
/|195,196
Adverse|197,204
Drug|205,209
Reactions|210,219
<EOL>|219,220
<EOL>|221,222
Attending|222,231
:|231,232
_|233,234
_|234,235
_|235,236
<EOL>|236,237
<EOL>|238,239
dyspnea|257,264
on|265,267
exertion|268,276
<EOL>|277,278
<EOL>|279,280
Major|280,285
Surgical|286,294
or|295,297
Invasive|298,306
Procedure|307,316
:|316,317
<EOL>|317,318
None|318,322
<EOL>|322,323
<EOL>|323,324
<EOL>|325,326
Patient|354,361
is|362,364
a|365,366
_|367,368
_|368,369
_|369,370
year|371,375
old|376,379
woman|380,385
s|386,387
/|387,388
p|388,389
robotic|390,397
radical|398,405
cystectomy|406,416
<EOL>|417,418
_|418,419
_|419,420
_|420,421
(|422,423
with|423,427
ileal|428,433
conduit|434,441
creation|442,450
)|450,451
with|452,456
postop|457,463
course|464,470
<EOL>|471,472
complicated|472,483
by|484,486
bacteremia|487,497
and|498,501
abscess|502,509
,|509,510
LLE|511,514
DVT|515,518
(|519,520
on|520,522
prophylactic|523,535
<EOL>|536,537
dosing|537,543
lovenox|544,551
)|551,552
who|553,556
presents|557,565
with|566,570
dyspnea|571,578
on|579,581
exertion|582,590
for|591,594
past|595,599
3|600,601
<EOL>|602,603
days|603,607
.|607,608
<EOL>|609,610
<EOL>|610,611
Briefly|611,618
,|618,619
patient|620,627
was|628,631
initially|632,641
admitted|642,650
to|651,653
the|654,657
Urology|658,665
service|666,673
<EOL>|674,675
from|675,679
_|680,681
_|681,682
_|682,683
for|684,687
robotic|688,695
anterior|696,704
exenteration|705,717
with|718,722
ileal|723,728
<EOL>|729,730
conduit|730,737
.|737,738
She|739,742
was|743,746
discharged|747,757
to|758,760
rehab|761,766
on|767,769
prophylactic|770,782
dosing|783,789
<EOL>|790,791
lovenox|791,798
for|799,802
1|803,804
month|805,810
.|810,811
She|812,815
was|816,819
then|820,824
readmitted|825,835
from|836,840
_|841,842
_|842,843
_|843,844
for|845,848
<EOL>|849,850
ileus|850,855
requiring|856,865
NGT|866,869
decompression|870,883
,|883,884
TPN|885,888
.|888,889
BCx|890,893
grew|894,898
Citrobacter|899,910
,|910,911
<EOL>|912,913
for|913,916
which|917,922
CTX|923,926
was|927,930
started|931,938
.|938,939
CT|940,942
showed|943,949
intra-abdominal|950,965
,|965,966
interloop|967,976
,|976,977
<EOL>|978,979
simple|979,985
fluid|986,991
collection|992,1002
and|1003,1006
LLQ|1007,1010
drain|1011,1016
was|1017,1020
placed|1021,1027
by|1028,1030
_|1031,1032
_|1032,1033
_|1033,1034
.|1034,1035
Patient|1036,1043
<EOL>|1044,1045
improved|1045,1053
,|1053,1054
passing|1055,1062
BMs|1063,1066
and|1067,1070
tolerating|1071,1081
PO|1082,1084
,|1084,1085
and|1086,1089
was|1090,1093
discharged|1094,1104
on|1105,1107
<EOL>|1108,1109
cipro|1109,1114
/|1114,1115
flagyl|1115,1121
.|1121,1122
She|1123,1126
was|1127,1130
also|1131,1135
discharged|1136,1146
on|1147,1149
PO|1150,1152
Bactrim|1153,1160
for|1161,1164
presumed|1165,1173
<EOL>|1174,1175
UTI|1175,1178
,|1178,1179
though|1180,1186
unclear|1187,1194
if|1195,1197
she|1198,1201
actually|1202,1210
took|1211,1215
this|1216,1220
.|1220,1221
During|1222,1228
this|1229,1233
<EOL>|1234,1235
admission|1235,1244
,|1244,1245
she|1246,1249
was|1250,1253
noted|1254,1259
to|1260,1262
have|1263,1267
new|1268,1271
bilateral|1272,1281
_|1282,1283
_|1283,1284
_|1284,1285
edema|1286,1291
.|1291,1292
LENIs|1293,1298
<EOL>|1299,1300
at|1300,1302
the|1303,1306
time|1307,1311
showed|1312,1318
aute|1319,1323
deep|1324,1328
vein|1329,1333
thrombosis|1334,1344
of|1345,1347
the|1348,1351
duplicated|1352,1362
<EOL>|1363,1364
mid|1364,1367
and|1368,1371
distal|1372,1378
left|1379,1383
femoral|1384,1391
veins|1392,1397
.|1397,1398
She|1399,1402
was|1403,1406
discharged|1407,1417
on|1418,1420
<EOL>|1422,1423
Enoxaparin|1423,1433
Sodium|1434,1440
40|1441,1443
mg|1444,1446
SC|1447,1449
daily|1450,1455
.|1455,1456
She|1457,1460
reports|1461,1468
that|1469,1473
her|1474,1477
PCP|1478,1481
<EOL>|1482,1483
started|1483,1490
PO|1491,1493
_|1494,1495
_|1495,1496
_|1496,1497
20mg|1498,1502
daily|1503,1508
and|1509,1512
since|1513,1518
then|1519,1523
there|1524,1529
has|1530,1533
been|1534,1538
<EOL>|1539,1540
improvement|1540,1551
of|1552,1554
the|1555,1558
swelling|1559,1567
.|1567,1568
Per|1569,1572
her|1573,1576
report|1577,1583
,|1583,1584
a|1585,1586
repeat|1587,1593
_|1594,1595
_|1595,1596
_|1596,1597
at|1598,1600
<EOL>|1601,1602
the|1602,1605
rehab|1606,1611
facility|1612,1620
(|1621,1622
_|1622,1623
_|1623,1624
_|1624,1625
)|1625,1626
was|1627,1630
negative|1631,1639
for|1640,1643
DVT|1644,1647
.|1647,1648
<EOL>|1648,1649
<EOL>|1649,1650
Patient|1650,1657
reports|1658,1665
that|1666,1670
she|1671,1674
recovered|1675,1684
well|1685,1689
post-operatively|1690,1706
and|1707,1710
was|1711,1714
<EOL>|1715,1716
doing|1716,1721
well|1722,1726
at|1727,1729
her|1730,1733
assisted|1734,1742
living|1743,1749
facility|1750,1758
up|1759,1761
until|1762,1767
a|1768,1769
week|1770,1774
ago|1775,1778
<EOL>|1779,1780
when|1780,1784
she|1785,1788
began|1789,1794
experiencing|1795,1807
dyspnea|1808,1815
on|1816,1818
exertion|1819,1827
.|1827,1828
She|1829,1832
states|1833,1839
that|1840,1844
<EOL>|1845,1846
she|1846,1849
typically|1850,1859
is|1860,1862
able|1863,1867
to|1868,1870
ambulate|1871,1879
a|1880,1881
block|1882,1887
before|1888,1894
stopping|1895,1903
to|1904,1906
<EOL>|1907,1908
catch|1908,1913
her|1914,1917
breath|1918,1924
,|1924,1925
however|1926,1933
in|1934,1936
the|1937,1940
past|1941,1945
week|1946,1950
she|1951,1954
has|1955,1958
been|1959,1963
unable|1964,1970
<EOL>|1971,1972
to|1972,1974
take|1975,1979
more|1980,1984
than|1985,1989
a|1990,1991
few|1992,1995
steps|1996,2001
.|2001,2002
She|2003,2006
states|2007,2013
that|2014,2018
it|2019,2021
has|2022,2025
become|2026,2032
<EOL>|2033,2034
increasingly|2034,2046
more|2047,2051
difficult|2052,2061
to|2062,2064
ambulate|2065,2073
from|2074,2078
her|2079,2082
bedroom|2083,2090
to|2091,2093
the|2094,2097
<EOL>|2098,2099
bathroom|2099,2107
.|2107,2108
When|2109,2113
visited|2114,2121
by|2122,2124
the|2125,2128
NP|2129,2131
her|2132,2135
ambulatory|2136,2146
saturation|2147,2157
was|2158,2161
<EOL>|2162,2163
noted|2163,2168
to|2169,2171
be|2172,2174
in|2175,2177
the|2178,2181
_|2182,2183
_|2183,2184
_|2184,2185
with|2186,2190
associated|2191,2201
tachycardia|2202,2213
to|2214,2216
110|2217,2220
,|2220,2221
<EOL>|2222,2223
pallor|2223,2229
and|2230,2233
diaphoresis|2234,2245
.|2245,2246
She|2247,2250
endorses|2251,2259
associated|2260,2270
leg|2271,2274
swelling|2275,2283
<EOL>|2284,2285
left|2285,2289
worse|2290,2295
than|2296,2300
right|2301,2306
,|2306,2307
and|2308,2311
she|2312,2315
states|2316,2322
that|2323,2327
her|2328,2331
thighs|2332,2338
"|2339,2340
feel|2340,2344
<EOL>|2345,2346
heavy|2346,2351
"|2351,2352
.|2352,2353
She|2354,2357
denies|2358,2364
any|2365,2368
associated|2369,2379
chest|2380,2385
pain|2386,2390
,|2390,2391
fever|2392,2397
,|2397,2398
chills|2399,2405
,|2405,2406
<EOL>|2407,2408
pain|2408,2412
with|2413,2417
deep|2418,2422
inspiration|2423,2434
,|2434,2435
abdominal|2436,2445
pain|2446,2450
,|2450,2451
rashes|2452,2458
,|2458,2459
dizziness|2460,2469
,|2469,2470
<EOL>|2471,2472
lightheadedness|2472,2487
.|2487,2488
<EOL>|2490,2491
<EOL>|2491,2492
In|2492,2494
the|2495,2498
ED|2499,2501
,|2501,2502
initial|2503,2510
VS|2511,2513
were|2514,2518
:|2518,2519
97.7|2520,2524
72|2525,2527
136|2528,2531
/|2531,2532
93|2532,2534
20|2535,2537
100|2538,2541
%|2541,2542
Nasal|2543,2548
Cannula|2549,2556
<EOL>|2557,2558
<EOL>|2558,2559
ED|2559,2561
physical|2562,2570
exam|2571,2575
was|2576,2579
recorded|2580,2588
as|2589,2591
patient|2592,2599
resting|2600,2607
comfortably|2608,2619
<EOL>|2620,2621
with|2621,2625
NC|2626,2628
,|2628,2629
pursed|2630,2636
lip|2637,2640
breathing|2641,2650
,|2650,2651
unable|2652,2658
to|2659,2661
speak|2662,2667
in|2668,2670
full|2671,2675
sentences|2676,2685
<EOL>|2686,2687
before|2687,2693
becoming|2694,2702
short|2703,2708
of|2709,2711
breath|2712,2718
,|2718,2719
urostomy|2720,2728
pouch|2729,2734
in|2735,2737
RLQ|2738,2741
,|2741,2742
stoma|2743,2748
<EOL>|2749,2750
pink|2750,2754
,|2754,2755
2|2756,2757
+|2757,2758
edema|2759,2764
to|2765,2767
bilateral|2768,2777
lower|2778,2783
extremities|2784,2795
L|2796,2797
>|2797,2798
R|2798,2799
.|2799,2800
<EOL>|2801,2802
<EOL>|2802,2803
ED|2803,2805
labs|2806,2810
were|2811,2815
notable|2816,2823
for|2824,2827
:|2827,2828
Hb|2829,2831
9|2832,2833
,|2833,2834
Hct|2835,2838
29|2839,2841
,|2841,2842
plt|2843,2846
479|2847,2850
,|2850,2851
UA|2852,2854
:|2854,2855
large|2856,2861
_|2862,2863
_|2863,2864
_|2864,2865
,|2865,2866
<EOL>|2867,2868
>|2868,2869
182|2869,2872
WBC|2873,2876
,|2876,2877
many|2878,2882
bact|2883,2887
0|2888,2889
epi|2890,2893
.|2893,2894
Trop|2895,2899
neg|2900,2903
x1|2904,2906
,|2906,2907
proBNP|2908,2914
normal|2915,2921
<EOL>|2921,2922
<EOL>|2922,2923
CTA|2923,2926
chest|2927,2932
showed|2933,2939
:|2939,2940
<EOL>|2940,2941
1.|2941,2943
Extensive|2944,2953
pulmonary|2954,2963
embolism|2964,2972
with|2973,2977
thrombus|2978,2986
seen|2987,2991
extending|2992,3001
<EOL>|3002,3003
from|3003,3007
the|3008,3011
right|3012,3017
main|3018,3022
pulmonary|3023,3032
artery|3033,3039
into|3040,3044
the|3045,3048
segmental|3049,3058
and|3059,3062
<EOL>|3063,3064
subsegmental|3064,3076
right|3077,3082
upper|3083,3088
,|3088,3089
middle|3090,3096
,|3096,3097
and|3098,3101
lower|3102,3107
lobe|3108,3112
pulmonary|3113,3122
<EOL>|3123,3124
arteries|3124,3132
.|3132,3133
No|3134,3136
right|3137,3142
heart|3143,3148
strain|3149,3155
identified|3156,3166
.|3166,3167
2.|3168,3170
Additionally|3171,3183
,|3183,3184
<EOL>|3185,3186
there|3186,3191
are|3192,3195
smaller|3196,3203
pulmonary|3204,3213
emboli|3214,3220
seen|3221,3225
in|3226,3228
the|3229,3232
segmental|3233,3242
and|3243,3246
<EOL>|3247,3248
subsegmental|3248,3260
branches|3261,3269
of|3270,3272
the|3273,3276
left|3277,3281
upper|3282,3287
and|3288,3291
lower|3292,3297
lobes|3298,3303
.|3303,3304
3|3305,3306
.|3306,3307
<EOL>|3308,3309
Several|3309,3316
pulmonary|3317,3326
nodules|3327,3334
are|3335,3338
noted|3339,3344
,|3344,3345
as|3346,3348
noted|3349,3354
previously|3355,3365
,|3365,3366
with|3367,3371
<EOL>|3372,3373
the|3373,3376
largest|3377,3384
appearing|3385,3394
spiculated|3395,3405
and|3406,3409
measuring|3410,3419
up|3420,3422
to|3423,3425
1|3426,3427
cm|3428,3430
in|3431,3433
the|3434,3437
<EOL>|3438,3439
right|3439,3444
middle|3445,3451
lobe|3452,3456
,|3456,3457
suspicious|3458,3468
for|3469,3472
malignancy|3473,3483
on|3484,3486
the|3487,3490
previous|3491,3499
<EOL>|3500,3501
PET|3501,3504
-|3504,3505
CT|3505,3507
.|3507,3508
4.|3509,3511
Re|3512,3514
-|3514,3515
demonstration|3516,3529
of|3530,3532
2|3533,3534
left|3535,3539
breast|3540,3546
nodules|3547,3554
for|3555,3558
which|3559,3564
<EOL>|3565,3566
correlation|3566,3577
with|3578,3582
mammography|3583,3594
and|3595,3598
ultrasound|3599,3609
is|3610,3612
suggested|3613,3622
.|3622,3623
<EOL>|3623,3624
<EOL>|3624,3625
EKG|3625,3628
showed|3629,3635
NSR|3636,3639
with|3640,3644
frequent|3645,3653
PAC|3654,3657
<EOL>|3657,3658
<EOL>|3658,3659
Patient|3659,3666
was|3667,3670
given|3671,3676
:|3676,3677
<EOL>|3677,3678
_|3678,3679
_|3679,3680
_|3680,3681
20|3682,3684
:|3684,3685
26|3685,3687
PO|3688,3690
/|3690,3691
NG|3691,3693
Ciprofloxacin|3694,3707
HCl|3708,3711
500|3712,3715
mg|3716,3718
<EOL>|3719,3720
_|3720,3721
_|3721,3722
_|3722,3723
20|3724,3726
:|3726,3727
26|3727,3729
IV|3730,3732
Heparin|3733,3740
6600|3741,3745
UNIT|3746,3750
<EOL>|3751,3752
_|3752,3753
_|3753,3754
_|3754,3755
20|3756,3758
:|3758,3759
26|3759,3761
IV|3762,3764
Heparin|3765,3772
<EOL>|3774,3775
<EOL>|3775,3776
Transfer|3776,3784
VS|3785,3787
were|3788,3792
:|3792,3793
98.1|3794,3798
77|3799,3801
145|3802,3805
/|3805,3806
63|3806,3808
20|3809,3811
99|3812,3814
%|3814,3815
Nasal|3816,3821
Cannula|3822,3829
<EOL>|3830,3831
When|3832,3836
seen|3837,3841
on|3842,3844
the|3845,3848
floor|3849,3854
,|3854,3855
she|3856,3859
reports|3860,3867
significant|3868,3879
dyspnea|3880,3887
with|3888,3892
<EOL>|3893,3894
minimal|3894,3901
exertion|3902,3910
.|3910,3911
Denies|3912,3918
chest|3919,3924
pain|3925,3929
,|3929,3930
palpitations|3931,3943
,|3943,3944
<EOL>|3945,3946
lightheadedness|3946,3961
.|3961,3962
<EOL>|3962,3963
A|3963,3964
ten|3965,3968
point|3969,3974
ROS|3975,3978
was|3979,3982
conducted|3983,3992
and|3993,3996
was|3997,4000
negative|4001,4009
except|4010,4016
as|4017,4019
above|4020,4025
<EOL>|4026,4027
in|4027,4029
the|4030,4033
HPI|4034,4037
.|4037,4038
<EOL>|4038,4039
<EOL>|4040,4041
Hypertension|4063,4075
,|4075,4076
laparoscopic|4077,4089
cholecystectomy|4090,4105
,|4105,4106
left|4107,4111
knee|4112,4116
<EOL>|4117,4118
replacement|4118,4129
six|4130,4133
to|4134,4136
_|4137,4138
_|4138,4139
_|4139,4140
years|4141,4146
ago|4147,4150
,|4150,4151
laminectomy|4152,4163
of|4164,4166
L5|4167,4169
-|4169,4170
S1|4170,4172
at|4173,4175
age|4176,4179
<EOL>|4180,4181
_|4181,4182
_|4182,4183
_|4183,4184
,|4184,4185
two|4186,4189
vaginal|4190,4197
deliveries|4198,4208
.|4208,4209
<EOL>|4209,4210
<EOL>|4210,4211
s|4211,4212
/|4212,4213
p|4213,4214
_|4215,4216
_|4216,4217
_|4217,4218
:|4218,4219
<EOL>|4220,4221
1.|4221,4223
Robot|4225,4230
-|4230,4231
assisted|4231,4239
laparoscopic|4240,4252
bilateral|4253,4262
pelvic|4263,4269
lymph|4270,4275
node|4276,4280
<EOL>|4281,4282
dissection|4282,4292
.|4292,4293
<EOL>|4293,4294
2.|4294,4296
Robot|4297,4302
-|4302,4303
assisted|4303,4311
hysterectomy|4312,4324
and|4325,4328
bilateral|4329,4338
oophorectomy|4339,4351
for|4352,4355
<EOL>|4356,4357
large|4357,4362
uterus|4363,4369
,|4369,4370
greater|4371,4378
than|4379,4383
300|4384,4387
grams|4388,4393
,|4393,4394
with|4395,4399
large|4400,4405
fibroid|4406,4413
.|4413,4414
<EOL>|4414,4415
3.|4415,4417
Laparoscopic|4418,4430
radical|4431,4438
cystectomy|4439,4449
and|4450,4453
anterior|4454,4462
vaginectomy|4463,4474
with|4475,4479
<EOL>|4480,4481
vaginal|4481,4488
reconstruction|4489,4503
.|4503,4504
<EOL>|4504,4505
<EOL>|4505,4506
<EOL>|4507,4508
:|4522,4523
<EOL>|4523,4524
_|4524,4525
_|4525,4526
_|4526,4527
<EOL>|4527,4528
:|4542,4543
<EOL>|4543,4544
Negative|4544,4552
for|4553,4556
bladder|4557,4564
CA|4565,4567
.|4567,4568
<EOL>|4568,4569
<EOL>|4569,4570
<EOL>|4571,4572
ADMISSION|4587,4596
EXAM|4597,4601
:|4601,4602
<EOL>|4602,4603
Gen|4604,4607
:|4607,4608
NAD|4609,4612
,|4612,4613
speaking|4614,4622
in|4623,4625
3|4626,4627
word|4628,4632
sentences|4633,4642
,|4642,4643
pursed|4644,4650
lip|4651,4654
breathing|4655,4664
,|4664,4665
<EOL>|4666,4667
no|4667,4669
accessory|4670,4679
muscle|4680,4686
use|4687,4690
,|4690,4691
lying|4692,4697
in|4698,4700
bed|4701,4704
<EOL>|4704,4705
Eyes|4706,4710
:|4710,4711
EOMI|4712,4716
,|4716,4717
sclerae|4718,4725
anicteric|4726,4735
<EOL>|4737,4738
ENT|4739,4742
:|4742,4743
MMM|4744,4747
,|4747,4748
OP|4749,4751
clear|4752,4757
<EOL>|4757,4758
Cardiovasc|4759,4769
:|4769,4770
RRR|4771,4774
,|4774,4775
no|4776,4778
MRG|4779,4782
,|4782,4783
full|4784,4788
pulses|4789,4795
,|4795,4796
1|4797,4798
+|4798,4799
edema|4800,4805
bilaterally|4806,4817
with|4818,4822
<EOL>|4823,4824
compression|4824,4835
stockings|4836,4845
in|4846,4848
place|4849,4854
,|4854,4855
no|4856,4858
JVD|4859,4862
<EOL>|4863,4864
Resp|4865,4869
:|4869,4870
normal|4871,4877
effort|4878,4884
,|4884,4885
no|4886,4888
accessory|4889,4898
muscle|4899,4905
use|4906,4909
,|4909,4910
lungs|4911,4916
CTA|4917,4920
_|4921,4922
_|4922,4923
_|4923,4924
to|4925,4927
<EOL>|4928,4929
anterior|4929,4937
auscultation|4938,4950
.|4950,4951
<EOL>|4951,4952
GI|4953,4955
:|4955,4956
soft|4957,4961
,|4961,4962
NT|4963,4965
,|4965,4966
ND|4967,4969
,|4969,4970
BS|4971,4973
+|4973,4974
.|4974,4975
Urostomy|4976,4984
site|4985,4989
does|4990,4994
not|4995,4998
appear|4999,5005
infected|5006,5014
<EOL>|5014,5015
MSK|5016,5019
:|5019,5020
No|5021,5023
significant|5024,5035
kyphosis|5036,5044
.|5044,5045
No|5046,5048
palpable|5049,5057
synovitis|5058,5067
.|5067,5068
<EOL>|5068,5069
Skin|5070,5074
:|5074,5075
No|5076,5078
visible|5079,5086
rash|5087,5091
.|5091,5092
No|5093,5095
jaundice|5096,5104
.|5104,5105
<EOL>|5105,5106
Neuro|5107,5112
:|5112,5113
AAOx3|5114,5119
.|5119,5120
No|5121,5123
facial|5124,5130
droop|5131,5136
.|5136,5137
<EOL>|5137,5138
Psych|5139,5144
:|5144,5145
Full|5146,5150
range|5151,5156
of|5157,5159
affect|5160,5166
<EOL>|5167,5168
<EOL>|5168,5169
DISCHARGE|5169,5178
EXAM|5179,5183
:|5183,5184
<EOL>|5184,5185
vitals|5185,5191
:|5191,5192
98.3|5193,5197
140|5198,5201
/|5201,5202
42|5202,5204
90|5205,5207
24|5208,5210
96|5211,5213
%|5213,5214
1L|5215,5217
<EOL>|5217,5218
Gen|5218,5221
:|5221,5222
Lying|5223,5228
in|5229,5231
bed|5232,5235
in|5236,5238
no|5239,5241
apparent|5242,5250
distress|5251,5259
<EOL>|5259,5260
HEENT|5260,5265
:|5265,5266
Anicteric|5267,5276
,|5276,5277
MMM|5278,5281
<EOL>|5281,5282
Cardiovascular|5282,5296
:|5296,5297
RRR|5298,5301
normal|5302,5308
S1|5309,5311
,|5311,5312
S2|5313,5315
,|5315,5316
no|5317,5319
right|5320,5325
sided|5326,5331
heave|5332,5337
,|5337,5338
_|5339,5340
_|5340,5341
_|5341,5342
<EOL>|5343,5344
systolic|5344,5352
murmur|5353,5359
<EOL>|5360,5361
Pulmonary|5361,5370
:|5370,5371
Lung|5372,5376
fields|5377,5383
clear|5384,5389
to|5390,5392
auscultation|5393,5405
throughout|5406,5416
.|5416,5417
No|5418,5420
<EOL>|5421,5422
crackles|5422,5430
or|5431,5433
wheezing|5434,5442
.|5442,5443
<EOL>|5444,5445
GI|5445,5447
:|5447,5448
Soft|5449,5453
,|5453,5454
distended|5455,5464
,|5464,5465
nontender|5466,5475
,|5475,5476
bowel|5477,5482
sounds|5483,5489
present|5490,5497
,|5497,5498
urostomy|5499,5507
<EOL>|5508,5509
in|5509,5511
place|5512,5517
.|5517,5518
<EOL>|5518,5519
Extremities|5519,5530
:|5530,5531
no|5532,5534
edema|5535,5540
,|5540,5541
though|5542,5548
left|5549,5553
leg|5554,5557
appears|5558,5565
larger|5566,5572
than|5573,5577
right|5578,5583
<EOL>|5584,5585
leg|5585,5588
,|5588,5589
warm|5590,5594
,|5594,5595
well|5596,5600
perfused|5601,5609
with|5610,5614
motor|5615,5620
function|5621,5629
intact|5630,5636
.|5636,5637
Her|5638,5641
left|5642,5646
<EOL>|5647,5648
lower|5648,5653
leg|5654,5657
is|5658,5660
wrapped|5661,5668
.|5668,5669
<EOL>|5670,5671
<EOL>|5671,5672
<EOL>|5673,5674
Pertinent|5674,5683
Results|5684,5691
:|5691,5692
<EOL>|5692,5693
LABS|5693,5697
:|5697,5698
<EOL>|5698,5699
=|5699,5700
=|5700,5701
=|5701,5702
=|5702,5703
=|5703,5704
=|5704,5705
=|5705,5706
=|5706,5707
=|5707,5708
=|5708,5709
=|5709,5710
=|5710,5711
=|5711,5712
=|5712,5713
=|5713,5714
=|5714,5715
=|5715,5716
=|5716,5717
=|5717,5718
=|5718,5719
=|5719,5720
=|5720,5721
=|5721,5722
=|5722,5723
=|5723,5724
=|5724,5725
<EOL>|5725,5726
Admission|5726,5735
labs|5736,5740
:|5740,5741
<EOL>|5741,5742
_|5742,5743
_|5743,5744
_|5744,5745
02|5746,5748
:|5748,5749
40PM|5749,5753
GLUCOSE|5756,5763
-|5763,5764
101|5764,5767
*|5767,5768
UREA|5769,5773
N|5774,5775
-|5775,5776
22|5776,5778
*|5778,5779
CREAT|5780,5785
-|5785,5786
0.7|5786,5789
SODIUM|5790,5796
-|5796,5797
136|5797,5800
<EOL>|5801,5802
POTASSIUM|5802,5811
-|5811,5812
4.1|5812,5815
CHLORIDE|5816,5824
-|5824,5825
98|5825,5827
TOTAL|5828,5833
CO2|5834,5837
-|5837,5838
22|5838,5840
ANION|5841,5846
GAP|5847,5850
-|5850,5851
20|5851,5853
<EOL>|5853,5854
_|5854,5855
_|5855,5856
_|5856,5857
02|5858,5860
:|5860,5861
40PM|5861,5865
cTropnT|5868,5875
-|5875,5876
<|5876,5877
0|5877,5878
.|5878,5879
01|5879,5881
<EOL>|5881,5882
_|5882,5883
_|5883,5884
_|5884,5885
02|5886,5888
:|5888,5889
40PM|5889,5893
proBNP|5896,5902
-|5902,5903
567|5903,5906
<EOL>|5906,5907
_|5907,5908
_|5908,5909
_|5909,5910
02|5911,5913
:|5913,5914
40PM|5914,5918
WBC|5921,5924
-|5924,5925
7.7|5925,5928
RBC|5929,5932
-|5932,5933
3|5933,5934
.|5934,5935
07|5935,5937
*|5937,5938
HGB|5939,5942
-|5942,5943
9|5943,5944
.|5944,5945
0|5945,5946
*|5946,5947
HCT|5948,5951
-|5951,5952
29|5952,5954
.|5954,5955
1|5955,5956
*|5956,5957
MCV|5958,5961
-|5961,5962
95|5962,5964
<EOL>|5965,5966
MCH|5966,5969
-|5969,5970
29.3|5970,5974
MCHC|5975,5979
-|5979,5980
30|5980,5982
.|5982,5983
9|5983,5984
*|5984,5985
RDW|5986,5989
-|5989,5990
14.9|5990,5994
RDWSD|5995,6000
-|6000,6001
52|6001,6003
.|6003,6004
1|6004,6005
*|6005,6006
<EOL>|6006,6007
_|6007,6008
_|6008,6009
_|6009,6010
02|6011,6013
:|6013,6014
40PM|6014,6018
PLT|6021,6024
COUNT|6025,6030
-|6030,6031
479|6031,6034
*|6034,6035
<EOL>|6035,6036
_|6036,6037
_|6037,6038
_|6038,6039
02|6040,6042
:|6042,6043
40PM|6043,6047
_|6050,6051
_|6051,6052
_|6052,6053
PTT|6054,6057
-|6057,6058
33.4|6058,6062
_|6063,6064
_|6064,6065
_|6065,6066
<EOL>|6066,6067
<EOL>|6067,6068
Discharge|6068,6077
labs|6078,6082
:|6082,6083
<EOL>|6083,6084
_|6084,6085
_|6085,6086
_|6086,6087
06|6088,6090
:|6090,6091
55AM|6091,6095
BLOOD|6096,6101
WBC|6102,6105
-|6105,6106
11|6106,6108
.|6108,6109
0|6109,6110
*|6110,6111
RBC|6112,6115
-|6115,6116
2|6116,6117
.|6117,6118
60|6118,6120
*|6120,6121
Hgb|6122,6125
-|6125,6126
7|6126,6127
.|6127,6128
5|6128,6129
*|6129,6130
Hct|6131,6134
-|6134,6135
24|6135,6137
.|6137,6138
5|6138,6139
*|6139,6140
<EOL>|6141,6142
MCV|6142,6145
-|6145,6146
94|6146,6148
MCH|6149,6152
-|6152,6153
28.8|6153,6157
MCHC|6158,6162
-|6162,6163
30|6163,6165
.|6165,6166
6|6166,6167
*|6167,6168
RDW|6169,6172
-|6172,6173
14.8|6173,6177
RDWSD|6178,6183
-|6183,6184
51|6184,6186
.|6186,6187
4|6187,6188
*|6188,6189
Plt|6190,6193
_|6194,6195
_|6195,6196
_|6196,6197
<EOL>|6197,6198
_|6198,6199
_|6199,6200
_|6200,6201
06|6202,6204
:|6204,6205
55AM|6205,6209
BLOOD|6210,6215
Glucose|6216,6223
-|6223,6224
99|6224,6226
UreaN|6227,6232
-|6232,6233
10|6233,6235
Creat|6236,6241
-|6241,6242
0.5|6242,6245
Na|6246,6248
-|6248,6249
141|6249,6252
<EOL>|6253,6254
K|6254,6255
-|6255,6256
4.3|6256,6259
Cl|6260,6262
-|6262,6263
105|6263,6266
HCO3|6267,6271
-|6271,6272
26|6272,6274
AnGap|6275,6280
-|6280,6281
14|6281,6283
<EOL>|6283,6284
_|6284,6285
_|6285,6286
_|6286,6287
06|6288,6290
:|6290,6291
55AM|6291,6295
BLOOD|6296,6301
Calcium|6302,6309
-|6309,6310
8|6310,6311
.|6311,6312
2|6312,6313
*|6313,6314
Phos|6315,6319
-|6319,6320
3.8|6320,6323
Mg|6324,6326
-|6326,6327
2.0|6327,6330
<EOL>|6330,6331
_|6331,6332
_|6332,6333
_|6333,6334
07|6335,6337
:|6337,6338
15AM|6338,6342
BLOOD|6343,6348
calTIBC|6349,6356
-|6356,6357
134|6357,6360
*|6360,6361
Ferritn|6362,6369
-|6369,6370
507|6370,6373
*|6373,6374
TRF|6375,6378
-|6378,6379
103|6379,6382
*|6382,6383
<EOL>|6383,6384
_|6384,6385
_|6385,6386
_|6386,6387
07|6388,6390
:|6390,6391
15AM|6391,6395
BLOOD|6396,6401
Iron|6402,6406
-|6406,6407
18|6407,6409
*|6409,6410
<EOL>|6410,6411
<EOL>|6411,6412
MICROBIOLOGY|6412,6424
<EOL>|6424,6425
=|6425,6426
=|6426,6427
=|6427,6428
=|6428,6429
=|6429,6430
=|6430,6431
=|6431,6432
=|6432,6433
=|6433,6434
=|6434,6435
=|6435,6436
=|6436,6437
=|6437,6438
=|6438,6439
=|6439,6440
=|6440,6441
=|6441,6442
=|6442,6443
=|6443,6444
=|6444,6445
=|6445,6446
=|6446,6447
=|6447,6448
=|6448,6449
=|6449,6450
=|6450,6451
<EOL>|6451,6452
_|6452,6453
_|6453,6454
_|6454,6455
4|6456,6457
:|6457,6458
30|6458,6460
pm|6461,6463
URINE|6464,6469
<EOL>|6469,6470
<EOL>|6470,6471
*|6499,6500
*|6500,6501
FINAL|6501,6506
REPORT|6507,6513
_|6514,6515
_|6515,6516
_|6516,6517
<EOL>|6517,6518
<EOL>|6518,6519
URINE|6522,6527
CULTURE|6528,6535
(|6536,6537
Final|6537,6542
_|6543,6544
_|6544,6545
_|6545,6546
:|6546,6547
<EOL>|6548,6549
MIXED|6555,6560
BACTERIAL|6561,6570
FLORA|6571,6576
(|6577,6578
>|6579,6580
=|6580,6581
3|6582,6583
COLONY|6584,6590
TYPES|6591,6596
)|6596,6597
,|6597,6598
CONSISTENT|6599,6609
<EOL>|6610,6611
WITH|6611,6615
SKIN|6616,6620
<EOL>|6620,6621
AND|6627,6630
/|6630,6631
OR|6631,6633
GENITAL|6634,6641
CONTAMINATION|6642,6655
.|6655,6656
<EOL>|6657,6658
ENTEROCOCCUS|6664,6676
SP|6677,6679
.|6679,6680
.|6680,6681
>|6685,6686
100,000|6686,6693
CFU|6694,6697
/|6697,6698
mL|6698,6700
.|6700,6701
<EOL>|6702,6703
PREDOMINATING|6712,6725
ORGANISM|6726,6734
INTERPRET|6735,6744
RESULTS|6745,6752
WITH|6753,6757
CAUTION|6758,6765
.|6765,6766
<EOL>|6767,6768
<EOL>|6768,6769
SENSITIVITIES|6799,6812
:|6812,6813
MIC|6814,6817
expressed|6818,6827
in|6828,6830
<EOL>|6831,6832
MCG|6832,6835
/|6835,6836
ML|6836,6838
<EOL>|6838,6839
<EOL>|6861,6862
_|6862,6863
_|6863,6864
_|6864,6865
_|6865,6866
_|6866,6867
_|6867,6868
_|6868,6869
_|6869,6870
_|6870,6871
_|6871,6872
_|6872,6873
_|6873,6874
_|6874,6875
_|6875,6876
_|6876,6877
_|6877,6878
_|6878,6879
_|6879,6880
_|6880,6881
_|6881,6882
_|6882,6883
_|6883,6884
_|6884,6885
_|6885,6886
_|6886,6887
_|6887,6888
_|6888,6889
_|6889,6890
_|6890,6891
_|6891,6892
_|6892,6893
_|6893,6894
_|6894,6895
_|6895,6896
_|6896,6897
_|6897,6898
_|6898,6899
_|6899,6900
_|6900,6901
_|6901,6902
_|6902,6903
_|6903,6904
_|6904,6905
_|6905,6906
_|6906,6907
_|6907,6908
_|6908,6909
_|6909,6910
_|6910,6911
_|6911,6912
_|6912,6913
_|6913,6914
_|6914,6915
_|6915,6916
_|6916,6917
_|6917,6918
_|6918,6919
<EOL>|6919,6920
ENTEROCOCCUS|6949,6961
SP|6962,6964
.|6964,6965
<EOL>|6965,6966
||6995,6996
<EOL>|6999,7000
AMPICILLIN|7000,7010
-|7010,7011
-|7011,7012
-|7012,7013
-|7013,7014
-|7014,7015
-|7015,7016
-|7016,7017
-|7017,7018
-|7018,7019
-|7019,7020
-|7020,7021
-|7021,7022
<|7025,7026
=|7026,7027
2|7027,7028
S|7029,7030
<EOL>|7030,7031
NITROFURANTOIN|7031,7045
-|7045,7046
-|7046,7047
-|7047,7048
-|7048,7049
-|7049,7050
-|7050,7051
-|7051,7052
-|7052,7053
<|7055,7056
=|7056,7057
16|7057,7059
S|7060,7061
<EOL>|7061,7062
TETRACYCLINE|7062,7074
-|7074,7075
-|7075,7076
-|7076,7077
-|7077,7078
-|7078,7079
-|7079,7080
-|7080,7081
-|7081,7082
-|7082,7083
-|7083,7084
<|7087,7088
=|7088,7089
1|7089,7090
S|7091,7092
<EOL>|7092,7093
VANCOMYCIN|7093,7103
-|7103,7104
-|7104,7105
-|7105,7106
-|7106,7107
-|7107,7108
-|7108,7109
-|7109,7110
-|7110,7111
-|7111,7112
-|7112,7113
-|7113,7114
-|7114,7115
1|7120,7121
S|7122,7123
<EOL>|7123,7124
<EOL>|7124,7125
IMAGING|7125,7132
<EOL>|7132,7133
=|7133,7134
=|7134,7135
=|7135,7136
=|7136,7137
=|7137,7138
=|7138,7139
=|7139,7140
=|7140,7141
=|7141,7142
=|7142,7143
=|7143,7144
=|7144,7145
=|7145,7146
=|7146,7147
=|7147,7148
=|7148,7149
=|7149,7150
=|7150,7151
=|7151,7152
=|7152,7153
=|7153,7154
=|7154,7155
=|7155,7156
=|7156,7157
=|7157,7158
=|7158,7159
<EOL>|7159,7160
_|7160,7161
_|7161,7162
_|7162,7163
CXR|7164,7167
<EOL>|7167,7168
IMPRESSION|7168,7178
:|7178,7179
Hilar|7180,7185
congestion|7186,7196
without|7197,7204
frank|7205,7210
edema|7211,7216
.|7216,7217
No|7219,7221
convincing|7222,7232
<EOL>|7233,7234
signs|7234,7239
of|7240,7242
pneumonia|7243,7252
.|7252,7253
<EOL>|7253,7254
<EOL>|7254,7255
_|7255,7256
_|7256,7257
_|7257,7258
CTA|7259,7262
chest|7263,7268
showed|7269,7275
:|7275,7276
<EOL>|7276,7277
1.|7277,7279
Extensive|7280,7289
pulmonary|7290,7299
embolism|7300,7308
with|7309,7313
thrombus|7314,7322
seen|7323,7327
extending|7328,7337
<EOL>|7338,7339
from|7339,7343
the|7344,7347
right|7348,7353
main|7354,7358
pulmonary|7359,7368
artery|7369,7375
into|7376,7380
the|7381,7384
segmental|7385,7394
and|7395,7398
<EOL>|7399,7400
subsegmental|7400,7412
right|7413,7418
upper|7419,7424
,|7424,7425
middle|7426,7432
,|7432,7433
and|7434,7437
lower|7438,7443
lobe|7444,7448
pulmonary|7449,7458
<EOL>|7459,7460
arteries|7460,7468
.|7468,7469
No|7470,7472
right|7473,7478
heart|7479,7484
strain|7485,7491
identified|7492,7502
.|7502,7503
2.|7504,7506
Additionally|7507,7519
,|7519,7520
<EOL>|7521,7522
there|7522,7527
are|7528,7531
smaller|7532,7539
pulmonary|7540,7549
emboli|7550,7556
seen|7557,7561
in|7562,7564
the|7565,7568
segmental|7569,7578
and|7579,7582
<EOL>|7583,7584
subsegmental|7584,7596
branches|7597,7605
of|7606,7608
the|7609,7612
left|7613,7617
upper|7618,7623
and|7624,7627
lower|7628,7633
lobes|7634,7639
.|7639,7640
3|7641,7642
.|7642,7643
<EOL>|7644,7645
Several|7645,7652
pulmonary|7653,7662
nodules|7663,7670
are|7671,7674
noted|7675,7680
,|7680,7681
as|7682,7684
noted|7685,7690
previously|7691,7701
,|7701,7702
with|7703,7707
<EOL>|7708,7709
the|7709,7712
largest|7713,7720
appearing|7721,7730
spiculated|7731,7741
and|7742,7745
measuring|7746,7755
up|7756,7758
to|7759,7761
1|7762,7763
cm|7764,7766
in|7767,7769
the|7770,7773
<EOL>|7774,7775
right|7775,7780
middle|7781,7787
lobe|7788,7792
,|7792,7793
suspicious|7794,7804
for|7805,7808
malignancy|7809,7819
on|7820,7822
the|7823,7826
previous|7827,7835
<EOL>|7836,7837
PET|7837,7840
-|7840,7841
CT|7841,7843
.|7843,7844
4.|7845,7847
Re|7848,7850
-|7850,7851
demonstration|7852,7865
of|7866,7868
2|7869,7870
left|7871,7875
breast|7876,7882
nodules|7883,7890
for|7891,7894
which|7895,7900
<EOL>|7901,7902
correlation|7902,7913
with|7914,7918
mammography|7919,7930
and|7931,7934
ultrasound|7935,7945
is|7946,7948
suggested|7949,7958
.|7958,7959
<EOL>|7959,7960
<EOL>|7960,7961
_|7961,7962
_|7962,7963
_|7963,7964
_|7965,7966
_|7966,7967
_|7967,7968
:|7968,7969
<EOL>|7969,7970
1.|7982,7984
Interval|7985,7993
progression|7994,8005
of|8006,8008
deep|8009,8013
vein|8014,8018
thrombosis|8019,8029
in|8030,8032
the|8033,8036
left|8037,8041
<EOL>|8042,8043
lower|8043,8048
extremity|8049,8058
,|8058,8059
with|8060,8064
occlusive|8065,8074
thrombus|8075,8083
involving|8084,8093
the|8094,8097
entire|8098,8104
<EOL>|8105,8106
femoral|8106,8113
vein|8114,8118
,|8118,8119
previously|8120,8130
only|8131,8135
involving|8136,8145
the|8146,8149
mid|8150,8153
and|8154,8157
distal|8158,8164
<EOL>|8165,8166
femoral|8166,8173
vein|8174,8178
.|8178,8179
There|8181,8186
is|8187,8189
additional|8190,8200
nonocclusive|8201,8213
thrombus|8214,8222
in|8223,8225
the|8226,8229
<EOL>|8230,8231
deep|8231,8235
femoral|8236,8243
vein|8244,8248
.|8248,8249
The|8251,8254
left|8255,8259
common|8260,8266
femoral|8267,8274
and|8275,8278
popliteal|8279,8288
veins|8289,8294
<EOL>|8295,8296
are|8296,8299
patent|8300,8306
.|8306,8307
<EOL>|8307,8308
2|8308,8309
.|8309,8310
The|8311,8314
bilateral|8315,8324
calf|8325,8329
veins|8330,8335
were|8336,8340
not|8341,8344
visualized|8345,8355
due|8356,8359
to|8360,8362
an|8363,8365
<EOL>|8366,8367
overlying|8367,8376
dressing|8377,8385
.|8385,8386
Otherwise|8387,8396
no|8397,8399
evidence|8400,8408
of|8409,8411
deep|8412,8416
venous|8417,8423
<EOL>|8424,8425
thrombosis|8425,8435
in|8436,8438
the|8439,8442
right|8443,8448
lower|8449,8454
extremity|8455,8464
.|8464,8465
<EOL>|8465,8466
<EOL>|8466,8467
_|8467,8468
_|8468,8469
_|8469,8470
TTE|8471,8474
:|8474,8475
<EOL>|8475,8476
Conclusions|8476,8487
<EOL>|8487,8488
The|8488,8491
left|8492,8496
atrium|8497,8503
is|8504,8506
normal|8507,8513
in|8514,8516
size|8517,8521
.|8521,8522
The|8523,8526
estimated|8527,8536
right|8537,8542
atrial|8543,8549
<EOL>|8550,8551
pressure|8551,8559
is|8560,8562
_|8563,8564
_|8564,8565
_|8565,8566
mmHg|8567,8571
.|8571,8572
Left|8573,8577
ventricular|8578,8589
wall|8590,8594
thickness|8595,8604
,|8604,8605
cavity|8606,8612
<EOL>|8613,8614
size|8614,8618
,|8618,8619
and|8620,8623
global|8624,8630
systolic|8631,8639
function|8640,8648
are|8649,8652
normal|8653,8659
(|8660,8661
LVEF|8661,8665
>|8665,8666
55|8666,8668
%|8668,8669
)|8669,8670
.|8670,8671
<EOL>|8672,8673
Doppler|8673,8680
parameters|8681,8691
are|8692,8695
most|8696,8700
consistent|8701,8711
with|8712,8716
Grade|8717,8722
I|8723,8724
(|8725,8726
mild|8726,8730
)|8730,8731
left|8732,8736
<EOL>|8737,8738
ventricular|8738,8749
diastolic|8750,8759
dysfunction|8760,8771
.|8771,8772
Right|8773,8778
ventricular|8779,8790
chamber|8791,8798
<EOL>|8799,8800
size|8800,8804
and|8805,8808
free|8809,8813
wall|8814,8818
motion|8819,8825
are|8826,8829
normal|8830,8836
.|8836,8837
The|8838,8841
aortic|8842,8848
valve|8849,8854
leaflets|8855,8863
<EOL>|8864,8865
are|8865,8868
mildly|8869,8875
thickened|8876,8885
(|8886,8887
?|8887,8888
#|8888,8889
)|8889,8890
.|8890,8891
There|8892,8897
is|8898,8900
no|8901,8903
aortic|8904,8910
valve|8911,8916
stenosis|8917,8925
.|8925,8926
<EOL>|8927,8928
Trivial|8928,8935
mitral|8936,8942
regurgitation|8943,8956
is|8957,8959
seen|8960,8964
.|8964,8965
There|8966,8971
is|8972,8974
mild|8975,8979
pulmonary|8980,8989
<EOL>|8990,8991
artery|8991,8997
systolic|8998,9006
hypertension|9007,9019
.|9019,9020
<EOL>|9021,9022
<EOL>|9022,9023
_|9023,9024
_|9024,9025
_|9025,9026
CXR|9027,9030
<EOL>|9030,9031
Compared|9044,9052
to|9053,9055
chest|9056,9061
radiographs|9062,9073
_|9074,9075
_|9075,9076
_|9076,9077
through|9078,9085
_|9086,9087
_|9087,9088
_|9088,9089
.|9089,9090
<EOL>|9091,9092
Heart|9092,9097
size|9098,9102
top|9103,9106
-|9106,9107
normal|9107,9113
.|9113,9114
Lungs|9116,9121
grossly|9122,9129
clear|9130,9135
.|9135,9136
No|9138,9140
pleural|9141,9148
<EOL>|9149,9150
abnormality|9150,9161
or|9162,9164
evidence|9165,9173
of|9174,9176
central|9177,9184
lymph|9185,9190
node|9191,9195
enlargement|9196,9207
.|9207,9208
<EOL>|9208,9209
<EOL>|9209,9210
<EOL>|9211,9212
Ms.|9235,9238
_|9239,9240
_|9240,9241
_|9241,9242
is|9243,9245
a|9246,9247
_|9248,9249
_|9249,9250
_|9250,9251
woman|9252,9257
s|9258,9259
/|9259,9260
p|9260,9261
robotic|9262,9269
radical|9270,9277
cystectomy|9278,9288
<EOL>|9289,9290
_|9290,9291
_|9291,9292
_|9292,9293
omplicated|9293,9303
by|9304,9306
bacteremia|9307,9317
and|9318,9321
<EOL>|9322,9323
abscess|9323,9330
,|9330,9331
LLE|9332,9335
DVT|9336,9339
,|9339,9340
currently|9341,9350
on|9351,9353
daily|9354,9359
lovenox|9360,9367
who|9368,9371
presents|9372,9380
with|9381,9385
<EOL>|9386,9387
dyspnea|9387,9394
on|9395,9397
exertion|9398,9406
and|9407,9410
dyspnea|9411,9418
on|9419,9421
exertion|9422,9430
and|9431,9434
found|9435,9440
to|9441,9443
have|9444,9448
<EOL>|9449,9450
large|9450,9455
PE|9456,9458
and|9459,9462
progression|9463,9474
of|9475,9477
DVT|9478,9481
.|9481,9482
<EOL>|9482,9483
<EOL>|9483,9484
#|9484,9485
PE|9486,9488
/|9488,9489
DVT|9489,9492
:|9492,9493
Likely|9494,9500
due|9501,9504
to|9505,9507
undertreatment|9508,9522
of|9523,9525
known|9526,9531
LLE|9532,9535
DVT|9536,9539
with|9540,9544
<EOL>|9545,9546
prophylactic|9546,9558
dosing|9559,9565
of|9566,9568
lovenox|9569,9576
.|9576,9577
Given|9578,9583
underdosing|9584,9595
of|9596,9598
lovenox|9599,9606
,|9606,9607
<EOL>|9608,9609
this|9609,9613
was|9614,9617
not|9618,9621
thought|9622,9629
to|9630,9632
be|9633,9635
treatment|9636,9645
failure|9646,9653
and|9654,9657
IVC|9658,9661
filter|9662,9668
was|9669,9672
<EOL>|9673,9674
deferred|9674,9682
.|9682,9683
She|9684,9687
had|9688,9691
no|9692,9694
signs|9695,9700
of|9701,9703
right|9704,9709
heart|9710,9715
strain|9716,9722
on|9723,9725
imaging|9726,9733
,|9733,9734
<EOL>|9735,9736
EKG|9736,9739
,|9739,9740
exam|9741,9745
.|9745,9746
TTE|9747,9750
showed|9751,9757
no|9758,9760
evidence|9761,9769
of|9770,9772
right|9773,9778
heart|9779,9784
strain|9785,9791
.|9791,9792
She|9793,9796
was|9797,9800
<EOL>|9801,9802
treated|9802,9809
with|9810,9814
a|9815,9816
heparin|9817,9824
gtt|9825,9828
,|9828,9829
then|9830,9834
transitioned|9835,9847
to|9848,9850
treatment|9851,9860
dose|9861,9865
<EOL>|9866,9867
lovenox|9867,9874
given|9875,9880
malignancy|9881,9891
associated|9892,9902
thrombosis|9903,9913
as|9914,9916
noted|9917,9922
in|9923,9925
CLOT|9926,9930
<EOL>|9931,9932
trial|9932,9937
.|9937,9938
She|9939,9942
is|9943,9945
quite|9946,9951
symptomatic|9952,9963
and|9964,9967
requires|9968,9976
oxygen|9977,9983
<EOL>|9984,9985
supplementation|9985,10000
,|10000,10001
though|10002,10008
improved|10009,10017
during|10018,10024
hospitalization|10025,10040
.|10040,10041
Please|10042,10048
<EOL>|10049,10050
wean|10050,10054
oxygen|10055,10061
as|10062,10064
tolerated|10065,10074
.|10074,10075
<EOL>|10075,10076
<EOL>|10076,10077
#|10077,10078
Pulmonary|10079,10088
nodules|10089,10096
:|10096,10097
Known|10098,10103
spiculated|10104,10114
masses|10115,10121
that|10122,10126
were|10127,10131
noted|10132,10137
on|10138,10140
<EOL>|10141,10142
CT|10142,10144
in|10145,10147
_|10148,10149
_|10149,10150
_|10150,10151
,|10151,10152
concerning|10153,10163
for|10164,10167
primary|10168,10175
lung|10176,10180
malignancy|10181,10191
vs|10192,10194
mets|10195,10199
.|10199,10200
<EOL>|10201,10202
Current|10202,10209
CT|10210,10212
showed|10213,10219
stable|10220,10226
nodules|10227,10234
still|10235,10240
concerning|10241,10251
for|10252,10255
<EOL>|10256,10257
malignancy|10257,10267
.|10267,10268
She|10269,10272
was|10273,10276
evaluated|10277,10286
by|10287,10289
the|10290,10293
thoracic|10294,10302
team|10303,10307
who|10308,10311
<EOL>|10312,10313
recommended|10313,10324
CT|10325,10327
biopsy|10328,10334
vs|10335,10337
.|10337,10338
surveillance|10339,10351
.|10351,10352
Given|10353,10358
her|10359,10362
current|10363,10370
<EOL>|10371,10372
PE|10372,10374
/|10374,10375
DVT|10375,10378
,|10378,10379
the|10380,10383
family|10384,10390
and|10391,10394
the|10395,10398
patient|10399,10406
decided|10407,10414
for|10415,10418
surveillance|10419,10431
at|10432,10434
<EOL>|10435,10436
this|10436,10440
time|10441,10445
.|10445,10446
They|10447,10451
will|10452,10456
follow|10457,10463
up|10464,10466
with|10467,10471
her|10472,10475
primary|10476,10483
care|10484,10488
provider|10489,10497
.|10497,10498
<EOL>|10499,10500
<EOL>|10500,10501
#|10501,10502
Enterococcal|10503,10515
UTI|10516,10519
<EOL>|10519,10520
She|10520,10523
was|10524,10527
noted|10528,10533
to|10534,10536
have|10537,10541
rising|10542,10548
WBC|10549,10552
in|10553,10555
the|10556,10559
setting|10560,10567
of|10568,10570
UCX|10571,10574
from|10575,10579
<EOL>|10580,10581
urostomy|10581,10589
growing|10590,10597
Enterococcus|10598,10610
.|10610,10611
Given|10612,10617
her|10618,10621
rising|10622,10628
leukocytosis|10629,10641
,|10641,10642
we|10643,10645
<EOL>|10646,10647
proceeded|10647,10656
with|10657,10661
treatment|10662,10671
.|10671,10672
She|10673,10676
was|10677,10680
started|10681,10688
on|10689,10691
IV|10692,10694
Ampicillin|10695,10705
and|10706,10709
<EOL>|10710,10711
transitioned|10711,10723
to|10724,10726
macrobid|10727,10735
,|10735,10736
based|10737,10742
on|10743,10745
sensitivies|10746,10757
.|10757,10758
Leukocytosis|10759,10771
<EOL>|10772,10773
improved|10773,10781
on|10782,10784
antibiotics|10785,10796
.|10796,10797
She|10798,10801
should|10802,10808
complete|10809,10817
a|10818,10819
7|10820,10821
day|10822,10825
course|10826,10832
(|10833,10834
day|10834,10837
<EOL>|10838,10839
1|10839,10840
:|10840,10841
_|10842,10843
_|10843,10844
_|10844,10845
,|10845,10846
day|10847,10850
7|10851,10852
:|10852,10853
_|10854,10855
_|10855,10856
_|10856,10857
.|10857,10858
<EOL>|10859,10860
<EOL>|10860,10861
#|10861,10862
Normocytic|10863,10873
Anemia|10874,10880
:|10880,10881
No|10882,10884
signs|10885,10890
of|10891,10893
bleeding|10894,10902
,|10902,10903
or|10904,10906
hemolysis|10907,10916
.|10916,10917
Hb|10918,10920
<EOL>|10921,10922
dropped|10922,10929
to|10930,10932
nadir|10933,10938
of|10939,10941
7.3|10942,10945
,|10945,10946
stable|10947,10953
at|10954,10956
discharge|10957,10966
at|10967,10969
7.5|10970,10973
.|10973,10974
Iron|10975,10979
<EOL>|10980,10981
studies|10981,10988
consistent|10989,10999
with|11000,11004
likely|11005,11011
combination|11012,11023
iron|11024,11028
deficiency|11029,11039
<EOL>|11040,11041
anemia|11041,11047
and|11048,11051
anemia|11052,11058
of|11059,11061
chronic|11062,11069
disease|11070,11077
with|11078,11082
low|11083,11086
iron|11087,11091
but|11092,11095
elevated|11096,11104
<EOL>|11105,11106
ferritin|11106,11114
and|11115,11118
low|11119,11122
TIBC|11123,11127
.|11127,11128
Would|11129,11134
recommend|11135,11144
checking|11145,11153
again|11154,11159
as|11160,11162
<EOL>|11163,11164
outpatient|11164,11174
and|11175,11178
work|11179,11183
-|11183,11184
up|11184,11186
as|11187,11189
needed|11190,11196
.|11196,11197
<EOL>|11197,11198
<EOL>|11198,11199
#|11199,11200
_|11201,11202
_|11202,11203
_|11203,11204
swelling|11205,11213
:|11213,11214
Likley|11215,11221
multifactorial|11222,11236
including|11237,11246
venous|11247,11253
<EOL>|11254,11255
insufficiency|11255,11268
,|11268,11269
as|11270,11272
well|11273,11277
as|11278,11280
known|11281,11286
LLE|11287,11290
DVT|11291,11294
.|11294,11295
She|11296,11299
responded|11300,11309
quite|11310,11315
<EOL>|11316,11317
well|11317,11321
with|11322,11326
compression|11327,11338
stockings|11339,11348
.|11348,11349
<EOL>|11349,11350
<EOL>|11350,11351
#|11351,11352
Hx|11353,11355
of|11356,11358
bladder|11359,11366
cancer|11367,11373
:|11373,11374
s|11375,11376
/|11376,11377
p|11377,11378
_|11379,11380
_|11380,11381
_|11381,11382
TURBT|11383,11388
,|11388,11389
high|11390,11394
-|11394,11395
grade|11395,11400
TCC|11401,11404
,|11404,11405
T1|11406,11408
<EOL>|11409,11410
(|11410,11411
no|11411,11413
muscle|11414,11420
identified|11421,11431
)|11431,11432
.|11432,11433
Then|11434,11438
in|11439,11441
_|11442,11443
_|11443,11444
_|11444,11445
,|11445,11446
pelvic|11447,11453
MRI|11454,11457
showed|11458,11464
<EOL>|11465,11466
bladder|11466,11473
mass|11474,11478
invasion|11479,11487
,|11487,11488
perivesical|11489,11500
soft|11501,11505
tissue|11506,11512
,|11512,11513
anterior|11514,11522
vaginal|11523,11530
<EOL>|11531,11532
wall|11532,11536
on|11537,11539
right|11540,11545
(|11546,11547
C|11547,11548
/|11548,11549
W|11549,11550
T4|11551,11553
lesion|11554,11560
)|11560,11561
.|11561,11562
In|11563,11565
_|11566,11567
_|11567,11568
_|11568,11569
,|11569,11570
underwent|11571,11580
robotic|11581,11588
<EOL>|11589,11590
TAH|11590,11593
-|11593,11594
BSO|11594,11597
,|11597,11598
lap|11599,11602
radical|11603,11610
cystectomy|11611,11621
and|11622,11625
anterior|11626,11634
vaginectomy|11635,11646
with|11647,11651
<EOL>|11652,11653
pathology|11653,11662
showing|11663,11670
pT2b|11671,11675
,|11675,11676
node|11677,11681
and|11682,11685
margins|11686,11693
negative|11694,11702
.|11702,11703
No|11704,11706
plan|11707,11711
for|11712,11715
<EOL>|11716,11717
any|11717,11720
further|11721,11728
therapy|11729,11736
at|11737,11739
this|11740,11744
time|11745,11749
per|11750,11753
Dr|11754,11756
_|11757,11758
_|11758,11759
_|11759,11760
.|11760,11761
<EOL>|11761,11762
<EOL>|11762,11763
The|11763,11766
patient|11767,11774
is|11775,11777
safe|11778,11782
to|11783,11785
discharge|11786,11795
today|11796,11801
,|11801,11802
and|11803,11806
>|11807,11808
30min|11808,11813
were|11814,11818
spent|11819,11824
on|11825,11827
<EOL>|11828,11829
discharge|11829,11838
day|11839,11842
management|11843,11853
services|11854,11862
.|11862,11863
<EOL>|11863,11864
<EOL>|11864,11865
Transitional|11865,11877
issues|11878,11884
:|11884,11885
<EOL>|11885,11886
-|11886,11887
She|11888,11891
will|11892,11896
need|11897,11901
follow|11902,11908
up|11909,11911
chest|11912,11917
CT|11918,11920
for|11921,11924
pulmonary|11925,11934
nodules|11935,11942
in|11943,11945
3|11946,11947
<EOL>|11948,11949
months|11949,11955
(|11956,11957
_|11957,11958
_|11958,11959
_|11959,11960
)|11960,11961
<EOL>|11961,11962
-|11962,11963
To|11964,11966
complete|11967,11975
7|11976,11977
day|11978,11981
course|11982,11988
for|11989,11992
UTI|11993,11996
with|11997,12001
macrobid|12002,12010
(|12011,12012
day|12012,12015
7|12016,12017
:|12017,12018
_|12019,12020
_|12020,12021
_|12021,12022
<EOL>|12022,12023
-|12023,12024
Continue|12025,12033
oxygen|12034,12040
therapy|12041,12048
and|12049,12052
wean|12053,12057
as|12058,12060
tolerated|12061,12070
to|12071,12073
maintain|12074,12082
O2|12083,12085
<EOL>|12086,12087
sat|12087,12090
>|12091,12092
92|12093,12095
%|12095,12096
<EOL>|12097,12098
-|12098,12099
Please|12100,12106
check|12107,12112
CBC|12113,12116
on|12117,12119
_|12120,12121
_|12121,12122
_|12122,12123
to|12124,12126
ensure|12127,12133
stability|12134,12143
of|12144,12146
h|12147,12148
/|12148,12149
h|12149,12150
<EOL>|12151,12152
and|12152,12155
demonstrate|12156,12167
resolution|12168,12178
of|12179,12181
leukocytosis|12182,12194
<EOL>|12194,12195
-|12195,12196
HCP|12197,12200
:|12200,12201
son|12202,12205
,|12205,12206
Dr.|12207,12210
_|12211,12212
_|12212,12213
_|12213,12214
_|12215,12216
_|12216,12217
_|12217,12218
<EOL>|12218,12219
<EOL>|12219,12220
<EOL>|12221,12222
Medications|12222,12233
on|12234,12236
Admission|12237,12246
:|12246,12247
<EOL>|12247,12248
The|12248,12251
Preadmission|12252,12264
Medication|12265,12275
list|12276,12280
may|12281,12284
be|12285,12287
inaccurate|12288,12298
and|12299,12302
requires|12303,12311
<EOL>|12312,12313
futher|12313,12319
investigation|12320,12333
.|12333,12334
<EOL>|12334,12335
1.|12335,12337
Acetaminophen|12338,12351
650|12352,12355
mg|12356,12358
PO|12359,12361
Q6H|12362,12365
<EOL>|12366,12367
2.|12367,12369
Docusate|12370,12378
Sodium|12379,12385
100|12386,12389
mg|12390,12392
PO|12393,12395
BID|12396,12399
<EOL>|12400,12401
3.|12401,12403
Enoxaparin|12404,12414
Sodium|12415,12421
40|12422,12424
mg|12425,12427
SC|12428,12430
DAILY|12431,12436
<EOL>|12437,12438
Start|12438,12443
:|12443,12444
_|12445,12446
_|12446,12447
_|12447,12448
,|12448,12449
First|12450,12455
Dose|12456,12460
:|12460,12461
Next|12462,12466
Routine|12467,12474
Administration|12475,12489
Time|12490,12494
<EOL>|12495,12496
4.|12496,12498
Levothyroxine|12499,12512
Sodium|12513,12519
175|12520,12523
mcg|12524,12527
PO|12528,12530
DAILY|12531,12536
<EOL>|12537,12538
5.|12538,12540
Atorvastatin|12541,12553
10|12554,12556
mg|12557,12559
PO|12560,12562
QPM|12563,12566
<EOL>|12567,12568
6.|12568,12570
Losartan|12571,12579
Potassium|12580,12589
50|12590,12592
mg|12593,12595
PO|12596,12598
DAILY|12599,12604
<EOL>|12605,12606
7.|12606,12608
OxyCODONE|12609,12618
(|12619,12620
Immediate|12620,12629
Release|12630,12637
)|12637,12638
5|12639,12640
mg|12641,12643
PO|12644,12646
Q4H|12647,12650
:|12650,12651
PRN|12651,12654
Pain|12655,12659
-|12660,12661
Moderate|12662,12670
<EOL>|12671,12672
<EOL>|12672,12673
8.|12673,12675
LORazepam|12676,12685
0.25|12686,12690
mg|12691,12693
PO|12694,12696
BID|12697,12700
:|12700,12701
PRN|12701,12704
anxiety|12705,12712
<EOL>|12713,12714
9.|12714,12716
Senna|12717,12722
8.6|12723,12726
mg|12727,12729
PO|12730,12732
BID|12733,12736
<EOL>|12737,12738
<EOL>|12738,12739
<EOL>|12740,12741
Discharge|12741,12750
Medications|12751,12762
:|12762,12763
<EOL>|12763,12764
1.|12764,12766
Nitrofurantoin|12768,12782
Monohyd|12783,12790
(|12791,12792
MacroBID|12792,12800
)|12800,12801
100|12802,12805
mg|12806,12808
PO|12809,12811
Q12H|12812,12816
<EOL>|12817,12818
Last|12818,12822
day|12823,12826
:|12826,12827
_|12828,12829
_|12829,12830
_|12830,12831
.|12831,12832
Enoxaparin|12834,12844
Sodium|12845,12851
90|12852,12854
mg|12855,12857
SC|12858,12860
Q12H|12861,12865
<EOL>|12866,12867
Start|12867,12872
:|12872,12873
Today|12874,12879
-|12880,12881
_|12882,12883
_|12883,12884
_|12884,12885
,|12885,12886
First|12887,12892
Dose|12893,12897
:|12897,12898
Next|12899,12903
Routine|12904,12911
Administration|12912,12926
<EOL>|12927,12928
Time|12928,12932
<EOL>|12934,12935
3.|12935,12937
LORazepam|12939,12948
0.25|12949,12953
mg|12954,12956
PO|12957,12959
QHS|12960,12963
:|12963,12964
PRN|12964,12967
insomnia|12968,12976
<EOL>|12977,12978
RX|12978,12980
*|12981,12982
lorazepam|12982,12991
0.5|12992,12995
mg|12996,12998
0.5|12999,13002
(|13003,13004
One|13004,13007
half|13008,13012
)|13012,13013
tab|13014,13017
by|13018,13020
mouth|13021,13026
QHS|13027,13030
:|13030,13031
prn|13031,13034
Disp|13035,13039
<EOL>|13040,13041
#|13041,13042
*|13042,13043
3|13043,13044
Tablet|13045,13051
Refills|13052,13059
:|13059,13060
*|13060,13061
0|13061,13062
<EOL>|13063,13064
4.|13064,13066
Acetaminophen|13068,13081
650|13082,13085
mg|13086,13088
PO|13089,13091
Q6H|13092,13095
<EOL>|13097,13098
5.|13098,13100
Atorvastatin|13102,13114
10|13115,13117
mg|13118,13120
PO|13121,13123
QPM|13124,13127
<EOL>|13129,13130
6.|13130,13132
Docusate|13134,13142
Sodium|13143,13149
100|13150,13153
mg|13154,13156
PO|13157,13159
BID|13160,13163
<EOL>|13165,13166
7.|13166,13168
Levothyroxine|13170,13183
Sodium|13184,13190
175|13191,13194
mcg|13195,13198
PO|13199,13201
DAILY|13202,13207
<EOL>|13209,13210
8.|13210,13212
OxyCODONE|13214,13223
(|13224,13225
Immediate|13225,13234
Release|13235,13242
)|13242,13243
5|13244,13245
mg|13246,13248
PO|13249,13251
Q4H|13252,13255
:|13255,13256
PRN|13256,13259
Pain|13260,13264
-|13265,13266
<EOL>|13267,13268
Moderate|13268,13276
<EOL>|13277,13278
RX|13278,13280
*|13281,13282
oxycodone|13282,13291
5|13292,13293
mg|13294,13296
1|13297,13298
tablet|13299,13305
(|13305,13306
s|13306,13307
)|13307,13308
by|13309,13311
mouth|13312,13317
Q8H|13318,13321
:|13321,13322
prn|13322,13325
Disp|13326,13330
#|13331,13332
*|13332,13333
3|13333,13334
Tablet|13335,13341
<EOL>|13342,13343
Refills|13343,13350
:|13350,13351
*|13351,13352
0|13352,13353
<EOL>|13354,13355
9.|13355,13357
Senna|13359,13364
8.6|13365,13368
mg|13369,13371
PO|13372,13374
BID|13375,13378
<EOL>|13380,13381
<EOL>|13381,13382
<EOL>|13383,13384
Discharge|13384,13393
Disposition|13394,13405
:|13405,13406
<EOL>|13406,13407
Extended|13407,13415
Care|13416,13420
<EOL>|13420,13421
<EOL>|13422,13423
Facility|13423,13431
:|13431,13432
<EOL>|13432,13433
_|13433,13434
_|13434,13435
_|13435,13436
<EOL>|13436,13437
<EOL>|13438,13439
Discharge|13439,13448
Diagnosis|13449,13458
:|13458,13459
<EOL>|13459,13460
PE|13460,13462
<EOL>|13462,13463
<EOL>|13464,13465
Mental|13486,13492
Status|13493,13499
:|13499,13500
Clear|13501,13506
and|13507,13510
coherent|13511,13519
.|13519,13520
<EOL>|13520,13521
Level|13521,13526
of|13527,13529
Consciousness|13530,13543
:|13543,13544
Alert|13545,13550
and|13551,13554
interactive|13555,13566
.|13566,13567
<EOL>|13567,13568
Activity|13568,13576
Status|13577,13583
:|13583,13584
Out|13585,13588
of|13589,13591
Bed|13592,13595
with|13596,13600
assistance|13601,13611
to|13612,13614
chair|13615,13620
or|13621,13623
<EOL>|13624,13625
wheelchair|13625,13635
.|13635,13636
<EOL>|13636,13637
<EOL>|13637,13638
<EOL>|13639,13640
Ms.|13664,13667
_|13668,13669
_|13669,13670
_|13670,13671
it|13672,13674
was|13675,13678
a|13679,13680
pleasure|13681,13689
taking|13690,13696
care|13697,13701
you|13702,13705
during|13706,13712
your|13713,13717
<EOL>|13718,13719
admission|13719,13728
to|13729,13731
_|13732,13733
_|13733,13734
_|13734,13735
.|13735,13736
You|13737,13740
were|13741,13745
admitted|13746,13754
for|13755,13758
a|13759,13760
clot|13761,13765
in|13766,13768
your|13769,13773
lungs|13774,13779
<EOL>|13780,13781
and|13781,13784
leg|13785,13788
.|13788,13789
You|13790,13793
were|13794,13798
treated|13799,13806
with|13807,13811
a|13812,13813
blood|13814,13819
thinner|13820,13827
.|13827,13828
You|13829,13832
will|13833,13837
need|13838,13842
to|13843,13845
<EOL>|13846,13847
continue|13847,13855
the|13856,13859
blood|13860,13865
thinner|13866,13873
.|13873,13874
You|13875,13878
were|13879,13883
also|13884,13888
treated|13889,13896
for|13897,13900
a|13901,13902
urinary|13903,13910
<EOL>|13911,13912
tract|13912,13917
infection|13918,13927
.|13927,13928
For|13929,13932
your|13933,13937
pulmonary|13938,13947
nodules|13948,13955
,|13955,13956
you|13957,13960
should|13961,13967
follow|13968,13974
<EOL>|13975,13976
up|13976,13978
with|13979,13983
your|13984,13988
primary|13989,13996
care|13997,14001
doctor|14002,14008
.|14008,14009
<EOL>|14010,14011
<EOL>|14012,14013
Followup|14013,14021
Instructions|14022,14034
:|14034,14035
<EOL>|14035,14036
_|14036,14037
_|14037,14038
_|14038,14039
<EOL>|14039,14040

