 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|42,51|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|42,51|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|42,56|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|76,85|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|76,85|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|76,85|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|76,85|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|76,85|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|76,90|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|108,113|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|108,113|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|108,113|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|132,135|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|143,150|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|143,150|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|152,160|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|SIMPLE_SEGMENT|163,172|false|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|163,172|false|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|163,172|false|false|false|C0020517|Hypersensitivity|Allergies
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|178,181|false|false|false|C0013343|Dyes|Dye
Event|Event|SIMPLE_SEGMENT|178,181|false|false|false|||Dye
Drug|Biologically Active Substance|SIMPLE_SEGMENT|183,189|false|false|false|C0021968;C0885449|Iodine, Homeopathic preparation;iodine|Iodine
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|183,189|false|false|false|C0021968;C0885449|Iodine, Homeopathic preparation;iodine|Iodine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|183,189|false|false|false|C0021968;C0885449|Iodine, Homeopathic preparation;iodine|Iodine
Event|Activity|SIMPLE_SEGMENT|190,200|false|false|false|C2700400|Contain (action)|Containing
Finding|Functional Concept|SIMPLE_SEGMENT|190,200|false|false|false|C0332256|Containing (qualifier value)|Containing
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|201,209|false|false|false|C0009924|Contrast Media|Contrast
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|201,215|false|false|false|C0009924|Contrast Media|Contrast Media
Anatomy|Tissue|SIMPLE_SEGMENT|210,215|false|false|false|C0162867;C1254021|Media layer;Tunica Media|Media
Finding|Intellectual Product|SIMPLE_SEGMENT|210,215|false|false|false|C0009458;C0677540|Communications Media;PAMS Media|Media
Drug|Organic Chemical|SIMPLE_SEGMENT|218,227|false|false|false|C0030049|oxycodone|Oxycodone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|218,227|false|false|false|C0030049|oxycodone|Oxycodone
Event|Event|SIMPLE_SEGMENT|218,227|false|false|false|||Oxycodone
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|218,227|false|false|false|C0524222|Oxycodone measurement|Oxycodone
Drug|Organic Chemical|SIMPLE_SEGMENT|231,241|false|false|false|C0055729|cilostazol|cilostazol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|231,241|false|false|false|C0055729|cilostazol|cilostazol
Event|Event|SIMPLE_SEGMENT|231,241|false|false|false|||cilostazol
Drug|Organic Chemical|SIMPLE_SEGMENT|244,255|false|false|false|C1569608|varenicline|Varenicline
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|244,255|false|false|false|C1569608|varenicline|Varenicline
Event|Event|SIMPLE_SEGMENT|244,255|false|false|false|||Varenicline
Event|Event|SIMPLE_SEGMENT|258,267|false|false|false|||Attending
Finding|Functional Concept|SIMPLE_SEGMENT|258,267|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|SIMPLE_SEGMENT|276,291|false|false|false|C0277786|Chief complaint (finding)|Chief Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|282,291|false|false|false|C3864418||Complaint
Event|Event|SIMPLE_SEGMENT|282,291|false|false|false|||Complaint
Finding|Finding|SIMPLE_SEGMENT|282,291|false|false|false|C5441521|Complaint (finding)|Complaint
Event|Event|SIMPLE_SEGMENT|293,302|false|false|false|||Shortness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|293,312|false|false|false|C2707305||Shortness of breath
Finding|Sign or Symptom|SIMPLE_SEGMENT|293,312|false|false|false|C0013404|Dyspnea|Shortness of breath
Finding|Body Substance|SIMPLE_SEGMENT|306,312|false|false|false|C0225386|Breath|breath
Finding|Classification|SIMPLE_SEGMENT|315,320|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|SIMPLE_SEGMENT|321,329|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|321,329|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|333,351|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|342,351|false|false|false|C0945766||Procedure
Event|Event|SIMPLE_SEGMENT|342,351|false|false|false|||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|342,351|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|342,351|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|342,351|false|false|false|C0184661|Interventional procedure|Procedure
Event|Event|SIMPLE_SEGMENT|361,368|true|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|361,368|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|361,368|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|361,368|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|361,371|true|false|false|C0262926|Medical History|History of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|361,387|true|false|false|C0488508||History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|361,387|true|false|false|C0262512|History of present illness (finding)|History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|372,379|true|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Idea or Concept|SIMPLE_SEGMENT|372,379|true|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Finding|SIMPLE_SEGMENT|372,387|true|false|false|C4264312|Present illness|Present Illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|380,387|true|false|false|C0221423|Illness (finding)|Illness
Event|Event|SIMPLE_SEGMENT|422,425|false|false|false|||PMH
Finding|Finding|SIMPLE_SEGMENT|422,425|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|PMH
Event|Event|SIMPLE_SEGMENT|426,433|false|false|false|||notable
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|438,442|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|438,442|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|SIMPLE_SEGMENT|438,442|false|false|false|||COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|438,442|false|false|false|C1412502|ARCN1 gene|COPD
Finding|Idea or Concept|SIMPLE_SEGMENT|447,451|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|447,451|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|447,451|false|false|false|C1553498|home health encounter|home
Event|Event|SIMPLE_SEGMENT|455,467|false|false|false|||hospitalized
Event|Event|SIMPLE_SEGMENT|492,498|false|false|false|||visits
Finding|Social Behavior|SIMPLE_SEGMENT|492,498|false|false|false|C0545082|Visit|visits
Procedure|Health Care Activity|SIMPLE_SEGMENT|492,498|false|false|false|C1512346|Patient Visit|visits
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|501,505|false|false|false|C0004238|Atrial Fibrillation|Afib
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|501,505|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Afib
Drug|Organic Chemical|SIMPLE_SEGMENT|510,518|false|false|false|C1831808|apixaban|apixaban
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|510,518|false|false|false|C1831808|apixaban|apixaban
Event|Event|SIMPLE_SEGMENT|510,518|false|false|false|||apixaban
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|520,523|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|SIMPLE_SEGMENT|520,523|false|false|false|||HTN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|525,528|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|525,528|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|525,528|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|525,528|false|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|525,528|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|525,528|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|525,528|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|525,528|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Event|Event|SIMPLE_SEGMENT|534,537|false|false|false|||HLD
Event|Event|SIMPLE_SEGMENT|542,550|false|false|false|||presents
Finding|Finding|SIMPLE_SEGMENT|556,568|false|false|false|C3845714|Several days|several days
Event|Event|SIMPLE_SEGMENT|573,582|false|false|false|||worsening
Event|Event|SIMPLE_SEGMENT|583,590|false|false|false|||dyspnea
Finding|Finding|SIMPLE_SEGMENT|583,590|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|583,590|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Body Substance|SIMPLE_SEGMENT|593,600|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|593,600|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|593,600|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Functional Concept|SIMPLE_SEGMENT|593,604|false|false|false|C0332310|Has patient|Patient has
Event|Event|SIMPLE_SEGMENT|620,626|false|false|false|||visits
Finding|Social Behavior|SIMPLE_SEGMENT|620,626|false|false|false|C0545082|Visit|visits
Procedure|Health Care Activity|SIMPLE_SEGMENT|620,626|false|false|false|C1512346|Patient Visit|visits
Event|Event|SIMPLE_SEGMENT|631,638|false|false|false|||dyspnea
Finding|Finding|SIMPLE_SEGMENT|631,638|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|631,638|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Event|Event|SIMPLE_SEGMENT|653,668|false|false|false|||hospitalization
Procedure|Health Care Activity|SIMPLE_SEGMENT|653,668|false|false|false|C0019993|Hospitalization|hospitalization
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|675,679|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|675,679|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|SIMPLE_SEGMENT|675,679|false|false|false|||COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|675,679|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|675,692|false|false|false|C0740304|COPD exacerbation|COPD exacerbation
Event|Event|SIMPLE_SEGMENT|680,692|false|false|false|||exacerbation
Finding|Finding|SIMPLE_SEGMENT|680,692|false|false|false|C4086268|Exacerbation|exacerbation
Drug|Organic Chemical|SIMPLE_SEGMENT|718,725|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|718,725|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|718,733|false|false|false|C0149783|Steroid therapy|steroid therapy
Event|Event|SIMPLE_SEGMENT|726,733|false|false|false|||therapy
Finding|Finding|SIMPLE_SEGMENT|726,733|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|SIMPLE_SEGMENT|726,733|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|726,733|false|false|false|C0087111|Therapeutic procedure|therapy
Event|Event|SIMPLE_SEGMENT|747,755|false|false|false|||attempts
Event|Event|SIMPLE_SEGMENT|759,764|false|false|false|||taper
Procedure|Health Care Activity|SIMPLE_SEGMENT|759,764|false|false|false|C0441640||taper
Event|Event|SIMPLE_SEGMENT|821,826|false|false|false|||visit
Finding|Social Behavior|SIMPLE_SEGMENT|821,826|false|false|false|C0545082|Visit|visit
Event|Event|SIMPLE_SEGMENT|846,852|false|false|false|||placed
Drug|Hormone|SIMPLE_SEGMENT|865,875|false|false|false|C0032952|prednisone|prednisone
Drug|Organic Chemical|SIMPLE_SEGMENT|865,875|false|false|false|C0032952|prednisone|prednisone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|865,875|false|false|false|C0032952|prednisone|prednisone
Event|Event|SIMPLE_SEGMENT|865,875|false|false|false|||prednisone
Event|Event|SIMPLE_SEGMENT|883,888|false|false|false|||taper
Procedure|Health Care Activity|SIMPLE_SEGMENT|883,888|false|false|false|C0441640||taper
Finding|Idea or Concept|SIMPLE_SEGMENT|909,912|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|909,912|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|918,921|false|false|false|||SOB
Finding|Sign or Symptom|SIMPLE_SEGMENT|918,921|false|false|false|C0013404|Dyspnea|SOB
Event|Event|SIMPLE_SEGMENT|922,930|false|false|false|||worsened
Event|Event|SIMPLE_SEGMENT|940,945|false|false|false|||taper
Procedure|Health Care Activity|SIMPLE_SEGMENT|940,945|false|false|false|C0441640||taper
Event|Event|SIMPLE_SEGMENT|958,962|false|false|false|||seen
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|978,981|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|978,981|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|978,981|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|978,981|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|SIMPLE_SEGMENT|978,981|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|978,981|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|SIMPLE_SEGMENT|978,981|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|978,981|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|SIMPLE_SEGMENT|978,981|false|false|false|||PCP
Finding|Gene or Genome|SIMPLE_SEGMENT|978,981|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|SIMPLE_SEGMENT|978,981|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Event|SIMPLE_SEGMENT|986,993|false|false|false|||started
Event|Event|SIMPLE_SEGMENT|1003,1009|false|false|false|||course
Drug|Hormone|SIMPLE_SEGMENT|1013,1023|false|false|false|C0032952|prednisone|prednisone
Drug|Organic Chemical|SIMPLE_SEGMENT|1013,1023|false|false|false|C0032952|prednisone|prednisone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1013,1023|false|false|false|C0032952|prednisone|prednisone
Event|Event|SIMPLE_SEGMENT|1013,1023|false|false|false|||prednisone
Event|Event|SIMPLE_SEGMENT|1040,1047|false|false|false|||tapered
Procedure|Health Care Activity|SIMPLE_SEGMENT|1084,1089|false|false|false|C0441640||taper
Drug|Hormone|SIMPLE_SEGMENT|1111,1121|false|false|false|C0032952|prednisone|prednisone
Drug|Organic Chemical|SIMPLE_SEGMENT|1111,1121|false|false|false|C0032952|prednisone|prednisone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1111,1121|false|false|false|C0032952|prednisone|prednisone
Event|Event|SIMPLE_SEGMENT|1111,1121|false|false|false|||prednisone
Event|Event|SIMPLE_SEGMENT|1137,1144|false|false|false|||reports
Event|Event|SIMPLE_SEGMENT|1154,1157|false|false|false|||SOB
Finding|Sign or Symptom|SIMPLE_SEGMENT|1154,1157|false|false|false|C0013404|Dyspnea|SOB
Event|Event|SIMPLE_SEGMENT|1158,1166|false|false|false|||improved
Event|Event|SIMPLE_SEGMENT|1182,1190|false|false|false|||starting
Drug|Organic Chemical|SIMPLE_SEGMENT|1196,1204|false|false|false|C0038317|Steroids|steroids
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1196,1204|false|false|false|C0038317|Steroids|steroids
Event|Event|SIMPLE_SEGMENT|1196,1204|false|false|false|||steroids
Event|Event|SIMPLE_SEGMENT|1244,1252|false|false|false|||worsened
Event|Event|SIMPLE_SEGMENT|1266,1272|false|false|false|||unable
Finding|Finding|SIMPLE_SEGMENT|1266,1272|false|false|false|C1299582|Unable|unable
Finding|Finding|SIMPLE_SEGMENT|1266,1281|false|false|false|C0424565|Cannot sleep at all|unable to sleep
Drug|Organic Chemical|SIMPLE_SEGMENT|1276,1281|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1276,1281|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Event|Event|SIMPLE_SEGMENT|1276,1281|false|false|false|||sleep
Finding|Organism Function|SIMPLE_SEGMENT|1276,1281|false|false|false|C0037313|Sleep|sleep
Finding|Finding|SIMPLE_SEGMENT|1287,1294|false|false|false|C3888388|Usually|usually
Event|Event|SIMPLE_SEGMENT|1302,1309|false|false|false|||pillows
Drug|Organic Chemical|SIMPLE_SEGMENT|1313,1318|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1313,1318|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Event|Event|SIMPLE_SEGMENT|1313,1318|false|false|false|||sleep
Finding|Organism Function|SIMPLE_SEGMENT|1313,1318|false|false|false|C0037313|Sleep|sleep
Event|Event|SIMPLE_SEGMENT|1333,1344|false|false|false|||comfortable
Finding|Finding|SIMPLE_SEGMENT|1333,1344|false|false|false|C5546696|Feeling comfortable|comfortable
Finding|Intellectual Product|SIMPLE_SEGMENT|1352,1359|false|false|false|C1550127|Special Handling Code - Upright|upright
Phenomenon|Human-caused Phenomenon or Process|SIMPLE_SEGMENT|1352,1359|false|false|false|C1550585|Entity Handling - upright|upright
Event|Event|SIMPLE_SEGMENT|1390,1399|false|false|false|||increased
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1404,1410|false|false|false|C0030054|oxygen|oxygen
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|1404,1410|false|false|false|C0030054|oxygen|oxygen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1404,1410|false|false|false|C0030054|oxygen|oxygen
Event|Event|SIMPLE_SEGMENT|1404,1410|false|false|false|||oxygen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1404,1410|false|false|false|C0184633|Oxygen Therapy Care|oxygen
Event|Event|SIMPLE_SEGMENT|1421,1425|false|false|false|||felt
Event|Event|SIMPLE_SEGMENT|1426,1432|false|false|false|||better
Finding|Idea or Concept|SIMPLE_SEGMENT|1426,1432|false|false|false|C1550462|Observation Interpretation - better|better
Finding|Finding|SIMPLE_SEGMENT|1441,1448|false|false|false|C3888388|Usually|usually
Finding|Finding|SIMPLE_SEGMENT|1459,1466|false|false|false|C4534363|At home|at home
Event|Event|SIMPLE_SEGMENT|1462,1466|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|1462,1466|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|1462,1466|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|1462,1466|false|false|false|C1553498|home health encounter|home
Event|Event|SIMPLE_SEGMENT|1472,1479|false|false|false|||reports
Event|Event|SIMPLE_SEGMENT|1527,1532|false|false|false|||using
Drug|Organic Chemical|SIMPLE_SEGMENT|1547,1556|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1547,1556|false|false|false|C0001927|albuterol|albuterol
Event|Event|SIMPLE_SEGMENT|1557,1565|false|false|false|||inhalers
Event|Event|SIMPLE_SEGMENT|1582,1587|false|false|false|||hours
Event|Event|SIMPLE_SEGMENT|1593,1598|false|false|false|||knows
Event|Event|SIMPLE_SEGMENT|1631,1641|false|false|false|||prescribed
Event|Event|SIMPLE_SEGMENT|1654,1659|false|false|false|||makes
Event|Event|SIMPLE_SEGMENT|1664,1675|false|false|false|||comfortable
Finding|Finding|SIMPLE_SEGMENT|1664,1675|false|false|false|C5546696|Feeling comfortable|comfortable
Finding|Idea or Concept|SIMPLE_SEGMENT|1681,1687|false|false|false|C0750554|MOSTLY|mostly
Event|Event|SIMPLE_SEGMENT|1688,1693|false|false|false|||stays
Event|Event|SIMPLE_SEGMENT|1705,1711|false|false|false|||second
Finding|Functional Concept|SIMPLE_SEGMENT|1705,1711|false|false|false|C1522484;C1561503;C1705190|Precision - second;Second Suffix;metastatic qualifier|second
Finding|Idea or Concept|SIMPLE_SEGMENT|1705,1711|false|false|false|C1522484;C1561503;C1705190|Precision - second;Second Suffix;metastatic qualifier|second
Finding|Intellectual Product|SIMPLE_SEGMENT|1705,1711|false|false|false|C1522484;C1561503;C1705190|Precision - second;Second Suffix;metastatic qualifier|second
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|1713,1718|false|false|false|C3714591|Floor (anatomic)|floor
Event|Event|SIMPLE_SEGMENT|1726,1730|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|1726,1730|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|1726,1730|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|1726,1730|false|false|false|C1553498|home health encounter|home
Event|Event|SIMPLE_SEGMENT|1736,1742|false|false|false|||states
Event|Event|SIMPLE_SEGMENT|1756,1760|true|false|false|||walk
Event|Event|SIMPLE_SEGMENT|1792,1797|true|false|false|||short
Finding|Sign or Symptom|SIMPLE_SEGMENT|1792,1807|true|false|false|C0013404|Dyspnea|short of breath
Finding|Body Substance|SIMPLE_SEGMENT|1801,1807|true|false|false|C0225386|Breath|breath
Event|Event|SIMPLE_SEGMENT|1822,1825|true|false|false|||use
Event|Event|SIMPLE_SEGMENT|1830,1836|true|false|false|||stairs
Finding|Finding|SIMPLE_SEGMENT|1830,1836|true|true|false|C4300351|Prior functioning.stairs|stairs
Event|Event|SIMPLE_SEGMENT|1856,1861|false|false|false|||leave
Event|Event|SIMPLE_SEGMENT|1883,1890|false|false|false|||worsens
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1896,1905|false|false|false|C5885990||breathing
Event|Event|SIMPLE_SEGMENT|1896,1905|false|false|false|||breathing
Finding|Finding|SIMPLE_SEGMENT|1896,1905|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|SIMPLE_SEGMENT|1896,1905|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|SIMPLE_SEGMENT|1896,1905|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|SIMPLE_SEGMENT|1896,1905|false|false|false|C1160636|respiratory system process|breathing
Event|Event|SIMPLE_SEGMENT|1911,1919|false|false|false|||endorses
Drug|Organic Chemical|SIMPLE_SEGMENT|1922,1927|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1922,1927|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|SIMPLE_SEGMENT|1922,1927|false|false|false|||cough
Finding|Sign or Symptom|SIMPLE_SEGMENT|1922,1927|false|false|false|C0010200|Coughing|cough
Event|Event|SIMPLE_SEGMENT|1941,1951|false|false|false|||productive
Event|Event|SIMPLE_SEGMENT|1960,1966|false|false|false|||sputum
Finding|Body Substance|SIMPLE_SEGMENT|1960,1966|false|false|false|C0038056;C1546789;C1576419|Specimen Type - Sputum;Sputum|sputum
Finding|Intellectual Product|SIMPLE_SEGMENT|1960,1966|false|false|false|C0038056;C1546789;C1576419|Specimen Type - Sputum;Sputum|sputum
Event|Event|SIMPLE_SEGMENT|1976,1986|false|false|false|||consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|1976,1986|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|1976,1991|false|false|false|C0332290|Consistent with|consistent with
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|1996,2004|false|true|false|C0168634|BaseLine dental cement|baseline
Event|Event|SIMPLE_SEGMENT|1996,2004|false|false|false|||baseline
Finding|Idea or Concept|SIMPLE_SEGMENT|1996,2004|false|true|false|C1552824|baseline - TableCellVerticalAlign|baseline
Event|Event|SIMPLE_SEGMENT|2010,2018|false|false|false|||endorses
Event|Event|SIMPLE_SEGMENT|2024,2031|false|false|false|||episode
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2050,2055|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|2050,2055|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2050,2060|false|true|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|2050,2060|false|true|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2056,2060|false|true|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|2056,2060|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|2056,2060|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|2056,2060|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|2087,2095|false|false|false|||resolved
Event|Event|SIMPLE_SEGMENT|2101,2107|false|false|false|||denies
Event|Event|SIMPLE_SEGMENT|2108,2113|true|false|false|||fever
Finding|Finding|SIMPLE_SEGMENT|2108,2113|true|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|2108,2113|true|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Event|Event|SIMPLE_SEGMENT|2115,2121|true|false|false|||chills
Finding|Sign or Symptom|SIMPLE_SEGMENT|2115,2121|true|false|false|C0085593|Chills|chills
Finding|Sign or Symptom|SIMPLE_SEGMENT|2130,2134|true|false|false|C0221423|Illness (finding)|sick
Event|Event|SIMPLE_SEGMENT|2135,2143|true|false|false|||contacts
Procedure|Health Care Activity|SIMPLE_SEGMENT|2135,2143|true|false|false|C4036459|Contacts|contacts
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2150,2155|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|2150,2155|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2150,2165|false|false|false|C0023216|Lower Extremity|lower extremity
Finding|Pathologic Function|SIMPLE_SEGMENT|2150,2171|false|false|false|C0239340|Edema of lower extremity|lower extremity edema
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2156,2165|false|false|false|C0015385|Limb structure|extremity
Finding|Pathologic Function|SIMPLE_SEGMENT|2156,2171|false|false|false|C0085649|Peripheral edema|extremity edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2166,2171|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|2166,2171|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|2166,2171|false|false|false|C0013604|Edema|edema
Finding|Idea or Concept|SIMPLE_SEGMENT|2185,2192|false|false|false|C1555582|Initial (abbreviation)|initial
Drug|Food|SIMPLE_SEGMENT|2193,2198|false|false|false|C1875856|Vital High Nitrogen Enteral Nutrition|vital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2193,2204|false|false|false|C0488614;C0518766|Vital signs|vital signs
Procedure|Health Care Activity|SIMPLE_SEGMENT|2193,2204|false|false|false|C0150404|Taking vital signs|vital signs
Event|Event|SIMPLE_SEGMENT|2199,2204|false|false|false|||signs
Finding|Finding|SIMPLE_SEGMENT|2199,2204|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|SIMPLE_SEGMENT|2199,2204|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Event|Event|SIMPLE_SEGMENT|2223,2225|false|false|false|||BP
Event|Event|SIMPLE_SEGMENT|2258,2262|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|2258,2262|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2258,2262|false|false|false|C0582103|Medical Examination|Exam
Event|Event|SIMPLE_SEGMENT|2263,2270|false|false|false|||notable
Finding|Organism Function|SIMPLE_SEGMENT|2284,2294|false|false|false|C0231800|Expiration, Respiratory|expiratory
Finding|Sign or Symptom|SIMPLE_SEGMENT|2284,2303|false|false|false|C0231875|Expiratory wheezing|expiratory wheezing
Event|Event|SIMPLE_SEGMENT|2295,2303|false|false|false|||wheezing
Finding|Sign or Symptom|SIMPLE_SEGMENT|2295,2303|false|false|false|C0043144|Wheezing|wheezing
Event|Event|SIMPLE_SEGMENT|2305,2314|false|false|false|||prolonged
Finding|Organism Function|SIMPLE_SEGMENT|2316,2326|false|false|false|C0231800|Expiration, Respiratory|expiratory
Event|Event|SIMPLE_SEGMENT|2327,2332|false|false|false|||phase
Finding|Functional Concept|SIMPLE_SEGMENT|2334,2338|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Finding|Organism Function|SIMPLE_SEGMENT|2339,2350|false|false|false|C0004048|Inspiration (function)|inspiratory
Finding|Finding|SIMPLE_SEGMENT|2339,2359|false|false|false|C0577961|Inspiratory crackles|inspiratory crackles
Event|Event|SIMPLE_SEGMENT|2351,2359|false|false|false|||crackles
Finding|Finding|SIMPLE_SEGMENT|2351,2359|false|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Event|Event|SIMPLE_SEGMENT|2384,2390|false|false|false|||rhthym
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2400,2405|false|false|false|C0016504;C0687080|Foot;Paw|pedal
Finding|Pathologic Function|SIMPLE_SEGMENT|2400,2411|false|false|false|C0239340;C0574002;C5700071|Edema of foot (finding);Edema of lower extremity;Foot swelling|pedal edema
Finding|Sign or Symptom|SIMPLE_SEGMENT|2400,2411|false|false|false|C0239340;C0574002;C5700071|Edema of foot (finding);Edema of lower extremity;Foot swelling|pedal edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2406,2411|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|2406,2411|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|2406,2411|false|false|false|C0013604|Edema|edema
Event|Event|SIMPLE_SEGMENT|2416,2420|false|false|false|||Labs
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2416,2420|false|false|false|C0587081|Laboratory test finding|Labs
Event|Event|SIMPLE_SEGMENT|2426,2433|false|false|false|||notable
Anatomy|Cell Component|SIMPLE_SEGMENT|2438,2441|false|false|false|C2263086|Nuclear cap binding complex location|CBC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2438,2441|false|false|false|C0009555|Complete Blood Count|CBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2447,2453|false|false|false|C5574646|Natriuretic Peptides B, human|proBNP
Drug|Hormone|SIMPLE_SEGMENT|2447,2453|false|false|false|C5574646|Natriuretic Peptides B, human|proBNP
Event|Event|SIMPLE_SEGMENT|2447,2453|false|false|false|||proBNP
Event|Event|SIMPLE_SEGMENT|2470,2474|false|false|false|||chem
Finding|Functional Concept|SIMPLE_SEGMENT|2470,2474|false|false|false|C0079107|chemical aspects|chem
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2470,2474|false|false|false|C0201682|Chemical procedure|chem
Event|Event|SIMPLE_SEGMENT|2476,2483|false|false|false|||notable
Drug|Organic Chemical|SIMPLE_SEGMENT|2488,2494|false|false|false|C0074722|sodium bicarbonate|bicarb
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2488,2494|false|false|false|C0074722|sodium bicarbonate|bicarb
Event|Event|SIMPLE_SEGMENT|2488,2494|false|false|false|||bicarb
Anatomy|Cell|SIMPLE_SEGMENT|2524,2528|false|false|false|C0014792|Erythrocytes|RBCs
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2524,2528|false|false|false|C0014792|Erythrocytes|RBCs
Event|Event|SIMPLE_SEGMENT|2533,2540|false|false|false|||Studies
Procedure|Research Activity|SIMPLE_SEGMENT|2533,2540|false|false|false|C0947630|Scientific Study|Studies
Event|Event|SIMPLE_SEGMENT|2559,2562|false|false|false|||CXR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2559,2562|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|SIMPLE_SEGMENT|2568,2574|false|false|false|||stable
Finding|Intellectual Product|SIMPLE_SEGMENT|2568,2574|false|false|false|C1547311|Patient Condition Code - Stable|stable
Finding|Intellectual Product|SIMPLE_SEGMENT|2575,2579|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Finding|SIMPLE_SEGMENT|2580,2588|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|SIMPLE_SEGMENT|2580,2588|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Event|Event|SIMPLE_SEGMENT|2590,2602|false|false|false|||cardiomegaly
Finding|Finding|SIMPLE_SEGMENT|2590,2602|false|false|false|C0018800|Cardiomegaly|cardiomegaly
Event|Event|SIMPLE_SEGMENT|2604,2615|false|false|false|||atelectasis
Finding|Pathologic Function|SIMPLE_SEGMENT|2604,2615|false|false|false|C0004144|Atelectasis|atelectasis
Drug|Chemical Viewed Functionally|SIMPLE_SEGMENT|2619,2624|false|false|false|C0178499|Base|bases
Finding|Idea or Concept|SIMPLE_SEGMENT|2636,2641|false|false|false|C1550016|Remote control command - Clear|clear
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2642,2646|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2642,2646|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2642,2646|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|SIMPLE_SEGMENT|2642,2646|false|false|false|C0740941|Lung Problem|lung
Event|Event|SIMPLE_SEGMENT|2647,2653|false|false|false|||fields
Finding|Body Substance|SIMPLE_SEGMENT|2656,2663|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|2656,2663|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|2656,2663|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|2668,2673|false|false|false|||given
Drug|Organic Chemical|SIMPLE_SEGMENT|2674,2683|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2674,2683|false|false|false|C0001927|albuterol|Albuterol
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2684,2687|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|neb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2684,2687|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|neb
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|2684,2687|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|neb
Event|Event|SIMPLE_SEGMENT|2684,2687|false|false|false|||neb
Finding|Cell Function|SIMPLE_SEGMENT|2684,2687|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|neb
Finding|Gene or Genome|SIMPLE_SEGMENT|2684,2687|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|neb
Drug|Organic Chemical|SIMPLE_SEGMENT|2693,2704|false|false|false|C0027235|ipratropium|ipratropium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2693,2704|false|false|false|C0027235|ipratropium|ipratropium
Event|Event|SIMPLE_SEGMENT|2693,2704|false|false|false|||ipratropium
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2705,2708|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|neb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2705,2708|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|neb
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|2705,2708|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|neb
Event|Event|SIMPLE_SEGMENT|2705,2708|false|false|false|||neb
Finding|Cell Function|SIMPLE_SEGMENT|2705,2708|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|neb
Finding|Gene or Genome|SIMPLE_SEGMENT|2705,2708|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|neb
Drug|Antibiotic|SIMPLE_SEGMENT|2715,2727|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|Azithromycin
Drug|Clinical Drug|SIMPLE_SEGMENT|2715,2727|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|Azithromycin
Drug|Organic Chemical|SIMPLE_SEGMENT|2715,2727|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|Azithromycin
Drug|Hormone|SIMPLE_SEGMENT|2739,2749|false|false|false|C0032952|prednisone|Prednisone
Drug|Organic Chemical|SIMPLE_SEGMENT|2739,2749|false|false|false|C0032952|prednisone|Prednisone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2739,2749|false|false|false|C0032952|prednisone|Prednisone
Event|Activity|SIMPLE_SEGMENT|2765,2772|false|false|false|C1706079||arrival
Event|Event|SIMPLE_SEGMENT|2765,2772|false|false|false|||arrival
Finding|Functional Concept|SIMPLE_SEGMENT|2765,2772|false|false|false|C1555577|arrival - ActRelationshipType|arrival
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|2780,2785|false|false|false|C3714591|Floor (anatomic)|floor
Finding|Body Substance|SIMPLE_SEGMENT|2791,2798|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|2791,2798|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|2791,2798|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|2799,2805|false|false|false|||states
Event|Event|SIMPLE_SEGMENT|2825,2829|false|false|false|||well
Finding|Finding|SIMPLE_SEGMENT|2825,2829|false|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|2835,2839|false|false|false|||says
Event|Event|SIMPLE_SEGMENT|2849,2852|false|false|false|||SOB
Finding|Sign or Symptom|SIMPLE_SEGMENT|2849,2852|false|false|false|C0013404|Dyspnea|SOB
Event|Event|SIMPLE_SEGMENT|2857,2865|false|false|false|||improved
Event|Event|SIMPLE_SEGMENT|2893,2899|false|false|false|||better
Finding|Idea or Concept|SIMPLE_SEGMENT|2893,2899|false|false|false|C1550462|Observation Interpretation - better|better
Event|Event|SIMPLE_SEGMENT|2935,2940|true|false|false|||sleep
Event|Event|SIMPLE_SEGMENT|2946,2952|false|false|false|||Review
Finding|Idea or Concept|SIMPLE_SEGMENT|2946,2952|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|Review
Finding|Intellectual Product|SIMPLE_SEGMENT|2946,2952|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|Review
Finding|Functional Concept|SIMPLE_SEGMENT|2946,2955|false|false|false|C0699752|Review of|Review of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2946,2963|false|false|false|C0488564;C0488565||Review of Systems
Procedure|Health Care Activity|SIMPLE_SEGMENT|2946,2963|false|false|false|C0489633|Review of systems (procedure)|Review of Systems
Event|Event|SIMPLE_SEGMENT|2956,2963|false|false|false|||Systems
Finding|Functional Concept|SIMPLE_SEGMENT|2956,2963|false|false|false|C0449913|System|Systems
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2976,2979|false|false|false|C0268529|Proline dehydrogenase deficiency|HPI
Event|Event|SIMPLE_SEGMENT|2976,2979|false|false|false|||HPI
Finding|Finding|SIMPLE_SEGMENT|2976,2979|false|false|false|C0262512;C1323983|History of present illness (finding);allene oxide synthase activity|HPI
Finding|Molecular Function|SIMPLE_SEGMENT|2976,2979|false|false|false|C0262512;C1323983|History of present illness (finding);allene oxide synthase activity|HPI
Event|Event|SIMPLE_SEGMENT|2987,2992|false|false|false|||fever
Finding|Finding|SIMPLE_SEGMENT|2987,2992|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|2987,2992|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Event|Event|SIMPLE_SEGMENT|2994,3000|false|false|false|||chills
Finding|Sign or Symptom|SIMPLE_SEGMENT|2994,3000|false|false|false|C0085593|Chills|chills
Finding|Sign or Symptom|SIMPLE_SEGMENT|3002,3014|false|false|false|C0028081|Night sweats|night sweats
Event|Event|SIMPLE_SEGMENT|3008,3014|false|false|false|||sweats
Finding|Body Substance|SIMPLE_SEGMENT|3008,3014|false|false|false|C0038984;C0038990|Sweat;Sweating|sweats
Finding|Finding|SIMPLE_SEGMENT|3008,3014|false|false|false|C0038984;C0038990|Sweat;Sweating|sweats
Event|Event|SIMPLE_SEGMENT|3016,3024|false|false|false|||headache
Finding|Sign or Symptom|SIMPLE_SEGMENT|3016,3024|false|false|false|C0018681|Headache|headache
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3026,3032|false|false|false|C2707266||vision
Finding|Organism Function|SIMPLE_SEGMENT|3026,3032|false|false|false|C0042789|Vision|vision
Event|Event|SIMPLE_SEGMENT|3033,3040|false|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|3033,3040|false|false|false|C0392747|Changing|changes
Event|Event|SIMPLE_SEGMENT|3043,3053|false|false|false|||rhinorrhea
Finding|Sign or Symptom|SIMPLE_SEGMENT|3043,3053|false|false|false|C1260880|Rhinorrhea|rhinorrhea
Event|Event|SIMPLE_SEGMENT|3055,3065|false|false|false|||congestion
Finding|Pathologic Function|SIMPLE_SEGMENT|3055,3065|false|false|false|C0700148|Congestion|congestion
Finding|Sign or Symptom|SIMPLE_SEGMENT|3067,3071|false|false|false|C0234233;C1442877|Sore skin;Sore to touch|sore
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3067,3078|false|false|false|C0031350|Pharyngitis|sore throat
Drug|Organic Chemical|SIMPLE_SEGMENT|3067,3078|false|false|false|C0723402;C3244654|Sore Throat brand of Phenol;Sore Throat brand of benzocaine & menthol|sore throat
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3067,3078|false|false|false|C0723402;C3244654|Sore Throat brand of Phenol;Sore Throat brand of benzocaine & menthol|sore throat
Finding|Sign or Symptom|SIMPLE_SEGMENT|3067,3078|false|false|false|C0242429|Sore Throat|sore throat
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3072,3078|false|false|false|C0031354;C0230069;C3665375|Anterior portion of neck;Pharyngeal structure;Throat|throat
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3072,3078|false|false|false|C0031354;C0230069;C3665375|Anterior portion of neck;Pharyngeal structure;Throat|throat
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3072,3078|false|false|false|C1950455|Throat Homeopathic Medication|throat
Event|Event|SIMPLE_SEGMENT|3072,3078|false|false|false|||throat
Finding|Body Substance|SIMPLE_SEGMENT|3072,3078|false|false|false|C1547926;C1550663|Specimen Type - Throat|throat
Finding|Intellectual Product|SIMPLE_SEGMENT|3072,3078|false|false|false|C1547926;C1550663|Specimen Type - Throat|throat
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3080,3089|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|SIMPLE_SEGMENT|3080,3094|false|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3090,3094|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|3090,3094|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|3090,3094|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|3090,3094|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3096,3102|false|false|false|C4255480||nausea
Event|Event|SIMPLE_SEGMENT|3096,3102|false|false|false|||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|3096,3102|false|false|false|C0027497|Nausea|nausea
Event|Event|SIMPLE_SEGMENT|3105,3113|false|false|false|||vomiting
Finding|Sign or Symptom|SIMPLE_SEGMENT|3105,3113|false|false|false|C0042963|Vomiting|vomiting
Event|Event|SIMPLE_SEGMENT|3115,3123|false|false|false|||diarrhea
Finding|Finding|SIMPLE_SEGMENT|3115,3123|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|SIMPLE_SEGMENT|3115,3123|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Event|Event|SIMPLE_SEGMENT|3125,3137|false|false|false|||constipation
Finding|Sign or Symptom|SIMPLE_SEGMENT|3125,3137|false|false|false|C0009806|Constipation|constipation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3139,3144|false|false|false|C0018932|Hematochezia|BRBPR
Event|Event|SIMPLE_SEGMENT|3139,3144|false|false|false|||BRBPR
Event|Event|SIMPLE_SEGMENT|3146,3152|false|false|false|||melena
Finding|Pathologic Function|SIMPLE_SEGMENT|3146,3152|false|false|false|C0025222|Melena|melena
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3154,3166|false|false|false|C0018932|Hematochezia|hematochezia
Event|Event|SIMPLE_SEGMENT|3154,3166|false|false|false|||hematochezia
Finding|Sign or Symptom|SIMPLE_SEGMENT|3154,3166|false|false|false|C1321898|Blood in stool|hematochezia
Event|Event|SIMPLE_SEGMENT|3169,3176|false|false|false|||dysuria
Finding|Sign or Symptom|SIMPLE_SEGMENT|3169,3176|false|false|false|C0013428|Dysuria|dysuria
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3178,3187|false|false|false|C0018965|Hematuria|hematuria
Event|Event|SIMPLE_SEGMENT|3178,3187|false|false|false|||hematuria
Finding|Finding|SIMPLE_SEGMENT|3193,3213|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Event|Event|SIMPLE_SEGMENT|3198,3205|false|false|false|||Medical
Finding|Functional Concept|SIMPLE_SEGMENT|3198,3205|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|3198,3205|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|3198,3205|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|3198,3205|false|false|false|C0199168|Medical service|Medical
Finding|Finding|SIMPLE_SEGMENT|3198,3213|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|3206,3213|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|3206,3213|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|3206,3213|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3215,3221|false|false|false|C0004096|Asthma|ASTHMA
Event|Event|SIMPLE_SEGMENT|3215,3221|false|false|false|||ASTHMA
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3222,3226|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3222,3226|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|SIMPLE_SEGMENT|3222,3226|false|false|false|||COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|3222,3226|false|false|false|C1412502|ARCN1 gene|COPD
Finding|Finding|SIMPLE_SEGMENT|3229,3237|false|false|false|C0741302|atypia morphology|ATYPICAL
Finding|Sign or Symptom|SIMPLE_SEGMENT|3229,3248|false|false|false|C0262384|Atypical chest pain|ATYPICAL CHEST PAIN
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3238,3243|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|CHEST
Finding|Finding|SIMPLE_SEGMENT|3238,3243|false|false|false|C0741025|Chest problem|CHEST
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3238,3248|false|false|false|C2926613||CHEST PAIN
Finding|Sign or Symptom|SIMPLE_SEGMENT|3238,3248|false|false|false|C0008031|Chest Pain|CHEST PAIN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3244,3248|false|true|false|C2598155||PAIN
Event|Event|SIMPLE_SEGMENT|3244,3248|false|false|false|||PAIN
Finding|Functional Concept|SIMPLE_SEGMENT|3244,3248|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|PAIN
Finding|Sign or Symptom|SIMPLE_SEGMENT|3244,3248|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|PAIN
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3251,3259|false|false|false|C0027530|Neck|CERVICAL
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3251,3271|false|false|false|C0263884|Cervical radiculitis|CERVICAL RADICULITIS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3260,3271|false|false|false|C0034544|Radiculitis|RADICULITIS
Event|Event|SIMPLE_SEGMENT|3260,3271|false|false|false|||RADICULITIS
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3274,3282|false|false|false|C0027530|Neck|CERVICAL
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3274,3294|false|false|false|C0158241;C1384641|Cervical spondylosis;Cervical spondylosis without myelopathy|CERVICAL SPONDYLOSIS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3283,3294|false|false|false|C0038019|Spondylosis|SPONDYLOSIS
Event|Event|SIMPLE_SEGMENT|3283,3294|false|false|false|||SPONDYLOSIS
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3297,3305|false|false|false|C0018787|Heart|CORONARY
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3297,3312|false|false|false|C0205042|Coronary artery|CORONARY ARTERY
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3297,3320|false|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|CORONARY ARTERY DISEASE
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3306,3312|false|false|false|C0003842;C0226004|Arterial system;Arteries|ARTERY
Anatomy|Body System|SIMPLE_SEGMENT|3306,3312|false|false|false|C0003842;C0226004|Arterial system;Arteries|ARTERY
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3306,3320|false|false|false|C0852949|Arteriopathic disease|ARTERY DISEASE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3313,3320|false|false|false|C0012634|Disease|DISEASE
Event|Event|SIMPLE_SEGMENT|3313,3320|false|false|false|||DISEASE
Finding|Sign or Symptom|SIMPLE_SEGMENT|3323,3331|false|false|false|C0018681|Headache|HEADACHE
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3334,3337|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|HIP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3334,3337|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|HIP
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3334,3337|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|HIP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3334,3337|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|HIP
Event|Event|SIMPLE_SEGMENT|3334,3337|false|false|false|||HIP
Finding|Gene or Genome|SIMPLE_SEGMENT|3334,3337|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|HIP
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3334,3337|false|false|false|C1292890|Procedure on hip|HIP
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3334,3349|false|false|false|C0392806|Prosthetic arthroplasty of hip (procedure)|HIP REPLACEMENT
Event|Event|SIMPLE_SEGMENT|3338,3349|false|false|false|||REPLACEMENT
Finding|Functional Concept|SIMPLE_SEGMENT|3338,3349|false|false|false|C0559956|Replacement|REPLACEMENT
Procedure|Health Care Activity|SIMPLE_SEGMENT|3338,3349|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|REPLACEMENT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3338,3349|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|REPLACEMENT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3352,3366|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|HYPERLIPIDEMIA
Event|Event|SIMPLE_SEGMENT|3352,3366|false|false|false|||HYPERLIPIDEMIA
Finding|Finding|SIMPLE_SEGMENT|3352,3366|false|false|false|C0428465|Serum lipids high (finding)|HYPERLIPIDEMIA
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3369,3381|false|false|false|C0020538|Hypertensive disease|HYPERTENSION
Event|Event|SIMPLE_SEGMENT|3369,3381|false|false|false|||HYPERTENSION
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3384,3398|false|false|false|C0029408|Degenerative polyarthritis|OSTEOARTHRITIS
Event|Event|SIMPLE_SEGMENT|3384,3398|false|false|false|||OSTEOARTHRITIS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3401,3407|false|false|false|C0019340;C0854331|Herpes simplex dermatitis|HERPES
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3401,3414|false|false|false|C0019360;C0042338|Herpes zoster (disorder);herpesvirus 3, human|HERPES ZOSTER
Disorder|Virus|SIMPLE_SEGMENT|3401,3414|false|false|false|C0019360;C0042338|Herpes zoster (disorder);herpesvirus 3, human|HERPES ZOSTER
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3408,3414|false|false|false|C0019360|Herpes zoster (disorder)|ZOSTER
Event|Event|SIMPLE_SEGMENT|3408,3414|false|false|false|||ZOSTER
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3417,3423|false|false|false|C0018792|Heart Atrium|ATRIAL
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3417,3436|false|false|false|C2926591||ATRIAL FIBRILLATION
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3417,3436|false|false|false|C0004238|Atrial Fibrillation|ATRIAL FIBRILLATION
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3417,3436|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|ATRIAL FIBRILLATION
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3424,3436|false|false|false|C0232197|Fibrillation|FIBRILLATION
Event|Event|SIMPLE_SEGMENT|3424,3436|false|false|false|||FIBRILLATION
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|3439,3446|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|ANXIETY
Event|Event|SIMPLE_SEGMENT|3439,3446|false|false|false|||ANXIETY
Finding|Sign or Symptom|SIMPLE_SEGMENT|3439,3446|false|false|false|C0860603|Anxiety symptoms|ANXIETY
Finding|Intellectual Product|SIMPLE_SEGMENT|3449,3465|false|false|false|C1314977|Gastrointestinal attachment|GASTROINTESTINAL
Finding|Pathologic Function|SIMPLE_SEGMENT|3449,3474|false|false|false|C0017181|Gastrointestinal Hemorrhage|GASTROINTESTINAL BLEEDING
Finding|Pathologic Function|SIMPLE_SEGMENT|3466,3474|false|false|false|C0019080|Hemorrhage|BLEEDING
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3477,3491|false|false|false|C0029408|Degenerative polyarthritis|OSTEOARTHRITIS
Event|Event|SIMPLE_SEGMENT|3477,3491|false|false|false|||OSTEOARTHRITIS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3496,3523|false|false|false|C0085096|Peripheral Vascular Diseases|PERIPHERAL VASCULAR DISEASE
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3507,3515|false|false|false|C0005847|Blood Vessel|VASCULAR
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3507,3523|false|false|false|C0042373|Vascular Diseases|VASCULAR DISEASE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3516,3523|false|false|false|C0012634|Disease|DISEASE
Event|Event|SIMPLE_SEGMENT|3516,3523|false|false|false|||DISEASE
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3539,3544|false|false|false|C0020889|Bone structure of ilium|iliac
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3539,3551|false|false|false|C0850459|iliac stents|iliac stents
Event|Event|SIMPLE_SEGMENT|3545,3551|false|false|false|||stents
Finding|Functional Concept|SIMPLE_SEGMENT|3555,3561|false|false|false|C0728831|Social|Social
Finding|Finding|SIMPLE_SEGMENT|3555,3569|false|false|false|C0424945;C3714536|Social History;Social and personal history|Social History
Event|Event|SIMPLE_SEGMENT|3562,3569|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|3562,3569|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|3562,3569|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|3562,3569|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Classification|SIMPLE_SEGMENT|3575,3581|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|SIMPLE_SEGMENT|3575,3581|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|SIMPLE_SEGMENT|3575,3581|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|SIMPLE_SEGMENT|3575,3581|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Finding|SIMPLE_SEGMENT|3575,3589|false|false|false|C0241889|Family Medical History|Family History
Event|Event|SIMPLE_SEGMENT|3582,3589|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|3582,3589|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|3582,3589|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|3582,3589|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Idea or Concept|SIMPLE_SEGMENT|3591,3597|false|false|false|C1546508|Relationship - Mother|Mother
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3604,3607|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|SIMPLE_SEGMENT|3604,3607|false|false|false|||HTN
Finding|Conceptual Entity|SIMPLE_SEGMENT|3610,3616|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Idea or Concept|SIMPLE_SEGMENT|3610,3616|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Event|Event|SIMPLE_SEGMENT|3627,3634|false|false|false|||Brother
Finding|Conceptual Entity|SIMPLE_SEGMENT|3627,3634|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Finding|Idea or Concept|SIMPLE_SEGMENT|3627,3634|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Event|Event|SIMPLE_SEGMENT|3642,3649|false|false|false|||Brother
Finding|Conceptual Entity|SIMPLE_SEGMENT|3642,3649|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Finding|Idea or Concept|SIMPLE_SEGMENT|3642,3649|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Event|Event|SIMPLE_SEGMENT|3658,3666|false|false|false|||Physical
Finding|Finding|SIMPLE_SEGMENT|3658,3666|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|3658,3666|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|3658,3666|false|false|false|C0031809|Physical Examination|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|3690,3699|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|SIMPLE_SEGMENT|3700,3704|false|false|false|||EXAM
Finding|Functional Concept|SIMPLE_SEGMENT|3700,3704|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|SIMPLE_SEGMENT|3700,3704|false|false|false|C0582103|Medical Examination|EXAM
Event|Event|SIMPLE_SEGMENT|3782,3789|false|false|false|||GENERAL
Finding|Classification|SIMPLE_SEGMENT|3782,3789|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|3782,3789|false|false|false|C3812897|General medical service|GENERAL
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3797,3800|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3797,3800|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3797,3800|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|3797,3800|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3797,3800|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|SIMPLE_SEGMENT|3797,3800|false|false|false|||NAD
Finding|Finding|SIMPLE_SEGMENT|3797,3800|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Event|Event|SIMPLE_SEGMENT|3802,3809|false|false|false|||sitting
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3816,3819|false|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Finding|Intellectual Product|SIMPLE_SEGMENT|3816,3819|false|false|false|C2346952|Bachelor of Education|bed
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3820,3825|false|false|false|C1512338|HEENT|HEENT
Event|Event|SIMPLE_SEGMENT|3827,3840|false|false|false|||Normocephalic
Event|Event|SIMPLE_SEGMENT|3842,3852|false|false|false|||atraumatic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3855,3861|false|false|false|C0034121|Pupil|Pupils
Finding|Finding|SIMPLE_SEGMENT|3855,3867|false|false|false|C0578617|Pupils equal|Pupils equal
Event|Event|SIMPLE_SEGMENT|3862,3867|false|false|false|||equal
Finding|Intellectual Product|SIMPLE_SEGMENT|3862,3867|false|false|false|C1549782|Relational Operator - Equal|equal
Event|Event|SIMPLE_SEGMENT|3881,3889|false|false|false|||reactive
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3881,3889|false|false|false|C4722408|Reactive Therapy|reactive
Finding|Functional Concept|SIMPLE_SEGMENT|3903,3914|false|false|false|C0241886|Extraocular|extraocular
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3903,3922|false|false|false|C0028863|Muscle of orbit|extraocular muscles
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3915,3922|false|false|false|C0026845;C1995013;C4083049|Muscle (organ);Muscle Tissue;Set of muscles|muscles
Anatomy|Tissue|SIMPLE_SEGMENT|3915,3922|false|false|false|C0026845;C1995013;C4083049|Muscle (organ);Muscle Tissue;Set of muscles|muscles
Event|Event|SIMPLE_SEGMENT|3923,3929|false|false|false|||intact
Finding|Finding|SIMPLE_SEGMENT|3923,3929|false|false|false|C1554187|Gender Status - Intact|intact
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3936,3948|true|false|false|C0009758|conjunctiva|conjunctival
Finding|Functional Concept|SIMPLE_SEGMENT|3936,3948|true|false|false|C1522483|Conjunctival Route of Administration|conjunctival
Finding|Finding|SIMPLE_SEGMENT|3936,3955|true|false|false|C2071267|Conjunctival pallor|conjunctival pallor
Event|Event|SIMPLE_SEGMENT|3949,3955|true|false|false|||pallor
Finding|Finding|SIMPLE_SEGMENT|3949,3955|true|false|false|C0241137|Pallor of skin|pallor
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3959,3968|true|false|false|C1272883|Injection|injection
Event|Event|SIMPLE_SEGMENT|3959,3968|true|false|false|||injection
Finding|Functional Concept|SIMPLE_SEGMENT|3959,3968|true|false|false|C1828121|Injection Route of Administration|injection
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3959,3968|true|false|false|C0021485;C1533685|Injection of therapeutic agent;Injection procedure|injection
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3970,3976|true|false|false|C0036410|Sclera|sclera
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3970,3976|true|false|false|C0036412|Scleral Diseases|sclera
Event|Event|SIMPLE_SEGMENT|3970,3976|true|false|false|||sclera
Procedure|Health Care Activity|SIMPLE_SEGMENT|3970,3976|true|false|false|C2228481|examination of sclera|sclera
Event|Event|SIMPLE_SEGMENT|3977,3986|true|false|false|||anicteric
Finding|Finding|SIMPLE_SEGMENT|3977,3986|true|false|false|C0205180|Anicteric|anicteric
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4000,4009|true|false|false|C1272883|Injection|injection
Event|Event|SIMPLE_SEGMENT|4000,4009|true|false|false|||injection
Finding|Functional Concept|SIMPLE_SEGMENT|4000,4009|true|false|false|C1828121|Injection Route of Administration|injection
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4000,4009|true|false|false|C0021485;C1533685|Injection of therapeutic agent;Injection procedure|injection
Finding|Finding|SIMPLE_SEGMENT|4011,4033|false|false|false|C0517391|Moist mucous membranes|Moist mucous membranes
Finding|Body Substance|SIMPLE_SEGMENT|4017,4023|false|false|false|C0026727;C2753459|Mucus (substance);mucus layer|mucous
Anatomy|Tissue|SIMPLE_SEGMENT|4017,4033|false|false|false|C0026724|Mucous Membrane|mucous membranes
Finding|Finding|SIMPLE_SEGMENT|4017,4033|false|false|false|C2230150|moisture of mucous membranes (physical finding)|mucous membranes
Anatomy|Tissue|SIMPLE_SEGMENT|4024,4033|false|false|false|C0025255|Membrane Tissue|membranes
Finding|Idea or Concept|SIMPLE_SEGMENT|4035,4039|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4040,4049|false|false|false|C0011443;C0040426|Dentition;Tooth structure|dentition
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4052,4062|false|false|false|C0521367|Oropharyngeal|Oropharynx
Event|Event|SIMPLE_SEGMENT|4067,4072|false|false|false|||clear
Finding|Idea or Concept|SIMPLE_SEGMENT|4067,4072|false|false|false|C1550016|Remote control command - Clear|clear
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4074,4078|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|SIMPLE_SEGMENT|4074,4078|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|SIMPLE_SEGMENT|4074,4078|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Event|Event|SIMPLE_SEGMENT|4080,4086|false|false|false|||Supple
Finding|Functional Concept|SIMPLE_SEGMENT|4080,4086|false|false|false|C0332254|Supple|Supple
Event|Event|SIMPLE_SEGMENT|4088,4091|true|false|false|||JVD
Finding|Finding|SIMPLE_SEGMENT|4088,4091|true|false|false|C0425687|Jugular venous engorgement|JVD
Event|Event|SIMPLE_SEGMENT|4096,4106|true|false|false|||visualized
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4108,4115|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|SIMPLE_SEGMENT|4108,4115|false|false|false|C1314974|Cardiac attachment|CARDIAC
Event|Event|SIMPLE_SEGMENT|4129,4138|false|false|false|||irregular
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|4144,4152|false|false|false|C0039155|Systole|systolic
Finding|Finding|SIMPLE_SEGMENT|4144,4159|true|false|false|C0232257|Systolic Murmurs|systolic murmur
Event|Event|SIMPLE_SEGMENT|4153,4159|true|false|false|||murmur
Finding|Finding|SIMPLE_SEGMENT|4153,4159|true|false|false|C0018808|Heart murmur|murmur
Event|Event|SIMPLE_SEGMENT|4160,4164|true|false|false|||best
Event|Event|SIMPLE_SEGMENT|4173,4176|true|false|false|||LSB
Event|Event|SIMPLE_SEGMENT|4181,4185|true|false|false|||rubs
Finding|Finding|SIMPLE_SEGMENT|4181,4185|true|false|false|C0232267|Pericardial friction rub|rubs
Event|Event|SIMPLE_SEGMENT|4189,4196|true|false|false|||gallops
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4198,4203|false|false|false|C0024109|Lung|LUNGS
Finding|Intellectual Product|SIMPLE_SEGMENT|4205,4209|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|Poor
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4210,4213|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4210,4213|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|SIMPLE_SEGMENT|4210,4213|false|false|false|C0001861;C3536832|Air (substance);air|air
Finding|Finding|SIMPLE_SEGMENT|4210,4213|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|SIMPLE_SEGMENT|4210,4213|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|SIMPLE_SEGMENT|4210,4213|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|4210,4222|false|false|false|C0001868|Air Movements|air movement
Event|Event|SIMPLE_SEGMENT|4214,4222|false|false|false|||movement
Finding|Organism Function|SIMPLE_SEGMENT|4214,4222|false|false|false|C0026649|Movement|movement
Finding|Intellectual Product|SIMPLE_SEGMENT|4235,4239|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Event|Event|SIMPLE_SEGMENT|4248,4259|false|false|false|||inspiratory
Finding|Organism Function|SIMPLE_SEGMENT|4248,4259|false|false|false|C0004048|Inspiration (function)|inspiratory
Finding|Organism Function|SIMPLE_SEGMENT|4265,4275|false|false|false|C0231800|Expiration, Respiratory|expiratory
Finding|Sign or Symptom|SIMPLE_SEGMENT|4265,4283|false|false|false|C0231875|Expiratory wheezing|expiratory wheezes
Event|Event|SIMPLE_SEGMENT|4276,4283|false|false|false|||wheezes
Finding|Sign or Symptom|SIMPLE_SEGMENT|4276,4283|false|false|false|C0043144|Wheezing|wheezes
Event|Event|SIMPLE_SEGMENT|4288,4291|true|false|false|||use
Finding|Functional Concept|SIMPLE_SEGMENT|4288,4291|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|SIMPLE_SEGMENT|4288,4291|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Functional Concept|SIMPLE_SEGMENT|4288,4294|true|false|false|C1524063|Use of|use of
Finding|Finding|SIMPLE_SEGMENT|4288,4312|true|false|false|C1821466|Use of accessory muscles|use of accessory muscles
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|4295,4312|true|false|false|C0158784|Accessory skeletal muscle|accessory muscles
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4305,4312|true|false|false|C0026845;C1995013;C4083049|Muscle (organ);Muscle Tissue;Set of muscles|muscles
Anatomy|Tissue|SIMPLE_SEGMENT|4305,4312|true|false|false|C0026845;C1995013;C4083049|Muscle (organ);Muscle Tissue;Set of muscles|muscles
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4317,4326|true|false|false|C5885990||breathing
Event|Event|SIMPLE_SEGMENT|4317,4326|true|false|false|||breathing
Finding|Finding|SIMPLE_SEGMENT|4317,4326|true|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|SIMPLE_SEGMENT|4317,4326|true|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|SIMPLE_SEGMENT|4317,4326|true|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|SIMPLE_SEGMENT|4317,4326|true|false|false|C1160636|respiratory system process|breathing
Event|Event|SIMPLE_SEGMENT|4331,4338|true|false|false|||rhonchi
Finding|Finding|SIMPLE_SEGMENT|4331,4338|true|false|false|C0035508|Rhonchi|rhonchi
Event|Event|SIMPLE_SEGMENT|4342,4347|true|false|false|||rales
Finding|Finding|SIMPLE_SEGMENT|4342,4347|true|false|false|C0034642;C0240859|Basilar Rales;Rales|rales
Event|Event|SIMPLE_SEGMENT|4349,4353|false|false|false|||BACK
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4358,4361|true|false|false|C0001365;C0038454|Acute ill-defined cerebrovascular disease;Cerebrovascular accident|CVA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4358,4361|true|false|false|C5779650|Cyclophosphamide/Doxorubicin/Vincristine|CVA
Event|Event|SIMPLE_SEGMENT|4358,4361|true|false|false|||CVA
Finding|Sign or Symptom|SIMPLE_SEGMENT|4358,4372|true|false|false|C0235634|Renal angle tenderness|CVA tenderness
Event|Event|SIMPLE_SEGMENT|4362,4372|true|false|false|||tenderness
Finding|Mental Process|SIMPLE_SEGMENT|4362,4372|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|SIMPLE_SEGMENT|4362,4372|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4374,4381|true|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4374,4381|true|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Event|Event|SIMPLE_SEGMENT|4374,4381|true|false|false|||ABDOMEN
Finding|Finding|SIMPLE_SEGMENT|4374,4381|true|false|false|C0941288|Abdomen problem|ABDOMEN
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4391,4397|false|false|false|C0021853|Intestines|bowels
Event|Event|SIMPLE_SEGMENT|4398,4404|false|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|4398,4404|false|false|false|C0037709||sounds
Event|Event|SIMPLE_SEGMENT|4410,4419|false|false|false|||distended
Finding|Finding|SIMPLE_SEGMENT|4410,4419|false|false|false|C0700124|Dilated|distended
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4436,4440|false|false|false|C4318566|Deep Resection Margin|deep
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4436,4450|false|false|false|C0278328|Deep palpation|deep palpation
Event|Event|SIMPLE_SEGMENT|4441,4450|false|false|false|||palpation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4441,4450|false|false|false|C0030247|Palpation|palpation
Event|Event|SIMPLE_SEGMENT|4477,4489|true|false|false|||organomegaly
Finding|Finding|SIMPLE_SEGMENT|4477,4489|true|false|false|C4054315|Organomegaly|organomegaly
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4491,4502|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|4507,4515|true|false|false|C0149651|Clubbing|clubbing
Event|Event|SIMPLE_SEGMENT|4507,4515|true|false|false|||clubbing
Event|Event|SIMPLE_SEGMENT|4519,4527|true|false|false|||cyanosis
Finding|Sign or Symptom|SIMPLE_SEGMENT|4519,4527|true|false|false|C0010520|Cyanosis|cyanosis
Finding|Finding|SIMPLE_SEGMENT|4529,4552|false|false|false|C2237594|bilateral pitting edema|Bilateral pitting edema
Finding|Functional Concept|SIMPLE_SEGMENT|4539,4546|false|false|false|C0205323|Pitting|pitting
Finding|Finding|SIMPLE_SEGMENT|4539,4552|false|false|false|C0333243|Pitting edema|pitting edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4547,4552|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|4547,4552|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|4547,4552|false|false|false|C0013604|Edema|edema
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4565,4569|false|false|false|C0230444|Shin|shin
Drug|Food|SIMPLE_SEGMENT|4571,4577|false|false|false|C5890763||Pulses
Event|Event|SIMPLE_SEGMENT|4571,4577|false|false|false|||Pulses
Finding|Physiologic Function|SIMPLE_SEGMENT|4571,4577|false|false|false|C0391850|Physiologic pulse|Pulses
Procedure|Health Care Activity|SIMPLE_SEGMENT|4571,4577|false|false|false|C0034107|Pulse taking|Pulses
Event|Event|SIMPLE_SEGMENT|4578,4580|false|false|false|||DP
Finding|Conceptual Entity|SIMPLE_SEGMENT|4581,4587|false|false|false|C0442038;C0920847|Circumpennate;Radial|Radial
Anatomy|Body System|SIMPLE_SEGMENT|4604,4608|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4604,4608|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4604,4608|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Event|Event|SIMPLE_SEGMENT|4604,4608|false|false|false|||SKIN
Finding|Body Substance|SIMPLE_SEGMENT|4604,4608|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|SIMPLE_SEGMENT|4604,4608|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4613,4617|true|false|false|C5779629|Eruption of skin (disorder)|rash
Event|Event|SIMPLE_SEGMENT|4613,4617|true|false|false|||rash
Finding|Pathologic Function|SIMPLE_SEGMENT|4613,4617|true|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Sign or Symptom|SIMPLE_SEGMENT|4613,4617|true|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Event|Event|SIMPLE_SEGMENT|4621,4627|true|false|false|||ulcers
Finding|Pathologic Function|SIMPLE_SEGMENT|4621,4627|true|false|false|C0041582|Ulcer|ulcers
Event|Event|SIMPLE_SEGMENT|4628,4638|true|false|false|||NEUROLOGIC
Finding|Gene or Genome|SIMPLE_SEGMENT|4640,4643|false|false|false|C1539110|CNDP2 gene|CN2
Event|Event|SIMPLE_SEGMENT|4647,4653|false|false|false|||intact
Finding|Finding|SIMPLE_SEGMENT|4647,4653|false|false|false|C1554187|Gender Status - Intact|intact
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4662,4677|false|false|false|C0278454|All extremities|all extremities
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4666,4677|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Event|Event|SIMPLE_SEGMENT|4702,4711|false|false|false|||sensation
Finding|Finding|SIMPLE_SEGMENT|4702,4711|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|4702,4711|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|SIMPLE_SEGMENT|4702,4711|false|false|false|C2229507|sensory exam|sensation
Finding|Body Substance|SIMPLE_SEGMENT|4732,4741|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|4732,4741|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|4732,4741|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|4732,4741|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|SIMPLE_SEGMENT|4742,4746|false|false|false|||EXAM
Finding|Functional Concept|SIMPLE_SEGMENT|4742,4746|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|SIMPLE_SEGMENT|4742,4746|false|false|false|C0582103|Medical Examination|EXAM
Event|Event|SIMPLE_SEGMENT|4824,4831|false|false|false|||GENERAL
Finding|Classification|SIMPLE_SEGMENT|4824,4831|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|4824,4831|false|false|false|C3812897|General medical service|GENERAL
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4839,4842|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4839,4842|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4839,4842|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|4839,4842|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4839,4842|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|SIMPLE_SEGMENT|4839,4842|false|false|false|||NAD
Finding|Finding|SIMPLE_SEGMENT|4839,4842|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Event|Event|SIMPLE_SEGMENT|4844,4851|false|false|false|||sitting
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4858,4861|false|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Finding|Intellectual Product|SIMPLE_SEGMENT|4858,4861|false|false|false|C2346952|Bachelor of Education|bed
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4862,4867|false|false|false|C1512338|HEENT|HEENT
Event|Event|SIMPLE_SEGMENT|4869,4873|false|false|false|||NCAT
Event|Event|SIMPLE_SEGMENT|4876,4881|false|false|false|||PERRL
Finding|Finding|SIMPLE_SEGMENT|4876,4881|false|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Event|Event|SIMPLE_SEGMENT|4883,4887|false|false|false|||EOMI
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4889,4895|true|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4889,4895|true|false|false|C0036412|Scleral Diseases|Sclera
Event|Event|SIMPLE_SEGMENT|4889,4895|true|false|false|||Sclera
Procedure|Health Care Activity|SIMPLE_SEGMENT|4889,4895|true|false|false|C2228481|examination of sclera|Sclera
Event|Event|SIMPLE_SEGMENT|4896,4905|true|false|false|||anicteric
Finding|Finding|SIMPLE_SEGMENT|4896,4905|true|false|false|C0205180|Anicteric|anicteric
Event|Event|SIMPLE_SEGMENT|4914,4922|true|false|false|||injected
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4925,4928|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4925,4928|false|false|false|C0026987|Myelofibrosis|MMM
Event|Event|SIMPLE_SEGMENT|4925,4928|false|false|false|||MMM
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4932,4942|false|false|false|C0521367|Oropharyngeal|Oropharynx
Event|Event|SIMPLE_SEGMENT|4946,4951|false|false|false|||clear
Finding|Idea or Concept|SIMPLE_SEGMENT|4946,4951|false|false|false|C1550016|Remote control command - Clear|clear
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4953,4957|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|SIMPLE_SEGMENT|4953,4957|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|SIMPLE_SEGMENT|4953,4957|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Event|Event|SIMPLE_SEGMENT|4959,4965|false|false|false|||Supple
Finding|Functional Concept|SIMPLE_SEGMENT|4959,4965|false|false|false|C0332254|Supple|Supple
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4970,4973|true|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4970,4973|true|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|SIMPLE_SEGMENT|4970,4973|true|false|false|||LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|4970,4973|true|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Event|Event|SIMPLE_SEGMENT|4975,4978|true|false|false|||JVP
Finding|Finding|SIMPLE_SEGMENT|4975,4978|true|false|false|C0428897|Jugular venous pressure|JVP
Event|Event|SIMPLE_SEGMENT|4983,4994|true|false|false|||appreciated
Event|Event|SIMPLE_SEGMENT|5001,5008|true|false|false|||degrees
Finding|Intellectual Product|SIMPLE_SEGMENT|5001,5008|true|false|false|C0542560|Academic degree|degrees
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5010,5017|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|SIMPLE_SEGMENT|5010,5017|false|false|false|C1314974|Cardiac attachment|CARDIAC
Event|Event|SIMPLE_SEGMENT|5031,5040|false|false|false|||irregular
Event|Activity|SIMPLE_SEGMENT|5049,5053|false|false|false|C0871208|Rating (action)|rate
Event|Event|SIMPLE_SEGMENT|5049,5053|false|false|false|||rate
Finding|Idea or Concept|SIMPLE_SEGMENT|5049,5053|false|false|false|C1549480|Amount type - Rate|rate
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|5059,5067|false|false|false|C0039155|Systole|systolic
Finding|Finding|SIMPLE_SEGMENT|5059,5074|false|false|false|C0232257|Systolic Murmurs|systolic murmur
Event|Event|SIMPLE_SEGMENT|5068,5074|false|false|false|||murmur
Finding|Finding|SIMPLE_SEGMENT|5068,5074|false|false|false|C0018808|Heart murmur|murmur
Event|Event|SIMPLE_SEGMENT|5083,5087|false|false|false|||RUSB
Event|Event|SIMPLE_SEGMENT|5092,5096|true|false|false|||rubs
Finding|Finding|SIMPLE_SEGMENT|5092,5096|true|false|false|C0232267|Pericardial friction rub|rubs
Event|Event|SIMPLE_SEGMENT|5100,5107|true|false|false|||gallops
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5109,5114|false|false|false|C0024109|Lung|LUNGS
Finding|Intellectual Product|SIMPLE_SEGMENT|5116,5120|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|Poor
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5121,5124|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5121,5124|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|SIMPLE_SEGMENT|5121,5124|false|false|false|C0001861;C3536832|Air (substance);air|air
Finding|Finding|SIMPLE_SEGMENT|5121,5124|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|SIMPLE_SEGMENT|5121,5124|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|SIMPLE_SEGMENT|5121,5124|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|5121,5133|false|false|false|C0001868|Air Movements|air movement
Event|Event|SIMPLE_SEGMENT|5125,5133|false|false|false|||movement
Finding|Organism Function|SIMPLE_SEGMENT|5125,5133|false|false|false|C0026649|Movement|movement
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5162,5167|false|false|false|C0024109|Lung|lungs
Event|Event|SIMPLE_SEGMENT|5173,5180|true|false|false|||wheezes
Finding|Sign or Symptom|SIMPLE_SEGMENT|5173,5180|true|false|false|C0043144|Wheezing|wheezes
Finding|Organism Function|SIMPLE_SEGMENT|5195,5205|true|false|false|C0231800|Expiration, Respiratory|expiratory
Event|Event|SIMPLE_SEGMENT|5206,5211|true|false|false|||phase
Event|Event|SIMPLE_SEGMENT|5216,5223|true|false|false|||rhonchi
Finding|Finding|SIMPLE_SEGMENT|5216,5223|true|false|false|C0035508|Rhonchi|rhonchi
Event|Event|SIMPLE_SEGMENT|5227,5232|true|false|false|||rales
Finding|Finding|SIMPLE_SEGMENT|5227,5232|true|false|false|C0034642;C0240859|Basilar Rales;Rales|rales
Event|Event|SIMPLE_SEGMENT|5235,5239|false|false|false|||Does
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5254,5259|false|false|false|C2936910|Cross syndrome|cross
Event|Event|SIMPLE_SEGMENT|5254,5259|false|false|false|||cross
Finding|Conceptual Entity|SIMPLE_SEGMENT|5254,5259|false|false|false|C2828360|Traverse|cross
Event|Event|SIMPLE_SEGMENT|5260,5266|false|false|false|||legged
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5274,5277|false|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Event|Event|SIMPLE_SEGMENT|5274,5277|false|false|false|||bed
Finding|Intellectual Product|SIMPLE_SEGMENT|5274,5277|false|false|false|C2346952|Bachelor of Education|bed
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5283,5291|false|false|false|C0016536|Forearm|forearms
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5300,5304|false|false|false|C1140621|Leg|legs
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5300,5304|false|false|false|C5781420||legs
Finding|Finding|SIMPLE_SEGMENT|5310,5325|false|false|false|C3875386|Tripod position|tripod position
Event|Event|SIMPLE_SEGMENT|5317,5325|false|false|false|||position
Event|Event|SIMPLE_SEGMENT|5327,5331|false|false|false|||BACK
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5336,5339|true|false|false|C0001365;C0038454|Acute ill-defined cerebrovascular disease;Cerebrovascular accident|CVA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5336,5339|true|false|false|C5779650|Cyclophosphamide/Doxorubicin/Vincristine|CVA
Event|Event|SIMPLE_SEGMENT|5336,5339|true|false|false|||CVA
Finding|Sign or Symptom|SIMPLE_SEGMENT|5336,5350|true|false|false|C0235634|Renal angle tenderness|CVA tenderness
Event|Event|SIMPLE_SEGMENT|5340,5350|true|false|false|||tenderness
Finding|Mental Process|SIMPLE_SEGMENT|5340,5350|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|SIMPLE_SEGMENT|5340,5350|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5353,5360|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5353,5360|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Event|Event|SIMPLE_SEGMENT|5353,5360|false|false|false|||ABDOMEN
Finding|Finding|SIMPLE_SEGMENT|5353,5360|false|false|false|C0941288|Abdomen problem|ABDOMEN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5368,5372|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|SIMPLE_SEGMENT|5368,5372|false|false|false|||soft
Event|Event|SIMPLE_SEGMENT|5374,5383|false|false|false|||nontender
Event|Event|SIMPLE_SEGMENT|5385,5397|false|false|false|||nondistended
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5398,5409|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Finding|Functional Concept|SIMPLE_SEGMENT|5411,5416|false|false|false|C1883002|Sequence Chromatogram|Trace
Event|Event|SIMPLE_SEGMENT|5417,5424|false|false|false|||pitting
Finding|Functional Concept|SIMPLE_SEGMENT|5417,5424|false|false|false|C0205323|Pitting|pitting
Finding|Finding|SIMPLE_SEGMENT|5417,5430|false|false|false|C0333243|Pitting edema|pitting edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5425,5430|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|5425,5430|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|5425,5430|false|false|false|C0013604|Edema|edema
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5442,5446|false|false|false|C0230444|Shin|shin
Drug|Food|SIMPLE_SEGMENT|5454,5460|false|false|false|C5890763||pulses
Event|Event|SIMPLE_SEGMENT|5454,5460|false|false|false|||pulses
Finding|Physiologic Function|SIMPLE_SEGMENT|5454,5460|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|SIMPLE_SEGMENT|5454,5460|false|false|false|C0034107|Pulse taking|pulses
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5478,5481|true|false|false|C0034155;C1268935|Congenital Thrombotic Thrombocytopenic Purpura;Purpura, Thrombotic Thrombocytopenic|TTP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5478,5481|true|false|false|C1506603;C4723973|ZFP36 protein, human;thiamine triphosphorate|TTP
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5478,5481|true|false|false|C1506603;C4723973|ZFP36 protein, human;thiamine triphosphorate|TTP
Drug|Organic Chemical|SIMPLE_SEGMENT|5478,5481|true|false|false|C1506603;C4723973|ZFP36 protein, human;thiamine triphosphorate|TTP
Drug|Vitamin|SIMPLE_SEGMENT|5478,5481|true|false|false|C1506603;C4723973|ZFP36 protein, human;thiamine triphosphorate|TTP
Event|Event|SIMPLE_SEGMENT|5478,5481|true|false|false|||TTP
Finding|Gene or Genome|SIMPLE_SEGMENT|5478,5481|true|false|false|C1413036;C1421571;C3539814|ADAMTS13 gene;ZFP36 gene;ZFP36 wt Allele|TTP
Anatomy|Body System|SIMPLE_SEGMENT|5483,5487|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5483,5487|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5483,5487|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Event|Event|SIMPLE_SEGMENT|5483,5487|false|false|false|||SKIN
Finding|Body Substance|SIMPLE_SEGMENT|5483,5487|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|SIMPLE_SEGMENT|5483,5487|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5492,5496|true|false|false|C5779629|Eruption of skin (disorder)|rash
Event|Event|SIMPLE_SEGMENT|5492,5496|true|false|false|||rash
Finding|Pathologic Function|SIMPLE_SEGMENT|5492,5496|true|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Sign or Symptom|SIMPLE_SEGMENT|5492,5496|true|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Event|Event|SIMPLE_SEGMENT|5500,5506|true|false|false|||ulcers
Finding|Pathologic Function|SIMPLE_SEGMENT|5500,5506|true|false|false|C0041582|Ulcer|ulcers
Event|Event|SIMPLE_SEGMENT|5508,5518|false|false|false|||NEUROLOGIC
Finding|Gene or Genome|SIMPLE_SEGMENT|5520,5523|false|false|false|C1539110|CNDP2 gene|CN2
Event|Event|SIMPLE_SEGMENT|5527,5533|false|false|false|||intact
Finding|Finding|SIMPLE_SEGMENT|5527,5533|false|false|false|C1554187|Gender Status - Intact|intact
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5542,5557|false|false|false|C0278454|All extremities|all extremities
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5546,5557|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Event|Event|SIMPLE_SEGMENT|5582,5591|false|false|false|||sensation
Finding|Finding|SIMPLE_SEGMENT|5582,5591|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|5582,5591|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|SIMPLE_SEGMENT|5582,5591|false|false|false|C2229507|sensory exam|sensation
Procedure|Health Care Activity|SIMPLE_SEGMENT|5634,5643|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|SIMPLE_SEGMENT|5644,5648|false|false|false|||LABS
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5644,5648|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5681,5686|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5681,5686|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5681,5686|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|5687,5690|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|5695,5698|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5695,5698|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5695,5698|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5704,5707|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5704,5707|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|5704,5707|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5704,5707|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5713,5716|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5713,5716|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|5722,5725|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|5722,5725|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5722,5725|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5722,5725|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5722,5725|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|5730,5733|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5730,5733|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|5730,5733|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|5730,5733|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|5730,5733|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5730,5733|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|SIMPLE_SEGMENT|5739,5743|false|false|false|||MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5739,5743|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5772,5775|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5792,5797|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5792,5797|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5792,5797|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5810,5816|false|false|false|C0024202|Lymph|Lymphs
Drug|Antibiotic|SIMPLE_SEGMENT|5822,5827|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5822,5827|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|SIMPLE_SEGMENT|5822,5827|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5833,5836|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|Eos
Event|Event|SIMPLE_SEGMENT|5833,5836|false|false|false|||Eos
Finding|Gene or Genome|SIMPLE_SEGMENT|5833,5836|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|Eos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5939,5944|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5939,5944|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5939,5944|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|5939,5952|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5939,5952|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5939,5952|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5945,5952|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|5945,5952|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5945,5952|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|5945,5952|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5945,5952|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5945,5952|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5998,6002|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5998,6002|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5998,6002|false|false|false|C0202059|Bicarbonate measurement|HCO3
Event|Event|SIMPLE_SEGMENT|6044,6051|false|false|false|||RESULTS
Event|Event|SIMPLE_SEGMENT|6072,6076|false|false|false|||LABS
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6072,6076|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6109,6114|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|6109,6114|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|6109,6114|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Event|Event|SIMPLE_SEGMENT|6119,6122|false|false|false|||pO2
Finding|Classification|SIMPLE_SEGMENT|6119,6122|false|false|false|C0391840;C4521535|Partial pressure of Oxygen;US Military enlisted E5|pO2
Finding|Molecular Function|SIMPLE_SEGMENT|6119,6122|false|false|false|C0391840;C4521535|Partial pressure of Oxygen;US Military enlisted E5|pO2
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6119,6122|false|false|false|C1283004|PO2 measurement|pO2
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6127,6131|false|false|false|C0391839|Carbon dioxide, partial pressure|pCO2
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6127,6131|false|false|false|C0201931|Carbon dioxide measurement, partial pressure|pCO2
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6157,6161|false|false|false|C2987514|Anatomical base|Base
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6157,6161|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|Base
Drug|Chemical Viewed Functionally|SIMPLE_SEGMENT|6157,6161|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|Base
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|6157,6161|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|Base
Finding|Gene or Genome|SIMPLE_SEGMENT|6157,6161|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|Base
Finding|Idea or Concept|SIMPLE_SEGMENT|6157,6161|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|Base
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6183,6188|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|6183,6188|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|6183,6188|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6203,6209|false|false|false|C5574646|Natriuretic Peptides B, human|proBNP
Drug|Hormone|SIMPLE_SEGMENT|6203,6209|false|false|false|C5574646|Natriuretic Peptides B, human|proBNP
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6226,6231|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|6226,6231|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|6226,6231|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6232,6237|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|SIMPLE_SEGMENT|6232,6237|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|SIMPLE_SEGMENT|6232,6237|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6232,6237|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6235,6239|false|false|false|C4722362|MB-6|MB-6
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6266,6271|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|6266,6271|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|6266,6271|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6272,6277|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|SIMPLE_SEGMENT|6272,6277|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|SIMPLE_SEGMENT|6272,6277|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6272,6277|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6275,6279|false|false|false|C4722362|MB-6|MB-6
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6310,6315|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|6310,6315|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|6310,6315|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|6316,6328|false|false|false|C0039771|theophylline|THEOPHYLLINE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6316,6328|false|false|false|C0039771|theophylline|THEOPHYLLINE
Event|Event|SIMPLE_SEGMENT|6316,6328|false|false|false|||THEOPHYLLINE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6316,6328|false|false|false|C0039773|Assay of theophylline|THEOPHYLLINE
Event|Event|SIMPLE_SEGMENT|6365,6372|false|false|false|||IMAGING
Finding|Finding|SIMPLE_SEGMENT|6365,6372|false|false|false|C0740845|Imaging problem|IMAGING
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6365,6372|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|IMAGING
Event|Event|SIMPLE_SEGMENT|6393,6396|false|false|false|||CXR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6393,6396|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|SIMPLE_SEGMENT|6404,6406|false|false|false|||PA
Event|Event|SIMPLE_SEGMENT|6419,6424|false|false|false|||views
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6429,6434|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|6429,6434|false|false|false|C0741025|Chest problem|chest
Event|Event|SIMPLE_SEGMENT|6435,6443|false|false|false|||provided
Anatomy|Tissue|SIMPLE_SEGMENT|6455,6462|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6455,6462|false|false|false|C0032226|Pleural Diseases|pleural
Event|Event|SIMPLE_SEGMENT|6475,6483|false|false|false|||scarring
Finding|Pathologic Function|SIMPLE_SEGMENT|6475,6483|false|false|false|C0008767;C2004491|Cicatrix;Cicatrization|scarring
Event|Event|SIMPLE_SEGMENT|6484,6489|false|false|false|||noted
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6501,6514|true|false|false|C0521530|Lung consolidation|consolidation
Event|Event|SIMPLE_SEGMENT|6501,6514|true|false|false|||consolidation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6531,6540|true|false|false|C0032285|Pneumonia|pneumonia
Event|Event|SIMPLE_SEGMENT|6531,6540|true|false|false|||pneumonia
Event|Event|SIMPLE_SEGMENT|6545,6553|true|false|false|||effusion
Finding|Body Substance|SIMPLE_SEGMENT|6545,6553|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|SIMPLE_SEGMENT|6545,6553|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|6545,6553|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6557,6569|true|false|false|C0032326|Pneumothorax|pneumothorax
Event|Event|SIMPLE_SEGMENT|6557,6569|true|false|false|||pneumothorax
Event|Event|SIMPLE_SEGMENT|6575,6580|true|false|false|||signs
Finding|Finding|SIMPLE_SEGMENT|6575,6580|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|SIMPLE_SEGMENT|6575,6580|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Event|Event|SIMPLE_SEGMENT|6585,6595|true|false|false|||congestion
Finding|Pathologic Function|SIMPLE_SEGMENT|6585,6595|true|false|false|C0700148|Congestion|congestion
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6599,6604|true|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|6599,6604|true|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|6599,6604|true|false|false|C0013604|Edema|edema
Event|Event|SIMPLE_SEGMENT|6624,6634|false|false|false|||silhouette
Event|Event|SIMPLE_SEGMENT|6638,6644|false|false|false|||stable
Finding|Intellectual Product|SIMPLE_SEGMENT|6638,6644|false|false|false|C1547311|Patient Condition Code - Stable|stable
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6663,6671|false|false|false|C0817096|Chest|thoracic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6663,6671|false|false|false|C5779551|Dissecting Thoracic Aortic Aneurysm|thoracic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6663,6677|false|false|false|C1522460;C4037977|Chest>Aorta.thoracic;Thoracic aorta|thoracic aorta
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6672,6677|false|false|false|C0003483;C4037978|Aorta;Chest+Abdomen>Aorta|aorta
Procedure|Health Care Activity|SIMPLE_SEGMENT|6672,6677|false|false|false|C0869784|Procedure on aorta|aorta
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6693,6698|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6693,6698|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|6693,6698|false|false|false|C0795691|HEART PROBLEM|heart
Finding|Finding|SIMPLE_SEGMENT|6693,6703|false|false|false|C0744689|heart size|heart size
Event|Event|SIMPLE_SEGMENT|6699,6703|false|false|false|||size
Finding|Functional Concept|SIMPLE_SEGMENT|6705,6709|false|false|false|C0443157|Bony|Bony
Event|Event|SIMPLE_SEGMENT|6711,6721|false|false|false|||structures
Event|Event|SIMPLE_SEGMENT|6726,6732|false|false|false|||intact
Finding|Finding|SIMPLE_SEGMENT|6726,6732|false|false|false|C1554187|Gender Status - Intact|intact
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6738,6746|false|false|false|C0881858||CT Chest
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6738,6746|false|false|false|C0202823|Chest CT|CT Chest
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6741,6746|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|SIMPLE_SEGMENT|6741,6746|false|false|false|C0741025|Chest problem|Chest
Finding|Finding|SIMPLE_SEGMENT|6758,6766|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Intellectual Product|SIMPLE_SEGMENT|6758,6766|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6767,6777|false|false|false|C0225756|Structure of upper lobe of lung|upper lobe
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6773,6777|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|SIMPLE_SEGMENT|6773,6777|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6820,6829|false|false|false|C0034067|Pulmonary Emphysema|emphysema
Event|Event|SIMPLE_SEGMENT|6820,6829|false|false|false|||emphysema
Finding|Pathologic Function|SIMPLE_SEGMENT|6820,6829|false|false|false|C0013990|Pathological accumulation of air in tissues|emphysema
Finding|Finding|SIMPLE_SEGMENT|6835,6838|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|New
Finding|Idea or Concept|SIMPLE_SEGMENT|6835,6838|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|New
Finding|Functional Concept|SIMPLE_SEGMENT|6839,6843|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6839,6854|false|false|false|C1261077|Structure of left lower lobe of lung|left lower lobe
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6844,6849|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|6844,6849|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6844,6854|false|false|false|C0225758|Structure of lower lobe of lung|lower lobe
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6850,6854|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|SIMPLE_SEGMENT|6850,6854|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Event|Event|SIMPLE_SEGMENT|6855,6861|false|false|false|||nodule
Event|Event|SIMPLE_SEGMENT|6875,6884|false|false|false|||measuring
Finding|Gene or Genome|SIMPLE_SEGMENT|6888,6893|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Event|Event|SIMPLE_SEGMENT|6908,6916|false|false|false|||warrants
Finding|Finding|SIMPLE_SEGMENT|6917,6922|false|false|false|C0587267;C3810854|Close;Closed|close
Finding|Functional Concept|SIMPLE_SEGMENT|6917,6922|false|false|false|C0587267;C3810854|Close;Closed|close
Event|Event|SIMPLE_SEGMENT|6923,6929|false|false|false|||follow
Finding|Functional Concept|SIMPLE_SEGMENT|6923,6929|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|SIMPLE_SEGMENT|6923,6929|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|SIMPLE_SEGMENT|6923,6932|false|false|false|C0589120|Follow-up status|follow-up
Procedure|Health Care Activity|SIMPLE_SEGMENT|6923,6932|false|false|false|C1522577|follow-up|follow-up
Event|Event|SIMPLE_SEGMENT|6930,6932|false|false|false|||up
Event|Event|SIMPLE_SEGMENT|6935,6941|false|false|false|||Stable
Finding|Intellectual Product|SIMPLE_SEGMENT|6935,6941|false|false|false|C1547311|Patient Condition Code - Stable|Stable
Finding|Functional Concept|SIMPLE_SEGMENT|6968,6973|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6968,6985|false|false|false|C4281590|Structure of middle lobe of right lung|right middle lobe
Finding|Intellectual Product|SIMPLE_SEGMENT|6974,6980|false|false|false|C1552826|Table Cell Vertical Align - middle|middle
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6974,6985|false|false|false|C4281590|Structure of middle lobe of right lung|middle lobe
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6981,6985|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|SIMPLE_SEGMENT|6981,6985|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Event|Event|SIMPLE_SEGMENT|6986,6992|false|false|false|||nodule
Finding|Finding|SIMPLE_SEGMENT|6998,7004|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|Severe
Finding|Intellectual Product|SIMPLE_SEGMENT|6998,7004|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|Severe
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7005,7013|false|false|false|C0018787|Heart|coronary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7005,7020|false|false|false|C0205042|Coronary artery|coronary artery
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7014,7020|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|SIMPLE_SEGMENT|7014,7020|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Event|Event|SIMPLE_SEGMENT|7021,7035|false|false|false|||calcifications
Finding|Finding|SIMPLE_SEGMENT|7021,7035|false|false|false|C0006660;C2242558|Pathologic calcification, calcified structure;Physiologic calcification|calcifications
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|7021,7035|false|false|false|C0006660;C2242558|Pathologic calcification, calcified structure;Physiologic calcification|calcifications
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7038,7044|false|false|false|C0003483|Aorta|Aortic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7038,7050|false|false|false|C0003501;C4533215|Aortic valve structure;Chest>Aortic valve|Aortic valve
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7045,7050|false|false|false|C1186983|Anatomical valve|valve
Event|Event|SIMPLE_SEGMENT|7052,7066|false|false|false|||calcifications
Finding|Finding|SIMPLE_SEGMENT|7052,7066|false|false|false|C0006660;C2242558|Pathologic calcification, calcified structure;Physiologic calcification|calcifications
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|7052,7066|false|false|false|C0006660;C2242558|Pathologic calcification, calcified structure;Physiologic calcification|calcifications
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|7073,7084|false|false|false|C2711450|Enlargement (morphologic abnormality)|Enlargement
Event|Event|SIMPLE_SEGMENT|7073,7084|false|false|false|||Enlargement
Finding|Pathologic Function|SIMPLE_SEGMENT|7073,7084|false|false|false|C0020564|Hypertrophy|Enlargement
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7073,7084|false|false|false|C1293134|Enlargement procedure|Enlargement
Finding|Functional Concept|SIMPLE_SEGMENT|7101,7106|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7101,7125|false|false|false|C0226054|Right pulmonary artery|right pulmonary arteries
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7107,7116|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7107,7116|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|7107,7116|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7107,7125|false|false|false|C0034052|Pulmonary artery structure|pulmonary arteries
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7117,7125|false|false|false|C0003842;C0226004|Arterial system;Arteries|arteries
Anatomy|Body System|SIMPLE_SEGMENT|7117,7125|false|false|false|C0003842;C0226004|Arterial system;Arteries|arteries
Procedure|Health Care Activity|SIMPLE_SEGMENT|7117,7125|false|false|false|C0397581|Procedure on artery|arteries
Event|Event|SIMPLE_SEGMENT|7130,7140|false|false|false|||suggestive
Finding|Functional Concept|SIMPLE_SEGMENT|7130,7140|false|false|false|C0332299|Suggestive of|suggestive
Finding|Functional Concept|SIMPLE_SEGMENT|7130,7143|false|false|false|C0332299|Suggestive of|suggestive of
Event|Event|SIMPLE_SEGMENT|7144,7151|false|false|false|||chronic
Finding|Intellectual Product|SIMPLE_SEGMENT|7144,7151|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|7144,7151|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7152,7161|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7152,7161|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|7152,7161|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7152,7183|false|false|false|C2973725;C3203102|Idiopathic pulmonary arterial hypertension;Pulmonary arterial hypertension|pulmonary arterial hypertension
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7162,7170|false|false|false|C0003842|Arteries|arterial
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7162,7183|false|false|false|C0020538|Hypertensive disease|arterial hypertension
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7171,7183|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|SIMPLE_SEGMENT|7171,7183|false|false|false|||hypertension
Finding|Pathologic Function|SIMPLE_SEGMENT|7199,7220|false|false|false|C0002940|Aneurysm|aneurysmal dilatation
Event|Event|SIMPLE_SEGMENT|7210,7220|false|false|false|||dilatation
Finding|Finding|SIMPLE_SEGMENT|7210,7220|false|false|false|C0012359;C0700124|Dilated;Pathological Dilatation|dilatation
Finding|Pathologic Function|SIMPLE_SEGMENT|7210,7220|false|false|false|C0012359;C0700124|Dilated;Pathological Dilatation|dilatation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7210,7220|false|false|false|C1322279|Dilate procedure|dilatation
Finding|Finding|SIMPLE_SEGMENT|7210,7243|false|true|false|C4025248|Dilatation of the abdominal aorta|dilatation of the abdominal aorta
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7228,7237|false|false|false|C0000726|Abdomen|abdominal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7228,7243|false|false|false|C0003484;C4037989|Abdomen>Aorta.abdominal;Abdominal aorta structure|abdominal aorta
Procedure|Health Care Activity|SIMPLE_SEGMENT|7228,7243|false|false|false|C2228415|examination of abdominal aorta|abdominal aorta
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7238,7243|false|false|false|C0003483;C4037978|Aorta;Chest+Abdomen>Aorta|aorta
Procedure|Health Care Activity|SIMPLE_SEGMENT|7238,7243|false|false|false|C0869784|Procedure on aorta|aorta
Event|Event|SIMPLE_SEGMENT|7245,7254|false|false|false|||measuring
Event|Event|SIMPLE_SEGMENT|7272,7282|false|false|false|||progressed
Event|Event|SIMPLE_SEGMENT|7283,7291|false|false|false|||compared
Event|Activity|SIMPLE_SEGMENT|7302,7313|false|false|false|C4321457|Examination|examination
Event|Event|SIMPLE_SEGMENT|7302,7313|false|false|false|||examination
Procedure|Health Care Activity|SIMPLE_SEGMENT|7302,7313|false|false|false|C0031809;C0582103|Medical Examination;Physical Examination|examination
Finding|Body Substance|SIMPLE_SEGMENT|7334,7343|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|7334,7343|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|7334,7343|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|7334,7343|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|SIMPLE_SEGMENT|7344,7348|false|false|false|||LABS
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|7344,7348|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7381,7386|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|7381,7386|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|7381,7386|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|7387,7390|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|7395,7398|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7395,7398|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7395,7398|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7404,7407|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7404,7407|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|7404,7407|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|7404,7407|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7413,7416|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7413,7416|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|7422,7425|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|7422,7425|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|7422,7425|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7422,7425|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7422,7425|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|7430,7433|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7430,7433|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|7430,7433|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|7430,7433|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|7430,7433|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7430,7433|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|SIMPLE_SEGMENT|7439,7443|false|false|false|||MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7439,7443|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7472,7475|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7492,7497|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|7492,7497|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|7492,7497|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|7492,7505|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|7492,7505|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7492,7505|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7498,7505|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|7498,7505|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7498,7505|false|false|false|C0017725|glucose|Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|7498,7505|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7498,7505|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|SIMPLE_SEGMENT|7549,7553|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7549,7553|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7549,7553|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7578,7583|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|7578,7583|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|7578,7583|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7578,7591|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7584,7591|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|7584,7591|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|7584,7591|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7584,7591|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|7584,7591|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|SIMPLE_SEGMENT|7584,7591|false|false|false|||Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|7584,7591|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7584,7591|false|false|false|C0201925|Calcium measurement|Calcium
Finding|Intellectual Product|SIMPLE_SEGMENT|7614,7619|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|Brief
Finding|Idea or Concept|SIMPLE_SEGMENT|7620,7628|false|false|false|C1547192|Organization unit type - Hospital|Hospital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7620,7635|false|false|false|C0488549||Hospital Course
Finding|Finding|SIMPLE_SEGMENT|7620,7635|false|false|false|C0489547|Hospital course|Hospital Course
Event|Event|SIMPLE_SEGMENT|7671,7674|false|false|false|||PMH
Finding|Finding|SIMPLE_SEGMENT|7671,7674|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|PMH
Event|Event|SIMPLE_SEGMENT|7675,7682|false|false|false|||notable
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7687,7691|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7687,7691|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|SIMPLE_SEGMENT|7687,7691|false|false|false|||COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|7687,7691|false|false|false|C1412502|ARCN1 gene|COPD
Finding|Idea or Concept|SIMPLE_SEGMENT|7696,7700|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|7696,7700|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|7696,7700|false|false|false|C1553498|home health encounter|home
Event|Event|SIMPLE_SEGMENT|7705,7717|false|false|false|||hospitalized
Event|Event|SIMPLE_SEGMENT|7742,7748|false|false|false|||visits
Finding|Social Behavior|SIMPLE_SEGMENT|7742,7748|false|false|false|C0545082|Visit|visits
Procedure|Health Care Activity|SIMPLE_SEGMENT|7742,7748|false|false|false|C1512346|Patient Visit|visits
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7751,7755|false|false|false|C0004238|Atrial Fibrillation|Afib
Event|Event|SIMPLE_SEGMENT|7751,7755|false|false|false|||Afib
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|7751,7755|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Afib
Drug|Organic Chemical|SIMPLE_SEGMENT|7760,7768|false|false|false|C1831808|apixaban|apixaban
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7760,7768|false|false|false|C1831808|apixaban|apixaban
Event|Event|SIMPLE_SEGMENT|7760,7768|false|false|false|||apixaban
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7770,7773|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|SIMPLE_SEGMENT|7770,7773|false|false|false|||HTN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7775,7778|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7775,7778|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|7775,7778|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|7775,7778|false|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|7775,7778|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7775,7778|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|7775,7778|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7775,7778|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Event|Event|SIMPLE_SEGMENT|7784,7787|false|false|false|||HLD
Event|Event|SIMPLE_SEGMENT|7792,7801|false|false|false|||presented
Event|Event|SIMPLE_SEGMENT|7807,7814|false|false|false|||dyspnea
Finding|Finding|SIMPLE_SEGMENT|7807,7814|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|7807,7814|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Event|Event|SIMPLE_SEGMENT|7820,7829|false|false|false|||orthopnea
Finding|Finding|SIMPLE_SEGMENT|7820,7829|false|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|7820,7829|false|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Finding|Mental Process|SIMPLE_SEGMENT|7837,7844|false|false|false|C0542559|contextual factors|setting
Drug|Organic Chemical|SIMPLE_SEGMENT|7850,7857|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7850,7857|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Event|Event|SIMPLE_SEGMENT|7858,7863|false|false|false|||taper
Procedure|Health Care Activity|SIMPLE_SEGMENT|7858,7863|false|false|false|C0441640||taper
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7875,7879|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7875,7879|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|SIMPLE_SEGMENT|7875,7879|false|false|false|||COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|7875,7879|false|false|false|C1412502|ARCN1 gene|COPD
Event|Event|SIMPLE_SEGMENT|7881,7893|false|false|false|||exacerbation
Finding|Finding|SIMPLE_SEGMENT|7881,7893|false|false|false|C4086268|Exacerbation|exacerbation
Event|Event|SIMPLE_SEGMENT|7899,7906|false|false|false|||dyspnea
Finding|Finding|SIMPLE_SEGMENT|7899,7906|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|7899,7906|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Event|Event|SIMPLE_SEGMENT|7911,7918|false|false|false|||thought
Finding|Finding|SIMPLE_SEGMENT|7925,7939|false|false|false|C1837655|Multifactorial|multifactorial
Event|Event|SIMPLE_SEGMENT|7940,7943|false|false|false|||due
Finding|Functional Concept|SIMPLE_SEGMENT|7940,7943|false|false|false|C0678226;C3146286|Due;Due to|due
Finding|Idea or Concept|SIMPLE_SEGMENT|7940,7943|false|false|false|C0678226;C3146286|Due;Due to|due
Finding|Finding|SIMPLE_SEGMENT|7952,7958|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|SIMPLE_SEGMENT|7952,7958|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7959,7963|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7959,7963|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|SIMPLE_SEGMENT|7959,7963|false|false|false|||COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|7959,7963|false|false|false|C1412502|ARCN1 gene|COPD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7975,7984|false|false|false|C1179435|Protein Component|component
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7975,7984|false|false|false|C1179435|Protein Component|component
Event|Event|SIMPLE_SEGMENT|7975,7984|false|false|false|||component
Finding|Conceptual Entity|SIMPLE_SEGMENT|7975,7984|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Finding|Idea or Concept|SIMPLE_SEGMENT|7975,7984|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Finding|Intellectual Product|SIMPLE_SEGMENT|7975,7984|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|7988,7995|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Event|Event|SIMPLE_SEGMENT|7988,7995|false|false|false|||anxiety
Finding|Sign or Symptom|SIMPLE_SEGMENT|7988,7995|false|false|false|C0860603|Anxiety symptoms|anxiety
Finding|Body Substance|SIMPLE_SEGMENT|8001,8008|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|8001,8008|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|8001,8008|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|8018,8025|true|false|false|||thought
Finding|Intellectual Product|SIMPLE_SEGMENT|8042,8047|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8042,8065|true|false|false|C0340044|Acute exacerbation of chronic obstructive pulmonary disease|acute COPD exacerbation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8048,8052|true|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8048,8052|true|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|SIMPLE_SEGMENT|8048,8052|true|false|false|||COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|8048,8052|true|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8048,8065|true|false|false|C0740304|COPD exacerbation|COPD exacerbation
Event|Event|SIMPLE_SEGMENT|8053,8065|false|false|false|||exacerbation
Finding|Finding|SIMPLE_SEGMENT|8053,8065|false|false|false|C4086268|Exacerbation|exacerbation
Event|Event|SIMPLE_SEGMENT|8092,8098|false|false|false|||ISSUES
Finding|Finding|SIMPLE_SEGMENT|8120,8127|false|false|false|C0013404;C2024878|Dyspnea|Dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|8120,8127|false|false|false|C0013404;C2024878|Dyspnea|Dyspnea
Finding|Body Substance|SIMPLE_SEGMENT|8129,8136|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|8129,8136|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|8129,8136|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|8141,8149|false|false|false|||admitted
Event|Event|SIMPLE_SEGMENT|8169,8177|false|false|false|||worsened
Finding|Finding|SIMPLE_SEGMENT|8169,8177|false|false|false|C1457868;C4084902|Got Worse;Worse|worsened
Finding|Intellectual Product|SIMPLE_SEGMENT|8169,8177|false|false|false|C1457868;C4084902|Got Worse;Worse|worsened
Event|Event|SIMPLE_SEGMENT|8179,8188|false|false|false|||orthopnea
Finding|Finding|SIMPLE_SEGMENT|8179,8188|false|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|8179,8188|false|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Event|Event|SIMPLE_SEGMENT|8193,8200|false|false|false|||dyspnea
Finding|Finding|SIMPLE_SEGMENT|8193,8200|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|8193,8200|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Mental Process|SIMPLE_SEGMENT|8208,8215|false|false|false|C0542559|contextual factors|setting
Drug|Organic Chemical|SIMPLE_SEGMENT|8221,8228|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8221,8228|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Event|Event|SIMPLE_SEGMENT|8229,8234|false|false|false|||taper
Procedure|Health Care Activity|SIMPLE_SEGMENT|8229,8234|false|false|false|C0441640||taper
Event|Event|SIMPLE_SEGMENT|8261,8268|false|false|false|||dyspnea
Finding|Finding|SIMPLE_SEGMENT|8261,8268|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|8261,8268|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Event|Event|SIMPLE_SEGMENT|8273,8280|false|false|false|||thought
Event|Event|SIMPLE_SEGMENT|8287,8301|false|false|false|||multifactorial
Finding|Finding|SIMPLE_SEGMENT|8287,8301|false|false|false|C1837655|Multifactorial|multifactorial
Finding|Finding|SIMPLE_SEGMENT|8314,8320|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|SIMPLE_SEGMENT|8314,8320|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8321,8325|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8321,8325|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|SIMPLE_SEGMENT|8321,8325|false|false|false|||COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|8321,8325|false|false|false|C1412502|ARCN1 gene|COPD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8337,8346|false|false|false|C1179435|Protein Component|component
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8337,8346|false|false|false|C1179435|Protein Component|component
Event|Event|SIMPLE_SEGMENT|8337,8346|false|false|false|||component
Finding|Conceptual Entity|SIMPLE_SEGMENT|8337,8346|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Finding|Idea or Concept|SIMPLE_SEGMENT|8337,8346|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Finding|Intellectual Product|SIMPLE_SEGMENT|8337,8346|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|8350,8357|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Event|Event|SIMPLE_SEGMENT|8350,8357|false|false|false|||anxiety
Finding|Sign or Symptom|SIMPLE_SEGMENT|8350,8357|false|false|false|C0860603|Anxiety symptoms|anxiety
Finding|Body Substance|SIMPLE_SEGMENT|8363,8370|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|8363,8370|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|8363,8370|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|8380,8387|true|false|false|||thought
Finding|Intellectual Product|SIMPLE_SEGMENT|8404,8409|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8404,8427|true|false|false|C0340044|Acute exacerbation of chronic obstructive pulmonary disease|acute COPD exacerbation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8410,8414|true|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8410,8414|true|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|SIMPLE_SEGMENT|8410,8414|true|false|false|||COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|8410,8414|true|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8410,8427|true|false|false|C0740304|COPD exacerbation|COPD exacerbation
Event|Event|SIMPLE_SEGMENT|8415,8427|false|false|false|||exacerbation
Finding|Finding|SIMPLE_SEGMENT|8415,8427|false|false|false|C4086268|Exacerbation|exacerbation
Finding|Body Substance|SIMPLE_SEGMENT|8433,8440|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|8433,8440|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|8433,8440|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|8446,8453|false|false|false|||treated
Event|Event|SIMPLE_SEGMENT|8470,8477|false|false|false|||duonebs
Drug|Organic Chemical|SIMPLE_SEGMENT|8482,8491|false|false|false|C0024002|lorazepam|lorazepam
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8482,8491|false|false|false|C0024002|lorazepam|lorazepam
Event|Event|SIMPLE_SEGMENT|8482,8491|false|false|false|||lorazepam
Event|Event|SIMPLE_SEGMENT|8499,8502|false|false|false|||PRN
Finding|Gene or Genome|SIMPLE_SEGMENT|8499,8502|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|SIMPLE_SEGMENT|8509,8515|false|false|false|||helped
Event|Event|SIMPLE_SEGMENT|8516,8523|false|false|false|||relieve
Event|Event|SIMPLE_SEGMENT|8528,8535|false|false|false|||dyspnea
Finding|Finding|SIMPLE_SEGMENT|8528,8535|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|8528,8535|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Event|Event|SIMPLE_SEGMENT|8537,8548|false|false|false|||Pulmonology
Event|Event|SIMPLE_SEGMENT|8553,8562|false|false|false|||consulted
Finding|Body Substance|SIMPLE_SEGMENT|8569,8576|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|8569,8576|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|8569,8576|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|8587,8589|false|false|false|||CT
Event|Event|SIMPLE_SEGMENT|8595,8601|false|false|false|||showed
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8602,8611|false|false|false|C0034067|Pulmonary Emphysema|emphysema
Event|Event|SIMPLE_SEGMENT|8602,8611|false|false|false|||emphysema
Finding|Pathologic Function|SIMPLE_SEGMENT|8602,8611|false|false|false|C0013990|Pathological accumulation of air in tissues|emphysema
Event|Event|SIMPLE_SEGMENT|8619,8627|true|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|8619,8627|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|8619,8630|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8632,8641|true|false|false|C0009450|Communicable Diseases|infection
Event|Event|SIMPLE_SEGMENT|8632,8641|true|false|false|||infection
Finding|Pathologic Function|SIMPLE_SEGMENT|8632,8641|true|false|false|C3714514|Infection|infection
Finding|Body Substance|SIMPLE_SEGMENT|8659,8666|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|8659,8666|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|8659,8666|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|8671,8680|false|false|false|||initiated
Drug|Organic Chemical|SIMPLE_SEGMENT|8686,8693|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8686,8693|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Event|Event|SIMPLE_SEGMENT|8686,8693|false|false|false|||steroid
Event|Event|SIMPLE_SEGMENT|8695,8700|false|false|false|||taper
Drug|Hormone|SIMPLE_SEGMENT|8711,8721|false|false|false|C0032952|prednisone|prednisone
Drug|Organic Chemical|SIMPLE_SEGMENT|8711,8721|false|false|false|C0032952|prednisone|prednisone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8711,8721|false|false|false|C0032952|prednisone|prednisone
Finding|Intellectual Product|SIMPLE_SEGMENT|8740,8744|false|false|false|C1720594|Then - dosing instruction fragment|then
Finding|Intellectual Product|SIMPLE_SEGMENT|8764,8768|false|false|false|C1720594|Then - dosing instruction fragment|then
Finding|Classification|SIMPLE_SEGMENT|8781,8791|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|8781,8791|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|SIMPLE_SEGMENT|8792,8798|false|false|false|||follow
Finding|Functional Concept|SIMPLE_SEGMENT|8792,8798|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|SIMPLE_SEGMENT|8792,8798|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|SIMPLE_SEGMENT|8792,8801|false|false|false|C0589120|Follow-up status|follow-up
Procedure|Health Care Activity|SIMPLE_SEGMENT|8792,8801|false|false|false|C1522577|follow-up|follow-up
Event|Event|SIMPLE_SEGMENT|8816,8827|false|false|false|||recommended
Event|Event|SIMPLE_SEGMENT|8828,8838|false|false|false|||increasing
Drug|Organic Chemical|SIMPLE_SEGMENT|8843,8849|false|false|false|C0965130|Advair|Advair
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8843,8849|false|false|false|C0965130|Advair|Advair
Event|Event|SIMPLE_SEGMENT|8850,8854|false|false|false|||dose
Event|Event|SIMPLE_SEGMENT|8893,8904|false|false|false|||recommended
Event|Event|SIMPLE_SEGMENT|8905,8914|false|false|false|||switching
Drug|Organic Chemical|SIMPLE_SEGMENT|8920,8932|false|false|false|C0039771|theophylline|theophylline
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8920,8932|false|false|false|C0039771|theophylline|theophylline
Event|Event|SIMPLE_SEGMENT|8920,8932|false|false|false|||theophylline
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8920,8932|false|false|false|C0039773|Assay of theophylline|theophylline
Drug|Organic Chemical|SIMPLE_SEGMENT|8937,8948|false|false|false|C0965618|roflumilast|roflumilast
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8937,8948|false|false|false|C0965618|roflumilast|roflumilast
Event|Event|SIMPLE_SEGMENT|8937,8948|false|false|false|||roflumilast
Event|Event|SIMPLE_SEGMENT|8953,8963|false|false|false|||initiation
Finding|Functional Concept|SIMPLE_SEGMENT|8953,8963|false|false|false|C0589507;C1158830;C1704686|Initiation;Transcription Initiation|initiation
Finding|Genetic Function|SIMPLE_SEGMENT|8953,8963|false|false|false|C0589507;C1158830;C1704686|Initiation;Transcription Initiation|initiation
Finding|Mental Process|SIMPLE_SEGMENT|8953,8963|false|false|false|C0589507;C1158830;C1704686|Initiation;Transcription Initiation|initiation
Finding|Idea or Concept|SIMPLE_SEGMENT|8972,8976|false|false|false|C0233324;C1705313|Term (lexical);Term Birth|term
Finding|Organism Function|SIMPLE_SEGMENT|8972,8976|false|false|false|C0233324;C1705313|Term (lexical);Term Birth|term
Drug|Antibiotic|SIMPLE_SEGMENT|8977,8989|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Clinical Drug|SIMPLE_SEGMENT|8977,8989|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Organic Chemical|SIMPLE_SEGMENT|8977,8989|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Event|Event|SIMPLE_SEGMENT|8990,8997|false|false|false|||therapy
Finding|Finding|SIMPLE_SEGMENT|8990,8997|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|SIMPLE_SEGMENT|8990,8997|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8990,8997|false|false|false|C0087111|Therapeutic procedure|therapy
Event|Event|SIMPLE_SEGMENT|8999,9007|true|false|false|||provided
Finding|Body Substance|SIMPLE_SEGMENT|9012,9019|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|9012,9019|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|9012,9019|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|9034,9043|true|false|false|||prolonged
Event|Event|SIMPLE_SEGMENT|9054,9062|false|false|false|||deferred
Finding|Classification|SIMPLE_SEGMENT|9071,9081|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|9071,9081|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|SIMPLE_SEGMENT|9082,9089|false|false|false|||setting
Finding|Mental Process|SIMPLE_SEGMENT|9082,9089|false|false|false|C0542559|contextual factors|setting
Event|Event|SIMPLE_SEGMENT|9106,9115|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|9106,9115|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9128,9132|false|false|false|C0312448|short-acting thyroid stimulator|sats
Drug|Hormone|SIMPLE_SEGMENT|9128,9132|false|false|false|C0312448|short-acting thyroid stimulator|sats
Event|Event|SIMPLE_SEGMENT|9128,9132|false|false|false|||sats
Event|Event|SIMPLE_SEGMENT|9156,9158|false|false|false|||NC
Event|Event|SIMPLE_SEGMENT|9172,9182|true|false|false|||desaturate
Event|Event|SIMPLE_SEGMENT|9187,9197|true|false|false|||ambulation
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|9187,9197|true|false|false|C0080331;C0945826|Ambulation;Walking (function)|ambulation
Finding|Functional Concept|SIMPLE_SEGMENT|9187,9197|true|false|false|C0080331;C0945826|Ambulation;Walking (function)|ambulation
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|9203,9210|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|Anxiety
Event|Event|SIMPLE_SEGMENT|9203,9210|false|false|false|||Anxiety
Finding|Sign or Symptom|SIMPLE_SEGMENT|9203,9210|false|false|false|C0860603|Anxiety symptoms|Anxiety
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9211,9219|false|false|false|C1950154|Insomnia homeopathic medication|Insomnia
Event|Event|SIMPLE_SEGMENT|9211,9219|false|false|false|||Insomnia
Finding|Sign or Symptom|SIMPLE_SEGMENT|9211,9219|false|false|false|C0917801|Sleeplessness|Insomnia
Finding|Body Substance|SIMPLE_SEGMENT|9221,9228|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|9221,9228|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|9221,9228|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|9236,9243|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|9236,9243|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|9236,9243|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|9236,9243|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|9236,9246|false|false|false|C0262926|Medical History|history of
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|9247,9254|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Event|Event|SIMPLE_SEGMENT|9247,9254|false|false|false|||anxiety
Finding|Sign or Symptom|SIMPLE_SEGMENT|9247,9254|false|false|false|C0860603|Anxiety symptoms|anxiety
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9260,9268|false|false|false|C1950154|Insomnia homeopathic medication|insomnia
Event|Event|SIMPLE_SEGMENT|9260,9268|false|false|false|||insomnia
Finding|Sign or Symptom|SIMPLE_SEGMENT|9260,9268|false|false|false|C0917801|Sleeplessness|insomnia
Event|Event|SIMPLE_SEGMENT|9270,9277|false|false|false|||thought
Finding|Idea or Concept|SIMPLE_SEGMENT|9270,9277|false|false|false|C0039869;C4319827|Thought|thought
Finding|Mental Process|SIMPLE_SEGMENT|9270,9277|false|false|false|C0039869;C4319827|Thought|thought
Event|Event|SIMPLE_SEGMENT|9284,9296|false|false|false|||contributing
Finding|Mental Process|SIMPLE_SEGMENT|9304,9314|false|false|false|C0237607;C0596545|Experience;Experience (Practice)|experience
Event|Event|SIMPLE_SEGMENT|9319,9326|false|false|false|||dyspnea
Finding|Finding|SIMPLE_SEGMENT|9319,9326|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|9319,9326|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Body Substance|SIMPLE_SEGMENT|9332,9339|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|9332,9339|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|9332,9339|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|9344,9354|false|false|false|||discharged
Drug|Organic Chemical|SIMPLE_SEGMENT|9360,9369|false|false|false|C0024002|lorazepam|lorazepam
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9360,9369|false|false|false|C0024002|lorazepam|lorazepam
Event|Event|SIMPLE_SEGMENT|9360,9369|false|false|false|||lorazepam
Event|Event|SIMPLE_SEGMENT|9377,9383|false|false|false|||needed
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|9389,9396|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Event|Event|SIMPLE_SEGMENT|9389,9396|false|false|false|||anxiety
Finding|Sign or Symptom|SIMPLE_SEGMENT|9389,9396|false|false|false|C0860603|Anxiety symptoms|anxiety
Finding|Body Substance|SIMPLE_SEGMENT|9402,9409|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|9402,9409|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|9402,9409|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Finding|SIMPLE_SEGMENT|9416,9422|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|9416,9422|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|SIMPLE_SEGMENT|9423,9430|false|false|false|||benefit
Event|Event|SIMPLE_SEGMENT|9436,9443|false|false|false|||therapy
Finding|Finding|SIMPLE_SEGMENT|9436,9443|false|true|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|SIMPLE_SEGMENT|9436,9443|false|true|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9436,9443|false|true|false|C0087111|Therapeutic procedure|therapy
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9453,9457|false|false|false|C0360105;C2911696|Selective Serotonin Reuptake Inhibitors;Serotonin Reuptake Inhibitor [EPC]|SSRI
Event|Event|SIMPLE_SEGMENT|9453,9457|false|false|false|||SSRI
Finding|Idea or Concept|SIMPLE_SEGMENT|9462,9468|false|false|false|C0699784|Economic demand|Demand
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9462,9468|false|false|false|C0441516|Demand (clinical)|Demand
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9462,9477|false|false|false|C4049375|Ischemia co-occurrent and due to increased oxygen demand|Demand Ischemia
Event|Event|SIMPLE_SEGMENT|9469,9477|false|false|false|||Ischemia
Finding|Pathologic Function|SIMPLE_SEGMENT|9469,9477|false|false|false|C0022116|Ischemia|Ischemia
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9469,9477|false|false|false|C4321499|Ischemia Procedure|Ischemia
Finding|Body Substance|SIMPLE_SEGMENT|9479,9486|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|9479,9486|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|9479,9486|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9492,9500|false|false|false|C0041199|Troponin|troponin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9492,9500|false|false|false|C0041199|Troponin|troponin
Event|Event|SIMPLE_SEGMENT|9492,9500|false|false|false|||troponin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9492,9500|false|false|false|C0523952|Troponin measurement|troponin
Finding|Intellectual Product|SIMPLE_SEGMENT|9514,9518|false|false|false|C1720594|Then - dosing instruction fragment|then
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9526,9529|true|false|false|C0018064|Equine Gonadotropins|ECG
Drug|Hormone|SIMPLE_SEGMENT|9526,9529|true|false|false|C0018064|Equine Gonadotropins|ECG
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9526,9529|true|false|false|C0018064|Equine Gonadotropins|ECG
Event|Event|SIMPLE_SEGMENT|9526,9529|true|false|false|||ECG
Finding|Intellectual Product|SIMPLE_SEGMENT|9526,9529|true|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|ECG
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|9526,9529|true|false|false|C1623258|Electrocardiography|ECG
Event|Event|SIMPLE_SEGMENT|9538,9543|true|false|false|||acute
Finding|Intellectual Product|SIMPLE_SEGMENT|9538,9543|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Functional Concept|SIMPLE_SEGMENT|9544,9552|true|false|false|C0475224|Ischemic|ischemic
Event|Event|SIMPLE_SEGMENT|9553,9560|true|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|9553,9560|true|false|false|C0392747|Changing|changes
Finding|Finding|SIMPLE_SEGMENT|9565,9586|false|false|false|C0239937|Microscopic hematuria|Microscopic hematuria
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9577,9586|false|false|false|C0018965|Hematuria|hematuria
Event|Event|SIMPLE_SEGMENT|9577,9586|false|false|false|||hematuria
Event|Event|SIMPLE_SEGMENT|9591,9600|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|9591,9600|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Body Substance|SIMPLE_SEGMENT|9605,9612|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|9605,9612|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|9605,9612|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|9619,9621|false|false|false|||UA
Anatomy|Cell|SIMPLE_SEGMENT|9631,9635|false|false|false|C0014792|Erythrocytes|RBCs
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9631,9635|false|false|false|C0014792|Erythrocytes|RBCs
Finding|Idea or Concept|SIMPLE_SEGMENT|9666,9670|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|SIMPLE_SEGMENT|9666,9670|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Event|Event|SIMPLE_SEGMENT|9674,9677|false|false|false|||OMR
Finding|Gene or Genome|SIMPLE_SEGMENT|9674,9677|false|false|false|C1412647|ATP5F1A gene|OMR
Finding|Finding|SIMPLE_SEGMENT|9684,9705|false|false|false|C0239937|Microscopic hematuria|microscopic hematuria
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9696,9705|false|false|false|C0018965|Hematuria|hematuria
Event|Event|SIMPLE_SEGMENT|9696,9705|false|false|false|||hematuria
Event|Event|SIMPLE_SEGMENT|9713,9722|false|false|false|||recommend
Event|Event|SIMPLE_SEGMENT|9723,9729|false|false|false|||repeat
Finding|Functional Concept|SIMPLE_SEGMENT|9723,9729|false|false|false|C0205341;C1705914|Repeat;Repeat Object|repeat
Event|Event|SIMPLE_SEGMENT|9740,9750|false|false|false|||outpatient
Finding|Classification|SIMPLE_SEGMENT|9740,9750|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|9740,9750|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|SIMPLE_SEGMENT|9754,9758|false|false|false|||work
Event|Occupational Activity|SIMPLE_SEGMENT|9754,9758|false|false|false|C0043227|Work|work
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|9754,9761|false|false|false|C0750430|Work-up|work-up
Event|Event|SIMPLE_SEGMENT|9759,9761|false|false|false|||up
Finding|Finding|SIMPLE_SEGMENT|9766,9787|false|false|false|C0239937|Microscopic hematuria|microscopic hematuria
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9778,9787|false|false|false|C0018965|Hematuria|hematuria
Event|Event|SIMPLE_SEGMENT|9778,9787|false|false|false|||hematuria
Event|Event|SIMPLE_SEGMENT|9807,9814|false|false|false|||CHRONIC
Finding|Intellectual Product|SIMPLE_SEGMENT|9807,9814|false|false|false|C1547296|Chronic - Admission Level of Care Code|CHRONIC
Procedure|Health Care Activity|SIMPLE_SEGMENT|9807,9814|false|false|false|C1555457|Provision of recurring care for chronic illness|CHRONIC
Finding|Individual Behavior|SIMPLE_SEGMENT|9843,9850|false|false|false|C0037369;C0453996;C1548578|Location characteristic ID - Smoking;Smoking;Tobacco smoking behavior|Smoking
Finding|Intellectual Product|SIMPLE_SEGMENT|9843,9850|false|false|false|C0037369;C0453996;C1548578|Location characteristic ID - Smoking;Smoking;Tobacco smoking behavior|Smoking
Finding|Body Substance|SIMPLE_SEGMENT|9852,9859|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|9852,9859|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|9852,9859|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|9869,9873|false|false|false|||quit
Event|Event|SIMPLE_SEGMENT|9874,9881|false|false|false|||smoking
Finding|Idea or Concept|SIMPLE_SEGMENT|9886,9891|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Intellectual Product|SIMPLE_SEGMENT|9886,9891|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Gene or Genome|SIMPLE_SEGMENT|9892,9895|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Finding|Body Substance|SIMPLE_SEGMENT|9897,9904|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|9897,9904|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|9897,9904|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|9910,9918|false|false|false|||provided
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|9926,9934|false|false|false|C0028040|nicotine|nicotine
Drug|Organic Chemical|SIMPLE_SEGMENT|9926,9934|false|false|false|C0028040|nicotine|nicotine
Drug|Clinical Drug|SIMPLE_SEGMENT|9926,9940|false|false|false|C0358855|Nicotine Transdermal Patch|nicotine patch
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9935,9940|false|false|false|C0445403;C1533128;C1707974|Body tissue patch material;Human patch material;Patch - Extended Release Film|patch
Event|Event|SIMPLE_SEGMENT|9935,9940|false|false|false|||patch
Finding|Finding|SIMPLE_SEGMENT|9935,9940|false|false|false|C0332461|Plaque (lesion)|patch
Event|Event|SIMPLE_SEGMENT|9969,9977|false|false|false|||consider
Event|Event|SIMPLE_SEGMENT|9978,9988|false|false|false|||continuing
Event|Event|SIMPLE_SEGMENT|9995,10005|false|false|false|||outpatient
Finding|Classification|SIMPLE_SEGMENT|9995,10005|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|9995,10005|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Body Substance|SIMPLE_SEGMENT|10009,10016|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|10009,10016|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|10009,10016|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|10027,10035|false|false|false|||cravings
Finding|Individual Behavior|SIMPLE_SEGMENT|10027,10035|false|false|false|C0870371|Craving|cravings
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10040,10046|false|false|false|C0018792|Heart Atrium|Atrial
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10040,10059|false|false|false|C2926591||Atrial fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10040,10059|false|false|false|C0004238|Atrial Fibrillation|Atrial fibrillation
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|10040,10059|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Atrial fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10047,10059|false|false|false|C0232197|Fibrillation|fibrillation
Event|Event|SIMPLE_SEGMENT|10047,10059|false|false|false|||fibrillation
Finding|Body Substance|SIMPLE_SEGMENT|10061,10068|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|10061,10068|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|10061,10068|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|10069,10078|false|false|false|||continued
Drug|Organic Chemical|SIMPLE_SEGMENT|10082,10091|false|false|false|C0012373|diltiazem|diltiazem
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10082,10091|false|false|false|C0012373|diltiazem|diltiazem
Event|Event|SIMPLE_SEGMENT|10082,10091|false|false|false|||diltiazem
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|10103,10106|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10103,10106|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|10103,10106|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|10103,10106|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|10103,10106|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|10111,10119|false|false|false|C1831808|apixaban|apixaban
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10111,10119|false|false|false|C1831808|apixaban|apixaban
Event|Event|SIMPLE_SEGMENT|10111,10119|false|false|false|||apixaban
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|10125,10128|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10125,10128|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|10125,10128|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|10125,10128|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|10125,10128|false|false|false|C1332410|BID gene|BID
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10133,10136|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|SIMPLE_SEGMENT|10133,10136|false|false|false|||HTN
Finding|Body Substance|SIMPLE_SEGMENT|10138,10145|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|10138,10145|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|10138,10145|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|10153,10160|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|10153,10160|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|10153,10160|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|10153,10160|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|10153,10163|false|false|false|C0262926|Medical History|history of
Finding|Finding|SIMPLE_SEGMENT|10153,10176|false|false|false|C0455527||history of hypertension
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10164,10176|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|SIMPLE_SEGMENT|10164,10176|false|false|false|||hypertension
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10178,10183|false|false|false|C0851353|Blood and lymphatic system disorders|Blood
Finding|Body Substance|SIMPLE_SEGMENT|10178,10183|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Finding|Finding|SIMPLE_SEGMENT|10178,10192|false|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|Blood pressure
Finding|Organism Function|SIMPLE_SEGMENT|10178,10192|false|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|Blood pressure
Procedure|Health Care Activity|SIMPLE_SEGMENT|10178,10192|false|false|false|C0005824|Blood pressure determination|Blood pressure
Event|Event|SIMPLE_SEGMENT|10184,10192|false|false|false|||pressure
Finding|Finding|SIMPLE_SEGMENT|10184,10192|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|SIMPLE_SEGMENT|10184,10192|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|10184,10192|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|10184,10192|false|false|false|C0033095||pressure
Finding|Finding|SIMPLE_SEGMENT|10194,10198|false|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|10199,10209|false|false|false|||controlled
Event|Event|SIMPLE_SEGMENT|10211,10220|false|false|false|||Continued
Drug|Organic Chemical|SIMPLE_SEGMENT|10224,10234|false|false|false|C0022251|isosorbide|isosorbide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10224,10234|false|false|false|C0022251|isosorbide|isosorbide
Drug|Organic Chemical|SIMPLE_SEGMENT|10224,10246|false|false|false|C0064079|isosorbide mononitrate|isosorbide mononitrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10224,10246|false|false|false|C0064079|isosorbide mononitrate|isosorbide mononitrate
Event|Event|SIMPLE_SEGMENT|10235,10246|false|false|false|||mononitrate
Drug|Organic Chemical|SIMPLE_SEGMENT|10271,10290|false|false|false|C0020261|hydrochlorothiazide|hydrochlorothiazide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10271,10290|false|false|false|C0020261|hydrochlorothiazide|hydrochlorothiazide
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10310,10313|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10310,10313|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|10310,10313|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|10310,10313|false|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|10310,10313|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10310,10313|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|10310,10313|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10310,10313|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10315,10322|true|false|false|C0018787|Heart|Cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|10315,10322|true|false|false|C1314974|Cardiac attachment|Cardiac
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|10315,10338|true|false|false|C0261588|Cardiac catheterisation as the cause of abnormal reaction of the patient, or of later complication, without mention of misadventure at the time of the procedure|Cardiac catheterization
Finding|Intellectual Product|SIMPLE_SEGMENT|10315,10338|true|false|false|C1547981|Diagnostic Service Section ID - Cardiac Catheterization|Cardiac catheterization
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10315,10338|true|false|false|C0018795;C1548828|Cardiac Catheterization Procedures;Consent Type - Cardiac Catheterization|Cardiac catheterization
Procedure|Health Care Activity|SIMPLE_SEGMENT|10315,10338|true|false|false|C0018795;C1548828|Cardiac Catheterization Procedures;Consent Type - Cardiac Catheterization|Cardiac catheterization
Event|Event|SIMPLE_SEGMENT|10323,10338|true|false|false|||catheterization
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10323,10338|true|false|false|C0007430|Catheterization|catheterization
Event|Event|SIMPLE_SEGMENT|10354,10362|true|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|10354,10362|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|10354,10365|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Finding|Idea or Concept|SIMPLE_SEGMENT|10367,10378|true|false|false|C0750502|Significant|significant
Event|Event|SIMPLE_SEGMENT|10379,10387|true|false|false|||stenosis
Finding|Pathologic Function|SIMPLE_SEGMENT|10379,10387|true|false|false|C1261287|Stenosis|stenosis
Event|Event|SIMPLE_SEGMENT|10391,10401|true|false|false|||coronaries
Event|Event|SIMPLE_SEGMENT|10403,10407|false|false|false|||ECHO
Procedure|Health Care Activity|SIMPLE_SEGMENT|10403,10407|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10403,10407|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10454,10465|true|false|false|C1980023|Wall motion|wall motion
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|10459,10465|true|false|false|C0026597|Motion|motion
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|10466,10479|true|false|false|C0000768|Congenital Abnormality|abnormalities
Event|Event|SIMPLE_SEGMENT|10466,10479|true|false|false|||abnormalities
Finding|Functional Concept|SIMPLE_SEGMENT|10466,10479|true|false|false|C0000769|teratologic|abnormalities
Finding|Body Substance|SIMPLE_SEGMENT|10485,10492|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|10485,10492|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|10485,10492|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|10498,10507|false|false|false|||continued
Drug|Organic Chemical|SIMPLE_SEGMENT|10511,10518|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10511,10518|false|false|false|C0004057|aspirin|aspirin
Event|Event|SIMPLE_SEGMENT|10511,10518|false|false|false|||aspirin
Drug|Organic Chemical|SIMPLE_SEGMENT|10535,10547|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10535,10547|false|false|false|C0286651|atorvastatin|atorvastatin
Event|Event|SIMPLE_SEGMENT|10535,10547|false|false|false|||atorvastatin
Finding|Idea or Concept|SIMPLE_SEGMENT|10580,10592|false|false|false|C1548597|Marketing basis - Transitional|TRANSITIONAL
Event|Event|SIMPLE_SEGMENT|10593,10599|false|false|false|||ISSUES
Finding|Finding|SIMPLE_SEGMENT|10622,10625|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|New
Finding|Idea or Concept|SIMPLE_SEGMENT|10622,10625|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|New
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10622,10637|false|false|false|C1718097|New medications|New Medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10626,10637|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10626,10637|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|10626,10637|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|10626,10637|false|false|false|C4284232|Medications|Medications
Drug|Hormone|SIMPLE_SEGMENT|10640,10650|false|false|false|C0032952|prednisone|Prednisone
Drug|Organic Chemical|SIMPLE_SEGMENT|10640,10650|false|false|false|C0032952|prednisone|Prednisone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10640,10650|false|false|false|C0032952|prednisone|Prednisone
Finding|Intellectual Product|SIMPLE_SEGMENT|10676,10680|false|false|false|C1720594|Then - dosing instruction fragment|then
Finding|Intellectual Product|SIMPLE_SEGMENT|10704,10708|false|false|false|C1720594|Then - dosing instruction fragment|then
Finding|Classification|SIMPLE_SEGMENT|10725,10735|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|10725,10735|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|SIMPLE_SEGMENT|10736,10742|false|false|false|||follow
Finding|Functional Concept|SIMPLE_SEGMENT|10736,10742|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|SIMPLE_SEGMENT|10736,10742|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|SIMPLE_SEGMENT|10736,10745|false|false|false|C0589120|Follow-up status|follow-up
Procedure|Health Care Activity|SIMPLE_SEGMENT|10736,10745|false|false|false|C1522577|follow-up|follow-up
Drug|Organic Chemical|SIMPLE_SEGMENT|10757,10763|false|false|false|C0965130|Advair|Advair
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10757,10763|false|false|false|C0965130|Advair|Advair
Event|Event|SIMPLE_SEGMENT|10757,10763|false|false|false|||Advair
Drug|Organic Chemical|SIMPLE_SEGMENT|10765,10776|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10765,10776|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10765,10787|false|false|false|C0939232|fluticasone / salmeterol|Fluticasone-Salmeterol
Drug|Organic Chemical|SIMPLE_SEGMENT|10777,10787|false|false|false|C0073992|salmeterol|Salmeterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10777,10787|false|false|false|C0073992|salmeterol|Salmeterol
Event|Event|SIMPLE_SEGMENT|10777,10787|false|false|false|||Salmeterol
Drug|Organic Chemical|SIMPLE_SEGMENT|10805,10814|false|false|false|C0024002|lorazepam|Lorazepam
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10805,10814|false|false|false|C0024002|lorazepam|Lorazepam
Event|Event|SIMPLE_SEGMENT|10829,10832|false|false|false|||PRN
Finding|Gene or Genome|SIMPLE_SEGMENT|10829,10832|false|false|false|C1422467|CIAO3 gene|PRN
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|10837,10844|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Event|Event|SIMPLE_SEGMENT|10837,10844|false|false|false|||anxiety
Finding|Sign or Symptom|SIMPLE_SEGMENT|10837,10844|false|false|false|C0860603|Anxiety symptoms|anxiety
Finding|Functional Concept|SIMPLE_SEGMENT|10847,10853|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|Follow
Finding|Intellectual Product|SIMPLE_SEGMENT|10847,10853|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|Follow
Finding|Finding|SIMPLE_SEGMENT|10847,10856|false|false|false|C0589120|Follow-up status|Follow-up
Procedure|Health Care Activity|SIMPLE_SEGMENT|10847,10856|false|false|false|C1522577|follow-up|Follow-up
Event|Activity|SIMPLE_SEGMENT|10859,10870|false|false|false|C0003629|Appointments|Appointment
Event|Event|SIMPLE_SEGMENT|10871,10879|false|false|false|||arranged
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10885,10888|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|10885,10888|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|10885,10888|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10885,10888|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|SIMPLE_SEGMENT|10885,10888|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|10885,10888|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|SIMPLE_SEGMENT|10885,10888|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10885,10888|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|SIMPLE_SEGMENT|10885,10888|false|false|false|||PCP
Finding|Gene or Genome|SIMPLE_SEGMENT|10885,10888|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|SIMPLE_SEGMENT|10885,10888|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Activity|SIMPLE_SEGMENT|10899,10910|false|false|false|C0003629|Appointments|Appointment
Event|Event|SIMPLE_SEGMENT|10899,10910|false|false|false|||Appointment
Event|Event|SIMPLE_SEGMENT|10911,10919|false|false|false|||arranged
Event|Event|SIMPLE_SEGMENT|10925,10938|false|false|false|||Pulmonologist
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10955,10959|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10955,10959|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|SIMPLE_SEGMENT|10955,10959|false|false|false|||COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|10955,10959|false|false|false|C1412502|ARCN1 gene|COPD
Finding|Body Substance|SIMPLE_SEGMENT|10961,10968|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|10961,10968|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|10961,10968|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|10973,10977|false|false|false|||seen
Event|Event|SIMPLE_SEGMENT|11000,11009|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|11000,11009|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|SIMPLE_SEGMENT|11033,11048|false|false|false|||recommendations
Finding|Idea or Concept|SIMPLE_SEGMENT|11033,11048|false|false|false|C0034866|Recommendation|recommendations
Event|Event|SIMPLE_SEGMENT|11052,11060|false|false|false|||consider
Event|Event|SIMPLE_SEGMENT|11067,11077|false|false|false|||outpatient
Finding|Classification|SIMPLE_SEGMENT|11067,11077|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|11067,11077|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|SIMPLE_SEGMENT|11080,11086|false|false|false|||Switch
Drug|Organic Chemical|SIMPLE_SEGMENT|11090,11101|false|false|false|C0965618|roflumilast|roflumilast
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11090,11101|false|false|false|C0965618|roflumilast|roflumilast
Event|Event|SIMPLE_SEGMENT|11090,11101|false|false|false|||roflumilast
Drug|Organic Chemical|SIMPLE_SEGMENT|11107,11119|false|false|false|C0039771|theophylline|theophylline
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11107,11119|false|false|false|C0039771|theophylline|theophylline
Event|Event|SIMPLE_SEGMENT|11107,11119|false|false|false|||theophylline
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|11107,11119|false|false|false|C0039773|Assay of theophylline|theophylline
Drug|Antibiotic|SIMPLE_SEGMENT|11127,11139|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Clinical Drug|SIMPLE_SEGMENT|11127,11139|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Organic Chemical|SIMPLE_SEGMENT|11127,11139|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Event|Event|SIMPLE_SEGMENT|11127,11139|false|false|false|||azithromycin
Event|Event|SIMPLE_SEGMENT|11144,11153|false|false|false|||treatment
Finding|Conceptual Entity|SIMPLE_SEGMENT|11144,11153|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|SIMPLE_SEGMENT|11144,11153|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|SIMPLE_SEGMENT|11144,11153|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11144,11153|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Finding|Intellectual Product|SIMPLE_SEGMENT|11157,11164|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|11157,11164|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Finding|Pathologic Function|SIMPLE_SEGMENT|11157,11177|false|false|false|C0021376|Chronic inflammation|chronic inflammation
Event|Event|SIMPLE_SEGMENT|11165,11177|false|false|false|||inflammation
Finding|Pathologic Function|SIMPLE_SEGMENT|11165,11177|false|false|false|C0021368|Inflammation|inflammation
Event|Event|SIMPLE_SEGMENT|11188,11191|false|false|false|||QTc
Finding|Finding|SIMPLE_SEGMENT|11192,11212|false|false|false|C0442816||within normal limits
Event|Event|SIMPLE_SEGMENT|11206,11212|false|false|false|||limits
Finding|Functional Concept|SIMPLE_SEGMENT|11206,11212|false|false|false|C0439801|Limited (extensiveness)|limits
Finding|Body Substance|SIMPLE_SEGMENT|11215,11222|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|11215,11222|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|11215,11222|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|11227,11234|false|false|false|||benefit
Event|Event|SIMPLE_SEGMENT|11240,11249|false|false|false|||treatment
Finding|Conceptual Entity|SIMPLE_SEGMENT|11240,11249|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|SIMPLE_SEGMENT|11240,11249|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|SIMPLE_SEGMENT|11240,11249|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11240,11249|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|11253,11260|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Event|Event|SIMPLE_SEGMENT|11253,11260|false|false|false|||anxiety
Finding|Sign or Symptom|SIMPLE_SEGMENT|11253,11260|false|false|false|C0860603|Anxiety symptoms|anxiety
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11269,11273|false|false|false|C0360105;C2911696|Selective Serotonin Reuptake Inhibitors;Serotonin Reuptake Inhibitor [EPC]|SSRI
Event|Event|SIMPLE_SEGMENT|11269,11273|false|false|false|||SSRI
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|11283,11290|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Event|Event|SIMPLE_SEGMENT|11283,11290|false|false|false|||anxiety
Finding|Sign or Symptom|SIMPLE_SEGMENT|11283,11290|false|false|false|C0860603|Anxiety symptoms|anxiety
Finding|Finding|SIMPLE_SEGMENT|11294,11300|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|11294,11300|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|SIMPLE_SEGMENT|11301,11313|false|false|false|||contributing
Event|Event|SIMPLE_SEGMENT|11321,11331|false|false|false|||experience
Finding|Mental Process|SIMPLE_SEGMENT|11321,11331|false|false|false|C0237607;C0596545|Experience;Experience (Practice)|experience
Event|Event|SIMPLE_SEGMENT|11335,11342|false|false|false|||dyspnea
Finding|Finding|SIMPLE_SEGMENT|11335,11342|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|11335,11342|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Finding|SIMPLE_SEGMENT|11360,11375|false|false|false|C0700049|Encounter due to palliative care|palliative care
Procedure|Health Care Activity|SIMPLE_SEGMENT|11360,11375|false|false|false|C0030231;C3816218|Palliative Care;Palliative Nursing|palliative care
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11360,11375|false|false|false|C0030231;C3816218|Palliative Care;Palliative Nursing|palliative care
Event|Activity|SIMPLE_SEGMENT|11371,11375|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|11371,11375|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|11371,11375|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|11371,11375|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Event|Event|SIMPLE_SEGMENT|11376,11383|false|false|false|||consult
Procedure|Health Care Activity|SIMPLE_SEGMENT|11376,11383|false|false|false|C0009818|Consultation|consult
Event|Event|SIMPLE_SEGMENT|11388,11401|false|false|false|||consideration
Finding|Finding|SIMPLE_SEGMENT|11388,11401|false|false|false|C0518609|Consideration|consideration
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|11406,11412|false|false|false|C0242402|Opioids|opioid
Drug|Organic Chemical|SIMPLE_SEGMENT|11406,11412|false|false|false|C0242402|Opioids|opioid
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11406,11412|false|false|false|C0242402|Opioids|opioid
Event|Event|SIMPLE_SEGMENT|11413,11422|false|false|false|||treatment
Finding|Conceptual Entity|SIMPLE_SEGMENT|11413,11422|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|SIMPLE_SEGMENT|11413,11422|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|SIMPLE_SEGMENT|11413,11422|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11413,11422|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Event|Event|SIMPLE_SEGMENT|11426,11433|false|false|false|||dyspnea
Finding|Finding|SIMPLE_SEGMENT|11426,11433|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|11426,11433|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Finding|SIMPLE_SEGMENT|11436,11457|false|false|false|C0239937|Microscopic hematuria|Microscopic hematuria
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11448,11457|false|false|false|C0018965|Hematuria|hematuria
Event|Event|SIMPLE_SEGMENT|11448,11457|false|false|false|||hematuria
Finding|Body Substance|SIMPLE_SEGMENT|11459,11466|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|11459,11466|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|11459,11466|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|11473,11475|false|false|false|||UA
Anatomy|Cell|SIMPLE_SEGMENT|11484,11488|false|false|false|C0014792|Erythrocytes|RBCs
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11484,11488|false|false|false|C0014792|Erythrocytes|RBCs
Event|Event|SIMPLE_SEGMENT|11493,11502|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|11493,11502|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|SIMPLE_SEGMENT|11515,11521|false|false|false|||repeat
Finding|Functional Concept|SIMPLE_SEGMENT|11515,11521|false|false|false|C0205341;C1705914|Repeat;Repeat Object|repeat
Event|Event|SIMPLE_SEGMENT|11531,11541|false|false|false|||outpatient
Finding|Classification|SIMPLE_SEGMENT|11531,11541|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|11531,11541|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|SIMPLE_SEGMENT|11545,11549|false|false|false|||work
Event|Occupational Activity|SIMPLE_SEGMENT|11545,11549|false|false|false|C0043227|Work|work
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|11545,11552|false|false|false|C0750430|Work-up|work-up
Event|Event|SIMPLE_SEGMENT|11550,11552|false|false|false|||up
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11570,11579|false|false|false|C0018965|Hematuria|hematuria
Event|Event|SIMPLE_SEGMENT|11570,11579|false|false|false|||hematuria
Anatomy|Body Location or Region|SIMPLE_SEGMENT|11582,11586|false|false|false|C0024109;C4037972|Chest>Lung;Lung|Lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11582,11586|false|false|false|C0024109;C4037972|Chest>Lung;Lung|Lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11582,11586|false|false|false|C0024115|Lung diseases|Lung
Finding|Finding|SIMPLE_SEGMENT|11582,11586|false|false|false|C0740941|Lung Problem|Lung
Finding|Finding|SIMPLE_SEGMENT|11582,11593|false|false|false|C0034079||Lung nodule
Event|Event|SIMPLE_SEGMENT|11587,11593|false|false|false|||nodule
Finding|Finding|SIMPLE_SEGMENT|11595,11598|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|New
Finding|Idea or Concept|SIMPLE_SEGMENT|11595,11598|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|New
Finding|Functional Concept|SIMPLE_SEGMENT|11599,11603|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11599,11614|false|false|false|C1261077|Structure of left lower lobe of lung|left lower lobe
Anatomy|Body Location or Region|SIMPLE_SEGMENT|11604,11609|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|11604,11609|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11604,11614|false|false|false|C0225758|Structure of lower lobe of lung|lower lobe
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11610,11614|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|SIMPLE_SEGMENT|11610,11614|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Event|Event|SIMPLE_SEGMENT|11615,11621|false|false|false|||nodule
Event|Event|SIMPLE_SEGMENT|11635,11644|false|false|false|||measuring
Finding|Gene or Genome|SIMPLE_SEGMENT|11649,11654|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Event|Event|SIMPLE_SEGMENT|11668,11676|false|false|false|||warrants
Finding|Finding|SIMPLE_SEGMENT|11677,11682|false|false|false|C0587267;C3810854|Close;Closed|close
Finding|Functional Concept|SIMPLE_SEGMENT|11677,11682|false|false|false|C0587267;C3810854|Close;Closed|close
Event|Event|SIMPLE_SEGMENT|11683,11689|false|false|false|||follow
Finding|Functional Concept|SIMPLE_SEGMENT|11683,11689|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|SIMPLE_SEGMENT|11683,11689|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|SIMPLE_SEGMENT|11683,11692|false|false|false|C0589120|Follow-up status|follow-up
Procedure|Health Care Activity|SIMPLE_SEGMENT|11683,11692|false|false|false|C1522577|follow-up|follow-up
Event|Event|SIMPLE_SEGMENT|11690,11692|false|false|false|||up
Event|Event|SIMPLE_SEGMENT|11695,11701|false|false|false|||Stable
Finding|Intellectual Product|SIMPLE_SEGMENT|11695,11701|false|false|false|C1547311|Patient Condition Code - Stable|Stable
Finding|Functional Concept|SIMPLE_SEGMENT|11728,11733|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11728,11745|false|false|false|C4281590|Structure of middle lobe of right lung|right middle lobe
Finding|Intellectual Product|SIMPLE_SEGMENT|11734,11740|false|false|false|C1552826|Table Cell Vertical Align - middle|middle
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11734,11745|false|false|false|C4281590|Structure of middle lobe of right lung|middle lobe
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11741,11745|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|SIMPLE_SEGMENT|11741,11745|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Event|Event|SIMPLE_SEGMENT|11746,11752|false|false|false|||nodule
Event|Event|SIMPLE_SEGMENT|11754,11760|false|false|false|||Follow
Event|Event|SIMPLE_SEGMENT|11793,11803|false|false|false|||guidelines
Finding|Intellectual Product|SIMPLE_SEGMENT|11793,11803|false|false|false|C0162791;C0220845;C0282423|Guideline (Publication Type);Guidelines;guiding characteristics|guidelines
Event|Event|SIMPLE_SEGMENT|11808,11818|false|false|false|||evaluation
Finding|Idea or Concept|SIMPLE_SEGMENT|11808,11818|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|SIMPLE_SEGMENT|11808,11818|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Finding|Finding|SIMPLE_SEGMENT|11823,11826|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|11823,11826|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Functional Concept|SIMPLE_SEGMENT|11827,11831|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11827,11842|false|false|false|C1261077|Structure of left lower lobe of lung|left lower lobe
Anatomy|Body Location or Region|SIMPLE_SEGMENT|11832,11837|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|11832,11837|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11832,11842|false|false|false|C0225758|Structure of lower lobe of lung|lower lobe
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11838,11842|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|SIMPLE_SEGMENT|11838,11842|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11838,11852|false|false|false|C0225752|Structure of lobe of lung|lobe pulmonary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11843,11852|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11843,11852|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|11843,11852|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Finding|SIMPLE_SEGMENT|11843,11859|false|false|false|C0034079||pulmonary nodule
Event|Event|SIMPLE_SEGMENT|11853,11859|false|false|false|||nodule
Event|Occupational Activity|SIMPLE_SEGMENT|11863,11867|false|false|false|C0009219|Coding|Code
Finding|Intellectual Product|SIMPLE_SEGMENT|11863,11867|false|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|Code
Procedure|Health Care Activity|SIMPLE_SEGMENT|11863,11874|false|false|false|C0742531|CODE STATUS|Code Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11868,11874|false|false|false|C5889824||Status
Event|Event|SIMPLE_SEGMENT|11868,11874|false|false|false|||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|11868,11874|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|11881,11885|false|false|false|||code
Event|Occupational Activity|SIMPLE_SEGMENT|11881,11885|false|false|false|C0009219|Coding|code
Finding|Intellectual Product|SIMPLE_SEGMENT|11881,11885|false|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|code
Event|Event|SIMPLE_SEGMENT|11887,11896|false|false|false|||Emergency
Finding|Finding|SIMPLE_SEGMENT|11887,11896|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Finding|Idea or Concept|SIMPLE_SEGMENT|11887,11896|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Finding|Intellectual Product|SIMPLE_SEGMENT|11887,11896|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Finding|Pathologic Function|SIMPLE_SEGMENT|11887,11896|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|11887,11896|false|false|false|C0013956|Emergency Situation|Emergency
Procedure|Health Care Activity|SIMPLE_SEGMENT|11887,11896|false|false|false|C1553500|emergency encounter|Emergency
Finding|Functional Concept|SIMPLE_SEGMENT|11887,11904|false|false|false|C1552023|emergency contact|Emergency Contact
Event|Activity|SIMPLE_SEGMENT|11897,11904|false|false|false|C3812666|Personal Contact|Contact
Finding|Functional Concept|SIMPLE_SEGMENT|11897,11904|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|Contact
Finding|Idea or Concept|SIMPLE_SEGMENT|11897,11904|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|Contact
Finding|Intellectual Product|SIMPLE_SEGMENT|11897,11904|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|Contact
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|11897,11904|false|false|false|C0392367|Physical contact|Contact
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11905,11908|false|false|false|C0162531|Hereditary Coproporphyria|HCP
Event|Event|SIMPLE_SEGMENT|11905,11908|false|false|false|||HCP
Finding|Gene or Genome|SIMPLE_SEGMENT|11905,11908|false|false|false|C1335283;C1412376;C1413681;C1705637;C5780748|AMBP gene;AMBP wt Allele;CPOX gene;PTPN6 gene;PTPN6 wt Allele|HCP
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11930,11941|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11930,11941|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|11930,11941|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|11930,11941|false|false|false|C4284232|Medications|Medications
Finding|Finding|SIMPLE_SEGMENT|11930,11954|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|SIMPLE_SEGMENT|11945,11954|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|11945,11954|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11973,11983|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|11973,11983|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|11973,11988|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|SIMPLE_SEGMENT|11984,11988|false|false|false|||list
Finding|Intellectual Product|SIMPLE_SEGMENT|11984,11988|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|SIMPLE_SEGMENT|11992,12000|false|false|false|||accurate
Drug|Organic Chemical|SIMPLE_SEGMENT|12005,12013|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12005,12013|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|SIMPLE_SEGMENT|12005,12013|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|SIMPLE_SEGMENT|12005,12013|false|false|false|||complete
Finding|Functional Concept|SIMPLE_SEGMENT|12005,12013|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|SIMPLE_SEGMENT|12005,12013|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Hormone|SIMPLE_SEGMENT|12018,12028|false|false|false|C0032952|prednisone|PredniSONE
Drug|Organic Chemical|SIMPLE_SEGMENT|12018,12028|false|false|false|C0032952|prednisone|PredniSONE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12018,12028|false|false|false|C0032952|prednisone|PredniSONE
Procedure|Health Care Activity|SIMPLE_SEGMENT|12044,12051|false|false|false|C0441640||Tapered
Event|Event|SIMPLE_SEGMENT|12059,12063|false|false|false|||DOWN
Drug|Organic Chemical|SIMPLE_SEGMENT|12068,12081|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12068,12081|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|SIMPLE_SEGMENT|12068,12081|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|12068,12081|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|SIMPLE_SEGMENT|12096,12099|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12100,12104|false|false|false|C2598155||Pain
Event|Event|SIMPLE_SEGMENT|12100,12104|false|false|false|||Pain
Finding|Functional Concept|SIMPLE_SEGMENT|12100,12104|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|12100,12104|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Drug|Organic Chemical|SIMPLE_SEGMENT|12109,12120|false|false|false|C0027235|ipratropium|Ipratropium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12109,12120|false|false|false|C0027235|ipratropium|Ipratropium
Event|Event|SIMPLE_SEGMENT|12109,12120|false|false|false|||Ipratropium
Drug|Organic Chemical|SIMPLE_SEGMENT|12109,12128|false|false|false|C0700580|ipratropium bromide|Ipratropium Bromide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12109,12128|false|false|false|C0700580|ipratropium bromide|Ipratropium Bromide
Drug|Inorganic Chemical|SIMPLE_SEGMENT|12121,12128|false|false|false|C0006222|Bromides|Bromide
Event|Event|SIMPLE_SEGMENT|12121,12128|false|false|false|||Bromide
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|12121,12128|false|false|false|C0202341|Bromides measurement|Bromide
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|12129,12132|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|12129,12132|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|12129,12132|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Event|Event|SIMPLE_SEGMENT|12129,12132|false|false|false|||Neb
Finding|Cell Function|SIMPLE_SEGMENT|12129,12132|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Finding|Gene or Genome|SIMPLE_SEGMENT|12129,12132|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|12135,12138|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biologically Active Substance|SIMPLE_SEGMENT|12135,12138|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|12135,12138|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Event|Event|SIMPLE_SEGMENT|12135,12138|false|false|false|||NEB
Finding|Cell Function|SIMPLE_SEGMENT|12135,12138|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|SIMPLE_SEGMENT|12135,12138|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|SIMPLE_SEGMENT|12146,12149|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|SIMPLE_SEGMENT|12150,12158|false|false|false|||Wheezing
Finding|Sign or Symptom|SIMPLE_SEGMENT|12150,12158|false|false|false|C0043144|Wheezing|Wheezing
Drug|Organic Chemical|SIMPLE_SEGMENT|12163,12173|false|false|false|C0213771|tiotropium|Tiotropium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12163,12173|false|false|false|C0213771|tiotropium|Tiotropium
Event|Event|SIMPLE_SEGMENT|12163,12173|false|false|false|||Tiotropium
Drug|Organic Chemical|SIMPLE_SEGMENT|12163,12181|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12163,12181|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Inorganic Chemical|SIMPLE_SEGMENT|12174,12181|false|false|false|C0006222|Bromides|Bromide
Event|Event|SIMPLE_SEGMENT|12174,12181|false|false|false|||Bromide
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|12174,12181|false|false|false|C0202341|Bromides measurement|Bromide
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|12184,12187|false|false|false|C1855179|CATARACT, ANTERIOR POLAR|CAP
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|12184,12187|false|false|false|C0006935|capsule (pharmacologic)|CAP
Event|Event|SIMPLE_SEGMENT|12184,12187|false|false|false|||CAP
Finding|Gene or Genome|SIMPLE_SEGMENT|12184,12187|false|false|false|C1416891;C1418551;C1419093;C1422073;C1422760;C2985259;C4522312|BRD4 gene;BRD4 wt Allele;CAP1 gene;HACD1 gene;LNPEP gene;SERPINB6 gene;SORBS1 gene|CAP
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|12184,12187|false|false|false|C0278651;C0280547;C1879916|CAP Regimen;cisplatin/cyclophosphamide/doxorubicin protocol;cyclophosphamide/doxorubicin/prednisone protocol|CAP
Drug|Organic Chemical|SIMPLE_SEGMENT|12201,12212|false|false|false|C0018305|guaifenesin|Guaifenesin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12201,12212|false|false|false|C0018305|guaifenesin|Guaifenesin
Finding|Gene or Genome|SIMPLE_SEGMENT|12231,12234|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Organic Chemical|SIMPLE_SEGMENT|12235,12240|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12235,12240|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|SIMPLE_SEGMENT|12235,12240|false|false|false|||cough
Finding|Sign or Symptom|SIMPLE_SEGMENT|12235,12240|false|false|false|C0010200|Coughing|cough
Drug|Organic Chemical|SIMPLE_SEGMENT|12245,12254|false|false|false|C0024002|lorazepam|Lorazepam
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12245,12254|false|false|false|C0024002|lorazepam|Lorazepam
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12269,12276|false|false|false|C1135208|Vertigo as late effect of cerebrovascular disease|vertigo
Event|Event|SIMPLE_SEGMENT|12269,12276|false|false|false|||vertigo
Finding|Sign or Symptom|SIMPLE_SEGMENT|12269,12276|false|false|false|C0042571|Vertigo|vertigo
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12277,12285|false|false|false|C1950154|Insomnia homeopathic medication|insomnia
Event|Event|SIMPLE_SEGMENT|12277,12285|false|false|false|||insomnia
Finding|Sign or Symptom|SIMPLE_SEGMENT|12277,12285|false|false|false|C0917801|Sleeplessness|insomnia
Drug|Organic Chemical|SIMPLE_SEGMENT|12290,12299|false|false|false|C0012373|diltiazem|Diltiazem
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12290,12299|false|false|false|C0012373|diltiazem|Diltiazem
Finding|Finding|SIMPLE_SEGMENT|12300,12308|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|SIMPLE_SEGMENT|12300,12308|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|SIMPLE_SEGMENT|12309,12316|false|false|false|||Release
Finding|Functional Concept|SIMPLE_SEGMENT|12309,12316|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|12309,12316|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|12309,12316|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|12327,12330|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|12327,12330|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|12327,12330|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|12327,12330|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|12327,12330|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|12335,12346|false|false|false|C0165590|dorzolamide|Dorzolamide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12335,12346|false|false|false|C0165590|dorzolamide|Dorzolamide
Finding|Functional Concept|SIMPLE_SEGMENT|12350,12355|false|false|false|C1522230|Ophthalmic Route of Administration|Ophth
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|12365,12369|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|SIMPLE_SEGMENT|12365,12369|false|false|false|C1705648|Dropping|DROP
Event|Event|SIMPLE_SEGMENT|12365,12369|false|false|false|||DROP
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|12370,12379|false|false|false|C0229118|Structure of both eyes|BOTH EYES
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|12375,12379|false|false|false|C0015392|Eye|EYES
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12375,12379|false|false|false|C5848506||EYES
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|12380,12383|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|12380,12383|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|12380,12383|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|12380,12383|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|12380,12383|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|12388,12396|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12388,12396|false|false|false|C1692318|docusate|Docusate
Event|Event|SIMPLE_SEGMENT|12388,12396|false|false|false|||Docusate
Drug|Organic Chemical|SIMPLE_SEGMENT|12388,12403|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12388,12403|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|12397,12403|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|12397,12403|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12397,12403|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|SIMPLE_SEGMENT|12397,12403|false|false|false|||Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|12397,12403|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|12397,12403|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|12414,12417|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|12414,12417|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|12414,12417|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|12414,12417|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|12414,12417|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|12423,12434|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12423,12434|false|false|false|C0082607|fluticasone|Fluticasone
Event|Event|SIMPLE_SEGMENT|12423,12434|false|false|false|||Fluticasone
Drug|Organic Chemical|SIMPLE_SEGMENT|12423,12445|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12423,12445|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Organic Chemical|SIMPLE_SEGMENT|12435,12445|false|false|false|C0033474;C0392214|Propionates;propionate|Propionate
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|12446,12451|false|false|false|C0028429||NASAL
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|12446,12451|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Drug|Organic Chemical|SIMPLE_SEGMENT|12446,12451|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12446,12451|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Finding|Finding|SIMPLE_SEGMENT|12446,12451|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|NASAL
Finding|Functional Concept|SIMPLE_SEGMENT|12446,12451|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|NASAL
Event|Event|SIMPLE_SEGMENT|12454,12458|false|false|false|||SPRY
Event|Event|SIMPLE_SEGMENT|12462,12467|false|false|false|||DAILY
Finding|Gene or Genome|SIMPLE_SEGMENT|12468,12471|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12472,12481|false|false|false|C1717415||allergies
Event|Event|SIMPLE_SEGMENT|12472,12481|false|false|false|||allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|12472,12481|false|false|false|C0020517|Hypersensitivity|allergies
Drug|Organic Chemical|SIMPLE_SEGMENT|12487,12495|false|false|false|C1831808|apixaban|Apixaban
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12487,12495|false|false|false|C1831808|apixaban|Apixaban
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|12504,12507|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|12504,12507|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|12504,12507|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|12504,12507|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|12504,12507|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|12513,12523|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12513,12523|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Organic Chemical|SIMPLE_SEGMENT|12545,12557|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12545,12557|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|12576,12583|false|false|false|C2346592|Ferrous|Ferrous
Drug|Inorganic Chemical|SIMPLE_SEGMENT|12576,12591|false|false|false|C0060282|ferrous sulfate|Ferrous Sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12576,12591|false|false|false|C0060282|ferrous sulfate|Ferrous Sulfate
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|12584,12591|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Inorganic Chemical|SIMPLE_SEGMENT|12584,12591|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12584,12591|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Event|Event|SIMPLE_SEGMENT|12584,12591|false|false|false|||Sulfate
Drug|Organic Chemical|SIMPLE_SEGMENT|12613,12626|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12613,12626|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|SIMPLE_SEGMENT|12613,12626|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Event|Event|SIMPLE_SEGMENT|12613,12626|false|false|false|||Multivitamins
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|12629,12632|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|SIMPLE_SEGMENT|12629,12632|false|false|false|||TAB
Drug|Organic Chemical|SIMPLE_SEGMENT|12647,12657|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12647,12657|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Organic Chemical|SIMPLE_SEGMENT|12647,12669|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12647,12669|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Event|Event|SIMPLE_SEGMENT|12658,12669|false|false|false|||Mononitrate
Finding|Finding|SIMPLE_SEGMENT|12671,12679|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|SIMPLE_SEGMENT|12671,12679|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|SIMPLE_SEGMENT|12680,12687|false|false|false|||Release
Finding|Functional Concept|SIMPLE_SEGMENT|12680,12687|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|12680,12687|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|12680,12687|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|SIMPLE_SEGMENT|12710,12721|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12710,12721|false|false|false|C0082607|fluticasone|Fluticasone
Event|Event|SIMPLE_SEGMENT|12710,12721|false|false|false|||Fluticasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12710,12732|false|false|false|C0939232|fluticasone / salmeterol|Fluticasone-Salmeterol
Drug|Organic Chemical|SIMPLE_SEGMENT|12710,12739|false|false|false|C4762496|Fluticasone-Salmeterol Diskus|Fluticasone-Salmeterol Diskus
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12710,12739|false|false|false|C4762496|Fluticasone-Salmeterol Diskus|Fluticasone-Salmeterol Diskus
Drug|Organic Chemical|SIMPLE_SEGMENT|12722,12732|false|false|false|C0073992|salmeterol|Salmeterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12722,12732|false|false|false|C0073992|salmeterol|Salmeterol
Event|Event|SIMPLE_SEGMENT|12733,12739|false|false|false|||Diskus
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|12752,12755|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Organic Chemical|SIMPLE_SEGMENT|12752,12755|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12752,12755|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Event|Event|SIMPLE_SEGMENT|12752,12755|false|false|false|||INH
Finding|Functional Concept|SIMPLE_SEGMENT|12752,12755|false|false|false|C0205535|Inhalation Route of Administration|INH
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|12759,12762|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|12759,12762|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|12759,12762|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|12759,12762|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|12759,12762|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|12768,12779|false|false|false|C0090306|latanoprost|Latanoprost
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12768,12779|false|false|false|C0090306|latanoprost|Latanoprost
Finding|Functional Concept|SIMPLE_SEGMENT|12787,12792|false|false|false|C1522230|Ophthalmic Route of Administration|Ophth
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|12802,12806|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|SIMPLE_SEGMENT|12802,12806|false|false|false|C1705648|Dropping|DROP
Event|Event|SIMPLE_SEGMENT|12802,12806|false|false|false|||DROP
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|12807,12816|false|false|false|C0229118|Structure of both eyes|BOTH EYES
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|12812,12816|false|false|false|C0015392|Eye|EYES
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12812,12816|false|false|false|C5848506||EYES
Drug|Organic Chemical|SIMPLE_SEGMENT|12826,12836|false|false|false|C3464797|Calcitrate|Calcitrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12826,12836|false|false|false|C3464797|Calcitrate|Calcitrate
Drug|Organic Chemical|SIMPLE_SEGMENT|12837,12844|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12837,12844|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|SIMPLE_SEGMENT|12837,12844|false|false|false|C0042890|Vitamins|Vitamin
Event|Event|SIMPLE_SEGMENT|12837,12844|false|false|false|||Vitamin
Drug|Hormone|SIMPLE_SEGMENT|12837,12846|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|SIMPLE_SEGMENT|12837,12846|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12837,12846|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|SIMPLE_SEGMENT|12837,12846|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|12837,12846|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Event|Event|SIMPLE_SEGMENT|12845,12846|false|false|false|||D
Drug|Biologically Active Substance|SIMPLE_SEGMENT|12848,12855|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|12848,12855|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|12848,12855|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12848,12855|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Vitamin|SIMPLE_SEGMENT|12848,12855|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Event|Event|SIMPLE_SEGMENT|12848,12855|false|false|false|||calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|12848,12855|false|false|false|C4553026|Calcium metabolic function|calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|12848,12855|false|false|false|C0201925|Calcium measurement|calcium
Drug|Organic Chemical|SIMPLE_SEGMENT|12848,12863|false|false|false|C0108101|calcium citrate|calcium citrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12848,12863|false|false|false|C0108101|calcium citrate|calcium citrate
Drug|Organic Chemical|SIMPLE_SEGMENT|12856,12863|false|false|false|C0008857;C0376259|Citrates;citrate|citrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12856,12863|false|false|false|C0008857;C0376259|Citrates;citrate|citrate
Event|Event|SIMPLE_SEGMENT|12856,12863|false|false|false|||citrate
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|12856,12863|false|false|false|C0201956|Citrate measurement|citrate
Drug|Organic Chemical|SIMPLE_SEGMENT|12864,12871|false|false|false|C0042890|Vitamins|vitamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12864,12871|false|false|false|C0042890|Vitamins|vitamin
Drug|Vitamin|SIMPLE_SEGMENT|12864,12871|false|false|false|C0042890|Vitamins|vitamin
Event|Event|SIMPLE_SEGMENT|12864,12871|false|false|false|||vitamin
Drug|Organic Chemical|SIMPLE_SEGMENT|12864,12874|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12864,12874|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Drug|Vitamin|SIMPLE_SEGMENT|12864,12874|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|12897,12901|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|12897,12901|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|12897,12901|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|12897,12901|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Event|Event|SIMPLE_SEGMENT|12902,12907|false|false|false|||DAILY
Drug|Organic Chemical|SIMPLE_SEGMENT|12913,12925|false|false|false|C0039771|theophylline|Theophylline
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12913,12925|false|false|false|C0039771|theophylline|Theophylline
Event|Event|SIMPLE_SEGMENT|12913,12925|false|false|false|||Theophylline
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|12913,12925|false|false|false|C0039773|Assay of theophylline|Theophylline
Drug|Organic Chemical|SIMPLE_SEGMENT|12913,12928|false|false|false|C0939729|Theophylline SR|Theophylline SR
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12913,12928|false|false|false|C0939729|Theophylline SR|Theophylline SR
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|12939,12942|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|12939,12942|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|12939,12942|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|12939,12942|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|12939,12942|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|12948,12955|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12948,12955|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|SIMPLE_SEGMENT|12976,12985|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12976,12985|false|false|false|C0001927|albuterol|albuterol
Event|Event|SIMPLE_SEGMENT|12976,12985|false|false|false|||albuterol
Drug|Organic Chemical|SIMPLE_SEGMENT|12976,12993|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12976,12993|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|12986,12993|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Inorganic Chemical|SIMPLE_SEGMENT|12986,12993|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12986,12993|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Event|Event|SIMPLE_SEGMENT|12986,12993|false|false|false|||sulfate
Finding|Functional Concept|SIMPLE_SEGMENT|13011,13021|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Finding|Organism Function|SIMPLE_SEGMENT|13011,13021|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Event|Event|SIMPLE_SEGMENT|13022,13025|false|false|false|||Q4H
Drug|Organic Chemical|SIMPLE_SEGMENT|13031,13050|false|false|false|C0020261|hydrochlorothiazide|Hydrochlorothiazide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13031,13050|false|false|false|C0020261|hydrochlorothiazide|Hydrochlorothiazide
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|13071,13074|false|false|false|C0056632;C0459207;C2702357;C3488428|Cyclophosphamide/Dacarbazine/Vincristine;cod, unspecified preparation;codfish allergenic extract|cod
Drug|Food|SIMPLE_SEGMENT|13071,13074|false|false|false|C0056632;C0459207;C2702357;C3488428|Cyclophosphamide/Dacarbazine/Vincristine;cod, unspecified preparation;codfish allergenic extract|cod
Drug|Immunologic Factor|SIMPLE_SEGMENT|13071,13074|false|false|false|C0056632;C0459207;C2702357;C3488428|Cyclophosphamide/Dacarbazine/Vincristine;cod, unspecified preparation;codfish allergenic extract|cod
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13071,13074|false|false|false|C0056632;C0459207;C2702357;C3488428|Cyclophosphamide/Dacarbazine/Vincristine;cod, unspecified preparation;codfish allergenic extract|cod
Event|Event|SIMPLE_SEGMENT|13071,13074|false|false|false|||cod
Finding|Finding|SIMPLE_SEGMENT|13071,13074|false|false|false|C0007465;C0457523;C1420285;C5444130|Cancerization of Pancreatic Ducts;Cause of Death;Cemento-osseous dysplasia;SNRPB gene|cod
Finding|Gene or Genome|SIMPLE_SEGMENT|13071,13074|false|false|false|C0007465;C0457523;C1420285;C5444130|Cancerization of Pancreatic Ducts;Cause of Death;Cemento-osseous dysplasia;SNRPB gene|cod
Finding|Pathologic Function|SIMPLE_SEGMENT|13071,13074|false|false|false|C0007465;C0457523;C1420285;C5444130|Cancerization of Pancreatic Ducts;Cause of Death;Cemento-osseous dysplasia;SNRPB gene|cod
Drug|Food|SIMPLE_SEGMENT|13071,13084|false|false|false|C0009213|cod liver oil|cod liver oil
Drug|Organic Chemical|SIMPLE_SEGMENT|13071,13084|false|false|false|C0009213|cod liver oil|cod liver oil
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13071,13084|false|false|false|C0009213|cod liver oil|cod liver oil
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|13075,13080|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13075,13080|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|SIMPLE_SEGMENT|13075,13080|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|SIMPLE_SEGMENT|13075,13080|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13075,13080|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|SIMPLE_SEGMENT|13075,13080|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|SIMPLE_SEGMENT|13075,13080|false|false|false|||liver
Finding|Finding|SIMPLE_SEGMENT|13075,13080|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|SIMPLE_SEGMENT|13075,13080|false|false|false|C0872387|Procedures on liver|liver
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|13081,13084|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|oil
Drug|Food|SIMPLE_SEGMENT|13081,13084|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|oil
Drug|Organic Chemical|SIMPLE_SEGMENT|13081,13084|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|oil
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13081,13084|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|oil
Event|Event|SIMPLE_SEGMENT|13081,13084|false|false|false|||oil
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|13087,13094|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Anatomy|Cell Component|SIMPLE_SEGMENT|13087,13094|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|13087,13094|false|false|false|C0006935|capsule (pharmacologic)|capsule
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|13096,13100|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|13096,13100|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|13096,13100|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|13096,13100|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|13101,13104|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|13101,13104|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|13101,13104|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|13101,13104|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|13101,13104|false|false|false|C1332410|BID gene|BID
Event|Event|SIMPLE_SEGMENT|13109,13118|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|13109,13118|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|13109,13118|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|13109,13118|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|13109,13118|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|13109,13130|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13119,13130|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13119,13130|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|13119,13130|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|13119,13130|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|SIMPLE_SEGMENT|13135,13148|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13135,13148|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|SIMPLE_SEGMENT|13135,13148|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|13135,13148|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|SIMPLE_SEGMENT|13163,13166|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13167,13171|false|false|false|C2598155||Pain
Event|Event|SIMPLE_SEGMENT|13167,13171|false|false|false|||Pain
Finding|Functional Concept|SIMPLE_SEGMENT|13167,13171|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|13167,13171|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Drug|Organic Chemical|SIMPLE_SEGMENT|13176,13184|false|false|false|C1831808|apixaban|Apixaban
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13176,13184|false|false|false|C1831808|apixaban|Apixaban
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|13193,13196|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|13193,13196|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|13193,13196|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|13193,13196|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|13193,13196|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|13201,13208|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13201,13208|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|SIMPLE_SEGMENT|13228,13240|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13228,13240|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|SIMPLE_SEGMENT|13258,13267|false|false|false|C0012373|diltiazem|Diltiazem
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13258,13267|false|false|false|C0012373|diltiazem|Diltiazem
Finding|Finding|SIMPLE_SEGMENT|13268,13276|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|SIMPLE_SEGMENT|13268,13276|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|SIMPLE_SEGMENT|13277,13284|false|false|false|||Release
Finding|Functional Concept|SIMPLE_SEGMENT|13277,13284|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|13277,13284|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|13277,13284|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|13295,13298|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|13295,13298|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|13295,13298|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|13295,13298|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|13295,13298|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|13303,13311|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13303,13311|false|false|false|C1692318|docusate|Docusate
Event|Event|SIMPLE_SEGMENT|13303,13311|false|false|false|||Docusate
Drug|Organic Chemical|SIMPLE_SEGMENT|13303,13318|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13303,13318|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|13312,13318|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|13312,13318|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13312,13318|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|SIMPLE_SEGMENT|13312,13318|false|false|false|||Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|13312,13318|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|13312,13318|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|13329,13332|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|13329,13332|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|13329,13332|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|13329,13332|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|13329,13332|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|13337,13348|false|false|false|C0165590|dorzolamide|Dorzolamide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13337,13348|false|false|false|C0165590|dorzolamide|Dorzolamide
Finding|Functional Concept|SIMPLE_SEGMENT|13352,13357|false|false|false|C1522230|Ophthalmic Route of Administration|Ophth
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|13367,13371|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|SIMPLE_SEGMENT|13367,13371|false|false|false|C1705648|Dropping|DROP
Event|Event|SIMPLE_SEGMENT|13367,13371|false|false|false|||DROP
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|13372,13381|false|false|false|C0229118|Structure of both eyes|BOTH EYES
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|13377,13381|false|false|false|C0015392|Eye|EYES
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13377,13381|false|false|false|C5848506||EYES
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|13382,13385|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|13382,13385|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|13382,13385|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|13382,13385|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|13382,13385|false|false|false|C1332410|BID gene|BID
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|13390,13397|false|false|false|C2346592|Ferrous|Ferrous
Drug|Inorganic Chemical|SIMPLE_SEGMENT|13390,13405|false|false|false|C0060282|ferrous sulfate|Ferrous Sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13390,13405|false|false|false|C0060282|ferrous sulfate|Ferrous Sulfate
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|13398,13405|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Inorganic Chemical|SIMPLE_SEGMENT|13398,13405|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13398,13405|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Event|Event|SIMPLE_SEGMENT|13398,13405|false|false|false|||Sulfate
Drug|Organic Chemical|SIMPLE_SEGMENT|13426,13437|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13426,13437|false|false|false|C0082607|fluticasone|Fluticasone
Event|Event|SIMPLE_SEGMENT|13426,13437|false|false|false|||Fluticasone
Drug|Organic Chemical|SIMPLE_SEGMENT|13426,13448|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13426,13448|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Organic Chemical|SIMPLE_SEGMENT|13438,13448|false|false|false|C0033474;C0392214|Propionates;propionate|Propionate
Event|Event|SIMPLE_SEGMENT|13438,13448|false|false|false|||Propionate
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|13449,13454|false|false|false|C0028429||NASAL
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|13449,13454|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Drug|Organic Chemical|SIMPLE_SEGMENT|13449,13454|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13449,13454|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Finding|Finding|SIMPLE_SEGMENT|13449,13454|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|NASAL
Finding|Functional Concept|SIMPLE_SEGMENT|13449,13454|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|NASAL
Event|Event|SIMPLE_SEGMENT|13457,13461|false|false|false|||SPRY
Event|Event|SIMPLE_SEGMENT|13465,13470|false|false|false|||DAILY
Finding|Gene or Genome|SIMPLE_SEGMENT|13471,13474|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13475,13484|false|false|false|C1717415||allergies
Event|Event|SIMPLE_SEGMENT|13475,13484|false|false|false|||allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|13475,13484|false|false|false|C0020517|Hypersensitivity|allergies
Drug|Organic Chemical|SIMPLE_SEGMENT|13490,13509|false|false|false|C0020261|hydrochlorothiazide|Hydrochlorothiazide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13490,13509|false|false|false|C0020261|hydrochlorothiazide|Hydrochlorothiazide
Drug|Organic Chemical|SIMPLE_SEGMENT|13530,13540|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13530,13540|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Organic Chemical|SIMPLE_SEGMENT|13530,13552|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13530,13552|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Event|Event|SIMPLE_SEGMENT|13541,13552|false|false|false|||Mononitrate
Finding|Finding|SIMPLE_SEGMENT|13554,13562|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|SIMPLE_SEGMENT|13554,13562|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|SIMPLE_SEGMENT|13563,13570|false|false|false|||Release
Finding|Functional Concept|SIMPLE_SEGMENT|13563,13570|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|13563,13570|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|13563,13570|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|SIMPLE_SEGMENT|13593,13604|false|false|false|C0090306|latanoprost|Latanoprost
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13593,13604|false|false|false|C0090306|latanoprost|Latanoprost
Finding|Functional Concept|SIMPLE_SEGMENT|13612,13617|false|false|false|C1522230|Ophthalmic Route of Administration|Ophth
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|13627,13631|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|SIMPLE_SEGMENT|13627,13631|false|false|false|C1705648|Dropping|DROP
Event|Event|SIMPLE_SEGMENT|13627,13631|false|false|false|||DROP
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|13632,13641|false|false|false|C0229118|Structure of both eyes|BOTH EYES
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|13637,13641|false|false|false|C0015392|Eye|EYES
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13637,13641|false|false|false|C5848506||EYES
Drug|Organic Chemical|SIMPLE_SEGMENT|13651,13664|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13651,13664|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|SIMPLE_SEGMENT|13651,13664|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Event|Event|SIMPLE_SEGMENT|13651,13664|false|false|false|||Multivitamins
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|13667,13670|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|SIMPLE_SEGMENT|13667,13670|false|false|false|||TAB
Drug|Hormone|SIMPLE_SEGMENT|13685,13695|false|false|false|C0032952|prednisone|PredniSONE
Drug|Organic Chemical|SIMPLE_SEGMENT|13685,13695|false|false|false|C0032952|prednisone|PredniSONE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13685,13695|false|false|false|C0032952|prednisone|PredniSONE
Drug|Hormone|SIMPLE_SEGMENT|13716,13726|false|false|false|C0032952|prednisone|prednisone
Drug|Organic Chemical|SIMPLE_SEGMENT|13716,13726|false|false|false|C0032952|prednisone|prednisone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13716,13726|false|false|false|C0032952|prednisone|prednisone
Event|Event|SIMPLE_SEGMENT|13716,13726|false|false|false|||prednisone
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|13735,13741|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|SIMPLE_SEGMENT|13745,13753|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|13748,13753|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|13748,13753|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|13770,13776|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|13770,13776|false|false|false|||Tablet
Event|Event|SIMPLE_SEGMENT|13778,13785|false|false|false|||Refills
Finding|Idea or Concept|SIMPLE_SEGMENT|13778,13785|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|13793,13803|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13793,13803|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Organic Chemical|SIMPLE_SEGMENT|13825,13837|false|false|false|C0039771|theophylline|Theophylline
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13825,13837|false|false|false|C0039771|theophylline|Theophylline
Event|Event|SIMPLE_SEGMENT|13825,13837|false|false|false|||Theophylline
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|13825,13837|false|false|false|C0039773|Assay of theophylline|Theophylline
Drug|Organic Chemical|SIMPLE_SEGMENT|13825,13840|false|false|false|C0939729|Theophylline SR|Theophylline SR
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13825,13840|false|false|false|C0939729|Theophylline SR|Theophylline SR
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|13851,13854|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|13851,13854|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|13851,13854|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|13851,13854|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|13851,13854|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|13860,13870|false|false|false|C0213771|tiotropium|Tiotropium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13860,13870|false|false|false|C0213771|tiotropium|Tiotropium
Event|Event|SIMPLE_SEGMENT|13860,13870|false|false|false|||Tiotropium
Drug|Organic Chemical|SIMPLE_SEGMENT|13860,13878|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13860,13878|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Inorganic Chemical|SIMPLE_SEGMENT|13871,13878|false|false|false|C0006222|Bromides|Bromide
Event|Event|SIMPLE_SEGMENT|13871,13878|false|false|false|||Bromide
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|13871,13878|false|false|false|C0202341|Bromides measurement|Bromide
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|13881,13884|false|false|false|C1855179|CATARACT, ANTERIOR POLAR|CAP
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|13881,13884|false|false|false|C0006935|capsule (pharmacologic)|CAP
Event|Event|SIMPLE_SEGMENT|13881,13884|false|false|false|||CAP
Finding|Gene or Genome|SIMPLE_SEGMENT|13881,13884|false|false|false|C1416891;C1418551;C1419093;C1422073;C1422760;C2985259;C4522312|BRD4 gene;BRD4 wt Allele;CAP1 gene;HACD1 gene;LNPEP gene;SERPINB6 gene;SORBS1 gene|CAP
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|13881,13884|false|false|false|C0278651;C0280547;C1879916|CAP Regimen;cisplatin/cyclophosphamide/doxorubicin protocol;cyclophosphamide/doxorubicin/prednisone protocol|CAP
Drug|Organic Chemical|SIMPLE_SEGMENT|13899,13910|false|false|false|C0018305|guaifenesin|Guaifenesin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13899,13910|false|false|false|C0018305|guaifenesin|Guaifenesin
Finding|Gene or Genome|SIMPLE_SEGMENT|13929,13932|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Organic Chemical|SIMPLE_SEGMENT|13933,13938|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13933,13938|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|SIMPLE_SEGMENT|13933,13938|false|false|false|||cough
Finding|Sign or Symptom|SIMPLE_SEGMENT|13933,13938|false|false|false|C0010200|Coughing|cough
Drug|Organic Chemical|SIMPLE_SEGMENT|13944,13955|false|false|false|C0027235|ipratropium|Ipratropium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13944,13955|false|false|false|C0027235|ipratropium|Ipratropium
Event|Event|SIMPLE_SEGMENT|13944,13955|false|false|false|||Ipratropium
Drug|Organic Chemical|SIMPLE_SEGMENT|13944,13963|false|false|false|C0700580|ipratropium bromide|Ipratropium Bromide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13944,13963|false|false|false|C0700580|ipratropium bromide|Ipratropium Bromide
Drug|Inorganic Chemical|SIMPLE_SEGMENT|13956,13963|false|false|false|C0006222|Bromides|Bromide
Event|Event|SIMPLE_SEGMENT|13956,13963|false|false|false|||Bromide
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|13956,13963|false|false|false|C0202341|Bromides measurement|Bromide
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|13964,13967|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|13964,13967|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|13964,13967|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Event|Event|SIMPLE_SEGMENT|13964,13967|false|false|false|||Neb
Finding|Cell Function|SIMPLE_SEGMENT|13964,13967|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Finding|Gene or Genome|SIMPLE_SEGMENT|13964,13967|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|13970,13973|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biologically Active Substance|SIMPLE_SEGMENT|13970,13973|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|13970,13973|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Event|Event|SIMPLE_SEGMENT|13970,13973|false|false|false|||NEB
Finding|Cell Function|SIMPLE_SEGMENT|13970,13973|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|SIMPLE_SEGMENT|13970,13973|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|SIMPLE_SEGMENT|13981,13984|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|SIMPLE_SEGMENT|13985,13993|false|false|false|||Wheezing
Finding|Sign or Symptom|SIMPLE_SEGMENT|13985,13993|false|false|false|C0043144|Wheezing|Wheezing
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|13999,14002|false|false|false|C0056632;C0459207;C2702357;C3488428|Cyclophosphamide/Dacarbazine/Vincristine;cod, unspecified preparation;codfish allergenic extract|cod
Drug|Food|SIMPLE_SEGMENT|13999,14002|false|false|false|C0056632;C0459207;C2702357;C3488428|Cyclophosphamide/Dacarbazine/Vincristine;cod, unspecified preparation;codfish allergenic extract|cod
Drug|Immunologic Factor|SIMPLE_SEGMENT|13999,14002|false|false|false|C0056632;C0459207;C2702357;C3488428|Cyclophosphamide/Dacarbazine/Vincristine;cod, unspecified preparation;codfish allergenic extract|cod
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13999,14002|false|false|false|C0056632;C0459207;C2702357;C3488428|Cyclophosphamide/Dacarbazine/Vincristine;cod, unspecified preparation;codfish allergenic extract|cod
Event|Event|SIMPLE_SEGMENT|13999,14002|false|false|false|||cod
Finding|Finding|SIMPLE_SEGMENT|13999,14002|false|false|false|C0007465;C0457523;C1420285;C5444130|Cancerization of Pancreatic Ducts;Cause of Death;Cemento-osseous dysplasia;SNRPB gene|cod
Finding|Gene or Genome|SIMPLE_SEGMENT|13999,14002|false|false|false|C0007465;C0457523;C1420285;C5444130|Cancerization of Pancreatic Ducts;Cause of Death;Cemento-osseous dysplasia;SNRPB gene|cod
Finding|Pathologic Function|SIMPLE_SEGMENT|13999,14002|false|false|false|C0007465;C0457523;C1420285;C5444130|Cancerization of Pancreatic Ducts;Cause of Death;Cemento-osseous dysplasia;SNRPB gene|cod
Drug|Food|SIMPLE_SEGMENT|13999,14012|false|false|false|C0009213|cod liver oil|cod liver oil
Drug|Organic Chemical|SIMPLE_SEGMENT|13999,14012|false|false|false|C0009213|cod liver oil|cod liver oil
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13999,14012|false|false|false|C0009213|cod liver oil|cod liver oil
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|14003,14008|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14003,14008|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|SIMPLE_SEGMENT|14003,14008|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|SIMPLE_SEGMENT|14003,14008|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14003,14008|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|SIMPLE_SEGMENT|14003,14008|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|SIMPLE_SEGMENT|14003,14008|false|false|false|||liver
Finding|Finding|SIMPLE_SEGMENT|14003,14008|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|SIMPLE_SEGMENT|14003,14008|false|false|false|C0872387|Procedures on liver|liver
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|14009,14012|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|oil
Drug|Food|SIMPLE_SEGMENT|14009,14012|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|oil
Drug|Organic Chemical|SIMPLE_SEGMENT|14009,14012|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|oil
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14009,14012|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|oil
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|14015,14022|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Anatomy|Cell Component|SIMPLE_SEGMENT|14015,14022|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|14015,14022|false|false|false|C0006935|capsule (pharmacologic)|capsule
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|14024,14028|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|14024,14028|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|14024,14028|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|14024,14028|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|14029,14032|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|14029,14032|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|14029,14032|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|14029,14032|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|14029,14032|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|14038,14048|false|false|false|C3464797|Calcitrate|Calcitrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14038,14048|false|false|false|C3464797|Calcitrate|Calcitrate
Drug|Organic Chemical|SIMPLE_SEGMENT|14049,14056|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14049,14056|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|SIMPLE_SEGMENT|14049,14056|false|false|false|C0042890|Vitamins|Vitamin
Event|Event|SIMPLE_SEGMENT|14049,14056|false|false|false|||Vitamin
Drug|Hormone|SIMPLE_SEGMENT|14049,14058|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|SIMPLE_SEGMENT|14049,14058|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14049,14058|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|SIMPLE_SEGMENT|14049,14058|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|14049,14058|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Event|Event|SIMPLE_SEGMENT|14057,14058|false|false|false|||D
Drug|Biologically Active Substance|SIMPLE_SEGMENT|14060,14067|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|14060,14067|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|14060,14067|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14060,14067|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Vitamin|SIMPLE_SEGMENT|14060,14067|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Event|Event|SIMPLE_SEGMENT|14060,14067|false|false|false|||calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|14060,14067|false|false|false|C4553026|Calcium metabolic function|calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|14060,14067|false|false|false|C0201925|Calcium measurement|calcium
Drug|Organic Chemical|SIMPLE_SEGMENT|14060,14075|false|false|false|C0108101|calcium citrate|calcium citrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14060,14075|false|false|false|C0108101|calcium citrate|calcium citrate
Drug|Organic Chemical|SIMPLE_SEGMENT|14068,14075|false|false|false|C0008857;C0376259|Citrates;citrate|citrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14068,14075|false|false|false|C0008857;C0376259|Citrates;citrate|citrate
Event|Event|SIMPLE_SEGMENT|14068,14075|false|false|false|||citrate
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|14068,14075|false|false|false|C0201956|Citrate measurement|citrate
Drug|Organic Chemical|SIMPLE_SEGMENT|14076,14083|false|false|false|C0042890|Vitamins|vitamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14076,14083|false|false|false|C0042890|Vitamins|vitamin
Drug|Vitamin|SIMPLE_SEGMENT|14076,14083|false|false|false|C0042890|Vitamins|vitamin
Event|Event|SIMPLE_SEGMENT|14076,14083|false|false|false|||vitamin
Drug|Organic Chemical|SIMPLE_SEGMENT|14076,14086|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14076,14086|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Drug|Vitamin|SIMPLE_SEGMENT|14076,14086|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|14109,14113|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|14109,14113|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|14109,14113|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|14109,14113|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Event|Event|SIMPLE_SEGMENT|14114,14119|false|false|false|||DAILY
Drug|Organic Chemical|SIMPLE_SEGMENT|14125,14134|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14125,14134|false|false|false|C0001927|albuterol|albuterol
Event|Event|SIMPLE_SEGMENT|14125,14134|false|false|false|||albuterol
Drug|Organic Chemical|SIMPLE_SEGMENT|14125,14142|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14125,14142|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|14135,14142|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Inorganic Chemical|SIMPLE_SEGMENT|14135,14142|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14135,14142|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Event|Event|SIMPLE_SEGMENT|14135,14142|false|false|false|||sulfate
Finding|Functional Concept|SIMPLE_SEGMENT|14160,14170|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Finding|Organism Function|SIMPLE_SEGMENT|14160,14170|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Event|Event|SIMPLE_SEGMENT|14171,14174|false|false|false|||Q4H
Drug|Organic Chemical|SIMPLE_SEGMENT|14180,14191|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14180,14191|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14180,14202|false|false|false|C0939232|fluticasone / salmeterol|Fluticasone-Salmeterol
Drug|Organic Chemical|SIMPLE_SEGMENT|14180,14209|false|false|false|C4762496|Fluticasone-Salmeterol Diskus|Fluticasone-Salmeterol Diskus
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14180,14209|false|false|false|C4762496|Fluticasone-Salmeterol Diskus|Fluticasone-Salmeterol Diskus
Drug|Organic Chemical|SIMPLE_SEGMENT|14192,14202|false|false|false|C0073992|salmeterol|Salmeterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14192,14202|false|false|false|C0073992|salmeterol|Salmeterol
Event|Event|SIMPLE_SEGMENT|14203,14209|false|false|false|||Diskus
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|14222,14225|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Organic Chemical|SIMPLE_SEGMENT|14222,14225|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14222,14225|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Event|Event|SIMPLE_SEGMENT|14222,14225|false|false|false|||INH
Finding|Functional Concept|SIMPLE_SEGMENT|14222,14225|false|false|false|C0205535|Inhalation Route of Administration|INH
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|14229,14232|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|14229,14232|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|14229,14232|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|14229,14232|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|14229,14232|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|14238,14249|false|false|false|C0082607|fluticasone|fluticasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14238,14249|false|false|false|C0082607|fluticasone|fluticasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14238,14260|false|false|false|C0939232|fluticasone / salmeterol|fluticasone-salmeterol
Drug|Organic Chemical|SIMPLE_SEGMENT|14250,14260|false|false|false|C0073992|salmeterol|salmeterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14250,14260|false|false|false|C0073992|salmeterol|salmeterol
Event|Event|SIMPLE_SEGMENT|14250,14260|false|false|false|||salmeterol
Drug|Organic Chemical|SIMPLE_SEGMENT|14262,14268|false|false|false|C0965130|Advair|Advair
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14262,14268|false|false|false|C0965130|Advair|Advair
Drug|Organic Chemical|SIMPLE_SEGMENT|14262,14275|false|false|false|C0939246|Advair Diskus|Advair Diskus
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14262,14275|false|false|false|C0939246|Advair Diskus|Advair Diskus
Event|Event|SIMPLE_SEGMENT|14269,14275|false|false|false|||Diskus
Event|Event|SIMPLE_SEGMENT|14300,14304|false|false|false|||dose
Event|Event|SIMPLE_SEGMENT|14305,14312|false|false|false|||Inhaled
Finding|Idea or Concept|SIMPLE_SEGMENT|14321,14324|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|14321,14324|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|14334,14338|false|false|false|C1556138|Disc - Body Part|Disk
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|14334,14338|false|false|false|C0993608|Disk Drug Form|Disk
Event|Event|SIMPLE_SEGMENT|14339,14346|false|false|false|||Refills
Finding|Idea or Concept|SIMPLE_SEGMENT|14339,14346|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|14354,14363|false|false|false|C0024002|lorazepam|Lorazepam
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14354,14363|false|false|false|C0024002|lorazepam|Lorazepam
Finding|Gene or Genome|SIMPLE_SEGMENT|14378,14381|false|false|false|C1422467|CIAO3 gene|PRN
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|14382,14389|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|Anxiety
Event|Event|SIMPLE_SEGMENT|14382,14389|false|false|false|||Anxiety
Finding|Sign or Symptom|SIMPLE_SEGMENT|14382,14389|false|false|false|C0860603|Anxiety symptoms|Anxiety
Event|Event|SIMPLE_SEGMENT|14391,14393|false|false|false|||RX
Drug|Organic Chemical|SIMPLE_SEGMENT|14395,14404|false|false|false|C0024002|lorazepam|lorazepam
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14395,14404|false|false|false|C0024002|lorazepam|lorazepam
Event|Event|SIMPLE_SEGMENT|14395,14404|false|false|false|||lorazepam
Drug|Organic Chemical|SIMPLE_SEGMENT|14406,14412|false|false|false|C0699194|Ativan|Ativan
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14406,14412|false|false|false|C0699194|Ativan|Ativan
Event|Event|SIMPLE_SEGMENT|14406,14412|false|false|false|||Ativan
Finding|Functional Concept|SIMPLE_SEGMENT|14439,14447|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|14442,14447|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|14442,14447|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Intellectual Product|SIMPLE_SEGMENT|14448,14453|false|false|false|C1720374|Every - dosing instruction fragment|Every
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|14473,14479|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|14480,14487|false|false|false|||Refills
Finding|Idea or Concept|SIMPLE_SEGMENT|14480,14487|false|false|false|C0807726|refill|Refills
Event|Event|SIMPLE_SEGMENT|14494,14503|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|14494,14503|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|14494,14503|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|14494,14503|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|14494,14503|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14494,14515|false|false|false|C4019243||Discharge Disposition
Finding|Finding|SIMPLE_SEGMENT|14494,14515|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14504,14515|false|false|false|C2926604||Disposition
Event|Event|SIMPLE_SEGMENT|14504,14515|false|false|false|||Disposition
Procedure|Health Care Activity|SIMPLE_SEGMENT|14504,14515|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|SIMPLE_SEGMENT|14517,14521|false|false|false|||Home
Finding|Idea or Concept|SIMPLE_SEGMENT|14517,14521|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|SIMPLE_SEGMENT|14517,14521|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|SIMPLE_SEGMENT|14517,14521|false|false|false|C1553498|home health encounter|Home
Event|Occupational Activity|SIMPLE_SEGMENT|14527,14534|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|14527,14534|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Event|Event|SIMPLE_SEGMENT|14537,14545|false|false|false|||Facility
Finding|Intellectual Product|SIMPLE_SEGMENT|14537,14545|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|SIMPLE_SEGMENT|14553,14562|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|14553,14562|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|14553,14562|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|14553,14562|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|14553,14562|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|14553,14572|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14563,14572|false|false|false|C0945731||Diagnosis
Event|Event|SIMPLE_SEGMENT|14563,14572|false|false|false|||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|14563,14572|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|14563,14572|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|14563,14572|false|false|false|C0011900|Diagnosis|Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14574,14591|false|false|false|C0801658||Primary Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14582,14591|false|false|false|C0945731||Diagnosis
Event|Event|SIMPLE_SEGMENT|14582,14591|false|false|false|||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|14582,14591|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|14582,14591|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|14582,14591|false|false|false|C0011900|Diagnosis|Diagnosis
Finding|Intellectual Product|SIMPLE_SEGMENT|14593,14600|false|false|false|C1547296|Chronic - Admission Level of Care Code|Chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|14593,14600|false|false|false|C1555457|Provision of recurring care for chronic illness|Chronic
Finding|Pathologic Function|SIMPLE_SEGMENT|14593,14612|false|false|false|C0333166|Chronic obstruction|Chronic obstruction
Finding|Finding|SIMPLE_SEGMENT|14601,14612|false|false|false|C0028778|Obstruction|obstruction
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|14613,14622|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14613,14622|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|14613,14622|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14613,14630|false|false|false|C0024115|Lung diseases|pulmonary disease
Finding|Finding|SIMPLE_SEGMENT|14613,14630|false|false|false|C0455540|History of - respiratory disease|pulmonary disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14623,14630|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|14623,14630|false|false|false|||disease
Finding|Finding|SIMPLE_SEGMENT|14623,14643|false|false|false|C0235874|Disease Exacerbation|disease exacerbation
Event|Event|SIMPLE_SEGMENT|14631,14643|false|false|false|||exacerbation
Finding|Finding|SIMPLE_SEGMENT|14631,14643|false|false|false|C4086268|Exacerbation|exacerbation
Disorder|Neoplastic Process|SIMPLE_SEGMENT|14645,14654|false|false|false|C0027627|Neoplasm Metastasis|Secondary
Event|Event|SIMPLE_SEGMENT|14645,14654|false|false|false|||Secondary
Finding|Functional Concept|SIMPLE_SEGMENT|14645,14654|false|false|false|C1522484|metastatic qualifier|Secondary
Event|Event|SIMPLE_SEGMENT|14655,14664|false|false|false|||Diagnoses
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|14655,14664|false|false|false|C0011900|Diagnosis|Diagnoses
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|14666,14673|true|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|Tobacco
Drug|Immunologic Factor|SIMPLE_SEGMENT|14666,14673|true|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|Tobacco
Drug|Organic Chemical|SIMPLE_SEGMENT|14666,14673|true|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|Tobacco
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14666,14673|true|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|Tobacco
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14666,14677|false|false|false|C4522050||Tobacco use
Finding|Finding|SIMPLE_SEGMENT|14666,14677|false|false|false|C0040335;C0543414;C0841002;C3853727|Encounter due to tobacco use;History of tobacco use;Tobacco use;Tobacco user|Tobacco use
Finding|Individual Behavior|SIMPLE_SEGMENT|14666,14677|false|false|false|C0040335;C0543414;C0841002;C3853727|Encounter due to tobacco use;History of tobacco use;Tobacco use;Tobacco user|Tobacco use
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|14666,14686|false|false|false|C0040336|Tobacco Use Disorder|Tobacco use disorder
Event|Event|SIMPLE_SEGMENT|14674,14677|false|false|false|||use
Finding|Functional Concept|SIMPLE_SEGMENT|14674,14677|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|SIMPLE_SEGMENT|14674,14677|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14678,14686|false|false|false|C0012634|Disease|disorder
Event|Event|SIMPLE_SEGMENT|14678,14686|false|false|false|||disorder
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|14687,14693|false|false|false|C0018792|Heart Atrium|Atrial
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14687,14706|false|false|false|C2926591||Atrial fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14687,14706|false|false|false|C0004238|Atrial Fibrillation|Atrial fibrillation
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|14687,14706|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Atrial fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14694,14706|false|false|false|C0232197|Fibrillation|fibrillation
Event|Event|SIMPLE_SEGMENT|14694,14706|false|false|false|||fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14707,14719|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|SIMPLE_SEGMENT|14707,14719|false|false|false|||Hypertension
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|14720,14727|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|Anxiety
Event|Event|SIMPLE_SEGMENT|14720,14727|false|false|false|||Anxiety
Finding|Sign or Symptom|SIMPLE_SEGMENT|14720,14727|false|false|false|C0860603|Anxiety symptoms|Anxiety
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|14728,14736|false|false|false|C0018787|Heart|Coronary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|14728,14743|false|false|false|C0205042|Coronary artery|Coronary Artery
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14728,14751|false|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|Coronary Artery Disease
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|14737,14743|false|false|false|C0003842;C0226004|Arterial system;Arteries|Artery
Anatomy|Body System|SIMPLE_SEGMENT|14737,14743|false|false|false|C0003842;C0226004|Arterial system;Arteries|Artery
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14737,14751|false|false|false|C0852949|Arteriopathic disease|Artery Disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14744,14751|false|false|false|C0012634|Disease|Disease
Event|Event|SIMPLE_SEGMENT|14744,14751|false|false|false|||Disease
Event|Event|SIMPLE_SEGMENT|14755,14764|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|14755,14764|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|14755,14764|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|14755,14764|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|14755,14764|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14765,14774|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14765,14774|false|false|false|C0012634|Disease|Condition
Event|Event|SIMPLE_SEGMENT|14765,14774|false|false|false|||Condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|14765,14774|false|false|false|C1705253|Logical Condition|Condition
Finding|Mental Process|SIMPLE_SEGMENT|14776,14782|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14776,14789|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|SIMPLE_SEGMENT|14776,14789|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14783,14789|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|14783,14789|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|14791,14796|false|false|false|||Clear
Finding|Idea or Concept|SIMPLE_SEGMENT|14791,14796|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|SIMPLE_SEGMENT|14801,14809|false|false|false|||coherent
Finding|Finding|SIMPLE_SEGMENT|14801,14809|false|false|false|C4068804|Coherent|coherent
Event|Event|SIMPLE_SEGMENT|14811,14816|false|false|false|||Level
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14811,14833|false|false|false|C4050479||Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|14811,14833|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|SIMPLE_SEGMENT|14820,14833|false|false|false|||Consciousness
Finding|Finding|SIMPLE_SEGMENT|14820,14833|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|SIMPLE_SEGMENT|14820,14833|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14835,14840|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|14835,14840|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14835,14840|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|SIMPLE_SEGMENT|14835,14840|false|false|false|||Alert
Finding|Finding|SIMPLE_SEGMENT|14835,14840|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|14835,14840|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|14835,14840|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|SIMPLE_SEGMENT|14845,14856|false|false|false|||interactive
Finding|Functional Concept|SIMPLE_SEGMENT|14845,14856|false|false|false|C1704675|Interaction|interactive
Event|Activity|SIMPLE_SEGMENT|14858,14866|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|14858,14866|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|SIMPLE_SEGMENT|14858,14866|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14867,14873|false|false|false|C5889824||Status
Event|Event|SIMPLE_SEGMENT|14867,14873|false|false|false|||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|14867,14873|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|14875,14885|false|false|false|||Ambulatory
Finding|Functional Concept|SIMPLE_SEGMENT|14875,14885|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|SIMPLE_SEGMENT|14875,14885|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|SIMPLE_SEGMENT|14875,14885|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|SIMPLE_SEGMENT|14875,14885|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|SIMPLE_SEGMENT|14888,14899|false|false|false|||Independent
Finding|Finding|SIMPLE_SEGMENT|14888,14899|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|SIMPLE_SEGMENT|14888,14899|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Event|Event|SIMPLE_SEGMENT|14904,14913|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|14904,14913|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|14904,14913|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|14904,14913|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|14904,14913|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14904,14926|false|false|false|C3669312||Discharge Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|14904,14926|false|false|false|C4282220|Discharge instructions|Discharge Instructions
Procedure|Health Care Activity|SIMPLE_SEGMENT|14904,14926|false|false|false|C2266673|hospital discharge instructions (treatment)|Discharge Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14914,14926|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|14914,14926|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|14914,14926|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Finding|Gene or Genome|SIMPLE_SEGMENT|14928,14932|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Event|Event|SIMPLE_SEGMENT|14952,14961|false|false|false|||privilege
Finding|Conceptual Entity|SIMPLE_SEGMENT|14952,14961|false|false|false|C1547898;C1706335;C1706336|Privilege;Role Privilege;User Privilege|privilege
Finding|Idea or Concept|SIMPLE_SEGMENT|14952,14961|false|false|false|C1547898;C1706335;C1706336|Privilege;Role Privilege;User Privilege|privilege
Event|Activity|SIMPLE_SEGMENT|14969,14973|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|14969,14973|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|14969,14973|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|14969,14973|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|14969,14976|false|false|false|C1555558|care of - AddressPartType|care of
Event|Event|SIMPLE_SEGMENT|14993,15002|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|14993,15002|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|SIMPLE_SEGMENT|15021,15029|false|false|false|||admitted
Finding|Idea or Concept|SIMPLE_SEGMENT|15037,15045|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|SIMPLE_SEGMENT|15051,15060|false|false|false|||shortness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|15051,15070|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|SIMPLE_SEGMENT|15051,15070|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|SIMPLE_SEGMENT|15064,15070|false|false|false|C0225386|Breath|breath
Event|Event|SIMPLE_SEGMENT|15075,15082|false|false|false|||concern
Finding|Idea or Concept|SIMPLE_SEGMENT|15075,15082|false|false|false|C2699424|Concern|concern
Event|Event|SIMPLE_SEGMENT|15106,15111|false|false|false|||flare
Finding|Finding|SIMPLE_SEGMENT|15106,15111|false|false|false|C1517205;C3540542|Exacerbation of cGVHD;Flare|flare
Finding|Sign or Symptom|SIMPLE_SEGMENT|15106,15111|false|false|false|C1517205;C3540542|Exacerbation of cGVHD;Flare|flare
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15121,15125|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|15121,15125|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|SIMPLE_SEGMENT|15121,15125|false|false|false|||COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|15121,15125|false|false|false|C1412502|ARCN1 gene|COPD
Finding|Idea or Concept|SIMPLE_SEGMENT|15141,15149|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|SIMPLE_SEGMENT|15153,15162|false|false|false|||increased
Event|Event|SIMPLE_SEGMENT|15168,15172|false|false|false|||dose
Drug|Organic Chemical|SIMPLE_SEGMENT|15176,15184|false|false|true|C0038317|Steroids|steroids
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|15176,15184|false|false|true|C0038317|Steroids|steroids
Event|Event|SIMPLE_SEGMENT|15176,15184|false|false|false|||steroids
Event|Event|SIMPLE_SEGMENT|15188,15192|false|false|false|||help
Finding|Intellectual Product|SIMPLE_SEGMENT|15188,15192|false|false|false|C1552861|Help document|help
Attribute|Clinical Attribute|SIMPLE_SEGMENT|15199,15208|false|false|false|C5885990||breathing
Event|Event|SIMPLE_SEGMENT|15199,15208|false|false|false|||breathing
Finding|Finding|SIMPLE_SEGMENT|15199,15208|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|SIMPLE_SEGMENT|15199,15208|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|SIMPLE_SEGMENT|15199,15208|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|SIMPLE_SEGMENT|15199,15208|false|false|false|C1160636|respiratory system process|breathing
Event|Event|SIMPLE_SEGMENT|15219,15227|false|false|false|||received
Event|Event|SIMPLE_SEGMENT|15246,15256|false|false|false|||treatments
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|15246,15256|false|false|false|C0087111|Therapeutic procedure|treatments
Event|Event|SIMPLE_SEGMENT|15263,15269|false|false|false|||helped
Attribute|Clinical Attribute|SIMPLE_SEGMENT|15275,15284|false|false|false|C5885990||breathing
Event|Event|SIMPLE_SEGMENT|15275,15284|false|false|false|||breathing
Finding|Finding|SIMPLE_SEGMENT|15275,15284|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|SIMPLE_SEGMENT|15275,15284|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|SIMPLE_SEGMENT|15275,15284|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|SIMPLE_SEGMENT|15275,15284|false|false|false|C1160636|respiratory system process|breathing
Event|Event|SIMPLE_SEGMENT|15300,15310|false|false|false|||expressing
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|15317,15324|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Event|Event|SIMPLE_SEGMENT|15317,15324|false|false|false|||anxiety
Finding|Sign or Symptom|SIMPLE_SEGMENT|15317,15324|false|false|false|C0860603|Anxiety symptoms|anxiety
Event|Event|SIMPLE_SEGMENT|15344,15356|false|false|false|||contributing
Event|Event|SIMPLE_SEGMENT|15365,15374|false|false|false|||shortness
Event|Event|SIMPLE_SEGMENT|15379,15385|false|false|false|||breath
Finding|Body Substance|SIMPLE_SEGMENT|15379,15385|false|false|false|C0225386|Breath|breath
Event|Event|SIMPLE_SEGMENT|15396,15401|false|false|false|||given
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|15404,15414|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|15404,15414|false|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|15404,15414|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|SIMPLE_SEGMENT|15415,15421|false|false|false|||called
Drug|Organic Chemical|SIMPLE_SEGMENT|15422,15428|false|false|false|C0699194|Ativan|Ativan
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|15422,15428|false|false|false|C0699194|Ativan|Ativan
Event|Event|SIMPLE_SEGMENT|15422,15428|false|false|false|||Ativan
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|15439,15446|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Event|Event|SIMPLE_SEGMENT|15439,15446|false|false|false|||anxiety
Finding|Sign or Symptom|SIMPLE_SEGMENT|15439,15446|false|false|false|C0860603|Anxiety symptoms|anxiety
Event|Event|SIMPLE_SEGMENT|15457,15463|false|false|false|||seemed
Event|Event|SIMPLE_SEGMENT|15467,15471|false|false|false|||help
Attribute|Clinical Attribute|SIMPLE_SEGMENT|15477,15486|false|false|false|C5885990||breathing
Event|Event|SIMPLE_SEGMENT|15477,15486|false|false|false|||breathing
Finding|Finding|SIMPLE_SEGMENT|15477,15486|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|SIMPLE_SEGMENT|15477,15486|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|SIMPLE_SEGMENT|15477,15486|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|SIMPLE_SEGMENT|15477,15486|false|false|false|C1160636|respiratory system process|breathing
Event|Event|SIMPLE_SEGMENT|15501,15510|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|15501,15510|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|SIMPLE_SEGMENT|15520,15524|false|false|false|||seen
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|15532,15541|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|15532,15541|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|15532,15541|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Event|Event|SIMPLE_SEGMENT|15543,15554|false|false|false|||specialists
Event|Event|SIMPLE_SEGMENT|15561,15572|false|false|false|||recommended
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|15575,15582|false|false|false|C0040405|X-Ray Computed Tomography|CT scan
Event|Event|SIMPLE_SEGMENT|15578,15582|false|false|false|||scan
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|15578,15582|false|false|false|C0034606;C0441633|Radionuclide Imaging;Scanning|scan
Event|Event|SIMPLE_SEGMENT|15588,15594|false|false|false|||showed
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15620,15624|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|15620,15624|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|SIMPLE_SEGMENT|15620,15624|false|false|false|||COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|15620,15624|false|false|false|C1412502|ARCN1 gene|COPD
Event|Event|SIMPLE_SEGMENT|15637,15641|true|false|false|||show
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15646,15655|true|false|false|C0009450|Communicable Diseases|infection
Event|Event|SIMPLE_SEGMENT|15646,15655|true|false|false|||infection
Finding|Pathologic Function|SIMPLE_SEGMENT|15646,15655|true|false|false|C3714514|Infection|infection
Event|Event|SIMPLE_SEGMENT|15668,15677|false|false|false|||suggested
Event|Event|SIMPLE_SEGMENT|15678,15688|false|false|false|||increasing
Event|Event|SIMPLE_SEGMENT|15693,15697|false|false|false|||dose
Drug|Organic Chemical|SIMPLE_SEGMENT|15706,15712|false|false|false|C0965130|Advair|Advair
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|15706,15712|false|false|false|C0965130|Advair|Advair
Event|Event|SIMPLE_SEGMENT|15713,15720|false|false|false|||inhaler
Finding|Functional Concept|SIMPLE_SEGMENT|15713,15720|false|false|false|C4319647|Inhaler (unit of presentation)|inhaler
Event|Event|SIMPLE_SEGMENT|15745,15749|false|false|false|||feel
Event|Event|SIMPLE_SEGMENT|15750,15755|false|false|false|||short
Finding|Sign or Symptom|SIMPLE_SEGMENT|15750,15765|false|false|false|C0013404|Dyspnea|short of breath
Finding|Body Substance|SIMPLE_SEGMENT|15759,15765|false|false|false|C0225386|Breath|breath
Event|Event|SIMPLE_SEGMENT|15780,15785|false|false|false|||check
Drug|Biologically Active Substance|SIMPLE_SEGMENT|15791,15797|false|false|false|C0030054|oxygen|oxygen
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|15791,15797|false|false|false|C0030054|oxygen|oxygen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|15791,15797|false|false|false|C0030054|oxygen|oxygen
Event|Event|SIMPLE_SEGMENT|15791,15797|false|false|false|||oxygen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|15791,15797|false|false|false|C0184633|Oxygen Therapy Care|oxygen
Drug|Biologically Active Substance|SIMPLE_SEGMENT|15841,15847|false|false|false|C0030054|oxygen|oxygen
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|15841,15847|false|false|false|C0030054|oxygen|oxygen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|15841,15847|false|false|false|C0030054|oxygen|oxygen
Event|Event|SIMPLE_SEGMENT|15841,15847|false|false|false|||oxygen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|15841,15847|false|false|false|C0184633|Oxygen Therapy Care|oxygen
Event|Event|SIMPLE_SEGMENT|15858,15865|false|false|false|||inhaler
Finding|Functional Concept|SIMPLE_SEGMENT|15858,15865|false|false|false|C4319647|Inhaler (unit of presentation)|inhaler
Event|Event|SIMPLE_SEGMENT|15882,15886|true|false|false|||wait
Attribute|Clinical Attribute|SIMPLE_SEGMENT|15913,15917|false|false|false|C4318566|Deep Resection Margin|deep
Event|Event|SIMPLE_SEGMENT|15919,15926|false|false|false|||breaths
Finding|Body Substance|SIMPLE_SEGMENT|15919,15926|false|false|false|C0225386|Breath|breaths
Event|Event|SIMPLE_SEGMENT|15931,15934|false|false|false|||see
Event|Event|SIMPLE_SEGMENT|15943,15952|false|false|false|||shortness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|15943,15962|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|SIMPLE_SEGMENT|15943,15962|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|SIMPLE_SEGMENT|15956,15962|false|false|false|C0225386|Breath|breath
Event|Event|SIMPLE_SEGMENT|15963,15971|false|false|false|||improves
Finding|Finding|SIMPLE_SEGMENT|15963,15971|false|false|false|C0184511|Improved|improves
Event|Event|SIMPLE_SEGMENT|15982,15985|false|false|false|||use
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|15990,16000|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|15990,16000|false|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|15990,16000|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|SIMPLE_SEGMENT|16001,16007|false|false|false|||called
Drug|Organic Chemical|SIMPLE_SEGMENT|16008,16014|false|false|false|C0699194|Ativan|Ativan
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|16008,16014|false|false|false|C0699194|Ativan|Ativan
Drug|Organic Chemical|SIMPLE_SEGMENT|16015,16024|false|false|false|C0024002|lorazepam|lorazepam
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|16015,16024|false|false|false|C0024002|lorazepam|lorazepam
Event|Event|SIMPLE_SEGMENT|16015,16024|false|false|false|||lorazepam
Event|Event|SIMPLE_SEGMENT|16029,16033|false|false|false|||help
Event|Event|SIMPLE_SEGMENT|16044,16053|true|false|false|||shortness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|16044,16063|true|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|SIMPLE_SEGMENT|16044,16063|true|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|SIMPLE_SEGMENT|16057,16063|true|false|false|C0225386|Breath|breath
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|16083,16088|true|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|SIMPLE_SEGMENT|16091,16094|true|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|16091,16094|true|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|16100,16105|true|false|false|C1410088|Still|still
Event|Event|SIMPLE_SEGMENT|16111,16119|true|false|false|||improved
Event|Event|SIMPLE_SEGMENT|16129,16132|true|false|false|||use
Drug|Biologically Active Substance|SIMPLE_SEGMENT|16153,16159|false|false|false|C0030054|oxygen|oxygen
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|16153,16159|false|false|false|C0030054|oxygen|oxygen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|16153,16159|false|false|false|C0030054|oxygen|oxygen
Event|Event|SIMPLE_SEGMENT|16153,16159|false|false|false|||oxygen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|16153,16159|false|false|false|C0184633|Oxygen Therapy Care|oxygen
Event|Event|SIMPLE_SEGMENT|16170,16176|false|false|false|||follow
Event|Activity|SIMPLE_SEGMENT|16194,16206|false|false|false|C0003629|Appointments|appointments
Event|Event|SIMPLE_SEGMENT|16194,16206|false|false|false|||appointments
Event|Event|SIMPLE_SEGMENT|16228,16236|false|false|false|||continue
Event|Event|SIMPLE_SEGMENT|16240,16244|false|false|false|||take
Attribute|Clinical Attribute|SIMPLE_SEGMENT|16257,16268|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|16257,16268|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|16257,16268|false|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|16257,16268|false|false|false|C4284232|Medications|medications
Event|Event|SIMPLE_SEGMENT|16272,16282|false|false|false|||prescribed
Event|Event|SIMPLE_SEGMENT|16292,16302|true|false|false|||experience
Finding|Gene or Genome|SIMPLE_SEGMENT|16314,16320|true|false|false|C1428845|ITPRIP gene|danger
Event|Event|SIMPLE_SEGMENT|16321,16326|true|false|false|||signs
Finding|Finding|SIMPLE_SEGMENT|16321,16326|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|SIMPLE_SEGMENT|16321,16326|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Event|Event|SIMPLE_SEGMENT|16345,16349|false|false|false|||call
Finding|Intellectual Product|SIMPLE_SEGMENT|16356,16362|false|false|false|C2348314|Doctor - Title|doctor
Event|Event|SIMPLE_SEGMENT|16378,16380|false|false|false|||go
Event|Event|SIMPLE_SEGMENT|16388,16397|false|false|false|||Emergency
Finding|Finding|SIMPLE_SEGMENT|16388,16397|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Finding|Idea or Concept|SIMPLE_SEGMENT|16388,16397|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Finding|Intellectual Product|SIMPLE_SEGMENT|16388,16397|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Finding|Pathologic Function|SIMPLE_SEGMENT|16388,16397|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|16388,16397|false|false|false|C0013956|Emergency Situation|Emergency
Procedure|Health Care Activity|SIMPLE_SEGMENT|16388,16397|false|false|false|C1553500|emergency encounter|Emergency
Finding|Idea or Concept|SIMPLE_SEGMENT|16388,16402|false|false|false|C1546435|Encounter Referral Source - emergency room|Emergency Room
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|16421,16425|false|false|false|C0339510|Vitelliform Macular Dystrophy|best
Event|Event|SIMPLE_SEGMENT|16421,16425|false|false|false|||best
Finding|Gene or Genome|SIMPLE_SEGMENT|16421,16425|false|false|false|C1826421;C5781213|BEST1 gene;BEST1 wt Allele|best
Event|Activity|SIMPLE_SEGMENT|16448,16452|false|false|false|C1947933|care activity|Care
Finding|Finding|SIMPLE_SEGMENT|16448,16452|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|SIMPLE_SEGMENT|16448,16452|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Attribute|Clinical Attribute|SIMPLE_SEGMENT|16448,16457|false|false|false|C4321316||Care Team
Finding|Finding|SIMPLE_SEGMENT|16448,16457|false|false|false|C4321315|Care team|Care Team
Procedure|Health Care Activity|SIMPLE_SEGMENT|16460,16468|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|16469,16481|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|16469,16481|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|16469,16481|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

