 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
.|12,13
Unit|23,27
No|28,30
:|30,31
_|34,35
_|35,36
_|36,37
<EOL>|37,38
<EOL>|39,40
Admission|40,49
Date|50,54
:|54,55
_|57,58
_|58,59
_|59,60
Discharge|74,83
Date|84,88
:|88,89
_|92,93
_|93,94
_|94,95
<EOL>|95,96
<EOL>|97,98
Date|98,102
of|103,105
Birth|106,111
:|111,112
_|114,115
_|115,116
_|116,117
Sex|130,133
:|133,134
F|137,138
<EOL>|138,139
<EOL>|140,141
Service|141,148
:|148,149
MEDICINE|150,158
<EOL>|158,159
<EOL>|160,161
Allergies|161,170
:|170,171
<EOL>|172,173
Patient|173,180
recorded|181,189
as|190,192
having|193,199
No|200,202
Known|203,208
Allergies|209,218
to|219,221
Drugs|222,227
<EOL>|227,228
<EOL>|229,230
Attending|230,239
:|239,240
_|241,242
_|242,243
_|243,244
<EOL>|244,245
<EOL>|246,247
Chief|247,252
Complaint|253,262
:|262,263
<EOL>|263,264
Abdominal|264,273
distention|274,284
.|284,285
<EOL>|285,286
<EOL>|287,288
Major|288,293
Surgical|294,302
or|303,305
Invasive|306,314
Procedure|315,324
:|324,325
<EOL>|325,326
Paracentesis|326,338
.|338,339
<EOL>|339,340
<EOL>|341,342
History|342,349
of|350,352
Present|353,360
Illness|361,368
:|368,369
<EOL>|369,370
This|370,374
is|375,377
a|378,379
very|380,384
nice|385,389
_|390,391
_|391,392
_|392,393
woman|394,399
with|400,404
ETOH|405,409
abuse|410,415
who|416,419
<EOL>|420,421
presents|421,429
with|430,434
constipation|435,447
,|447,448
abdominal|449,458
distention|459,469
x|470,471
10|472,474
days|475,479
.|479,480
<EOL>|482,483
Patient|483,490
drinks|491,497
about|498,503
_|504,505
_|505,506
_|506,507
glasses|508,515
of|516,518
wine|519,523
per|524,527
night|528,533
and|534,537
went|538,542
on|543,545
a|546,547
<EOL>|548,549
2|549,550
month|551,556
binge|557,562
drinking|563,571
~|572,573
10|573,575
/|575,576
day|576,579
,|579,580
which|581,586
ended|587,592
about|593,598
1|599,600
month|601,606
ago|607,610
.|610,611
<EOL>|613,614
She|614,617
noted|618,623
abdominal|624,633
distension|634,644
progressive|645,656
over|657,661
the|662,665
past|666,670
week|671,675
<EOL>|676,677
and|677,680
has|681,684
also|685,689
not|690,693
had|694,697
a|698,699
solid|700,705
stool|706,711
x|712,713
7|714,715
days|716,720
.|720,721
She|723,726
denies|727,733
any|734,737
<EOL>|738,739
f|739,740
/|740,741
C|741,742
/|742,743
NS|743,745
,|745,746
CP|747,749
/|749,750
SOB|750,753
/|753,754
DOE|754,757
or|758,760
decrease|761,769
in|770,772
her|773,776
excercise|777,786
tolerance|787,796
.|796,797
No|799,801
<EOL>|802,803
recent|803,809
travel|810,816
but|817,820
has|821,824
traveled|825,833
to|834,836
_|837,838
_|838,839
_|839,840
and|841,844
_|845,846
_|846,847
_|847,848
<EOL>|849,850
previously|850,860
.|860,861
No|863,865
NSAIDs|866,872
,|872,873
Tylenol|874,881
or|882,884
OTC|885,888
medications|889,900
other|901,906
than|907,911
<EOL>|912,913
occasional|913,923
peptobismol|924,935
.|935,936
She|938,941
notes|942,947
that|948,952
she|953,956
has|957,960
missed|961,967
her|968,971
past|972,976
<EOL>|977,978
two|978,981
periods|982,989
.|989,990
<EOL>|992,993
<EOL>|993,994
In|994,996
ED|997,999
,|999,1000
bedside|1001,1008
US|1009,1011
with|1012,1016
ascites|1017,1024
.|1024,1025
CT|1027,1029
with|1030,1034
fatty|1035,1040
liver|1041,1046
,|1046,1047
good|1048,1052
<EOL>|1053,1054
portal|1054,1060
flow|1061,1065
.|1065,1066
Patient|1068,1075
with|1076,1080
HR|1081,1083
110|1084,1087
in|1088,1090
ED|1091,1093
,|1093,1094
for|1095,1098
IV|1099,1101
5mg|1102,1105
valium|1106,1112
.|1112,1113
Got|1115,1118
<EOL>|1119,1120
NS|1120,1122
IVF|1123,1126
at|1127,1129
100cc|1130,1135
/|1135,1136
hr|1136,1138
and|1139,1142
thiamine|1143,1151
100mg|1152,1157
IV|1158,1160
.|1160,1161
<EOL>|1161,1162
<EOL>|1163,1164
Past|1164,1168
Medical|1169,1176
History|1177,1184
:|1184,1185
<EOL>|1185,1186
-|1186,1187
-|1187,1188
Alcohol|1188,1195
abuse|1196,1201
<EOL>|1201,1202
-|1202,1203
-|1203,1204
Chronic|1204,1211
back|1212,1216
pain|1217,1221
<EOL>|1221,1222
<EOL>|1223,1224
Social|1224,1230
History|1231,1238
:|1238,1239
<EOL>|1239,1240
_|1240,1241
_|1241,1242
_|1242,1243
<EOL>|1243,1244
Family|1244,1250
History|1251,1258
:|1258,1259
<EOL>|1259,1260
Breast|1260,1266
Ca|1267,1269
in|1270,1272
mother|1273,1279
age|1280,1283
_|1284,1285
_|1285,1286
_|1286,1287
,|1287,1288
No|1289,1291
IBD|1292,1295
,|1295,1296
liver|1297,1302
failure|1303,1310
.|1310,1311
Multiple|1313,1321
<EOL>|1322,1323
relatives|1323,1332
with|1333,1337
alcoholism|1338,1348
.|1348,1349
<EOL>|1349,1350
<EOL>|1351,1352
Physical|1352,1360
Exam|1361,1365
:|1365,1366
<EOL>|1366,1367
VS|1367,1369
:|1369,1370
97.9|1371,1375
,|1375,1376
103|1377,1380
/|1380,1381
73|1381,1383
,|1383,1384
86|1385,1387
,|1387,1388
18|1389,1391
,|1391,1392
96|1393,1395
%|1395,1396
RA|1397,1399
<EOL>|1401,1402
GEN|1402,1405
:|1405,1406
A|1407,1408
/|1408,1409
Ox3|1409,1412
,|1412,1413
pleasant|1414,1422
,|1422,1423
appropriate|1424,1435
,|1435,1436
well|1437,1441
appearing|1442,1451
<EOL>|1453,1454
HEENT|1454,1459
:|1459,1460
No|1461,1463
temporal|1464,1472
wasting|1473,1480
,|1480,1481
JVD|1482,1485
not|1486,1489
elevated|1490,1498
,|1498,1499
neck|1500,1504
veins|1505,1510
fill|1511,1515
<EOL>|1516,1517
from|1517,1521
above|1522,1527
.|1527,1528
<EOL>|1530,1531
CV|1531,1533
:|1533,1534
RRR|1535,1538
,|1538,1539
No|1540,1542
MRG|1543,1546
<EOL>|1548,1549
PULM|1549,1553
:|1553,1554
CTAB|1555,1559
but|1560,1563
decreased|1564,1573
BS|1574,1576
in|1577,1579
R|1580,1581
base|1582,1586
.|1586,1587
<EOL>|1589,1590
ABD|1590,1593
:|1593,1594
Distended|1595,1604
and|1605,1608
tight|1609,1614
,|1614,1615
diffusely|1616,1625
tender|1626,1632
to|1633,1635
palpation|1636,1645
,|1645,1646
BS|1647,1649
+|1649,1650
,|1650,1651
+|1652,1653
<EOL>|1654,1655
passing|1655,1662
flatulence|1663,1673
.|1673,1674
<EOL>|1676,1677
LIMBS|1677,1682
:|1682,1683
2|1684,1685
+|1685,1686
edema|1687,1692
of|1693,1695
the|1696,1699
LEs|1700,1703
to|1704,1706
knee|1707,1711
bilaterally|1712,1723
_|1724,1725
_|1725,1726
_|1726,1727
pulses|1728,1734
2|1735,1736
+|1736,1737
<EOL>|1738,1739
bilaterally|1739,1750
<EOL>|1752,1753
NEURO|1753,1758
:|1758,1759
No|1760,1762
asterixis|1763,1772
,|1772,1773
very|1774,1778
mild|1779,1783
general|1784,1791
tremor|1792,1798
.|1798,1799
<EOL>|1801,1802
<EOL>|1802,1803
<EOL>|1804,1805
Pertinent|1805,1814
Results|1815,1822
:|1822,1823
<EOL>|1823,1824
_|1824,1825
_|1825,1826
_|1826,1827
04|1828,1830
:|1830,1831
50AM|1831,1835
BLOOD|1836,1841
WBC|1842,1845
-|1845,1846
12|1846,1848
.|1848,1849
2|1849,1850
*|1850,1851
RBC|1852,1855
-|1855,1856
3|1856,1857
.|1857,1858
37|1858,1860
*|1860,1861
Hgb|1862,1865
-|1865,1866
12.0|1866,1870
Hct|1871,1874
-|1874,1875
37.2|1875,1879
<EOL>|1880,1881
MCV|1881,1884
-|1884,1885
110|1885,1888
*|1888,1889
MCH|1890,1893
-|1893,1894
35|1894,1896
.|1896,1897
5|1897,1898
*|1898,1899
MCHC|1900,1904
-|1904,1905
32.2|1905,1909
RDW|1910,1913
-|1913,1914
13.9|1914,1918
Plt|1919,1922
_|1923,1924
_|1924,1925
_|1925,1926
<EOL>|1926,1927
_|1927,1928
_|1928,1929
_|1929,1930
04|1931,1933
:|1933,1934
50AM|1934,1938
BLOOD|1939,1944
WBC|1945,1948
-|1948,1949
11|1949,1951
.|1951,1952
5|1952,1953
*|1953,1954
RBC|1955,1958
-|1958,1959
3|1959,1960
.|1960,1961
52|1961,1963
*|1963,1964
Hgb|1965,1968
-|1968,1969
12.2|1969,1973
Hct|1974,1977
-|1977,1978
37.7|1978,1982
<EOL>|1983,1984
MCV|1984,1987
-|1987,1988
107|1988,1991
*|1991,1992
MCH|1993,1996
-|1996,1997
34|1997,1999
.|1999,2000
6|2000,2001
*|2001,2002
MCHC|2003,2007
-|2007,2008
32.3|2008,2012
RDW|2013,2016
-|2016,2017
13.3|2017,2021
Plt|2022,2025
_|2026,2027
_|2027,2028
_|2028,2029
<EOL>|2029,2030
_|2030,2031
_|2031,2032
_|2032,2033
04|2034,2036
:|2036,2037
55AM|2037,2041
BLOOD|2042,2047
WBC|2048,2051
-|2051,2052
11|2052,2054
.|2054,2055
6|2055,2056
*|2056,2057
RBC|2058,2061
-|2061,2062
3|2062,2063
.|2063,2064
67|2064,2066
*|2066,2067
Hgb|2068,2071
-|2071,2072
12.8|2072,2076
Hct|2077,2080
-|2080,2081
39.0|2081,2085
<EOL>|2086,2087
MCV|2087,2090
-|2090,2091
106|2091,2094
*|2094,2095
MCH|2096,2099
-|2099,2100
34|2100,2102
.|2102,2103
8|2103,2104
*|2104,2105
MCHC|2106,2110
-|2110,2111
32.7|2111,2115
RDW|2116,2119
-|2119,2120
13.2|2120,2124
Plt|2125,2128
_|2129,2130
_|2130,2131
_|2131,2132
<EOL>|2132,2133
_|2133,2134
_|2134,2135
_|2135,2136
06|2137,2139
:|2139,2140
35AM|2140,2144
BLOOD|2145,2150
WBC|2151,2154
-|2154,2155
12|2155,2157
.|2157,2158
2|2158,2159
*|2159,2160
RBC|2161,2164
-|2164,2165
3|2165,2166
.|2166,2167
37|2167,2169
*|2169,2170
Hgb|2171,2174
-|2174,2175
12.0|2175,2179
Hct|2180,2183
-|2183,2184
36.4|2184,2188
<EOL>|2189,2190
MCV|2190,2193
-|2193,2194
108|2194,2197
*|2197,2198
MCH|2199,2202
-|2202,2203
35|2203,2205
.|2205,2206
7|2206,2207
*|2207,2208
MCHC|2209,2213
-|2213,2214
33.1|2214,2218
RDW|2219,2222
-|2222,2223
13.3|2223,2227
Plt|2228,2231
_|2232,2233
_|2233,2234
_|2234,2235
<EOL>|2235,2236
_|2236,2237
_|2237,2238
_|2238,2239
09|2240,2242
:|2242,2243
00AM|2243,2247
BLOOD|2248,2253
WBC|2254,2257
-|2257,2258
13|2258,2260
.|2260,2261
7|2261,2262
*|2262,2263
RBC|2264,2267
-|2267,2268
3|2268,2269
.|2269,2270
35|2270,2272
*|2272,2273
Hgb|2274,2277
-|2277,2278
11|2278,2280
.|2280,2281
6|2281,2282
*|2282,2283
Hct|2284,2287
-|2287,2288
35|2288,2290
.|2290,2291
6|2291,2292
*|2292,2293
<EOL>|2294,2295
MCV|2295,2298
-|2298,2299
106|2299,2302
*|2302,2303
MCH|2304,2307
-|2307,2308
34|2308,2310
.|2310,2311
5|2311,2312
*|2312,2313
MCHC|2314,2318
-|2318,2319
32.5|2319,2323
RDW|2324,2327
-|2327,2328
13.1|2328,2332
Plt|2333,2336
_|2337,2338
_|2338,2339
_|2339,2340
<EOL>|2340,2341
_|2341,2342
_|2342,2343
_|2343,2344
11|2345,2347
:|2347,2348
30AM|2348,2352
BLOOD|2353,2358
WBC|2359,2362
-|2362,2363
14|2363,2365
.|2365,2366
4|2366,2367
*|2367,2368
RBC|2369,2372
-|2372,2373
3|2373,2374
.|2374,2375
80|2375,2377
*|2377,2378
Hgb|2379,2382
-|2382,2383
13.2|2383,2387
Hct|2388,2391
-|2391,2392
40.3|2392,2396
<EOL>|2397,2398
MCV|2398,2401
-|2401,2402
106|2402,2405
*|2405,2406
MCH|2407,2410
-|2410,2411
34|2411,2413
.|2413,2414
8|2414,2415
*|2415,2416
MCHC|2417,2421
-|2421,2422
32.8|2422,2426
RDW|2427,2430
-|2430,2431
13.6|2431,2435
Plt|2436,2439
_|2440,2441
_|2441,2442
_|2442,2443
<EOL>|2443,2444
_|2444,2445
_|2445,2446
_|2446,2447
11|2448,2450
:|2450,2451
30AM|2451,2455
BLOOD|2456,2461
Neuts|2462,2467
-|2467,2468
80|2468,2470
.|2470,2471
6|2471,2472
*|2472,2473
Lymphs|2474,2480
-|2480,2481
11|2481,2483
.|2483,2484
7|2484,2485
*|2485,2486
Monos|2487,2492
-|2492,2493
5.5|2493,2496
<EOL>|2497,2498
Eos|2498,2501
-|2501,2502
0.5|2502,2505
Baso|2506,2510
-|2510,2511
1.7|2511,2514
<EOL>|2514,2515
_|2515,2516
_|2516,2517
_|2517,2518
04|2519,2521
:|2521,2522
50AM|2522,2526
BLOOD|2527,2532
Plt|2533,2536
_|2537,2538
_|2538,2539
_|2539,2540
<EOL>|2540,2541
_|2541,2542
_|2542,2543
_|2543,2544
04|2545,2547
:|2547,2548
50AM|2548,2552
BLOOD|2553,2558
_|2559,2560
_|2560,2561
_|2561,2562
PTT|2563,2566
-|2566,2567
35.0|2567,2571
_|2572,2573
_|2573,2574
_|2574,2575
<EOL>|2575,2576
_|2576,2577
_|2577,2578
_|2578,2579
:|2579,2580
50AM|2580,2584
BLOOD|2585,2590
Plt|2591,2594
_|2595,2596
_|2596,2597
_|2597,2598
<EOL>|2598,2599
_|2599,2600
_|2600,2601
_|2601,2602
04|2603,2605
:|2605,2606
50AM|2606,2610
BLOOD|2611,2616
_|2617,2618
_|2618,2619
_|2619,2620
PTT|2621,2624
-|2624,2625
36|2625,2627
.|2627,2628
3|2628,2629
*|2629,2630
_|2631,2632
_|2632,2633
_|2633,2634
<EOL>|2634,2635
_|2635,2636
_|2636,2637
_|2637,2638
04|2639,2641
:|2641,2642
55AM|2642,2646
BLOOD|2647,2652
Plt|2653,2656
_|2657,2658
_|2658,2659
_|2659,2660
<EOL>|2660,2661
_|2661,2662
_|2662,2663
_|2663,2664
04|2665,2667
:|2667,2668
55AM|2668,2672
BLOOD|2673,2678
_|2679,2680
_|2680,2681
_|2681,2682
PTT|2683,2686
-|2686,2687
32.4|2687,2691
_|2692,2693
_|2693,2694
_|2694,2695
<EOL>|2695,2696
_|2696,2697
_|2697,2698
_|2698,2699
06|2700,2702
:|2702,2703
35AM|2703,2707
BLOOD|2708,2713
Plt|2714,2717
_|2718,2719
_|2719,2720
_|2720,2721
<EOL>|2721,2722
_|2722,2723
_|2723,2724
_|2724,2725
06|2726,2728
:|2728,2729
35AM|2729,2733
BLOOD|2734,2739
_|2740,2741
_|2741,2742
_|2742,2743
PTT|2744,2747
-|2747,2748
32.5|2748,2752
_|2753,2754
_|2754,2755
_|2755,2756
<EOL>|2756,2757
_|2757,2758
_|2758,2759
_|2759,2760
09|2761,2763
:|2763,2764
00AM|2764,2768
BLOOD|2769,2774
Plt|2775,2778
_|2779,2780
_|2780,2781
_|2781,2782
<EOL>|2782,2783
_|2783,2784
_|2784,2785
_|2785,2786
11|2787,2789
:|2789,2790
30AM|2790,2794
BLOOD|2795,2800
_|2801,2802
_|2802,2803
_|2803,2804
PTT|2805,2808
-|2808,2809
26.0|2809,2813
_|2814,2815
_|2815,2816
_|2816,2817
<EOL>|2817,2818
_|2818,2819
_|2819,2820
_|2820,2821
11|2822,2824
:|2824,2825
30AM|2825,2829
BLOOD|2830,2835
Plt|2836,2839
_|2840,2841
_|2841,2842
_|2842,2843
<EOL>|2843,2844
_|2844,2845
_|2845,2846
_|2846,2847
04|2848,2850
:|2850,2851
50AM|2851,2855
BLOOD|2856,2861
Glucose|2862,2869
-|2869,2870
156|2870,2873
*|2873,2874
UreaN|2875,2880
-|2880,2881
5|2881,2882
*|2882,2883
Creat|2884,2889
-|2889,2890
0|2890,2891
.|2891,2892
3|2892,2893
*|2893,2894
Na|2895,2897
-|2897,2898
129|2898,2901
*|2901,2902
<EOL>|2903,2904
K|2904,2905
-|2905,2906
3.6|2906,2909
Cl|2910,2912
-|2912,2913
95|2913,2915
*|2915,2916
HCO3|2917,2921
-|2921,2922
25|2922,2924
AnGap|2925,2930
-|2930,2931
13|2931,2933
<EOL>|2933,2934
_|2934,2935
_|2935,2936
_|2936,2937
04|2938,2940
:|2940,2941
50AM|2941,2945
BLOOD|2946,2951
Glucose|2952,2959
-|2959,2960
113|2960,2963
*|2963,2964
UreaN|2965,2970
-|2970,2971
4|2971,2972
*|2972,2973
Creat|2974,2979
-|2979,2980
0|2980,2981
.|2981,2982
3|2982,2983
*|2983,2984
Na|2985,2987
-|2987,2988
131|2988,2991
*|2991,2992
<EOL>|2993,2994
K|2994,2995
-|2995,2996
3|2996,2997
.|2997,2998
2|2998,2999
*|2999,3000
Cl|3001,3003
-|3003,3004
96|3004,3006
HCO3|3007,3011
-|3011,3012
27|3012,3014
AnGap|3015,3020
-|3020,3021
11|3021,3023
<EOL>|3023,3024
_|3024,3025
_|3025,3026
_|3026,3027
04|3028,3030
:|3030,3031
55AM|3031,3035
BLOOD|3036,3041
Glucose|3042,3049
-|3049,3050
105|3050,3053
*|3053,3054
UreaN|3055,3060
-|3060,3061
5|3061,3062
*|3062,3063
Creat|3064,3069
-|3069,3070
0.4|3070,3073
Na|3074,3076
-|3076,3077
134|3077,3080
<EOL>|3081,3082
K|3082,3083
-|3083,3084
3.3|3084,3087
Cl|3088,3090
-|3090,3091
96|3091,3093
HCO3|3094,3098
-|3098,3099
30|3099,3101
AnGap|3102,3107
-|3107,3108
11|3108,3110
<EOL>|3110,3111
_|3111,3112
_|3112,3113
_|3113,3114
06|3115,3117
:|3117,3118
35AM|3118,3122
BLOOD|3123,3128
Glucose|3129,3136
-|3136,3137
101|3137,3140
*|3140,3141
UreaN|3142,3147
-|3147,3148
4|3148,3149
*|3149,3150
Creat|3151,3156
-|3156,3157
0.4|3157,3160
Na|3161,3163
-|3163,3164
132|3164,3167
*|3167,3168
<EOL>|3169,3170
K|3170,3171
-|3171,3172
3.6|3172,3175
Cl|3176,3178
-|3178,3179
94|3179,3181
*|3181,3182
HCO3|3183,3187
-|3187,3188
30|3188,3190
AnGap|3191,3196
-|3196,3197
12|3197,3199
<EOL>|3199,3200
_|3200,3201
_|3201,3202
_|3202,3203
04|3204,3206
:|3206,3207
24AM|3207,3211
BLOOD|3212,3217
Glucose|3218,3225
-|3225,3226
100|3226,3229
UreaN|3230,3235
-|3235,3236
3|3236,3237
*|3237,3238
Creat|3239,3244
-|3244,3245
0.4|3245,3248
Na|3249,3251
-|3251,3252
135|3252,3255
<EOL>|3256,3257
K|3257,3258
-|3258,3259
3.4|3259,3262
Cl|3263,3265
-|3265,3266
95|3266,3268
*|3268,3269
HCO3|3270,3274
-|3274,3275
30|3275,3277
AnGap|3278,3283
-|3283,3284
13|3284,3286
<EOL>|3286,3287
_|3287,3288
_|3288,3289
_|3289,3290
11|3291,3293
:|3293,3294
30AM|3294,3298
BLOOD|3299,3304
Glucose|3305,3312
-|3312,3313
141|3313,3316
*|3316,3317
UreaN|3318,3323
-|3323,3324
4|3324,3325
*|3325,3326
Creat|3327,3332
-|3332,3333
0.4|3333,3336
Na|3337,3339
-|3339,3340
138|3340,3343
<EOL>|3344,3345
K|3345,3346
-|3346,3347
3.6|3347,3350
Cl|3351,3353
-|3353,3354
98|3354,3356
HCO3|3357,3361
-|3361,3362
26|3362,3364
AnGap|3365,3370
-|3370,3371
18|3371,3373
<EOL>|3373,3374
_|3374,3375
_|3375,3376
_|3376,3377
04|3378,3380
:|3380,3381
50AM|3381,3385
BLOOD|3386,3391
ALT|3392,3395
-|3395,3396
45|3396,3398
*|3398,3399
AST|3400,3403
-|3403,3404
144|3404,3407
*|3407,3408
AlkPhos|3409,3416
-|3416,3417
275|3417,3420
*|3420,3421
<EOL>|3422,3423
TotBili|3423,3430
-|3430,3431
1|3431,3432
.|3432,3433
6|3433,3434
*|3434,3435
<EOL>|3435,3436
_|3436,3437
_|3437,3438
_|3438,3439
04|3440,3442
:|3442,3443
50AM|3443,3447
BLOOD|3448,3453
ALT|3454,3457
-|3457,3458
41|3458,3460
*|3460,3461
AST|3462,3465
-|3465,3466
158|3466,3469
*|3469,3470
LD|3471,3473
(|3473,3474
_|3474,3475
_|3475,3476
_|3476,3477
)|3477,3478
-|3478,3479
260|3479,3482
*|3482,3483
<EOL>|3484,3485
AlkPhos|3485,3492
-|3492,3493
277|3493,3496
*|3496,3497
TotBili|3498,3505
-|3505,3506
2|3506,3507
.|3507,3508
3|3508,3509
*|3509,3510
<EOL>|3510,3511
_|3511,3512
_|3512,3513
_|3513,3514
04|3515,3517
:|3517,3518
55AM|3518,3522
BLOOD|3523,3528
ALT|3529,3532
-|3532,3533
46|3533,3535
*|3535,3536
AST|3537,3540
-|3540,3541
187|3541,3544
*|3544,3545
AlkPhos|3546,3553
-|3553,3554
299|3554,3557
*|3557,3558
<EOL>|3559,3560
TotBili|3560,3567
-|3567,3568
2|3568,3569
.|3569,3570
1|3570,3571
*|3571,3572
<EOL>|3572,3573
_|3573,3574
_|3574,3575
_|3575,3576
06|3577,3579
:|3579,3580
35AM|3580,3584
BLOOD|3585,3590
ALT|3591,3594
-|3594,3595
46|3595,3597
*|3597,3598
AST|3599,3602
-|3602,3603
223|3603,3606
*|3606,3607
AlkPhos|3608,3615
-|3615,3616
297|3616,3619
*|3619,3620
<EOL>|3621,3622
TotBili|3622,3629
-|3629,3630
2|3630,3631
.|3631,3632
1|3632,3633
*|3633,3634
<EOL>|3634,3635
_|3635,3636
_|3636,3637
_|3637,3638
04|3639,3641
:|3641,3642
24AM|3642,3646
BLOOD|3647,3652
ALT|3653,3656
-|3656,3657
56|3657,3659
*|3659,3660
AST|3661,3664
-|3664,3665
335|3665,3668
*|3668,3669
LD|3670,3672
(|3672,3673
LDH|3673,3676
)|3676,3677
-|3677,3678
370|3678,3681
*|3681,3682
<EOL>|3683,3684
AlkPhos|3684,3691
-|3691,3692
313|3692,3695
*|3695,3696
TotBili|3697,3704
-|3704,3705
1|3705,3706
.|3706,3707
7|3707,3708
*|3708,3709
<EOL>|3709,3710
_|3710,3711
_|3711,3712
_|3712,3713
11|3714,3716
:|3716,3717
30AM|3717,3721
BLOOD|3722,3727
ALT|3728,3731
-|3731,3732
71|3732,3734
*|3734,3735
AST|3736,3739
-|3739,3740
401|3740,3743
*|3743,3744
LD|3745,3747
(|3747,3748
_|3748,3749
_|3749,3750
_|3750,3751
)|3751,3752
-|3752,3753
470|3753,3756
*|3756,3757
CK|3758,3760
(|3760,3761
CPK|3761,3764
)|3764,3765
-|3765,3766
87|3766,3768
<EOL>|3769,3770
AlkPhos|3770,3777
-|3777,3778
325|3778,3781
*|3781,3782
TotBili|3783,3790
-|3790,3791
1.5|3791,3794
<EOL>|3794,3795
_|3795,3796
_|3796,3797
_|3797,3798
04|3799,3801
:|3801,3802
24AM|3802,3806
BLOOD|3807,3812
Lipase|3813,3819
-|3819,3820
33|3820,3822
<EOL>|3822,3823
_|3823,3824
_|3824,3825
_|3825,3826
11|3827,3829
:|3829,3830
30AM|3830,3834
BLOOD|3835,3840
Lipase|3841,3847
-|3847,3848
40|3848,3850
GGT|3851,3854
-|3854,3855
2266|3855,3859
*|3859,3860
<EOL>|3860,3861
_|3861,3862
_|3862,3863
_|3863,3864
04|3865,3867
:|3867,3868
50AM|3868,3872
BLOOD|3873,3878
Calcium|3879,3886
-|3886,3887
7|3887,3888
.|3888,3889
5|3889,3890
*|3890,3891
Phos|3892,3896
-|3896,3897
2|3897,3898
.|3898,3899
6|3899,3900
*|3900,3901
Mg|3902,3904
-|3904,3905
1.7|3905,3908
<EOL>|3908,3909
_|3909,3910
_|3910,3911
_|3911,3912
04|3913,3915
:|3915,3916
50AM|3916,3920
BLOOD|3921,3926
Calcium|3927,3934
-|3934,3935
7|3935,3936
.|3936,3937
3|3937,3938
*|3938,3939
Phos|3940,3944
-|3944,3945
2|3945,3946
.|3946,3947
4|3947,3948
*|3948,3949
Mg|3950,3952
-|3952,3953
1.6|3953,3956
<EOL>|3956,3957
_|3957,3958
_|3958,3959
_|3959,3960
04|3961,3963
:|3963,3964
55AM|3964,3968
BLOOD|3969,3974
Albumin|3975,3982
-|3982,3983
2|3983,3984
.|3984,3985
7|3985,3986
*|3986,3987
Calcium|3988,3995
-|3995,3996
7|3996,3997
.|3997,3998
7|3998,3999
*|3999,4000
Phos|4001,4005
-|4005,4006
2|4006,4007
.|4007,4008
1|4008,4009
*|4009,4010
<EOL>|4011,4012
Mg|4012,4014
-|4014,4015
1.7|4015,4018
Iron|4019,4023
-|4023,4024
47|4024,4026
<EOL>|4026,4027
_|4027,4028
_|4028,4029
_|4029,4030
06|4031,4033
:|4033,4034
35AM|4034,4038
BLOOD|4039,4044
Calcium|4045,4052
-|4052,4053
7|4053,4054
.|4054,4055
4|4055,4056
*|4056,4057
Phos|4058,4062
-|4062,4063
2|4063,4064
.|4064,4065
6|4065,4066
*|4066,4067
Mg|4068,4070
-|4070,4071
1.9|4071,4074
<EOL>|4074,4075
_|4075,4076
_|4076,4077
_|4077,4078
04|4079,4081
:|4081,4082
24AM|4082,4086
BLOOD|4087,4092
Albumin|4093,4100
-|4100,4101
3|4101,4102
.|4102,4103
0|4103,4104
*|4104,4105
Calcium|4106,4113
-|4113,4114
7|4114,4115
.|4115,4116
1|4116,4117
*|4117,4118
Phos|4119,4123
-|4123,4124
3.3|4124,4127
<EOL>|4128,4129
Mg|4129,4131
-|4131,4132
1|4132,4133
.|4133,4134
5|4134,4135
*|4135,4136
Iron|4137,4141
-|4141,4142
65|4142,4144
<EOL>|4144,4145
_|4145,4146
_|4146,4147
_|4147,4148
11|4149,4151
:|4151,4152
30AM|4152,4156
BLOOD|4157,4162
Albumin|4163,4170
-|4170,4171
3|4171,4172
.|4172,4173
2|4173,4174
*|4174,4175
<EOL>|4175,4176
_|4176,4177
_|4177,4178
_|4178,4179
04|4180,4182
:|4182,4183
24AM|4183,4187
BLOOD|4188,4193
calTIBC|4194,4201
-|4201,4202
151|4202,4205
*|4205,4206
VitB12|4207,4213
-|4213,4214
1059|4214,4218
*|4218,4219
Folate|4220,4226
-|4226,4227
11.1|4227,4231
<EOL>|4232,4233
Ferritn|4233,4240
-|4240,4241
GREATER|4241,4248
TH|4249,4251
TRF|4252,4255
-|4255,4256
116|4256,4259
*|4259,4260
<EOL>|4260,4261
_|4261,4262
_|4262,4263
_|4263,4264
06|4265,4267
:|4267,4268
35AM|4268,4272
BLOOD|4273,4278
TSH|4279,4282
-|4282,4283
5|4283,4284
.|4284,4285
6|4285,4286
*|4286,4287
<EOL>|4287,4288
_|4288,4289
_|4289,4290
_|4290,4291
04|4292,4294
:|4294,4295
55AM|4295,4299
BLOOD|4300,4305
Free|4306,4310
T4|4311,4313
-|4313,4314
1.2|4314,4317
<EOL>|4317,4318
_|4318,4319
_|4319,4320
_|4320,4321
11|4322,4324
:|4324,4325
30AM|4325,4329
BLOOD|4330,4335
HBsAg|4336,4341
-|4341,4342
NEGATIVE|4342,4350
HBsAb|4351,4356
-|4356,4357
POSITIVE|4357,4365
<EOL>|4366,4367
HBcAb|4367,4372
-|4372,4373
NEGATIVE|4373,4381
HAV|4382,4385
Ab|4386,4388
-|4388,4389
POSITIVE|4389,4397
IgM|4398,4401
HAV|4402,4405
-|4405,4406
NEGATIVE|4406,4414
<EOL>|4414,4415
_|4415,4416
_|4416,4417
_|4417,4418
11|4419,4421
:|4421,4422
30AM|4422,4426
BLOOD|4427,4432
HCG|4433,4436
-|4436,4437
<|4437,4438
5|4438,4439
<EOL>|4439,4440
_|4440,4441
_|4441,4442
_|4442,4443
04|4444,4446
:|4446,4447
24AM|4447,4451
BLOOD|4452,4457
AMA|4458,4461
-|4461,4462
NEGATIVE|4462,4470
Smooth|4471,4477
-|4477,4478
NEGATIVE|4478,4486
<EOL>|4486,4487
_|4487,4488
_|4488,4489
_|4489,4490
04|4491,4493
:|4493,4494
24AM|4494,4498
BLOOD|4499,4504
_|4505,4506
_|4506,4507
_|4507,4508
<EOL>|4508,4509
_|4509,4510
_|4510,4511
_|4511,4512
04|4513,4515
:|4515,4516
24AM|4516,4520
BLOOD|4521,4526
HIV|4527,4530
Ab|4531,4533
-|4533,4534
NEGATIVE|4534,4542
<EOL>|4542,4543
_|4543,4544
_|4544,4545
_|4545,4546
11|4547,4549
:|4549,4550
30AM|4550,4554
BLOOD|4555,4560
ASA|4561,4564
-|4564,4565
NEG|4565,4568
_|4569,4570
_|4570,4571
_|4571,4572
Acetmnp|4573,4580
-|4580,4581
NEG|4581,4584
<EOL>|4585,4586
Bnzodzp|4586,4593
-|4593,4594
NEG|4594,4597
Barbitr|4598,4605
-|4605,4606
NEG|4606,4609
Tricycl|4610,4617
-|4617,4618
NEG|4618,4621
<EOL>|4621,4622
_|4622,4623
_|4623,4624
_|4624,4625
11|4626,4628
:|4628,4629
30AM|4629,4633
BLOOD|4634,4639
HoldBLu|4640,4647
-|4647,4648
HOLD|4648,4652
<EOL>|4652,4653
_|4653,4654
_|4654,4655
_|4655,4656
11|4657,4659
:|4659,4660
30AM|4660,4664
BLOOD|4665,4670
LtGrnHD|4671,4678
-|4678,4679
HOLD|4679,4683
<EOL>|4683,4684
_|4684,4685
_|4685,4686
_|4686,4687
11|4688,4690
:|4690,4691
30AM|4691,4695
BLOOD|4696,4701
HCV|4702,4705
Ab|4706,4708
-|4708,4709
NEGATIVE|4709,4717
<EOL>|4717,4718
_|4718,4719
_|4719,4720
_|4720,4721
11|4722,4724
:|4724,4725
49AM|4725,4729
BLOOD|4730,4735
Glucose|4736,4743
-|4743,4744
125|4744,4747
*|4747,4748
Lactate|4749,4756
-|4756,4757
2|4757,4758
.|4758,4759
3|4759,4760
*|4760,4761
<EOL>|4761,4762
_|4762,4763
_|4763,4764
_|4764,4765
04|4766,4768
:|4768,4769
55AM|4769,4773
BLOOD|4774,4779
CERULOPLASMIN|4780,4793
-|4793,4794
PND|4794,4797
<EOL>|4797,4798
_|4798,4799
_|4799,4800
_|4800,4801
04|4802,4804
:|4804,4805
55AM|4805,4809
BLOOD|4810,4815
ALPHA|4816,4821
-|4821,4822
1|4822,4823
-|4823,4824
ANTITRYPSIN|4824,4835
-|4835,4836
PND|4836,4839
<EOL>|4839,4840
<EOL>|4840,4841
Imaging|4841,4848
<EOL>|4848,4849
_|4849,4850
_|4850,4851
_|4851,4852
US|4853,4855
abd|4856,4859
/|4859,4860
pelvis|4860,4866
<EOL>|4866,4867
IMPRESSION|4867,4877
:|4877,4878
<EOL>|4879,4880
1.|4880,4882
Diffusely|4883,4892
echogenic|4893,4902
liver|4903,4908
,|4908,4909
suggestive|4910,4920
of|4921,4923
fatty|4924,4929
infiltration|4930,4942
.|4942,4943
<EOL>|4944,4945
Other|4945,4950
forms|4951,4956
of|4957,4959
liver|4960,4965
disease|4966,4973
and|4974,4977
more|4978,4982
advanced|4983,4991
liver|4992,4997
disease|4998,5005
<EOL>|5006,5007
including|5007,5016
fibrosis|5017,5025
and|5026,5029
cirrhosis|5030,5039
can|5040,5043
not|5043,5046
be|5047,5049
excluded|5050,5058
.|5058,5059
<EOL>|5060,5061
2.|5061,5063
Layering|5064,5072
sludge|5073,5079
within|5080,5086
the|5087,5090
gallbladder|5091,5102
,|5102,5103
with|5104,5108
mild|5109,5113
gallbladder|5114,5125
<EOL>|5126,5127
wall|5127,5131
<EOL>|5132,5133
thickening|5133,5143
,|5143,5144
which|5145,5150
may|5151,5154
relate|5155,5161
to|5162,5164
underlying|5165,5175
liver|5176,5181
disease|5182,5189
.|5189,5190
<EOL>|5192,5193
3.|5193,5195
Patent|5196,5202
portal|5203,5209
venous|5210,5216
system|5217,5223
.|5223,5224
<EOL>|5225,5226
4.|5226,5228
Moderate|5229,5237
ascites|5238,5245
.|5245,5246
<EOL>|5247,5248
The|5248,5251
study|5252,5257
and|5258,5261
the|5262,5265
report|5266,5272
were|5273,5277
reviewed|5278,5286
by|5287,5289
the|5290,5293
staff|5294,5299
radiologist|5300,5311
.|5311,5312
<EOL>|5313,5314
<EOL>|5314,5315
<EOL>|5315,5316
CT|5316,5318
abd|5319,5322
/|5322,5323
pelvis|5323,5329
_|5330,5331
_|5331,5332
_|5332,5333
<EOL>|5333,5334
IMPRESSION|5334,5344
:|5344,5345
<EOL>|5346,5347
1.|5347,5349
Large|5350,5355
volume|5356,5362
ascites|5363,5370
and|5371,5374
enlarged|5375,5383
edematous|5384,5393
liver|5394,5399
.|5399,5400
The|5401,5404
<EOL>|5405,5406
findings|5406,5414
are|5415,5418
<EOL>|5419,5420
suggestive|5420,5430
of|5431,5433
acute|5434,5439
hepatitis|5440,5449
.|5449,5450
<EOL>|5452,5453
2.|5453,5455
Small|5456,5461
bilateral|5462,5471
pleural|5472,5479
effusions|5480,5489
.|5489,5490
<EOL>|5490,5491
<EOL>|5491,5492
ECHO|5492,5496
_|5497,5498
_|5498,5499
_|5499,5500
:|5500,5501
<EOL>|5501,5502
The|5502,5505
left|5506,5510
atrium|5511,5517
and|5518,5521
right|5522,5527
atrium|5528,5534
are|5535,5538
normal|5539,5545
in|5546,5548
cavity|5549,5555
size|5556,5560
.|5560,5561
Left|5562,5566
<EOL>|5567,5568
ventricular|5568,5579
wall|5580,5584
thickness|5585,5594
,|5594,5595
cavity|5596,5602
size|5603,5607
and|5608,5611
regional|5612,5620
/|5620,5621
global|5621,5627
<EOL>|5628,5629
systolic|5629,5637
function|5638,5646
are|5647,5650
normal|5651,5657
(|5658,5659
LVEF|5659,5663
>|5664,5665
55|5665,5667
%|5667,5668
)|5668,5669
.|5669,5670
Transmitral|5671,5682
and|5683,5686
tissue|5687,5693
<EOL>|5694,5695
Doppler|5695,5702
imaging|5703,5710
suggests|5711,5719
normal|5720,5726
diastolic|5727,5736
function|5737,5745
,|5745,5746
and|5747,5750
a|5751,5752
normal|5753,5759
<EOL>|5760,5761
left|5761,5765
ventricular|5766,5777
filling|5778,5785
pressure|5786,5794
(|5795,5796
PCWP|5796,5800
<|5800,5801
12mmHg|5801,5807
)|5807,5808
.|5808,5809
There|5810,5815
is|5816,5818
no|5819,5821
<EOL>|5822,5823
ventricular|5823,5834
septal|5835,5841
defect|5842,5848
.|5848,5849
Right|5850,5855
ventricular|5856,5867
chamber|5868,5875
size|5876,5880
and|5881,5884
<EOL>|5885,5886
free|5886,5890
wall|5891,5895
motion|5896,5902
are|5903,5906
normal|5907,5913
.|5913,5914
The|5915,5918
diameters|5919,5928
of|5929,5931
aorta|5932,5937
at|5938,5940
the|5941,5944
<EOL>|5945,5946
sinus|5946,5951
,|5951,5952
ascending|5953,5962
and|5963,5966
arch|5967,5971
levels|5972,5978
are|5979,5982
normal|5983,5989
.|5989,5990
The|5991,5994
aortic|5995,6001
valve|6002,6007
<EOL>|6008,6009
leaflets|6009,6017
(|6018,6019
3|6019,6020
)|6020,6021
appear|6022,6028
structurally|6029,6041
normal|6042,6048
with|6049,6053
good|6054,6058
leaflet|6059,6066
<EOL>|6067,6068
excursion|6068,6077
and|6078,6081
no|6082,6084
aortic|6085,6091
regurgitation|6092,6105
.|6105,6106
The|6107,6110
mitral|6111,6117
valve|6118,6123
appears|6124,6131
<EOL>|6132,6133
structurally|6133,6145
normal|6146,6152
with|6153,6157
trivial|6158,6165
mitral|6166,6172
regurgitation|6173,6186
.|6186,6187
There|6188,6193
is|6194,6196
<EOL>|6197,6198
no|6198,6200
mitral|6201,6207
valve|6208,6213
prolapse|6214,6222
.|6222,6223
There|6224,6229
is|6230,6232
no|6233,6235
pericardial|6236,6247
effusion|6248,6256
.|6256,6257
<EOL>|6258,6259
<EOL>|6259,6260
IMPRESSION|6260,6270
:|6270,6271
Normal|6272,6278
global|6279,6285
and|6286,6289
regional|6290,6298
biventricular|6299,6312
systolic|6313,6321
<EOL>|6322,6323
function|6323,6331
.|6331,6332
No|6333,6335
diastolic|6336,6345
dysfunction|6346,6357
,|6357,6358
pulmonary|6359,6368
hypertension|6369,6381
or|6382,6384
<EOL>|6385,6386
pathologic|6386,6396
valvular|6397,6405
disease|6406,6413
seen|6414,6418
.|6418,6419
<EOL>|6419,6420
<EOL>|6421,6422
Brief|6422,6427
Hospital|6428,6436
Course|6437,6443
:|6443,6444
<EOL>|6444,6445
This|6445,6449
is|6450,6452
a|6453,6454
_|6455,6456
_|6456,6457
_|6457,6458
woman|6459,6464
with|6465,6469
history|6470,6477
of|6478,6480
EtOH|6481,6485
_|6486,6487
_|6487,6488
_|6488,6489
years|6490,6495
,|6495,6496
<EOL>|6497,6498
heavy|6498,6503
at|6504,6506
times|6507,6512
,|6512,6513
with|6514,6518
new|6519,6522
onset|6523,6528
liver|6529,6534
failure|6535,6542
and|6543,6546
ascites|6547,6554
.|6554,6555
<EOL>|6557,6558
<EOL>|6560,6561
#|6561,6562
ASCITES|6564,6571
/|6571,6572
LFTs|6572,6576
:|6576,6577
New|6579,6582
onset|6583,6588
ascites|6589,6596
with|6597,6601
SAAG|6602,6606
supportive|6607,6617
of|6618,6620
<EOL>|6621,6622
portal|6622,6628
hypertension|6629,6641
.|6641,6642
Likely|6644,6650
alcoholic|6651,6660
hepatitis|6661,6670
with|6671,6675
ascites|6676,6683
<EOL>|6684,6685
and|6685,6688
possibility|6689,6700
of|6701,6703
cirrhosis|6704,6713
.|6713,6714
Steroids|6716,6724
and|6725,6728
pentoxyphyline|6729,6743
were|6744,6748
<EOL>|6749,6750
deferred|6750,6758
given|6759,6764
her|6765,6768
low|6769,6772
discriminate|6773,6785
factor|6786,6792
.|6792,6793
In|6795,6797
terms|6798,6803
of|6804,6806
other|6807,6812
<EOL>|6813,6814
etiologies|6814,6824
of|6825,6827
liver|6828,6833
disease|6834,6841
,|6841,6842
iron|6843,6847
panel|6848,6853
was|6854,6857
not|6858,6861
consistent|6862,6872
with|6873,6877
<EOL>|6878,6879
hemochromatosis|6879,6894
,|6894,6895
and|6896,6899
_|6900,6901
_|6901,6902
_|6902,6903
,|6903,6904
AMA|6905,6908
,|6908,6909
_|6910,6911
_|6911,6912
_|6912,6913
were|6914,6918
negative|6919,6927
,|6927,6928
making|6929,6935
<EOL>|6936,6937
autoimmune|6937,6947
causes|6948,6954
unlikely.|6955,6964
Alpha|6966,6971
1|6972,6973
antitrypsin|6974,6985
and|6986,6989
<EOL>|6990,6991
ceruloplasmin|6991,7004
were|7005,7009
normal|7010,7016
.|7016,7017
Viral|7019,7024
studies|7025,7032
show|7033,7037
immunity|7038,7046
to|7047,7049
Hep|7050,7053
B|7054,7055
<EOL>|7056,7057
and|7057,7060
A.|7061,7063
HIV|7065,7068
was|7069,7072
negative|7073,7081
.|7081,7082
U|7084,7085
/|7085,7086
S|7086,7087
and|7088,7091
CT|7092,7094
abd|7095,7098
/|7098,7099
pelvis|7099,7105
were|7106,7110
not|7111,7114
<EOL>|7115,7116
suggestive|7116,7126
of|7127,7129
mass|7130,7134
or|7135,7137
obstructive|7138,7149
lesions|7150,7157
.|7157,7158
Patient|7160,7167
received|7168,7176
a|7177,7178
<EOL>|7179,7180
2.5|7180,7183
L|7183,7184
paracentesis|7185,7197
on|7198,7200
_|7201,7202
_|7202,7203
_|7203,7204
,|7204,7205
day|7206,7209
prior|7210,7215
to|7216,7218
discharge|7219,7228
.|7228,7229
Low|7231,7234
-|7234,7235
dose|7235,7239
<EOL>|7240,7241
spironolactone|7241,7255
was|7256,7259
started|7260,7267
.|7267,7268
Ms.|7270,7273
_|7274,7275
_|7275,7276
_|7276,7277
will|7278,7282
follow|7283,7289
-|7289,7290
up|7290,7292
with|7293,7297
<EOL>|7298,7299
Dr.|7299,7302
_|7303,7304
_|7304,7305
_|7305,7306
in|7307,7309
1|7310,7311
week|7312,7316
.|7316,7317
<EOL>|7317,7318
<EOL>|7320,7321
#|7321,7322
ALCOHOLISM|7324,7334
:|7334,7335
On|7337,7339
admission|7340,7349
,|7349,7350
alcohol|7351,7358
level|7359,7364
was|7365,7368
336|7369,7372
though|7373,7379
<EOL>|7380,7381
patient|7381,7388
was|7389,7392
clinically|7393,7403
sober|7404,7409
.|7409,7410
Patient|7412,7419
was|7420,7423
monitored|7424,7433
on|7434,7436
a|7437,7438
CIWA|7439,7443
<EOL>|7444,7445
scale|7445,7450
and|7451,7454
treated|7455,7462
with|7463,7467
MVI|7468,7471
,|7471,7472
thiamine|7473,7481
,|7481,7482
and|7483,7486
folate|7487,7493
.|7493,7494
She|7496,7499
was|7500,7503
seen|7504,7508
<EOL>|7509,7510
by|7510,7512
social|7513,7519
work|7520,7524
and|7525,7528
given|7529,7534
the|7535,7538
contact|7539,7546
information|7547,7558
for|7559,7562
rehab|7563,7568
<EOL>|7569,7570
facilities|7570,7580
.|7580,7581
Although|7583,7591
patient|7592,7599
was|7600,7603
encouraged|7604,7614
to|7615,7617
enter|7618,7623
_|7624,7625
_|7625,7626
_|7626,7627
<EOL>|7628,7629
rehab|7629,7634
,|7634,7635
she|7636,7639
refused|7640,7647
.|7647,7648
She|7650,7653
will|7654,7658
seek|7659,7663
outpatient|7664,7674
treatment|7675,7684
for|7685,7688
her|7689,7692
<EOL>|7693,7694
addiction|7694,7703
.|7703,7704
Ms.|7706,7709
_|7710,7711
_|7711,7712
_|7712,7713
was|7714,7717
warned|7718,7724
on|7725,7727
multiple|7728,7736
occasions|7737,7746
that|7747,7751
<EOL>|7752,7753
if|7753,7755
she|7756,7759
continues|7760,7769
to|7770,7772
drink|7773,7778
she|7779,7782
will|7783,7787
irreperably|7788,7799
destroy|7800,7807
her|7808,7811
liver|7812,7817
<EOL>|7818,7819
and|7819,7822
could|7823,7828
even|7829,7833
die|7834,7837
.|7837,7838
<EOL>|7838,7839
<EOL>|7839,7840
#|7840,7841
BACK|7843,7847
PAIN|7848,7852
:|7852,7853
Patient|7855,7862
was|7863,7866
started|7867,7874
on|7875,7877
a|7878,7879
lidocaine|7880,7889
patch|7890,7895
and|7896,7899
<EOL>|7900,7901
given|7901,7906
oxycodone|7907,7916
for|7917,7920
breakthrough|7921,7933
pain|7934,7938
while|7939,7944
in|7945,7947
the|7948,7951
hospital|7952,7960
.|7960,7961
<EOL>|7961,7962
<EOL>|7964,7965
#|7965,7966
LEUKOCYTOSIS|7968,7980
:|7980,7981
Likely|7983,7989
a|7990,7991
combination|7992,8003
of|8004,8006
alcoholic|8007,8016
hepatitis|8017,8026
<EOL>|8027,8028
and|8028,8031
UTI|8032,8035
;|8035,8036
patient|8037,8044
was|8045,8048
started|8049,8056
on|8057,8059
ciprofloxacin|8060,8073
.|8073,8074
Other|8076,8081
infectious|8082,8092
<EOL>|8093,8094
work|8094,8098
-|8098,8099
up|8099,8101
was|8102,8105
unrevealing|8106,8117
.|8117,8118
On|8120,8122
day|8123,8126
prior|8127,8132
to|8133,8135
discharge|8136,8145
,|8145,8146
patient|8147,8154
<EOL>|8155,8156
spiked|8156,8162
a|8163,8164
fever|8165,8170
to|8171,8173
101|8174,8177
and|8178,8181
was|8182,8185
pan|8186,8189
cultured|8190,8198
.|8198,8199
CXR|8201,8204
was|8205,8208
unrevealing|8209,8220
<EOL>|8221,8222
and|8222,8225
urine|8226,8231
was|8232,8235
negative|8236,8244
for|8245,8248
infection|8249,8258
after|8259,8264
the|8265,8268
Cipro|8269,8274
.|8274,8275
Ms|8277,8279
.|8279,8280
<EOL>|8281,8282
_|8282,8283
_|8283,8284
_|8284,8285
was|8286,8289
discharged|8290,8300
on|8301,8303
levofloxacin|8304,8316
for|8317,8320
a|8321,8322
5|8323,8324
day|8325,8328
course|8329,8335
.|8335,8336
<EOL>|8336,8337
<EOL>|8339,8340
#|8340,8341
MACROCYTIC|8343,8353
ANEMIA|8354,8360
:|8360,8361
Likely|8363,8369
from|8370,8374
folate|8375,8381
and|8382,8385
nutritional|8386,8397
<EOL>|8398,8399
deficiency|8399,8409
in|8410,8412
setting|8413,8420
of|8421,8423
alcoholism|8424,8434
.|8434,8435
Patient|8437,8444
was|8445,8448
started|8449,8456
on|8457,8459
MV|8460,8462
,|8462,8463
<EOL>|8464,8465
thiamine|8465,8473
,|8473,8474
and|8475,8478
folate|8479,8485
supplementation|8486,8501
.|8501,8502
HCT|8504,8507
was|8508,8511
monitored|8512,8521
<EOL>|8522,8523
throughout|8523,8533
admission|8534,8543
.|8543,8544
<EOL>|8544,8545
<EOL>|8545,8546
#|8546,8547
ANXIETY|8549,8556
:|8556,8557
Patient|8559,8566
with|8567,8571
marked|8572,8578
anxiety|8579,8586
.|8586,8587
She|8589,8592
would|8593,8598
likely|8599,8605
<EOL>|8606,8607
benefit|8607,8614
from|8615,8619
outpatient|8620,8630
therapy|8631,8638
and|8639,8642
/|8642,8643
or|8643,8645
SSRI|8646,8650
treatment|8651,8660
.|8660,8661
<EOL>|8661,8662
<EOL>|8662,8663
#|8663,8664
SINUS|8666,8671
TACHYCARDIA|8672,8683
:|8683,8684
Likely|8686,8692
in|8693,8695
context|8696,8703
of|8704,8706
decompensated|8707,8720
liver|8721,8726
<EOL>|8727,8728
disease|8728,8735
.|8735,8736
ECHO|8738,8742
was|8743,8746
within|8747,8753
normal|8754,8760
limits|8761,8767
.|8767,8768
Patient|8770,8777
was|8778,8781
monitred|8782,8790
<EOL>|8791,8792
on|8792,8794
telemetry|8795,8804
throughout|8805,8815
hospitalization|8816,8831
.|8831,8832
<EOL>|8832,8833
<EOL>|8833,8834
#|8834,8835
CONSTIPATION|8837,8849
:|8849,8850
Patient|8852,8859
was|8860,8863
maintained|8864,8874
on|8875,8877
senna|8878,8883
and|8884,8887
colace|8888,8894
.|8894,8895
<EOL>|8895,8896
<EOL>|8897,8898
Medications|8898,8909
on|8910,8912
Admission|8913,8922
:|8922,8923
<EOL>|8923,8924
None|8924,8928
.|8928,8929
<EOL>|8929,8930
<EOL>|8931,8932
Discharge|8932,8941
Medications|8942,8953
:|8953,8954
<EOL>|8954,8955
1.|8955,8957
Multivitamin|8958,8970
Tablet|8975,8981
Sig|8982,8985
:|8985,8986
One|8987,8990
(|8991,8992
1|8992,8993
)|8993,8994
Tablet|8995,9001
PO|9002,9004
DAILY|9005,9010
(|9011,9012
Daily|9012,9017
)|9017,9018
.|9018,9019
<EOL>|9019,9020
Disp|9020,9024
:|9024,9025
*|9025,9026
30|9026,9028
Tablet|9029,9035
(|9035,9036
s|9036,9037
)|9037,9038
*|9038,9039
Refills|9040,9047
:|9047,9048
*|9048,9049
2|9049,9050
*|9050,9051
<EOL>|9051,9052
2.|9052,9054
Folic|9055,9060
Acid|9061,9065
1|9066,9067
mg|9068,9070
Tablet|9071,9077
Sig|9078,9081
:|9081,9082
One|9083,9086
(|9087,9088
1|9088,9089
)|9089,9090
Tablet|9091,9097
PO|9098,9100
DAILY|9101,9106
(|9107,9108
Daily|9108,9113
)|9113,9114
.|9114,9115
<EOL>|9115,9116
Disp|9116,9120
:|9120,9121
*|9121,9122
30|9122,9124
Tablet|9125,9131
(|9131,9132
s|9132,9133
)|9133,9134
*|9134,9135
Refills|9136,9143
:|9143,9144
*|9144,9145
2|9145,9146
*|9146,9147
<EOL>|9147,9148
3.|9148,9150
Thiamine|9151,9159
HCl|9160,9163
100|9164,9167
mg|9168,9170
Tablet|9171,9177
Sig|9178,9181
:|9181,9182
One|9183,9186
(|9187,9188
1|9188,9189
)|9189,9190
Tablet|9191,9197
PO|9198,9200
DAILY|9201,9206
<EOL>|9207,9208
(|9208,9209
Daily|9209,9214
)|9214,9215
.|9215,9216
<EOL>|9216,9217
Disp|9217,9221
:|9221,9222
*|9222,9223
30|9223,9225
Tablet|9226,9232
(|9232,9233
s|9233,9234
)|9234,9235
*|9235,9236
Refills|9237,9244
:|9244,9245
*|9245,9246
2|9246,9247
*|9247,9248
<EOL>|9248,9249
4.|9249,9251
Lidocaine|9252,9261
5|9262,9263
%|9264,9265
(|9265,9266
700|9266,9269
mg|9270,9272
/|9272,9273
patch|9273,9278
)|9278,9279
Adhesive|9280,9288
Patch|9289,9294
,|9294,9295
Medicated|9296,9305
Sig|9306,9309
:|9309,9310
<EOL>|9311,9312
One|9312,9315
(|9316,9317
1|9317,9318
)|9318,9319
Adhesive|9320,9328
Patch|9329,9334
,|9334,9335
Medicated|9336,9345
Topical|9346,9353
DAILY|9354,9359
(|9360,9361
Daily|9361,9366
)|9366,9367
:|9367,9368
Apply|9369,9374
<EOL>|9375,9376
to|9376,9378
affected|9379,9387
area|9388,9392
once|9393,9397
daily|9398,9403
as|9404,9406
directed|9407,9415
.|9415,9416
<EOL>|9416,9417
Disp|9417,9421
:|9421,9422
*|9422,9423
30|9423,9425
Adhesive|9426,9434
Patch|9435,9440
,|9440,9441
Medicated|9442,9451
(|9451,9452
s|9452,9453
)|9453,9454
*|9454,9455
Refills|9456,9463
:|9463,9464
*|9464,9465
2|9465,9466
*|9466,9467
<EOL>|9467,9468
5.|9468,9470
Nicotine|9471,9479
14|9480,9482
mg|9483,9485
/|9485,9486
24|9486,9488
hr|9489,9491
Patch|9492,9497
24|9498,9500
hr|9501,9503
Sig|9504,9507
:|9507,9508
One|9509,9512
(|9513,9514
1|9514,9515
)|9515,9516
Patch|9517,9522
24|9523,9525
hr|9526,9528
<EOL>|9529,9530
Transdermal|9530,9541
DAILY|9542,9547
(|9548,9549
Daily|9549,9554
)|9554,9555
:|9555,9556
Apply|9557,9562
once|9563,9567
daily|9568,9573
as|9574,9576
directed|9577,9585
.|9585,9586
<EOL>|9586,9587
Disp|9587,9591
:|9591,9592
*|9592,9593
30|9593,9595
Patch|9596,9601
24|9602,9604
hr|9605,9607
(|9607,9608
s|9608,9609
)|9609,9610
*|9610,9611
Refills|9612,9619
:|9619,9620
*|9620,9621
2|9621,9622
*|9622,9623
<EOL>|9623,9624
6.|9624,9626
Spironolactone|9627,9641
25|9642,9644
mg|9645,9647
Tablet|9648,9654
Sig|9655,9658
:|9658,9659
One|9660,9663
(|9664,9665
1|9665,9666
)|9666,9667
Tablet|9668,9674
PO|9675,9677
once|9678,9682
a|9683,9684
<EOL>|9685,9686
day|9686,9689
.|9689,9690
<EOL>|9690,9691
Disp|9691,9695
:|9695,9696
*|9696,9697
30|9697,9699
Tablet|9700,9706
(|9706,9707
s|9707,9708
)|9708,9709
*|9709,9710
Refills|9711,9718
:|9718,9719
*|9719,9720
0|9720,9721
*|9721,9722
<EOL>|9722,9723
7.|9723,9725
Levofloxacin|9726,9738
750|9739,9742
mg|9743,9745
Tablet|9746,9752
Sig|9753,9756
:|9756,9757
One|9758,9761
(|9762,9763
1|9763,9764
)|9764,9765
Tablet|9766,9772
PO|9773,9775
once|9776,9780
a|9781,9782
day|9783,9786
<EOL>|9787,9788
for|9788,9791
5|9792,9793
days|9794,9798
.|9798,9799
<EOL>|9799,9800
Disp|9800,9804
:|9804,9805
*|9805,9806
5|9806,9807
Tablet|9808,9814
(|9814,9815
s|9815,9816
)|9816,9817
*|9817,9818
Refills|9819,9826
:|9826,9827
*|9827,9828
0|9828,9829
*|9829,9830
<EOL>|9830,9831
8.|9831,9833
Outpatient|9834,9844
Lab|9845,9848
Work|9849,9853
<EOL>|9853,9854
Please|9854,9860
draw|9861,9865
blood|9866,9871
samples|9872,9879
for|9880,9883
CBC|9884,9887
with|9888,9892
differential|9893,9905
,|9905,9906
AST|9907,9910
/|9910,9911
ALT|9911,9914
,|9914,9915
<EOL>|9916,9917
total|9917,9922
bilirubin|9923,9932
,|9932,9933
alkaline|9934,9942
phosphatase|9943,9954
,|9954,9955
albumin|9956,9963
,|9963,9964
LDH|9965,9968
,|9968,9969
INR|9970,9973
/|9973,9974
PTT|9974,9977
,|9977,9978
<EOL>|9979,9980
and|9980,9983
chem10|9984,9990
(|9991,9992
K|9992,9993
,|9993,9994
Na|9995,9997
,|9997,9998
P|9999,10000
,|10000,10001
Ca|10002,10004
,|10004,10005
Mg|10006,10008
,|10008,10009
Cl|10010,10012
,|10012,10013
CO3|10014,10017
,|10017,10018
renal|10019,10024
function|10025,10033
,|10033,10034
glucose|10035,10042
)|10042,10043
<EOL>|10043,10044
<EOL>|10045,10046
Discharge|10046,10055
Disposition|10056,10067
:|10067,10068
<EOL>|10068,10069
Home|10069,10073
<EOL>|10073,10074
<EOL>|10075,10076
Discharge|10076,10085
Diagnosis|10086,10095
:|10095,10096
<EOL>|10096,10097
Primary|10097,10104
Diagnoses|10105,10114
:|10114,10115
<EOL>|10115,10116
-|10116,10117
alcohol|10118,10125
-|10125,10126
related|10126,10133
hepatitis|10134,10143
<EOL>|10143,10144
-|10144,10145
ascites|10146,10153
<EOL>|10153,10154
<EOL>|10155,10156
Discharge|10156,10165
Condition|10166,10175
:|10175,10176
<EOL>|10176,10177
Mental|10177,10183
Status|10184,10190
:|10190,10191
Clear|10192,10197
and|10198,10201
coherent|10202,10210
.|10210,10211
<EOL>|10211,10212
Level|10212,10217
of|10218,10220
Consciousness|10221,10234
:|10234,10235
Alert|10236,10241
and|10242,10245
interactive|10246,10257
.|10257,10258
<EOL>|10258,10259
Activity|10259,10267
Status|10268,10274
:|10274,10275
Ambulatory|10276,10286
-|10287,10288
Independent|10289,10300
.|10300,10301
<EOL>|10301,10302
<EOL>|10303,10304
Discharge|10304,10313
Instructions|10314,10326
:|10326,10327
<EOL>|10327,10328
You|10328,10331
were|10332,10336
admitted|10337,10345
to|10346,10348
the|10349,10352
hospital|10353,10361
for|10362,10365
inflammation|10366,10378
in|10379,10381
the|10382,10385
liver|10386,10391
<EOL>|10392,10393
that|10393,10397
was|10398,10401
likely|10402,10408
due|10409,10412
to|10413,10415
alcohol|10416,10423
consumption|10424,10435
.|10435,10436
You|10437,10440
were|10441,10445
treated|10446,10453
<EOL>|10454,10455
supportively|10455,10467
with|10468,10472
nutrition|10473,10482
and|10483,10486
also|10487,10491
treated|10492,10499
with|10500,10504
medicines|10505,10514
for|10515,10518
<EOL>|10519,10520
alcohol|10520,10527
withdrawal|10528,10538
.|10538,10539
We|10540,10542
monitored|10543,10552
your|10553,10557
liver|10558,10563
function|10564,10572
daily|10573,10578
with|10579,10583
<EOL>|10584,10585
blood|10585,10590
tests|10591,10596
and|10597,10600
found|10601,10606
that|10607,10611
the|10612,10615
liver|10616,10621
function|10622,10630
was|10631,10634
improving|10635,10644
at|10645,10647
<EOL>|10648,10649
time|10649,10653
of|10654,10656
discharge|10657,10666
.|10666,10667
During|10668,10674
this|10675,10679
admission|10680,10689
,|10689,10690
you|10691,10694
were|10695,10699
also|10700,10704
found|10705,10710
to|10711,10713
<EOL>|10714,10715
have|10715,10719
a|10720,10721
urinary|10722,10729
tract|10730,10735
infection|10736,10745
and|10746,10749
a|10750,10751
pneumonia|10752,10761
.|10761,10762
Please|10763,10769
complete|10770,10778
<EOL>|10779,10780
five|10780,10784
more|10785,10789
days|10790,10794
of|10795,10797
antibiotics|10798,10809
(|10810,10811
levofloxacin|10811,10823
)|10823,10824
to|10825,10827
treat|10828,10833
these|10834,10839
<EOL>|10840,10841
infections|10841,10851
.|10851,10852
<EOL>|10852,10853
<EOL>|10853,10854
We|10854,10856
have|10857,10861
started|10862,10869
a|10870,10871
new|10872,10875
medicine|10876,10884
that|10885,10889
will|10890,10894
help|10895,10899
remove|10900,10906
fluid|10907,10912
from|10913,10917
<EOL>|10918,10919
the|10919,10922
abdomen|10923,10930
and|10931,10934
legs|10935,10939
.|10939,10940
This|10941,10945
medicine|10946,10954
is|10955,10957
called|10958,10964
spironolactone|10965,10979
.|10979,10980
<EOL>|10981,10982
Since|10982,10987
this|10988,10992
medicine|10993,11001
can|11002,11005
raise|11006,11011
potassium|11012,11021
levels|11022,11028
in|11029,11031
the|11032,11035
blood|11036,11041
,|11041,11042
we|11043,11045
<EOL>|11046,11047
would|11047,11052
like|11053,11057
you|11058,11061
to|11062,11064
have|11065,11069
your|11070,11074
blood|11075,11080
-|11080,11081
work|11081,11085
checked|11086,11093
next|11094,11098
_|11099,11100
_|11100,11101
_|11101,11102
.|11102,11103
<EOL>|11104,11105
You|11105,11108
can|11109,11112
have|11113,11117
this|11118,11122
done|11123,11127
at|11128,11130
_|11131,11132
_|11132,11133
_|11133,11134
in|11135,11137
the|11138,11141
Atrium|11142,11148
Suite|11149,11154
on|11155,11157
the|11158,11161
first|11162,11167
floor|11168,11173
or|11174,11176
on|11177,11179
<EOL>|11180,11181
the|11181,11184
sixth|11185,11190
floor|11191,11196
,|11196,11197
anytime|11198,11205
from|11206,11210
8am|11211,11214
to|11215,11217
6pm|11218,11221
.|11221,11222
<EOL>|11222,11223
<EOL>|11223,11224
We|11224,11226
made|11227,11231
the|11232,11235
following|11236,11245
changes|11246,11253
to|11254,11256
your|11257,11261
medicines|11262,11271
:|11271,11272
<EOL>|11272,11273
-|11273,11274
we|11275,11277
ADDED|11278,11283
folate|11284,11290
,|11290,11291
thiamine|11292,11300
,|11300,11301
and|11302,11305
multivitamin|11306,11318
(|11319,11320
for|11320,11323
general|11324,11331
<EOL>|11332,11333
nutrition|11333,11342
)|11342,11343
<EOL>|11343,11344
-|11344,11345
we|11346,11348
ADDED|11349,11354
lidocaine|11355,11364
patch|11365,11370
(|11371,11372
for|11372,11375
pain|11376,11380
)|11380,11381
<EOL>|11381,11382
-|11382,11383
we|11384,11386
ADDED|11387,11392
nicotine|11393,11401
patch|11402,11407
<EOL>|11407,11408
-|11408,11409
we|11410,11412
ADDED|11413,11418
levofloxacin|11419,11431
(|11432,11433
antibiotic|11433,11443
for|11444,11447
pneumonia|11448,11457
)|11457,11458
<EOL>|11458,11459
-|11459,11460
we|11461,11463
ADDED|11464,11469
spironolactone|11470,11484
(|11485,11486
diuretic|11486,11494
to|11495,11497
prevent|11498,11505
fluid|11506,11511
<EOL>|11512,11513
accumulation|11513,11525
)|11525,11526
<EOL>|11526,11527
There|11527,11532
were|11533,11537
no|11538,11540
other|11541,11546
changes|11547,11554
to|11555,11557
your|11558,11562
medicines|11563,11572
.|11572,11573
<EOL>|11573,11574
<EOL>|11574,11575
Please|11575,11581
see|11582,11585
the|11586,11589
appointments|11590,11602
that|11603,11607
we|11608,11610
have|11611,11615
scheduled|11616,11625
for|11626,11629
you|11630,11633
<EOL>|11634,11635
below|11635,11640
.|11640,11641
<EOL>|11641,11642
<EOL>|11643,11644
Followup|11644,11652
Instructions|11653,11665
:|11665,11666
<EOL>|11666,11667
_|11667,11668
_|11668,11669
_|11669,11670
<EOL>|11670,11671

