 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Procedure|Health Care Activity|SIMPLE_SEGMENT|49,58|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|49,63|false|false|false|C2598112||Admission Date
Finding|Body Substance|SIMPLE_SEGMENT|83,92|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|83,92|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|83,92|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|83,92|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|83,97|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|115,120|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|115,120|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|115,120|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|139,142|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|139,142|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|139,142|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|139,142|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|139,142|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|150,157|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|150,157|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|159,167|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|SIMPLE_SEGMENT|170,179|false|false|false|C1717415||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|170,179|false|false|false|C0020517|Hypersensitivity|Allergies
Attribute|Clinical Attribute|SIMPLE_SEGMENT|191,200|false|false|false|C1717415||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|191,200|false|false|false|C0020517|Hypersensitivity|Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|203,225|true|false|false|C0041755|Adverse reaction to drug|Adverse Drug Reactions
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|211,215|false|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|Drug
Finding|Finding|SIMPLE_SEGMENT|211,215|false|false|false|C0740721|Drug problem|Drug
Finding|Pathologic Function|SIMPLE_SEGMENT|211,225|true|false|false|C0041755|Adverse reaction to drug|Drug Reactions
Finding|Functional Concept|SIMPLE_SEGMENT|228,237|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|SIMPLE_SEGMENT|246,261|false|false|false|C0277786|Chief complaint (finding)|Chief Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|252,261|false|false|false|C3864418||Complaint
Finding|Finding|SIMPLE_SEGMENT|252,261|false|false|false|C5441521|Complaint (finding)|Complaint
Finding|Functional Concept|SIMPLE_SEGMENT|263,269|false|false|false|C0234621|Visual|Visual
Finding|Sign or Symptom|SIMPLE_SEGMENT|263,284|false|false|false|C0233763|Hallucinations, Visual|Visual hallucinations
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|270,284|false|false|false|C0018524|Hallucinations|hallucinations
Finding|Classification|SIMPLE_SEGMENT|287,292|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|SIMPLE_SEGMENT|293,301|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|293,301|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|305,323|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|314,323|false|false|false|C0945766||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|314,323|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|314,323|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|314,323|false|false|false|C0184661|Interventional procedure|Procedure
Finding|Conceptual Entity|SIMPLE_SEGMENT|332,339|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|332,339|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|332,339|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|332,342|false|false|false|C0262926|Medical History|History of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|332,358|false|false|false|C0488508||History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|332,358|false|false|false|C0262512|History of present illness (finding)|History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|343,350|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Idea or Concept|SIMPLE_SEGMENT|343,350|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Finding|SIMPLE_SEGMENT|343,358|false|false|false|C4264312|Present illness|Present Illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|351,358|false|false|false|C0221423|Illness (finding)|Illness
Finding|Finding|SIMPLE_SEGMENT|364,368|false|false|false|C1706180|Male Gender|male
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|378,385|false|false|false|C0012634|Disease|disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|387,399|false|false|false|C0242339|Dyslipidemias|dyslipidemia
Finding|Conceptual Entity|SIMPLE_SEGMENT|407,414|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|407,414|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|407,414|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|407,417|false|false|false|C0262926|Medical History|history of
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|418,426|false|false|false|C0033572;C4266527|Prostate;Structure of prostate (body structure)|prostate
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|418,426|false|false|false|C0033575;C0154009;C0154088;C0496923|Benign neoplasm of prostate;Carcinoma in situ of prostate;Neoplasm of uncertain or unknown behavior of prostate;Prostatic Diseases|prostate
Disorder|Neoplastic Process|SIMPLE_SEGMENT|418,426|false|false|false|C0033575;C0154009;C0154088;C0496923|Benign neoplasm of prostate;Carcinoma in situ of prostate;Neoplasm of uncertain or unknown behavior of prostate;Prostatic Diseases|prostate
Disorder|Neoplastic Process|SIMPLE_SEGMENT|418,433|false|false|false|C0376358;C0600139|Malignant neoplasm of prostate;Prostate carcinoma|prostate cancer
Disorder|Neoplastic Process|SIMPLE_SEGMENT|427,433|false|false|false|C0006826|Malignant Neoplasms|cancer
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|439,452|false|false|false|C0033573|Prostatectomy|prostatectomy
Finding|Finding|SIMPLE_SEGMENT|514,518|false|false|false|C0016928|Gait|gait
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|520,525|false|false|false|C0000921|Accidental Falls|falls
Finding|Finding|SIMPLE_SEGMENT|520,525|false|false|false|C0085639|Falls|falls
Finding|Functional Concept|SIMPLE_SEGMENT|531,537|false|false|false|C0234621|Visual|visual
Finding|Sign or Symptom|SIMPLE_SEGMENT|531,552|false|false|false|C0233763|Hallucinations, Visual|visual hallucinations
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|538,552|false|false|false|C0018524|Hallucinations|hallucinations
Finding|Conceptual Entity|SIMPLE_SEGMENT|570,577|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|570,577|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|570,577|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Intellectual Product|SIMPLE_SEGMENT|592,597|false|false|false|C0684240|Charts (publication)|chart
Procedure|Health Care Activity|SIMPLE_SEGMENT|592,604|false|false|false|C0541653|Chart evaluation by healthcare professional|chart review
Finding|Idea or Concept|SIMPLE_SEGMENT|598,604|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Finding|Intellectual Product|SIMPLE_SEGMENT|598,604|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Finding|Body Substance|SIMPLE_SEGMENT|612,619|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|612,619|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|612,619|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Finding|SIMPLE_SEGMENT|664,668|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|664,668|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|664,668|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Functional Concept|SIMPLE_SEGMENT|690,696|false|false|false|C0234621|Visual|visual
Finding|Sign or Symptom|SIMPLE_SEGMENT|690,711|false|false|false|C0233763|Hallucinations, Visual|visual hallucinations
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|697,711|false|false|false|C0018524|Hallucinations|hallucinations
Finding|Idea or Concept|SIMPLE_SEGMENT|716,725|false|false|false|C1546960|Patient Outcome - Worsening|worsening
Finding|Finding|SIMPLE_SEGMENT|726,730|false|false|false|C0016928|Gait|gait
Finding|Functional Concept|SIMPLE_SEGMENT|731,739|false|false|false|C0677542|Frozen behavior|freezing
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|731,739|false|false|false|C0016701|Freezing|freezing
Finding|Finding|SIMPLE_SEGMENT|749,753|false|false|false|C0016928|Gait|gait
Finding|Functional Concept|SIMPLE_SEGMENT|754,762|false|false|false|C0677542|Frozen behavior|freezing
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|754,762|false|false|false|C0016701|Freezing|freezing
Drug|Organic Chemical|SIMPLE_SEGMENT|768,775|false|false|false|C0721754|Mirapex|mirapex
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|768,775|false|false|false|C0721754|Mirapex|mirapex
Finding|Intellectual Product|SIMPLE_SEGMENT|808,812|false|false|false|C1561540|Transaction counts and value totals - week|week
Finding|Idea or Concept|SIMPLE_SEGMENT|818,822|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Finding|Intellectual Product|SIMPLE_SEGMENT|818,822|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|878,886|false|false|false|C0013227|Pharmaceutical Preparations|medicine
Finding|Functional Concept|SIMPLE_SEGMENT|925,931|false|false|false|C0234621|Visual|visual
Finding|Sign or Symptom|SIMPLE_SEGMENT|925,946|false|false|false|C0233763|Hallucinations, Visual|visual hallucinations
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|932,946|false|false|false|C0018524|Hallucinations|hallucinations
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|951,960|false|false|false|C0009676|Confusion|confusion
Finding|Finding|SIMPLE_SEGMENT|951,960|false|false|false|C0683369|Clouded consciousness|confusion
Finding|Functional Concept|SIMPLE_SEGMENT|1046,1053|false|false|false|C0392747|Changing|changes
Drug|Organic Chemical|SIMPLE_SEGMENT|1061,1068|false|false|false|C0721754|Mirapex|Mirapex
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1061,1068|false|false|false|C0721754|Mirapex|Mirapex
Finding|Body Substance|SIMPLE_SEGMENT|1074,1081|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1074,1081|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1074,1081|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|SIMPLE_SEGMENT|1103,1114|false|false|false|C0205329|Progressive|progressive
Finding|Finding|SIMPLE_SEGMENT|1115,1119|false|false|false|C0016928|Gait|gait
Finding|Sign or Symptom|SIMPLE_SEGMENT|1120,1129|false|false|false|C0427008|Stiffness|stiffness
Finding|Finding|SIMPLE_SEGMENT|1144,1154|false|false|false|C1299586|Has difficulty doing (qualifier value)|difficulty
Finding|Finding|SIMPLE_SEGMENT|1186,1196|false|false|false|C1299586|Has difficulty doing (qualifier value)|difficulty
Finding|Finding|SIMPLE_SEGMENT|1186,1201|false|false|false|C0332218|Difficult (qualifier value)|difficulty with
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1256,1268|false|false|false|C0021167|Incontinence|incontinence
Procedure|Health Care Activity|SIMPLE_SEGMENT|1296,1306|false|false|false|C0557055|Reassuring (procedure)|reassuring
Finding|Idea or Concept|SIMPLE_SEGMENT|1317,1320|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|1317,1320|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Idea or Concept|SIMPLE_SEGMENT|1324,1336|false|false|false|C0449450|Presentation|presentation
Finding|Idea or Concept|SIMPLE_SEGMENT|1344,1352|false|false|false|C1547192|Organization unit type - Hospital|hospital
Finding|Body Substance|SIMPLE_SEGMENT|1358,1365|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1358,1365|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1358,1365|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Mental Process|SIMPLE_SEGMENT|1375,1385|false|false|false|C0237607;C0596545|Experience;Experience (Practice)|experience
Finding|Functional Concept|SIMPLE_SEGMENT|1386,1392|false|false|false|C0234621|Visual|visual
Finding|Sign or Symptom|SIMPLE_SEGMENT|1386,1407|false|false|false|C0233763|Hallucinations, Visual|visual hallucinations
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|1393,1407|false|false|false|C0018524|Hallucinations|hallucinations
Finding|Functional Concept|SIMPLE_SEGMENT|1413,1418|false|false|false|C1513492|motor movement|motor
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1419,1424|false|false|false|C2936910|Cross syndrome|cross
Finding|Conceptual Entity|SIMPLE_SEGMENT|1419,1424|false|false|false|C2828360|Traverse|cross
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1425,1429|false|false|false|C1315098||race
Finding|Gene or Genome|SIMPLE_SEGMENT|1425,1429|false|false|false|C1412374;C1706779|AMACR gene;AMACR wt Allele|race
Procedure|Molecular Biology Research Technique|SIMPLE_SEGMENT|1425,1429|false|false|false|C5551096|Rapid Amplification of cDNA Ends|race
Finding|Finding|SIMPLE_SEGMENT|1467,1473|false|false|false|C1561668|History of fall|a fall
Finding|Finding|SIMPLE_SEGMENT|1469,1473|false|false|false|C0085639|Falls|fall
Finding|Finding|SIMPLE_SEGMENT|1533,1539|false|false|false|C1299582|Unable|unable
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|1559,1564|false|false|false|C3714591|Floor (anatomic)|floor
Finding|Finding|SIMPLE_SEGMENT|1570,1574|false|false|false|C0085639|Falls|fall
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1606,1610|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1606,1610|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1606,1610|false|false|false|C0362076|Problems with head|head
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1606,1610|false|false|false|C0876917|Procedure on head|head
Event|Occupational Activity|SIMPLE_SEGMENT|1611,1617|true|false|false|C0038452|Strikes, Employee|strike
Finding|Body Substance|SIMPLE_SEGMENT|1627,1634|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1627,1634|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1627,1634|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Finding|SIMPLE_SEGMENT|1647,1651|false|false|false|C0016928|Gait|gait
Finding|Finding|SIMPLE_SEGMENT|1727,1733|false|false|false|C1299582|Unable|unable
Finding|Finding|SIMPLE_SEGMENT|1737,1745|false|false|false|C4036205|Ambulate|ambulate
Finding|Finding|SIMPLE_SEGMENT|1753,1756|false|false|false|C5939094|Own|own
Finding|Body Substance|SIMPLE_SEGMENT|1762,1769|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1762,1769|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1762,1769|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1820,1832|false|false|false|C0449450|Presentation|presentation
Finding|Body Substance|SIMPLE_SEGMENT|1861,1868|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1861,1868|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1861,1868|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Finding|SIMPLE_SEGMENT|1873,1881|false|false|false|C0277797|Apyrexial|afebrile
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1883,1886|false|false|false|C0751781|Dentatorubral-Pallidoluysian Atrophy|HRs
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1883,1886|false|false|false|C1568891|HGS protein, human|HRs
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1883,1886|false|false|false|C1568891|HGS protein, human|HRs
Finding|Gene or Genome|SIMPLE_SEGMENT|1883,1886|false|false|false|C1366514;C1415473;C1419996;C1708271;C5575450;C5780798|ATN1 wt Allele;HARS1 gene;HARS1 wt Allele;HGS gene;HGS wt Allele;SRSF5 gene|HRs
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1910,1914|false|false|false|C2317096|Saturation of Peripheral Oxygen|SpO2
Finding|Functional Concept|SIMPLE_SEGMENT|1927,1931|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|1927,1931|false|false|false|C0582103|Medical Examination|exam
Finding|Sign or Symptom|SIMPLE_SEGMENT|1953,1964|false|false|false|C0151564|Cogwheel Rigidity|cogwheeling
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1974,1985|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Finding|Finding|SIMPLE_SEGMENT|1990,1998|false|false|false|C0392756|Reduced|decrease
Finding|Idea or Concept|SIMPLE_SEGMENT|2003,2011|false|false|false|C0808080|Strength (attribute)|strength
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2013,2017|false|false|false|C0587081|Laboratory test finding|Labs
Finding|Classification|SIMPLE_SEGMENT|2040,2048|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|2040,2048|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2040,2048|false|false|false|C5237010|Expression Negative|negative
Finding|Body Substance|SIMPLE_SEGMENT|2049,2054|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Functional Concept|SIMPLE_SEGMENT|2049,2054|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Intellectual Product|SIMPLE_SEGMENT|2049,2054|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|2059,2064|false|false|false|C5575602|Cell Culture Serum|serum
Finding|Body Substance|SIMPLE_SEGMENT|2059,2064|false|false|false|C0229671;C1546774;C1550100|Serum;Serum specimen|serum
Finding|Intellectual Product|SIMPLE_SEGMENT|2059,2064|false|false|false|C0229671;C1546774;C1550100|Serum;Serum specimen|serum
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2065,2068|false|false|false|C3177193|TOX protein, human|tox
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2065,2068|false|false|false|C3177193|TOX protein, human|tox
Finding|Gene or Genome|SIMPLE_SEGMENT|2065,2068|false|false|false|C1847320|TOX gene|tox
Finding|Intellectual Product|SIMPLE_SEGMENT|2103,2106|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2103,2106|false|false|false|C1623258|Electrocardiography|EKG
Finding|Functional Concept|SIMPLE_SEGMENT|2107,2114|false|false|false|C0392747|Changing|changes
Finding|Classification|SIMPLE_SEGMENT|2117,2125|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|2117,2125|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2117,2125|false|false|false|C5237010|Expression Negative|negative
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2126,2134|false|false|false|C0041199|Troponin|troponin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2126,2134|false|false|false|C0041199|Troponin|troponin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2126,2134|false|false|false|C0523952|Troponin measurement|troponin
Anatomy|Cell Component|SIMPLE_SEGMENT|2162,2165|false|false|false|C2263086|Nuclear cap binding complex location|CBC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2162,2165|false|false|false|C0009555|Complete Blood Count|CBC
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2168,2173|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|SIMPLE_SEGMENT|2168,2173|false|false|false|C0741025|Chest problem|Chest
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|2174,2178|false|false|false|C0043309|Roentgen Rays|Xray
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2174,2178|false|false|false|C0043299|Diagnostic radiologic examination|Xray
Finding|Intellectual Product|SIMPLE_SEGMENT|2189,2194|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2195,2202|false|false|false|C1184743|bony process|process
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2195,2202|false|false|false|C1951340|Process Pharmacologic Substance|process
Finding|Functional Concept|SIMPLE_SEGMENT|2195,2202|false|false|false|C4521054|Process (qualifier value)|process
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|2195,2202|false|false|false|C1522240|Process|process
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2207,2210|false|false|false|C5849006|CTH protein, human|CTH
Drug|Enzyme|SIMPLE_SEGMENT|2207,2210|false|false|false|C5849006|CTH protein, human|CTH
Finding|Gene or Genome|SIMPLE_SEGMENT|2207,2210|false|false|false|C1413792;C1538070|CTH gene;VSIG2 gene|CTH
Procedure|Health Care Activity|SIMPLE_SEGMENT|2215,2225|false|false|false|C0557055|Reassuring (procedure)|reassuring
Procedure|Health Care Activity|SIMPLE_SEGMENT|2273,2282|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2286,2294|false|false|false|C0013227|Pharmaceutical Preparations|medicine
Finding|Functional Concept|SIMPLE_SEGMENT|2299,2306|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|SIMPLE_SEGMENT|2299,2306|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|SIMPLE_SEGMENT|2299,2306|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Body Substance|SIMPLE_SEGMENT|2334,2341|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|2334,2341|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|2334,2341|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|2344,2348|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|2344,2348|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|2344,2348|false|false|false|C1553498|home health encounter|home
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2349,2360|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2349,2360|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|SIMPLE_SEGMENT|2349,2360|false|false|false|C4284232|Medications|medications
Finding|Cell Function|SIMPLE_SEGMENT|2382,2391|false|false|false|C0311400;C1524026|Metabolic;Metabolic Process, Cellular|metabolic
Finding|Functional Concept|SIMPLE_SEGMENT|2382,2391|false|false|false|C0311400;C1524026|Metabolic;Metabolic Process, Cellular|metabolic
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2382,2391|false|false|false|C4263342|Multisection metabolic|metabolic
Finding|Body Substance|SIMPLE_SEGMENT|2404,2411|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|2404,2411|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|2404,2411|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|2426,2430|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|2426,2430|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|2426,2430|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|2431,2442|false|false|false|C0074710|pramipexole|pramipexole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2431,2442|false|false|false|C0074710|pramipexole|pramipexole
Drug|Organic Chemical|SIMPLE_SEGMENT|2447,2458|false|false|false|C0085542|pravastatin|pravastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2447,2458|false|false|false|C0085542|pravastatin|pravastatin
Event|Activity|SIMPLE_SEGMENT|2489,2496|false|false|false|C1706079||arrival
Finding|Functional Concept|SIMPLE_SEGMENT|2489,2496|false|false|false|C1555577|arrival - ActRelationshipType|arrival
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|2504,2509|false|false|false|C3714591|Floor (anatomic)|floor
Finding|Body Substance|SIMPLE_SEGMENT|2515,2522|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|2515,2522|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|2515,2522|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Finding|SIMPLE_SEGMENT|2526,2537|false|false|false|C5546696|Feeling comfortable|comfortable
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2541,2544|false|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Finding|Intellectual Product|SIMPLE_SEGMENT|2541,2544|false|false|false|C2346952|Bachelor of Education|bed
Finding|Classification|SIMPLE_SEGMENT|2572,2578|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|2572,2578|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|2572,2578|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|2572,2578|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Event|Activity|SIMPLE_SEGMENT|2585,2594|false|false|false|C0021822|Interview|interview
Finding|Intellectual Product|SIMPLE_SEGMENT|2585,2594|false|false|false|C0935630|Published Interview|interview
Finding|Idea or Concept|SIMPLE_SEGMENT|2624,2632|false|false|false|C1547192|Organization unit type - Hospital|hospital
Finding|Intellectual Product|SIMPLE_SEGMENT|2663,2667|true|false|false|C4724437|SURE Test|sure
Finding|Conceptual Entity|SIMPLE_SEGMENT|2713,2718|false|false|true|C1518904|Party|party
Finding|Functional Concept|SIMPLE_SEGMENT|2739,2744|false|false|true|C1513492|motor movement|motor
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2745,2750|false|false|false|C2936910|Cross syndrome|cross
Finding|Conceptual Entity|SIMPLE_SEGMENT|2745,2750|false|false|false|C2828360|Traverse|cross
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2751,2755|false|false|false|C1315098||race
Finding|Gene or Genome|SIMPLE_SEGMENT|2751,2755|false|false|false|C1412374;C1706779|AMACR gene;AMACR wt Allele|race
Procedure|Molecular Biology Research Technique|SIMPLE_SEGMENT|2751,2755|false|false|false|C5551096|Rapid Amplification of cDNA Ends|race
Finding|Finding|SIMPLE_SEGMENT|2800,2804|false|false|true|C0085639|Falls|fall
Finding|Finding|SIMPLE_SEGMENT|2838,2844|false|false|true|C1561668|History of fall|a fall
Finding|Finding|SIMPLE_SEGMENT|2840,2844|false|false|true|C0085639|Falls|fall
Finding|Sign or Symptom|SIMPLE_SEGMENT|2874,2880|false|false|false|C0015967|Fever|fevers
Finding|Sign or Symptom|SIMPLE_SEGMENT|2882,2888|false|false|false|C0085593|Chills|chills
Drug|Organic Chemical|SIMPLE_SEGMENT|2890,2895|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2890,2895|false|false|false|C3815497|Cough (guaifenesin)|cough
Finding|Sign or Symptom|SIMPLE_SEGMENT|2890,2895|false|false|false|C0010200|Coughing|cough
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2897,2902|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|2897,2902|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2897,2907|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|2897,2907|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2903,2907|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|2903,2907|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|2903,2907|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|2903,2918|false|false|false|C0000737|Abdominal Pain|pain, abdominal
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2909,2918|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|SIMPLE_SEGMENT|2909,2923|false|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2919,2923|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|2919,2923|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|2919,2923|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2925,2931|false|false|false|C4255480||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|2925,2931|false|false|false|C0027497|Nausea|nausea
Finding|Finding|SIMPLE_SEGMENT|2933,2941|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|SIMPLE_SEGMENT|2933,2941|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|SIMPLE_SEGMENT|2946,2953|false|false|false|C0013428|Dysuria|dysuria
Finding|Idea or Concept|SIMPLE_SEGMENT|2957,2963|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|REVIEW
Finding|Intellectual Product|SIMPLE_SEGMENT|2957,2963|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|REVIEW
Finding|Functional Concept|SIMPLE_SEGMENT|2957,2966|false|false|false|C0699752|Review of|REVIEW OF
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2957,2974|false|false|false|C0488564;C0488565||REVIEW OF SYSTEMS
Procedure|Health Care Activity|SIMPLE_SEGMENT|2957,2974|false|false|false|C0489633|Review of systems (procedure)|REVIEW OF SYSTEMS
Finding|Functional Concept|SIMPLE_SEGMENT|2967,2974|false|false|false|C0449913|System|SYSTEMS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2999,3002|false|false|false|C0268529|Proline dehydrogenase deficiency|HPI
Finding|Finding|SIMPLE_SEGMENT|2999,3002|false|false|false|C0262512;C1323983|History of present illness (finding);allene oxide synthase activity|HPI
Finding|Molecular Function|SIMPLE_SEGMENT|2999,3002|false|false|false|C0262512;C1323983|History of present illness (finding);allene oxide synthase activity|HPI
Finding|Idea or Concept|SIMPLE_SEGMENT|3024,3030|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Finding|Intellectual Product|SIMPLE_SEGMENT|3024,3030|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Finding|Functional Concept|SIMPLE_SEGMENT|3024,3033|false|false|false|C0699752|Review of|review of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3024,3041|false|false|false|C0488564;C0488565||review of systems
Procedure|Health Care Activity|SIMPLE_SEGMENT|3024,3041|false|false|false|C0489633|Review of systems (procedure)|review of systems
Finding|Functional Concept|SIMPLE_SEGMENT|3034,3041|false|false|false|C0449913|System|systems
Finding|Functional Concept|SIMPLE_SEGMENT|3060,3066|false|false|false|C0439801|Limited (extensiveness)|limits
Finding|Finding|SIMPLE_SEGMENT|3071,3091|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Finding|Functional Concept|SIMPLE_SEGMENT|3076,3083|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|3076,3083|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|3076,3083|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|3076,3083|false|false|false|C0199168|Medical service|Medical
Finding|Finding|SIMPLE_SEGMENT|3076,3091|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|3084,3091|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|3084,3091|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|3084,3091|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3097,3104|false|false|false|C0012634|Disease|disease
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|3109,3113|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|Body
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3109,3113|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|Body
Finding|Intellectual Product|SIMPLE_SEGMENT|3109,3113|false|false|false|C1551342|Document Body|Body
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|3114,3122|false|false|false|C0011265;C0497327|Dementia;Presenile dementia|Dementia
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3124,3136|false|false|false|C0242339|Dyslipidemias|dyslipidemia
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3138,3146|false|false|false|C0033572;C4266527|Prostate;Structure of prostate (body structure)|prostate
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3138,3146|false|false|false|C0033575;C0154009;C0154088;C0496923|Benign neoplasm of prostate;Carcinoma in situ of prostate;Neoplasm of uncertain or unknown behavior of prostate;Prostatic Diseases|prostate
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3138,3146|false|false|false|C0033575;C0154009;C0154088;C0496923|Benign neoplasm of prostate;Carcinoma in situ of prostate;Neoplasm of uncertain or unknown behavior of prostate;Prostatic Diseases|prostate
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3138,3153|false|false|false|C0376358;C0600139|Malignant neoplasm of prostate;Prostate carcinoma|prostate cancer
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3147,3153|false|false|false|C0006826|Malignant Neoplasms|cancer
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3159,3172|false|false|false|C0033573|Prostatectomy|prostatectomy
Finding|Functional Concept|SIMPLE_SEGMENT|3176,3182|false|false|false|C0728831|Social|Social
Finding|Finding|SIMPLE_SEGMENT|3176,3190|false|false|false|C0424945;C3714536|Social History;Social and personal history|Social History
Finding|Conceptual Entity|SIMPLE_SEGMENT|3183,3190|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|3183,3190|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|3183,3190|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Classification|SIMPLE_SEGMENT|3196,3202|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|SIMPLE_SEGMENT|3196,3202|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|SIMPLE_SEGMENT|3196,3202|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|SIMPLE_SEGMENT|3196,3202|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Finding|SIMPLE_SEGMENT|3196,3210|false|false|false|C0241889|Family Medical History|Family History
Finding|Conceptual Entity|SIMPLE_SEGMENT|3203,3210|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|3203,3210|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|3203,3210|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Idea or Concept|SIMPLE_SEGMENT|3216,3222|false|false|false|C1546508|Relationship - Mother|mother
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3231,3234|false|false|false|C1114365||age
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3231,3234|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|SIMPLE_SEGMENT|3231,3234|false|false|false|C0162574|Glycation End Products, Advanced|age
Finding|Finding|SIMPLE_SEGMENT|3243,3250|false|false|false|C0231337|Senility|old age
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3247,3250|false|false|false|C1114365||age
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3247,3250|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|SIMPLE_SEGMENT|3247,3250|false|false|false|C0162574|Glycation End Products, Advanced|age
Finding|Conceptual Entity|SIMPLE_SEGMENT|3257,3263|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|father
Finding|Idea or Concept|SIMPLE_SEGMENT|3257,3263|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|father
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3272,3280|false|false|false|C0033572;C4266527|Prostate;Structure of prostate (body structure)|prostate
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3272,3280|false|false|false|C0033575;C0154009;C0154088;C0496923|Benign neoplasm of prostate;Carcinoma in situ of prostate;Neoplasm of uncertain or unknown behavior of prostate;Prostatic Diseases|prostate
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3272,3280|false|false|false|C0033575;C0154009;C0154088;C0496923|Benign neoplasm of prostate;Carcinoma in situ of prostate;Neoplasm of uncertain or unknown behavior of prostate;Prostatic Diseases|prostate
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3272,3287|false|false|false|C0376358;C0600139|Malignant neoplasm of prostate;Prostate carcinoma|prostate cancer
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3281,3287|false|false|false|C0006826|Malignant Neoplasms|cancer
Finding|Conceptual Entity|SIMPLE_SEGMENT|3314,3320|false|false|false|C1546515;C1704647|Relationship - Sister;Sister - courtesy title|sister
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3322,3325|false|false|false|C1114365||age
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3322,3325|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|SIMPLE_SEGMENT|3322,3325|false|false|false|C0162574|Glycation End Products, Advanced|age
Finding|Conceptual Entity|SIMPLE_SEGMENT|3344,3350|false|false|false|C1546515;C1704647|Relationship - Sister;Sister - courtesy title|sister
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3352,3355|false|false|false|C1114365||age
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3352,3355|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|SIMPLE_SEGMENT|3352,3355|false|false|false|C0162574|Glycation End Products, Advanced|age
Finding|Conceptual Entity|SIMPLE_SEGMENT|3380,3387|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|brother
Finding|Idea or Concept|SIMPLE_SEGMENT|3380,3387|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|brother
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3389,3392|false|false|false|C1114365||age
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3389,3392|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|SIMPLE_SEGMENT|3389,3392|false|false|false|C0162574|Glycation End Products, Advanced|age
Finding|Classification|SIMPLE_SEGMENT|3442,3448|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|3442,3448|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|3442,3448|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|3442,3448|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|3449,3456|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|3449,3456|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|3449,3456|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|3449,3459|false|false|false|C0262926|Medical History|history of
Finding|Sign or Symptom|SIMPLE_SEGMENT|3471,3478|false|false|false|C0221423|Illness (finding)|illness
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|3482,3490|false|false|false|C0011265;C0497327|Dementia;Presenile dementia|dementia
Finding|Classification|SIMPLE_SEGMENT|3505,3511|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|3505,3511|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|3505,3511|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|3505,3511|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|3512,3519|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|3512,3519|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|3512,3519|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|3512,3522|false|false|false|C0262926|Medical History|history of
Finding|Mental Process|SIMPLE_SEGMENT|3542,3548|false|false|false|C0229992|Psyche structure|mental
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|3542,3558|false|false|false|C0004936|Mental disorders|mental disorders
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3549,3558|false|false|false|C0012634|Disease|disorders
Finding|Mental Process|SIMPLE_SEGMENT|3567,3575|false|false|false|C0023185|Learning|learning
Procedure|Educational Activity|SIMPLE_SEGMENT|3567,3575|false|false|false|C0013621|Knowledge acquisition|learning
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3576,3586|false|false|false|C5240435||disability
Finding|Finding|SIMPLE_SEGMENT|3576,3586|false|false|false|C0231170|Disability|disability
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|3590,3594|false|false|false|C1263846|Attention deficit hyperactivity disorder|ADHD
Finding|Classification|SIMPLE_SEGMENT|3609,3615|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|3609,3615|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|3609,3615|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|3609,3615|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Finding|SIMPLE_SEGMENT|3609,3623|true|false|false|C0241889|Family Medical History|family history
Finding|Finding|SIMPLE_SEGMENT|3609,3626|true|false|false|C0241889|Family Medical History|family history of
Finding|Conceptual Entity|SIMPLE_SEGMENT|3616,3623|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|3616,3623|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|3616,3623|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|3616,3626|true|false|false|C0262926|Medical History|history of
Finding|Finding|SIMPLE_SEGMENT|3627,3638|true|false|false|C0205487;C1548428|Psychiatric;Referral type - Psychiatric|psychiatric
Finding|Functional Concept|SIMPLE_SEGMENT|3627,3638|true|false|false|C0205487;C1548428|Psychiatric;Referral type - Psychiatric|psychiatric
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3627,3638|true|false|false|C3526598|Psychiatric service|psychiatric
Finding|Idea or Concept|SIMPLE_SEGMENT|3639,3647|false|false|false|C1546466|Problems - What subject filter|problems
Finding|Finding|SIMPLE_SEGMENT|3651,3659|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|3651,3659|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|3651,3659|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|3651,3664|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|3651,3664|false|false|false|C0031809|Physical Examination|Physical Exam
Finding|Functional Concept|SIMPLE_SEGMENT|3660,3664|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|3660,3664|false|false|false|C0582103|Medical Examination|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|3666,3675|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Finding|Finding|SIMPLE_SEGMENT|3676,3684|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|SIMPLE_SEGMENT|3676,3684|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|3676,3684|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|SIMPLE_SEGMENT|3676,3689|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAM
Procedure|Health Care Activity|SIMPLE_SEGMENT|3676,3689|false|false|false|C0031809|Physical Examination|PHYSICAL EXAM
Finding|Functional Concept|SIMPLE_SEGMENT|3685,3689|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|SIMPLE_SEGMENT|3685,3689|false|false|false|C0582103|Medical Examination|EXAM
Finding|Gene or Genome|SIMPLE_SEGMENT|3736,3739|false|false|false|C1412647|ATP5F1A gene|OMR
Finding|Classification|SIMPLE_SEGMENT|3741,3748|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|3741,3748|false|false|false|C3812897|General medical service|GENERAL
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3750,3755|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|3750,3755|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3750,3755|false|false|false|C0718338|Alert brand of caffeine|Alert
Finding|Finding|SIMPLE_SEGMENT|3750,3755|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|3750,3755|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|3750,3755|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|3760,3771|false|false|false|C1704675|Interaction|interactive
Finding|Finding|SIMPLE_SEGMENT|3773,3793|false|false|false|C2051415|patient appears in no acute distress (physical finding)|In no acute distress
Finding|Intellectual Product|SIMPLE_SEGMENT|3779,3784|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Finding|SIMPLE_SEGMENT|3785,3793|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|SIMPLE_SEGMENT|3785,3793|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3795,3800|false|false|false|C1512338|HEENT|HEENT
Finding|Finding|SIMPLE_SEGMENT|3802,3807|false|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3815,3821|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3815,3821|false|false|false|C0036412|Scleral Diseases|Sclera
Procedure|Health Care Activity|SIMPLE_SEGMENT|3815,3821|false|false|false|C2228481|examination of sclera|Sclera
Finding|Finding|SIMPLE_SEGMENT|3822,3831|false|false|false|C0205180|Anicteric|anicteric
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3844,3853|true|false|false|C1272883|Injection|injection
Finding|Functional Concept|SIMPLE_SEGMENT|3844,3853|true|false|false|C1828121|Injection Route of Administration|injection
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3844,3853|true|false|false|C0021485;C1533685|Injection of therapeutic agent;Injection procedure|injection
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3855,3858|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3855,3858|false|false|false|C0026987|Myelofibrosis|MMM
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3860,3864|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|SIMPLE_SEGMENT|3860,3864|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|SIMPLE_SEGMENT|3860,3864|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3869,3877|false|false|false|C0027530|Neck|cervical
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3869,3893|true|false|false|C0235592|Cervical lymphadenopathy|cervical lymphadenopathy
Finding|Finding|SIMPLE_SEGMENT|3869,3893|true|false|false|C4551446|Swollen lymph nodes in the neck|cervical lymphadenopathy
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3878,3893|true|false|false|C0497156|Lymphadenopathy|lymphadenopathy
Finding|Sign or Symptom|SIMPLE_SEGMENT|3878,3893|true|false|false|C4282165|Swollen Lymph Node|lymphadenopathy
Finding|Finding|SIMPLE_SEGMENT|3898,3901|true|false|false|C0425687|Jugular venous engorgement|JVD
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3903,3910|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|SIMPLE_SEGMENT|3903,3910|false|false|false|C1314974|Cardiac attachment|CARDIAC
Finding|Finding|SIMPLE_SEGMENT|3920,3926|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|SIMPLE_SEGMENT|3920,3926|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Event|Activity|SIMPLE_SEGMENT|3935,3939|false|false|false|C0871208|Rating (action)|rate
Finding|Idea or Concept|SIMPLE_SEGMENT|3935,3939|false|false|false|C1549480|Amount type - Rate|rate
Finding|Finding|SIMPLE_SEGMENT|3963,3970|false|false|false|C0018808|Heart murmur|murmurs
Finding|Finding|SIMPLE_SEGMENT|3971,3975|false|false|false|C0232267|Pericardial friction rub|rubs
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3985,3990|false|false|false|C0024109|Lung|LUNGS
Finding|Idea or Concept|SIMPLE_SEGMENT|3992,3997|false|false|false|C1550016|Remote control command - Clear|Clear
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4001,4013|false|false|false|C0004339|Auscultation|auscultation
Finding|Sign or Symptom|SIMPLE_SEGMENT|4030,4037|true|false|false|C0043144|Wheezing|wheezes
Finding|Finding|SIMPLE_SEGMENT|4039,4046|true|false|false|C0035508|Rhonchi|rhonchi
Finding|Finding|SIMPLE_SEGMENT|4050,4055|false|false|false|C0034642;C0240859|Basilar Rales;Rales|rales
Finding|Finding|SIMPLE_SEGMENT|4060,4069|true|false|false|C0442805;C5236002|Increase;Increased (finding)|increased
Finding|Functional Concept|SIMPLE_SEGMENT|4060,4069|true|false|false|C0442805;C5236002|Increase;Increased (finding)|increased
Finding|Sign or Symptom|SIMPLE_SEGMENT|4060,4087|true|false|false|C0859927|Increased work of breathing|increased work of breathing
Event|Occupational Activity|SIMPLE_SEGMENT|4070,4074|true|false|false|C0043227|Work|work
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|4070,4087|true|false|false|C0043229|Work of Breathing|work of breathing
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4078,4087|false|false|false|C5885990||breathing
Finding|Finding|SIMPLE_SEGMENT|4078,4087|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|SIMPLE_SEGMENT|4078,4087|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|SIMPLE_SEGMENT|4078,4087|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|SIMPLE_SEGMENT|4078,4087|false|false|false|C1160636|respiratory system process|breathing
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4098,4101|false|false|false|C0001365;C0038454|Acute ill-defined cerebrovascular disease;Cerebrovascular accident|CVA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4098,4101|false|false|false|C5779650|Cyclophosphamide/Doxorubicin/Vincristine|CVA
Finding|Sign or Symptom|SIMPLE_SEGMENT|4098,4112|true|false|false|C0235634|Renal angle tenderness|CVA tenderness
Finding|Mental Process|SIMPLE_SEGMENT|4102,4112|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|SIMPLE_SEGMENT|4102,4112|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4114,4121|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4114,4121|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Finding|Finding|SIMPLE_SEGMENT|4114,4121|false|false|false|C0941288|Abdomen problem|ABDOMEN
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4130,4136|false|false|false|C0021853|Intestines|bowels
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|4137,4143|false|false|false|C0037709||sounds
Finding|Finding|SIMPLE_SEGMENT|4149,4158|false|false|false|C0700124|Dilated|distended
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4174,4178|false|false|false|C4318566|Deep Resection Margin|deep
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4179,4188|false|false|false|C0030247|Palpation|palpation
Finding|Finding|SIMPLE_SEGMENT|4215,4227|true|false|false|C4054315|Organomegaly|organomegaly
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4229,4240|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|4245,4253|true|false|false|C0149651|Clubbing|clubbing
Finding|Sign or Symptom|SIMPLE_SEGMENT|4255,4263|true|false|false|C0010520|Cyanosis|cyanosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4268,4273|true|false|false|C1717255||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|4268,4273|true|false|false|C0013604|Edema|edema
Drug|Food|SIMPLE_SEGMENT|4275,4281|false|false|false|C5890763||Pulses
Finding|Physiologic Function|SIMPLE_SEGMENT|4275,4281|false|false|false|C0391850|Physiologic pulse|Pulses
Procedure|Health Care Activity|SIMPLE_SEGMENT|4275,4281|false|false|false|C0034107|Pulse taking|Pulses
Finding|Conceptual Entity|SIMPLE_SEGMENT|4285,4291|false|false|false|C0442038;C0920847|Circumpennate;Radial|Radial
Anatomy|Body System|SIMPLE_SEGMENT|4309,4313|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4309,4313|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4309,4313|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Finding|Body Substance|SIMPLE_SEGMENT|4309,4313|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|SIMPLE_SEGMENT|4309,4313|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Finding|SIMPLE_SEGMENT|4315,4319|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|4315,4319|false|false|false|C0687712|warming process|Warm
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|4321,4324|false|false|false|C1855179|CATARACT, ANTERIOR POLAR|Cap
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4321,4324|false|false|false|C0006935|capsule (pharmacologic)|Cap
Finding|Gene or Genome|SIMPLE_SEGMENT|4321,4324|false|false|false|C1416891;C1418551;C1419093;C1422073;C1422760;C2985259;C4522312|BRD4 gene;BRD4 wt Allele;CAP1 gene;HACD1 gene;LNPEP gene;SERPINB6 gene;SORBS1 gene|Cap
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4321,4324|false|false|false|C0278651;C0280547;C1879916|CAP Regimen;cisplatin/cyclophosphamide/doxorubicin protocol;cyclophosphamide/doxorubicin/prednisone protocol|Cap
Finding|Idea or Concept|SIMPLE_SEGMENT|4325,4331|false|false|false|C0807726|refill|refill
Finding|Sign or Symptom|SIMPLE_SEGMENT|4340,4346|true|false|false|C0015230;C5779628|Exanthema;Skin rash|rashes
Finding|Gene or Genome|SIMPLE_SEGMENT|4366,4369|false|false|false|C1539110|CNDP2 gene|CN2
Finding|Finding|SIMPLE_SEGMENT|4373,4379|false|false|false|C1554187|Gender Status - Intact|intact
Finding|Finding|SIMPLE_SEGMENT|4398,4412|false|false|false|C0026826|Muscle Hypertonia|Increased tone
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4416,4419|false|false|false|C0227192|Inferior esophageal sphincter structure|LEs
Finding|Classification|SIMPLE_SEGMENT|4416,4419|false|false|false|C0023595|Lewis Blood-Group System|LEs
Finding|Idea or Concept|SIMPLE_SEGMENT|4425,4433|false|false|false|C0808080|Strength (attribute)|strength
Finding|Finding|SIMPLE_SEGMENT|4450,4459|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|4450,4459|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|SIMPLE_SEGMENT|4450,4459|false|false|false|C2229507|sensory exam|sensation
Finding|Body Substance|SIMPLE_SEGMENT|4462,4471|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|4462,4471|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|4462,4471|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|4462,4471|false|false|false|C0030685|Patient Discharge|DISCHARGE
Finding|Finding|SIMPLE_SEGMENT|4472,4480|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|SIMPLE_SEGMENT|4472,4480|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|4472,4480|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|SIMPLE_SEGMENT|4472,4485|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAM
Procedure|Health Care Activity|SIMPLE_SEGMENT|4472,4485|false|false|false|C0031809|Physical Examination|PHYSICAL EXAM
Finding|Functional Concept|SIMPLE_SEGMENT|4481,4485|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|SIMPLE_SEGMENT|4481,4485|false|false|false|C0582103|Medical Examination|EXAM
Finding|Idea or Concept|SIMPLE_SEGMENT|4515,4519|false|false|false|C1511726|Data|Data
Finding|Gene or Genome|SIMPLE_SEGMENT|4550,4554|false|false|false|C1823816|C1orf210 gene|Temp
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4550,4554|false|false|false|C0279848|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Temp
Finding|Finding|SIMPLE_SEGMENT|4657,4665|false|false|false|C1314680;C1705822;C2053584|Transfer Technique;delivery (history)|delivery
Finding|Functional Concept|SIMPLE_SEGMENT|4657,4665|false|false|false|C1314680;C1705822;C2053584|Transfer Technique;delivery (history)|delivery
Finding|Organism Function|SIMPLE_SEGMENT|4657,4665|false|false|false|C1314680;C1705822;C2053584|Transfer Technique;delivery (history)|delivery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4657,4665|false|false|false|C0011209|Obstetric Delivery|delivery
Finding|Classification|SIMPLE_SEGMENT|4673,4680|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|4673,4680|false|false|false|C3812897|General medical service|GENERAL
Finding|Finding|SIMPLE_SEGMENT|4682,4702|false|false|false|C2051415|patient appears in no acute distress (physical finding)|In no acute distress
Finding|Intellectual Product|SIMPLE_SEGMENT|4688,4693|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Finding|SIMPLE_SEGMENT|4694,4702|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|SIMPLE_SEGMENT|4694,4702|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4726,4733|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|SIMPLE_SEGMENT|4726,4733|false|false|false|C1314974|Cardiac attachment|CARDIAC
Finding|Finding|SIMPLE_SEGMENT|4743,4749|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|SIMPLE_SEGMENT|4743,4749|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Event|Activity|SIMPLE_SEGMENT|4758,4762|false|false|false|C0871208|Rating (action)|rate
Finding|Idea or Concept|SIMPLE_SEGMENT|4758,4762|false|false|false|C1549480|Amount type - Rate|rate
Finding|Finding|SIMPLE_SEGMENT|4786,4793|false|false|false|C0018808|Heart murmur|murmurs
Finding|Finding|SIMPLE_SEGMENT|4794,4798|false|false|false|C0232267|Pericardial friction rub|rubs
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4808,4813|false|false|false|C0024109|Lung|LUNGS
Finding|Idea or Concept|SIMPLE_SEGMENT|4815,4820|false|false|false|C1550016|Remote control command - Clear|Clear
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4824,4836|false|false|false|C0004339|Auscultation|auscultation
Finding|Sign or Symptom|SIMPLE_SEGMENT|4853,4860|true|false|false|C0043144|Wheezing|wheezes
Finding|Finding|SIMPLE_SEGMENT|4862,4869|true|false|false|C0035508|Rhonchi|rhonchi
Finding|Finding|SIMPLE_SEGMENT|4873,4878|false|false|false|C0034642;C0240859|Basilar Rales;Rales|rales
Finding|Finding|SIMPLE_SEGMENT|4883,4892|true|false|false|C0442805;C5236002|Increase;Increased (finding)|increased
Finding|Functional Concept|SIMPLE_SEGMENT|4883,4892|true|false|false|C0442805;C5236002|Increase;Increased (finding)|increased
Finding|Sign or Symptom|SIMPLE_SEGMENT|4883,4910|true|false|false|C0859927|Increased work of breathing|increased work of breathing
Event|Occupational Activity|SIMPLE_SEGMENT|4893,4897|true|false|false|C0043227|Work|work
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|4893,4910|true|false|false|C0043229|Work of Breathing|work of breathing
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4901,4910|false|false|false|C5885990||breathing
Finding|Finding|SIMPLE_SEGMENT|4901,4910|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|SIMPLE_SEGMENT|4901,4910|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|SIMPLE_SEGMENT|4901,4910|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|SIMPLE_SEGMENT|4901,4910|false|false|false|C1160636|respiratory system process|breathing
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4912,4919|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4912,4919|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Finding|Finding|SIMPLE_SEGMENT|4912,4919|false|false|false|C0941288|Abdomen problem|ABDOMEN
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4928,4934|false|false|false|C0021853|Intestines|bowels
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|4935,4941|false|false|false|C0037709||sounds
Finding|Finding|SIMPLE_SEGMENT|4947,4956|false|false|false|C0700124|Dilated|distended
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4972,4976|false|false|false|C4318566|Deep Resection Margin|deep
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4977,4986|false|false|false|C0030247|Palpation|palpation
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5010,5021|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|5026,5034|true|false|false|C0149651|Clubbing|clubbing
Finding|Sign or Symptom|SIMPLE_SEGMENT|5036,5044|true|false|false|C0010520|Cyanosis|cyanosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5049,5054|true|false|false|C1717255||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|5049,5054|true|false|false|C0013604|Edema|edema
Drug|Food|SIMPLE_SEGMENT|5056,5062|false|false|false|C5890763||Pulses
Finding|Physiologic Function|SIMPLE_SEGMENT|5056,5062|false|false|false|C0391850|Physiologic pulse|Pulses
Procedure|Health Care Activity|SIMPLE_SEGMENT|5056,5062|false|false|false|C0034107|Pulse taking|Pulses
Finding|Conceptual Entity|SIMPLE_SEGMENT|5066,5072|false|false|false|C0442038;C0920847|Circumpennate;Radial|Radial
Anatomy|Body System|SIMPLE_SEGMENT|5090,5094|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5090,5094|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5090,5094|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Finding|Body Substance|SIMPLE_SEGMENT|5090,5094|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|SIMPLE_SEGMENT|5090,5094|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Finding|SIMPLE_SEGMENT|5096,5100|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|5096,5100|false|false|false|C0687712|warming process|Warm
Finding|Gene or Genome|SIMPLE_SEGMENT|5120,5123|false|false|false|C1539110|CNDP2 gene|CN2
Finding|Finding|SIMPLE_SEGMENT|5127,5133|false|false|false|C1554187|Gender Status - Intact|intact
Finding|Finding|SIMPLE_SEGMENT|5152,5166|false|false|false|C0026826|Muscle Hypertonia|Increased tone
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5170,5173|false|false|false|C0227192|Inferior esophageal sphincter structure|LEs
Finding|Classification|SIMPLE_SEGMENT|5170,5173|false|false|false|C0023595|Lewis Blood-Group System|LEs
Finding|Idea or Concept|SIMPLE_SEGMENT|5179,5187|false|false|false|C0808080|Strength (attribute)|strength
Finding|Finding|SIMPLE_SEGMENT|5204,5213|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|5204,5213|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|SIMPLE_SEGMENT|5204,5213|false|false|false|C2229507|sensory exam|sensation
Procedure|Health Care Activity|SIMPLE_SEGMENT|5237,5246|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5247,5251|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5281,5286|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5281,5286|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|5287,5290|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|5295,5298|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5295,5298|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5295,5298|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5305,5308|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5305,5308|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|5305,5308|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5305,5308|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5315,5318|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5315,5318|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|5326,5329|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5326,5329|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5326,5329|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5326,5329|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|5333,5336|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5333,5336|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|5333,5336|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|5333,5336|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5333,5336|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5342,5346|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5372,5375|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5392,5397|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5392,5397|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Antibiotic|SIMPLE_SEGMENT|5413,5418|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5413,5418|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|SIMPLE_SEGMENT|5413,5418|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5426,5429|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|Eos
Finding|Gene or Genome|SIMPLE_SEGMENT|5426,5429|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|Eos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5528,5533|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5528,5533|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5538,5541|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5538,5541|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5564,5569|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5564,5569|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|5564,5577|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5564,5577|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5564,5577|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5570,5577|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|5570,5577|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5570,5577|false|false|false|C0017725|glucose|Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5570,5577|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5570,5577|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5623,5627|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5623,5627|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5623,5627|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5653,5658|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5653,5658|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5659,5662|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5659,5662|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|SIMPLE_SEGMENT|5659,5662|false|false|false|C0001899|Alanine Transaminase|ALT
Finding|Gene or Genome|SIMPLE_SEGMENT|5659,5662|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|SIMPLE_SEGMENT|5659,5662|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|SIMPLE_SEGMENT|5659,5662|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5659,5662|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5666,5669|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5666,5669|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5666,5669|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5666,5669|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|SIMPLE_SEGMENT|5666,5669|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Finding|Gene or Genome|SIMPLE_SEGMENT|5666,5669|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5673,5680|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|SIMPLE_SEGMENT|5673,5680|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5709,5714|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5709,5714|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5715,5721|false|false|false|C0023764|lipase|Lipase
Drug|Enzyme|SIMPLE_SEGMENT|5715,5721|false|false|false|C0023764|lipase|Lipase
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5715,5721|false|false|false|C0023764|lipase|Lipase
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5715,5721|false|false|false|C0373670|Lipase measurement|Lipase
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5737,5742|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5737,5742|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5769,5774|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5769,5774|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5769,5782|false|false|false|C0853248|Blood albumin|BLOOD Albumin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5775,5782|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5775,5782|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5775,5782|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Finding|Gene or Genome|SIMPLE_SEGMENT|5775,5782|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Finding|Physiologic Function|SIMPLE_SEGMENT|5775,5782|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5775,5782|false|false|false|C0201838|Albumin measurement|Albumin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5787,5794|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|5787,5794|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5787,5794|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5787,5794|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|5787,5794|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|5787,5794|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5787,5794|false|false|false|C0201925|Calcium measurement|Calcium
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5827,5832|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5827,5832|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5856,5861|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5856,5861|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5862,5865|false|false|false|C2708739||TSH
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5862,5865|false|false|false|C0040160|thyrotropin|TSH
Drug|Hormone|SIMPLE_SEGMENT|5862,5865|false|false|false|C0040160|thyrotropin|TSH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5862,5865|false|false|false|C0040160|thyrotropin|TSH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5862,5865|false|false|false|C0202230|Thyroid stimulating hormone measurement|TSH
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5882,5887|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5882,5887|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Finding|Finding|SIMPLE_SEGMENT|5896,5899|false|false|false|C5848551|Neg - answer|NEG
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5912,5917|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5912,5917|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5918,5921|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Enzyme|SIMPLE_SEGMENT|5918,5921|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Organic Chemical|SIMPLE_SEGMENT|5918,5921|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5918,5921|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Finding|Gene or Genome|SIMPLE_SEGMENT|5918,5921|false|false|false|C1412553|ARSA gene|ASA
Finding|Finding|SIMPLE_SEGMENT|5922,5925|false|false|false|C5848551|Neg - answer|NEG
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|5926,5933|false|false|false|C0161679|Toxic effect of ethyl alcohol|Ethanol
Drug|Organic Chemical|SIMPLE_SEGMENT|5926,5933|false|false|false|C0001962;C3854029;C3854030|CNS depressants ethanol;antiseptics ethanol;ethanol|Ethanol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5926,5933|false|false|false|C0001962;C3854029;C3854030|CNS depressants ethanol;antiseptics ethanol;ethanol|Ethanol
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5926,5933|false|false|false|C0202304|Ethanol measurement|Ethanol
Finding|Finding|SIMPLE_SEGMENT|5934,5937|false|false|false|C5848551|Neg - answer|NEG
Finding|Finding|SIMPLE_SEGMENT|5946,5949|false|false|false|C5848551|Neg - answer|NEG
Finding|Finding|SIMPLE_SEGMENT|5959,5962|false|false|false|C5848551|Neg - answer|NEG
Finding|Finding|SIMPLE_SEGMENT|5964,5971|false|false|false|C0740845|Imaging problem|IMAGING
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5964,5971|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|IMAGING
Finding|Finding|SIMPLE_SEGMENT|5986,5993|false|false|false|C0740845|Imaging problem|Imaging
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5986,5993|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|Imaging
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5994,6001|false|false|false|C0881943||CT HEAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5994,6001|false|false|false|C0202691|CAT scan of head|CT HEAD
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5997,6001|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|HEAD
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5997,6001|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|HEAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5997,6001|false|false|false|C0362076|Problems with head|HEAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5997,6001|false|false|false|C0876917|Procedure on head|HEAD
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|6006,6014|false|false|false|C0009924|Contrast Media|CONTRAST
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6017,6025|false|false|false|C2926606||FINDINGS
Finding|Functional Concept|SIMPLE_SEGMENT|6017,6025|false|false|false|C2607943|findings aspects|FINDINGS
Finding|Idea or Concept|SIMPLE_SEGMENT|6041,6049|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|6041,6052|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Finding|Pathologic Function|SIMPLE_SEGMENT|6053,6063|true|false|false|C0021308|Infarction|infarction
Finding|Pathologic Function|SIMPLE_SEGMENT|6065,6075|true|false|false|C0019080|Hemorrhage|hemorrhage
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6077,6082|true|false|false|C1717255||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|6077,6082|true|false|false|C0013604|Edema|edema
Finding|Finding|SIMPLE_SEGMENT|6087,6091|true|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|SIMPLE_SEGMENT|6087,6091|true|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|SIMPLE_SEGMENT|6087,6091|true|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6123,6133|false|false|false|C0018827|Heart Ventricle|ventricles
Finding|Functional Concept|SIMPLE_SEGMENT|6144,6154|false|false|false|C0332299|Suggestive of|suggestive
Finding|Functional Concept|SIMPLE_SEGMENT|6144,6157|false|false|false|C0332299|Suggestive of|suggestive of
Finding|Functional Concept|SIMPLE_SEGMENT|6172,6179|false|false|false|C0392747|Changing|changes
Finding|Idea or Concept|SIMPLE_SEGMENT|6194,6202|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|6194,6205|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|6206,6214|true|false|false|C0016658|Fracture|fracture
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|6259,6276|false|false|false|C0030471|Nasal sinus|paranasal sinuses
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|6269,6276|false|false|false|C0030471;C4071871|Head>Sinuses;Nasal sinus|sinuses
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|6269,6276|false|false|false|C0016169|pathologic fistula|sinuses
Finding|Intellectual Product|SIMPLE_SEGMENT|6281,6287|false|false|false|C1552826|Table Cell Vertical Align - middle|middle
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|6281,6291|false|false|false|C0013455|middle ear|middle ear
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6281,6291|false|false|false|C0271428;C0496788|Disorder of middle ear;Malignant neoplasm of middle ear|middle ear
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6281,6291|false|false|false|C0271428;C0496788|Disorder of middle ear;Malignant neoplasm of middle ear|middle ear
Procedure|Health Care Activity|SIMPLE_SEGMENT|6281,6291|false|false|false|C2228461|examination of middle ear|middle ear
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6288,6291|false|false|false|C0013443;C0521421|Ear structure|ear
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6288,6291|false|false|false|C0851354|Ear and labyrinth disorders|ear
Finding|Body Substance|SIMPLE_SEGMENT|6288,6291|false|false|false|C1546608;C1550629|SpecimenType - Ear|ear
Finding|Intellectual Product|SIMPLE_SEGMENT|6288,6291|false|false|false|C1546608;C1550629|SpecimenType - Ear|ear
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|6292,6300|false|false|false|C0333343|Body cavities|cavities
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|6292,6300|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavities
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6292,6300|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavities
Finding|Idea or Concept|SIMPLE_SEGMENT|6305,6310|false|false|false|C1550016|Remote control command - Clear|clear
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|6344,6350|false|false|false|C0029180|Ocular orbit|orbits
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6390,6394|false|false|false|C0023317|Lens, Crystalline|lens
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6390,6394|false|false|false|C0023308|Lens Diseases|lens
Procedure|Health Care Activity|SIMPLE_SEGMENT|6390,6394|false|false|false|C2239142|examination of lens|lens
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6395,6407|false|false|false|C0035139|Surgical Replantation|replacements
Finding|Intellectual Product|SIMPLE_SEGMENT|6410,6420|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|6410,6420|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|6429,6434|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6435,6447|false|false|false|C0524466|Intracranial|intracranial
Finding|Functional Concept|SIMPLE_SEGMENT|6435,6447|false|false|false|C1522213|Intracranial Route of Administration|intracranial
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|6448,6459|true|false|false|C0000768|Congenital Abnormality|abnormality
Finding|Finding|SIMPLE_SEGMENT|6448,6459|true|false|false|C1704258|Abnormality|abnormality
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6465,6478|true|false|false|C0020255|Hydrocephalus|hydrocephalus
Finding|Finding|SIMPLE_SEGMENT|6486,6493|false|false|false|C0740845|Imaging problem|Imaging
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6486,6493|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|Imaging
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6494,6499|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|CHEST
Finding|Finding|SIMPLE_SEGMENT|6494,6499|false|false|false|C0741025|Chest problem|CHEST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6506,6509|false|false|false|C1366678;C1433371;C4049852|L-Type Amino Acid Transporter;LAT protein, human;ORC3 protein, human|LAT
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6506,6509|false|false|false|C1366678;C1433371;C4049852|L-Type Amino Acid Transporter;LAT protein, human;ORC3 protein, human|LAT
Drug|Immunologic Factor|SIMPLE_SEGMENT|6506,6509|false|false|false|C1366678;C1433371;C4049852|L-Type Amino Acid Transporter;LAT protein, human;ORC3 protein, human|LAT
Finding|Gene or Genome|SIMPLE_SEGMENT|6506,6509|false|false|false|C1335085;C1425844;C1705279;C2240043|LAT gene;ORC3 gene;ORC3 wt Allele;SPNS1 gene|LAT
Finding|Intellectual Product|SIMPLE_SEGMENT|6512,6522|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|6512,6522|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|6526,6530|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Finding|Pathologic Function|SIMPLE_SEGMENT|6531,6542|false|false|false|C0004144|Atelectasis|atelectasis
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6550,6554|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6550,6554|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6550,6554|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|SIMPLE_SEGMENT|6550,6554|false|false|false|C0740941|Lung Problem|lung
Drug|Chemical Viewed Functionally|SIMPLE_SEGMENT|6555,6560|false|false|false|C0178499|Base|bases
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6575,6588|true|false|false|C0521530|Lung consolidation|consolidation
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6593,6596|false|false|false|C1114365||Age
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6593,6596|false|false|false|C0162574|Glycation End Products, Advanced|Age
Drug|Organic Chemical|SIMPLE_SEGMENT|6593,6596|false|false|false|C0162574|Glycation End Products, Advanced|Age
Finding|Finding|SIMPLE_SEGMENT|6611,6619|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|SIMPLE_SEGMENT|6611,6619|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Finding|SIMPLE_SEGMENT|6623,6629|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|SIMPLE_SEGMENT|6623,6629|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Functional Concept|SIMPLE_SEGMENT|6630,6641|false|false|false|C0332459;C4551657|Compressed structure|compression
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|6630,6641|false|false|false|C0728907|Compression|compression
Procedure|Machine Activity|SIMPLE_SEGMENT|6630,6641|false|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6630,6641|false|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|6642,6651|false|false|false|C0000768;C0302142|Congenital Abnormality;Deformity|deformity
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|6642,6651|false|false|false|C0000768;C0302142|Congenital Abnormality;Deformity|deformity
Finding|Finding|SIMPLE_SEGMENT|6642,6651|false|false|false|C2117111||deformity
Finding|Finding|SIMPLE_SEGMENT|6658,6661|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|SIMPLE_SEGMENT|6658,6661|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6662,6670|false|false|false|C0817096|Chest|thoracic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6662,6670|false|false|false|C5779551|Dissecting Thoracic Aortic Aneurysm|thoracic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6662,6685|false|false|false|C0223199;C1305451|Structure of body of thoracic vertebra|thoracic vertebral body
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6671,6680|false|false|false|C0549207|Bone structure of spine|vertebral
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6671,6685|false|false|false|C0223084|Body of vertebra|vertebral body
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|6681,6685|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6681,6685|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Finding|Intellectual Product|SIMPLE_SEGMENT|6681,6685|false|false|false|C1551342|Document Body|body
Finding|Body Substance|SIMPLE_SEGMENT|6689,6698|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|6689,6698|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|6689,6698|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|6689,6698|false|false|false|C0030685|Patient Discharge|DISCHARGE
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6699,6703|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6733,6738|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|6733,6738|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|6739,6742|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|6747,6750|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6747,6750|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6747,6750|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6757,6760|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6757,6760|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|6757,6760|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6757,6760|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6767,6770|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6767,6770|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|6778,6781|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6778,6781|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6778,6781|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6778,6781|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|6785,6788|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6785,6788|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|6785,6788|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|6785,6788|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6785,6788|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6795,6799|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6825,6828|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6845,6850|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|6845,6850|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|6845,6858|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6845,6858|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6845,6858|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6851,6858|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|6851,6858|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6851,6858|false|false|false|C0017725|glucose|Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6851,6858|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6851,6858|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|SIMPLE_SEGMENT|6902,6906|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6902,6906|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6902,6906|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6931,6936|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|6931,6936|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6931,6944|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6937,6944|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|6937,6944|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|6937,6944|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6937,6944|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|6937,6944|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|6937,6944|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6937,6944|false|false|false|C0201925|Calcium measurement|Calcium
Finding|Finding|SIMPLE_SEGMENT|6967,6971|false|false|false|C1706180|Male Gender|male
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6981,6988|false|false|false|C0012634|Disease|disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6990,7002|false|false|false|C0242339|Dyslipidemias|dyslipidemia
Finding|Conceptual Entity|SIMPLE_SEGMENT|7010,7017|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|7010,7017|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|7010,7017|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|7010,7020|false|false|false|C0262926|Medical History|history of
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7021,7029|false|false|false|C0033572;C4266527|Prostate;Structure of prostate (body structure)|prostate
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7021,7029|false|false|false|C0033575;C0154009;C0154088;C0496923|Benign neoplasm of prostate;Carcinoma in situ of prostate;Neoplasm of uncertain or unknown behavior of prostate;Prostatic Diseases|prostate
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7021,7029|false|false|false|C0033575;C0154009;C0154088;C0496923|Benign neoplasm of prostate;Carcinoma in situ of prostate;Neoplasm of uncertain or unknown behavior of prostate;Prostatic Diseases|prostate
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7021,7036|false|false|false|C0376358;C0600139|Malignant neoplasm of prostate;Prostate carcinoma|prostate cancer
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7030,7036|false|false|false|C0006826|Malignant Neoplasms|cancer
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7042,7055|false|false|false|C0033573|Prostatectomy|prostatectomy
Finding|Finding|SIMPLE_SEGMENT|7117,7121|false|false|false|C0016928|Gait|gait
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|7123,7128|false|false|false|C0000921|Accidental Falls|falls
Finding|Finding|SIMPLE_SEGMENT|7123,7128|false|false|false|C0085639|Falls|falls
Finding|Functional Concept|SIMPLE_SEGMENT|7134,7140|false|false|false|C0234621|Visual|visual
Finding|Sign or Symptom|SIMPLE_SEGMENT|7134,7155|false|false|false|C0233763|Hallucinations, Visual|visual hallucinations
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|7141,7155|false|false|false|C0018524|Hallucinations|hallucinations
Finding|Functional Concept|SIMPLE_SEGMENT|7171,7182|false|false|false|C0242656;C0449258|Disease Progression;Progression|progression
Finding|Pathologic Function|SIMPLE_SEGMENT|7171,7182|false|false|false|C0242656;C0449258|Disease Progression;Progression|progression
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7190,7209|false|false|false|C0027765|nervous system disorder|neurologic disorder
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7201,7209|false|false|false|C0012634|Disease|disorder
Finding|Intellectual Product|SIMPLE_SEGMENT|7213,7218|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|ACUTE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7259,7266|false|false|false|C0012634|Disease|disease
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|7271,7275|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|Body
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7271,7275|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|Body
Finding|Intellectual Product|SIMPLE_SEGMENT|7271,7275|false|false|false|C1551342|Document Body|Body
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|7276,7284|false|false|false|C0011265;C0497327|Dementia;Presenile dementia|Dementia
Finding|Functional Concept|SIMPLE_SEGMENT|7287,7293|false|false|false|C0234621|Visual|Visual
Finding|Sign or Symptom|SIMPLE_SEGMENT|7287,7308|false|false|false|C0233763|Hallucinations, Visual|Visual Hallucinations
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|7294,7308|false|false|false|C0018524|Hallucinations|Hallucinations
Finding|Body Substance|SIMPLE_SEGMENT|7314,7321|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|7314,7321|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|7314,7321|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|7338,7343|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Intellectual Product|SIMPLE_SEGMENT|7347,7354|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|7347,7354|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Finding|Functional Concept|SIMPLE_SEGMENT|7355,7366|false|false|false|C0242656;C0449258|Disease Progression;Progression|progression
Finding|Pathologic Function|SIMPLE_SEGMENT|7355,7366|false|false|false|C0242656;C0449258|Disease Progression;Progression|progression
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7378,7385|false|false|false|C0012634|Disease|disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7406,7413|false|false|false|C0012634|Disease|disease
Finding|Pathologic Function|SIMPLE_SEGMENT|7406,7425|false|false|false|C0242656|Disease Progression|disease progression
Finding|Functional Concept|SIMPLE_SEGMENT|7414,7425|false|false|false|C0242656;C0449258|Disease Progression;Progression|progression
Finding|Pathologic Function|SIMPLE_SEGMENT|7414,7425|false|false|false|C0242656;C0449258|Disease Progression;Progression|progression
Finding|Functional Concept|SIMPLE_SEGMENT|7440,7447|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Idea or Concept|SIMPLE_SEGMENT|7440,7447|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Intellectual Product|SIMPLE_SEGMENT|7440,7447|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|7440,7447|false|false|false|C0199168|Medical service|medical
Finding|Conceptual Entity|SIMPLE_SEGMENT|7448,7453|false|false|false|C0015127;C1524003|Etiology aspects;Science of Etiology|cause
Finding|Functional Concept|SIMPLE_SEGMENT|7448,7453|false|false|false|C0015127;C1524003|Etiology aspects;Science of Etiology|cause
Drug|Organic Chemical|SIMPLE_SEGMENT|7465,7472|false|false|false|C0721754|Mirapex|mirapex
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7465,7472|false|false|false|C0721754|Mirapex|mirapex
Drug|Organic Chemical|SIMPLE_SEGMENT|7474,7484|false|false|false|C0525678|rasagiline|rasagiline
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7474,7484|false|false|false|C0525678|rasagiline|rasagiline
Drug|Organic Chemical|SIMPLE_SEGMENT|7491,7503|false|false|false|C0649350|rivastigmine|rivastigmine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7491,7503|false|false|false|C0649350|rivastigmine|rivastigmine
Drug|Organic Chemical|SIMPLE_SEGMENT|7535,7543|false|false|false|C0287163|Seroquel|Seroquel
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7535,7543|false|false|false|C0287163|Seroquel|Seroquel
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|7553,7567|false|false|false|C0018524|Hallucinations|hallucinations
Finding|Finding|SIMPLE_SEGMENT|7590,7598|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Finding|Functional Concept|SIMPLE_SEGMENT|7590,7598|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|7590,7598|false|false|false|C0031809|Physical Examination|physical
Finding|Intellectual Product|SIMPLE_SEGMENT|7590,7606|false|false|false|C1547999|Diagnostic Service Section ID - Physical Therapy|physical therapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7590,7606|false|false|false|C0949766|Physical therapy|physical therapy
Finding|Finding|SIMPLE_SEGMENT|7599,7606|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|SIMPLE_SEGMENT|7599,7606|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7599,7606|false|false|false|C0087111|Therapeutic procedure|therapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7623,7628|false|false|false|C0034991|Rehabilitation therapy|rehab
Finding|Idea or Concept|SIMPLE_SEGMENT|7636,7650|false|false|false|C0034866|Recommendation|recommendation
Finding|Classification|SIMPLE_SEGMENT|7674,7680|false|false|true|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|7674,7680|false|false|true|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|7674,7680|false|false|true|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|7674,7680|false|false|true|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Body Substance|SIMPLE_SEGMENT|7696,7705|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|7696,7705|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|7696,7705|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|7696,7705|false|false|false|C0030685|Patient Discharge|discharge
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7696,7713|false|false|false|C0184713|Discharge to home|discharge to home
Finding|Idea or Concept|SIMPLE_SEGMENT|7709,7713|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|7709,7713|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|7709,7713|false|false|false|C1553498|home health encounter|home
Finding|Idea or Concept|SIMPLE_SEGMENT|7719,7723|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|7719,7723|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|7719,7723|false|false|false|C1553498|home health encounter|home
Finding|Finding|SIMPLE_SEGMENT|7724,7732|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Finding|Functional Concept|SIMPLE_SEGMENT|7724,7732|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|7724,7732|false|false|false|C0031809|Physical Examination|physical
Finding|Intellectual Product|SIMPLE_SEGMENT|7724,7740|false|false|false|C1547999|Diagnostic Service Section ID - Physical Therapy|physical therapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7724,7740|false|false|false|C0949766|Physical therapy|physical therapy
Finding|Finding|SIMPLE_SEGMENT|7733,7740|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|SIMPLE_SEGMENT|7733,7740|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7733,7740|false|false|false|C0087111|Therapeutic procedure|therapy
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7756,7760|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|7756,7760|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Substance|SIMPLE_SEGMENT|7756,7760|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Finding|Intellectual Product|SIMPLE_SEGMENT|7756,7760|false|false|false|C1546701|line source specimen code|line
Finding|Body Substance|SIMPLE_SEGMENT|7771,7778|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|7771,7778|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|7771,7778|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7781,7786|false|false|false|C2979882||goals
Finding|Idea or Concept|SIMPLE_SEGMENT|7781,7786|false|false|false|C0018017;C0679840;C1546459|What subject filter - Goals;objective (goal);treatment goals|goals
Finding|Intellectual Product|SIMPLE_SEGMENT|7781,7786|false|false|false|C0018017;C0679840;C1546459|What subject filter - Goals;objective (goal);treatment goals|goals
Procedure|Health Care Activity|SIMPLE_SEGMENT|7781,7794|false|false|false|C2930505|Goals of Care|goals of care
Event|Activity|SIMPLE_SEGMENT|7790,7794|false|false|false|C1947933|care activity|care
Finding|Finding|SIMPLE_SEGMENT|7790,7794|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|7790,7794|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Idea or Concept|SIMPLE_SEGMENT|7797,7809|false|false|false|C1548597|Marketing basis - Transitional|TRANSITIONAL
Finding|Functional Concept|SIMPLE_SEGMENT|7825,7831|false|false|false|C0234621|Visual|visual
Finding|Sign or Symptom|SIMPLE_SEGMENT|7825,7845|false|false|false|C0233763|Hallucinations, Visual|visual hallucination
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|7832,7845|false|false|false|C0018524|Hallucinations|hallucination
Finding|Functional Concept|SIMPLE_SEGMENT|7846,7854|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|7846,7854|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Drug|Organic Chemical|SIMPLE_SEGMENT|7858,7866|false|false|false|C0287163|Seroquel|Seroquel
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7858,7866|false|false|false|C0287163|Seroquel|Seroquel
Finding|Finding|SIMPLE_SEGMENT|7874,7882|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Finding|Functional Concept|SIMPLE_SEGMENT|7874,7882|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|7874,7882|false|false|false|C0031809|Physical Examination|physical
Finding|Intellectual Product|SIMPLE_SEGMENT|7874,7890|false|false|false|C1547999|Diagnostic Service Section ID - Physical Therapy|physical therapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7874,7890|false|false|false|C0949766|Physical therapy|physical therapy
Finding|Finding|SIMPLE_SEGMENT|7883,7890|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|SIMPLE_SEGMENT|7883,7890|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7883,7890|false|false|false|C0087111|Therapeutic procedure|therapy
Finding|Finding|SIMPLE_SEGMENT|7891,7898|false|false|false|C4534363|At home|at home
Finding|Idea or Concept|SIMPLE_SEGMENT|7894,7898|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|7894,7898|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|7894,7898|false|false|false|C1553498|home health encounter|home
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7901,7912|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7901,7912|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|7901,7912|false|false|false|C4284232|Medications|Medications
Finding|Finding|SIMPLE_SEGMENT|7901,7925|false|false|false|C1627937|Medications on admission|Medications on Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|7916,7925|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7944,7954|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|7944,7954|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|7944,7959|false|false|false|C0746470|MEDICATION LIST|Medication list
Finding|Intellectual Product|SIMPLE_SEGMENT|7955,7959|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Finding|Intellectual Product|SIMPLE_SEGMENT|7999,8012|false|false|false|C1552578|Act Class - investigation|investigation
Procedure|Health Care Activity|SIMPLE_SEGMENT|7999,8012|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|investigation
Drug|Organic Chemical|SIMPLE_SEGMENT|8017,8027|false|false|false|C0525678|rasagiline|Rasagiline
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8017,8027|false|false|false|C0525678|rasagiline|Rasagiline
Drug|Organic Chemical|SIMPLE_SEGMENT|8046,8057|false|false|false|C0074710|pramipexole|Pramipexole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8046,8057|false|false|false|C0074710|pramipexole|Pramipexole
Drug|Organic Chemical|SIMPLE_SEGMENT|8078,8090|false|false|false|C0649350|rivastigmine|rivastigmine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8078,8090|false|false|false|C0649350|rivastigmine|rivastigmine
Finding|Finding|SIMPLE_SEGMENT|8104,8115|false|false|false|C0040652;C0694643;C4521342|Transdermal (intended site);Transdermal Route of Administration;transdermal|transdermal
Finding|Functional Concept|SIMPLE_SEGMENT|8104,8115|false|false|false|C0040652;C0694643;C4521342|Transdermal (intended site);Transdermal Route of Administration;transdermal|transdermal
Drug|Organic Chemical|SIMPLE_SEGMENT|8126,8137|false|false|false|C0085542|pravastatin|Pravastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8126,8137|false|false|false|C0085542|pravastatin|Pravastatin
Drug|Organic Chemical|SIMPLE_SEGMENT|8155,8169|false|false|false|C0042845;C3714801|Cyanocobalamin Drug Class;vitamin B12|Cyanocobalamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8155,8169|false|false|false|C0042845;C3714801|Cyanocobalamin Drug Class;vitamin B12|Cyanocobalamin
Drug|Vitamin|SIMPLE_SEGMENT|8155,8169|false|false|false|C0042845;C3714801|Cyanocobalamin Drug Class;vitamin B12|Cyanocobalamin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8178,8185|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|Unknown
Drug|Immunologic Factor|SIMPLE_SEGMENT|8178,8185|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|Unknown
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8178,8185|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|Unknown
Finding|Finding|SIMPLE_SEGMENT|8178,8185|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|Unknown
Finding|Functional Concept|SIMPLE_SEGMENT|8178,8185|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|Unknown
Finding|Idea or Concept|SIMPLE_SEGMENT|8178,8185|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|Unknown
Finding|Intellectual Product|SIMPLE_SEGMENT|8178,8185|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|Unknown
Drug|Organic Chemical|SIMPLE_SEGMENT|8200,8210|false|false|false|C0065180|loratadine|Loratadine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8200,8210|false|false|false|C0065180|loratadine|Loratadine
Finding|Body Substance|SIMPLE_SEGMENT|8230,8239|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|8230,8239|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|8230,8239|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|8230,8239|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|8230,8251|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8240,8251|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8240,8251|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|8240,8251|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|SIMPLE_SEGMENT|8257,8267|false|false|false|C0123091|quetiapine|QUEtiapine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8257,8267|false|false|false|C0123091|quetiapine|QUEtiapine
Drug|Organic Chemical|SIMPLE_SEGMENT|8257,8276|false|false|false|C0724680|quetiapine fumarate|QUEtiapine Fumarate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8257,8276|false|false|false|C0724680|quetiapine fumarate|QUEtiapine Fumarate
Drug|Organic Chemical|SIMPLE_SEGMENT|8268,8276|false|false|false|C0220833|fumarate|Fumarate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8268,8276|false|false|false|C0220833|fumarate|Fumarate
Drug|Organic Chemical|SIMPLE_SEGMENT|8295,8305|false|false|false|C0123091|quetiapine|quetiapine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8295,8305|false|false|false|C0123091|quetiapine|quetiapine
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8314,8320|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|SIMPLE_SEGMENT|8324,8332|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|8327,8332|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|8327,8332|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8353,8359|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|SIMPLE_SEGMENT|8360,8367|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|8376,8386|false|false|false|C0065180|loratadine|Loratadine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8376,8386|false|false|false|C0065180|loratadine|Loratadine
Drug|Organic Chemical|SIMPLE_SEGMENT|8408,8419|false|false|false|C0074710|pramipexole|Pramipexole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8408,8419|false|false|false|C0074710|pramipexole|Pramipexole
Drug|Organic Chemical|SIMPLE_SEGMENT|8442,8453|false|false|false|C0085542|pravastatin|Pravastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8442,8453|false|false|false|C0085542|pravastatin|Pravastatin
Drug|Organic Chemical|SIMPLE_SEGMENT|8473,8483|false|false|false|C0525678|rasagiline|Rasagiline
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8473,8483|false|false|false|C0525678|rasagiline|Rasagiline
Drug|Organic Chemical|SIMPLE_SEGMENT|8504,8516|false|false|false|C0649350|rivastigmine|rivastigmine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8504,8516|false|false|false|C0649350|rivastigmine|rivastigmine
Finding|Finding|SIMPLE_SEGMENT|8530,8541|false|false|false|C0040652;C0694643;C4521342|Transdermal (intended site);Transdermal Route of Administration;transdermal|transdermal
Finding|Functional Concept|SIMPLE_SEGMENT|8530,8541|false|false|false|C0040652;C0694643;C4521342|Transdermal (intended site);Transdermal Route of Administration;transdermal|transdermal
Finding|Body Substance|SIMPLE_SEGMENT|8553,8562|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|8553,8562|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|8553,8562|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|8553,8562|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8553,8574|false|false|false|C4019243||Discharge Disposition
Finding|Finding|SIMPLE_SEGMENT|8553,8574|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8563,8574|false|false|false|C2926604||Disposition
Procedure|Health Care Activity|SIMPLE_SEGMENT|8563,8574|false|false|false|C0184758|Patient disposition|Disposition
Finding|Idea or Concept|SIMPLE_SEGMENT|8576,8580|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|SIMPLE_SEGMENT|8576,8580|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|SIMPLE_SEGMENT|8576,8580|false|false|false|C1553498|home health encounter|Home
Event|Occupational Activity|SIMPLE_SEGMENT|8586,8593|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|8586,8593|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Finding|Intellectual Product|SIMPLE_SEGMENT|8596,8604|false|false|false|C4695111|ADMIN.FACILITY|Facility
Finding|Body Substance|SIMPLE_SEGMENT|8612,8621|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|8612,8621|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|8612,8621|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|8612,8621|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|8612,8631|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8622,8631|false|false|false|C0945731||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|8622,8631|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|8622,8631|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8622,8631|false|false|false|C0011900|Diagnosis|Diagnosis
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|8637,8645|false|false|false|C0011265;C0497327|Dementia;Presenile dementia|Dementia
Finding|Body Substance|SIMPLE_SEGMENT|8648,8657|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|8648,8657|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|8648,8657|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|8648,8657|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8658,8667|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8658,8667|false|false|false|C0012634|Disease|Condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|8658,8667|false|false|false|C1705253|Logical Condition|Condition
Finding|Mental Process|SIMPLE_SEGMENT|8669,8675|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8669,8682|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|SIMPLE_SEGMENT|8669,8682|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8676,8682|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|8676,8682|false|false|false|C1546481|What subject filter - Status|Status
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|8684,8692|false|false|false|C0009676|Confusion|Confused
Finding|Finding|SIMPLE_SEGMENT|8684,8692|false|false|false|C0683369;C1547301|Clouded consciousness;Precaution Code - Confused|Confused
Finding|Intellectual Product|SIMPLE_SEGMENT|8684,8692|false|false|false|C0683369;C1547301|Clouded consciousness;Precaution Code - Confused|Confused
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8706,8728|false|false|false|C4050479||Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|8706,8728|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|8715,8728|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|SIMPLE_SEGMENT|8715,8728|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8730,8735|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|8730,8735|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8730,8735|false|false|false|C0718338|Alert brand of caffeine|Alert
Finding|Finding|SIMPLE_SEGMENT|8730,8735|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|8730,8735|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|8730,8735|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|8740,8751|false|false|false|C1704675|Interaction|interactive
Finding|Body Substance|SIMPLE_SEGMENT|8756,8765|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|8756,8765|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|8756,8765|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|8756,8765|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8756,8778|false|false|false|C3669312||Discharge Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|8756,8778|false|false|false|C4282220|Discharge instructions|Discharge Instructions
Procedure|Health Care Activity|SIMPLE_SEGMENT|8756,8778|false|false|false|C2266673|hospital discharge instructions (treatment)|Discharge Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8766,8778|false|false|false|C3263700||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|8766,8778|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Finding|Gene or Genome|SIMPLE_SEGMENT|8780,8784|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Finding|Conceptual Entity|SIMPLE_SEGMENT|8805,8814|false|false|false|C1547898;C1706335;C1706336|Privilege;Role Privilege;User Privilege|privilege
Finding|Idea or Concept|SIMPLE_SEGMENT|8805,8814|false|false|false|C1547898;C1706335;C1706336|Privilege;Role Privilege;User Privilege|privilege
Finding|Idea or Concept|SIMPLE_SEGMENT|8857,8865|false|false|false|C1547192|Organization unit type - Hospital|HOSPITAL
Finding|Finding|SIMPLE_SEGMENT|8891,8900|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Idea or Concept|SIMPLE_SEGMENT|8891,8900|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Intellectual Product|SIMPLE_SEGMENT|8891,8900|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Pathologic Function|SIMPLE_SEGMENT|8891,8900|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|8891,8900|false|false|false|C0013956|Emergency Situation|emergency
Procedure|Health Care Activity|SIMPLE_SEGMENT|8891,8900|false|false|false|C1553500|emergency encounter|emergency
Finding|Idea or Concept|SIMPLE_SEGMENT|8891,8905|false|false|false|C1546435|Encounter Referral Source - emergency room|emergency room
Finding|Functional Concept|SIMPLE_SEGMENT|8966,8972|false|false|false|C0234621|Visual|visual
Finding|Sign or Symptom|SIMPLE_SEGMENT|8966,8987|false|false|false|C0233763|Hallucinations, Visual|visual hallucinations
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|8973,8987|false|false|false|C0018524|Hallucinations|hallucinations
Finding|Idea or Concept|SIMPLE_SEGMENT|9017,9025|false|false|false|C1547192|Organization unit type - Hospital|HOSPITAL
Finding|Finding|SIMPLE_SEGMENT|9052,9055|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|9052,9055|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9056,9066|false|false|false|C0013227|Pharmaceutical Preparations|medication
Finding|Intellectual Product|SIMPLE_SEGMENT|9056,9066|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Finding|Functional Concept|SIMPLE_SEGMENT|9087,9095|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|9087,9095|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Idea or Concept|SIMPLE_SEGMENT|9133,9141|false|false|false|C1547192|Organization unit type - Hospital|HOSPITAL
Finding|Idea or Concept|SIMPLE_SEGMENT|9146,9154|false|false|false|C0549178|Continuous|Continue
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9172,9181|false|false|false|C0013227|Pharmaceutical Preparations|medicines
Event|Activity|SIMPLE_SEGMENT|9197,9209|false|false|false|C0003629|Appointments|appointments
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9229,9233|false|false|false|C0339510|Vitelliform Macular Dystrophy|best
Finding|Gene or Genome|SIMPLE_SEGMENT|9229,9233|false|false|false|C1826421;C5781213|BEST1 gene;BEST1 wt Allele|best
Procedure|Health Care Activity|SIMPLE_SEGMENT|9266,9274|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9275,9287|false|false|false|C3263700||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|9275,9287|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

