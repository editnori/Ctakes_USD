 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|28,32
No|33,35
:|35,36
_|39,40
_|40,41
_|41,42
<EOL>|42,43
<EOL>|44,45
Admission|45,54
Date|55,59
:|59,60
_|62,63
_|63,64
_|64,65
Discharge|79,88
Date|89,93
:|93,94
_|97,98
_|98,99
_|99,100
<EOL>|100,101
<EOL>|102,103
Date|103,107
of|108,110
Birth|111,116
:|116,117
_|119,120
_|120,121
_|121,122
Sex|135,138
:|138,139
F|142,143
<EOL>|143,144
<EOL>|145,146
Service|146,153
:|153,154
ORTHOPAEDICS|155,167
<EOL>|167,168
<EOL>|169,170
Allergies|170,179
:|179,180
<EOL>|181,182
Codeine|182,189
/|190,191
Augmentin|192,201
/|202,203
Topamax|204,211
<EOL>|211,212
<EOL>|213,214
Attending|214,223
:|223,224
_|225,226
_|226,227
_|227,228
.|228,229
<EOL>|229,230
<EOL>|231,232
Chief|232,237
Complaint|238,247
:|247,248
<EOL>|248,249
Low|249,252
back|253,257
pain|258,262
with|263,267
radiation|268,277
down|278,282
the|283,286
right|287,292
leg|293,296
<EOL>|297,298
<EOL>|299,300
Major|300,305
Surgical|306,314
or|315,317
Invasive|318,326
Procedure|327,336
:|336,337
<EOL>|337,338
DECOMPRESSION|338,351
L2|352,354
-|354,355
S1|355,357
,|357,358
FUSION|359,365
L4|366,368
-|368,369
L5|369,371
,|371,372
DURAPLASTY|373,383
on|384,386
_|387,388
_|388,389
_|389,390
<EOL>|390,391
<EOL>|392,393
History|393,400
of|401,403
Present|404,411
Illness|412,419
:|419,420
<EOL>|420,421
Ms.|421,424
_|425,426
_|426,427
_|427,428
is|429,431
a|432,433
_|434,435
_|435,436
_|436,437
female|438,444
with|445,449
a|450,451
past|452,456
medical|457,464
<EOL>|465,466
history|466,473
significant|474,485
for|486,489
cerebral|490,498
aneurysm|499,507
,|507,508
abdominal|509,518
aortic|519,525
<EOL>|526,527
aneurysm|527,535
,|535,536
antiphospholipid|537,553
syndrome|554,562
w|563,564
/|564,565
multiple|566,574
DVTs|575,579
and|580,583
one|584,587
<EOL>|588,589
event|589,594
of|595,597
bilateral|598,607
large|608,613
PEs|614,617
on|618,620
warfarin|621,629
,|629,630
BRCA1|631,636
mutation|637,645
w|646,647
/|647,648
<EOL>|649,650
L|650,651
-|651,652
sided|652,657
breast|658,664
cancer|665,671
s|672,673
/|673,674
p|674,675
lumpectomy|676,686
,|686,687
who|688,691
presents|692,700
with|701,705
over|706,710
one|711,714
<EOL>|715,716
month|716,721
of|722,724
right|725,730
lower|731,736
back|737,741
pain|742,746
with|747,751
radicular|752,761
pain|762,766
down|767,771
the|772,775
<EOL>|776,777
right|777,782
leg|783,786
pain|787,791
.|791,792
She|793,796
had|797,800
recent|801,807
admission|808,817
_|818,819
_|819,820
_|820,821
for|822,825
acute|826,831
<EOL>|832,833
worsening|833,842
of|843,845
RLE|846,849
pain|850,854
and|855,858
swelling|859,867
in|868,870
background|871,881
of|882,884
about|885,890
4|891,892
<EOL>|893,894
months|894,900
right|901,906
leg|907,910
pain|911,915
.|915,916
RLE|917,920
US|921,923
did|924,927
not|928,931
show|932,936
evidence|937,945
of|946,948
DVT|949,952
.|952,953
Exam|954,958
<EOL>|959,960
was|960,963
most|964,968
consistent|969,979
with|980,984
right|985,990
trochanteric|991,1003
bursitis|1004,1012
and|1013,1016
pt|1017,1019
<EOL>|1020,1021
received|1021,1029
a|1030,1031
steroid|1032,1039
injection|1040,1049
.|1049,1050
Her|1051,1054
right|1055,1060
tibia|1061,1066
pain|1067,1071
was|1072,1075
felt|1076,1080
to|1081,1083
<EOL>|1084,1085
be|1085,1087
_|1088,1089
_|1089,1090
_|1090,1091
to|1092,1094
her|1095,1098
varicose|1099,1107
veins|1108,1113
.|1113,1114
On|1115,1117
this|1118,1122
admission|1123,1132
Imaging|1133,1140
notable|1141,1148
<EOL>|1149,1150
for|1150,1153
:|1153,1154
Normal|1156,1162
CT|1163,1165
A|1166,1167
/|1167,1168
P|1168,1169
with|1170,1174
no|1175,1177
e|1178,1179
/|1179,1180
o|1180,1181
nephrolithiasis|1182,1197
,|1197,1198
MR|1199,1201
_|1202,1203
_|1203,1204
_|1204,1205
spine|1206,1211
with|1212,1216
<EOL>|1217,1218
disc|1218,1222
bulge|1223,1228
at|1229,1231
L2|1232,1234
-|1234,1235
L3|1235,1237
and|1238,1241
L3|1242,1244
-|1244,1245
4|1245,1246
cause|1247,1252
severe|1253,1259
narrowing|1260,1269
of|1270,1272
the|1273,1276
<EOL>|1277,1278
spinal|1278,1284
canal|1285,1290
with|1291,1295
crowding|1296,1304
of|1305,1307
the|1308,1311
traversing|1312,1322
cauda|1323,1328
equina|1329,1335
.|1335,1336
<EOL>|1336,1337
<EOL>|1337,1338
<EOL>|1339,1340
Past|1340,1344
Medical|1345,1352
History|1353,1360
:|1360,1361
<EOL>|1361,1362
Dyslipidemia|1362,1374
,|1374,1375
<EOL>|1376,1377
Varicose|1377,1385
veins|1386,1391
(|1392,1393
R|1393,1394
>|1394,1395
L|1395,1396
)|1396,1397
s|1398,1399
/|1399,1400
p|1400,1401
ligation|1402,1410
,|1410,1411
<EOL>|1412,1413
COPD|1413,1417
,|1417,1418
<EOL>|1419,1420
OSA|1420,1423
(|1424,1425
+|1425,1426
CPap|1426,1430
)|1430,1431
,|1431,1432
<EOL>|1433,1434
recent|1434,1440
URI|1441,1444
(|1445,1446
received|1446,1454
course|1455,1461
of|1462,1464
Zithromax|1465,1474
)|1474,1475
,|1475,1476
<EOL>|1477,1478
bilateral|1478,1487
PEs|1488,1491
(|1492,1493
_|1493,1494
_|1494,1495
_|1495,1496
)|1496,1497
,|1497,1498
<EOL>|1499,1500
antiphospholipid|1500,1516
antibody|1517,1525
syndrome|1526,1534
(|1535,1536
on|1536,1538
lifelong|1539,1547
<EOL>|1548,1549
anticoagulation|1549,1564
)|1564,1565
,|1565,1566
<EOL>|1566,1567
<EOL>|1567,1568
T2DM|1568,1572
(|1573,1574
last|1574,1578
A1C|1579,1582
6.2|1583,1586
on|1587,1589
_|1590,1591
_|1591,1592
_|1592,1593
,|1593,1594
<EOL>|1595,1596
cerebral|1596,1604
aneurysm|1605,1613
(|1614,1615
followed|1615,1623
by|1624,1626
Dr.|1627,1630
_|1631,1632
_|1632,1633
_|1633,1634
,|1634,1635
unchanged|1636,1645
)|1645,1646
,|1646,1647
<EOL>|1648,1649
GERD|1649,1653
,|1653,1654
<EOL>|1655,1656
diverticulosis|1656,1670
,|1670,1671
<EOL>|1672,1673
h|1673,1674
/|1674,1675
o|1675,1676
colon|1677,1682
polyps|1683,1689
,|1689,1690
<EOL>|1691,1692
depression|1692,1702
,|1702,1703
<EOL>|1704,1705
s|1705,1706
/|1706,1707
p|1707,1708
right|1709,1714
CMC|1715,1718
joint|1719,1724
arthroplasty|1725,1737
,|1737,1738
<EOL>|1739,1740
b|1740,1741
/|1741,1742
l|1742,1743
rotator|1744,1751
cuff|1752,1756
repair|1757,1763
,|1763,1764
<EOL>|1765,1766
excision|1766,1774
right|1775,1780
_|1781,1782
_|1782,1783
_|1783,1784
digit|1785,1790
mass|1791,1795
,|1795,1796
<EOL>|1797,1798
CCY|1798,1801
w|1802,1803
/|1803,1804
stone|1804,1809
&|1810,1811
pancreatic|1812,1822
duct|1823,1827
exploration|1828,1839
(|1840,1841
_|1841,1842
_|1842,1843
_|1843,1844
)|1844,1845
,|1845,1846
<EOL>|1847,1848
hysterectomy|1848,1860
,|1860,1861
<EOL>|1862,1863
tonsillectomy|1863,1876
<EOL>|1877,1878
<EOL>|1878,1879
<EOL>|1880,1881
Social|1881,1887
History|1888,1895
:|1895,1896
<EOL>|1896,1897
_|1897,1898
_|1898,1899
_|1899,1900
<EOL>|1900,1901
Family|1901,1907
History|1908,1915
:|1915,1916
<EOL>|1916,1917
Mother|1917,1923
_|1924,1925
_|1925,1926
_|1926,1927
_|1928,1929
_|1929,1930
_|1930,1931
OVARIAN|1932,1939
CANCER|1940,1946
dx|1947,1949
age|1950,1953
_|1954,1955
_|1955,1956
_|1956,1957
<EOL>|1958,1959
Father|1959,1965
_|1966,1967
_|1967,1968
_|1968,1969
_|1970,1971
_|1971,1972
_|1972,1973
BRAIN|1974,1979
CANCER|1980,1986
<EOL>|1987,1988
PGM|1988,1991
OVARIAN|1992,1999
CANCER|2000,2006
<EOL>|2007,2008
Aunt|2008,2012
OVARIAN|2013,2020
CANCER|2021,2027
paternal|2028,2036
aunt|2037,2041
in|2042,2044
<EOL>|2045,2046
_|2047,2048
_|2048,2049
_|2049,2050
<EOL>|2051,2052
MGM|2052,2055
ENDOMETRIAL|2056,2067
CANCER|2068,2074
<EOL>|2075,2076
MGF|2076,2079
PROSTATE|2080,2088
CANCER|2089,2095
<EOL>|2096,2097
Brother|2097,2104
_|2105,2106
_|2106,2107
_|2107,2108
_|2109,2110
_|2110,2111
_|2111,2112
KIDNEY|2113,2119
CANCER|2120,2126
<EOL>|2127,2128
RENAL|2129,2134
FAILURE|2135,2142
<EOL>|2143,2144
CONGESTIVE|2145,2155
HEART|2156,2161
<EOL>|2162,2163
FAILURE|2164,2171
<EOL>|2172,2173
DIABETES|2174,2182
MELLITUS|2183,2191
<EOL>|2192,2193
TOBACCO|2194,2201
ABUSE|2202,2207
<EOL>|2208,2209
ALCOHOL|2210,2217
ABUSE|2218,2223
<EOL>|2224,2225
Sister|2225,2231
_|2232,2233
_|2233,2234
_|2234,2235
_|2236,2237
_|2237,2238
_|2238,2239
OVARIAN|2240,2247
CANCER|2248,2254
dx|2255,2257
age|2258,2261
_|2262,2263
_|2263,2264
_|2264,2265
<EOL>|2266,2267
Brother|2267,2274
_|2275,2276
_|2276,2277
_|2277,2278
THROAT|2279,2285
CANCER|2286,2292
dx|2293,2295
age|2296,2299
_|2300,2301
_|2301,2302
_|2302,2303
,|2303,2304
died|2305,2309
in|2310,2312
<EOL>|2313,2314
_|2315,2316
_|2316,2317
_|2317,2318
<EOL>|2319,2320
Sister|2320,2326
BRCA1|2327,2332
MUTATION|2333,2341
,|2341,2342
BREAST|2343,2349
CANCER|2350,2356
<EOL>|2357,2358
Daughter|2358,2366
Living|2367,2373
40|2374,2376
ABNORMAL|2377,2385
PAP|2386,2389
SMEAR|2390,2395
_|2396,2397
_|2397,2398
_|2398,2399
<EOL>|2399,2400
SUBSTANCE|2401,2410
ABUSE|2411,2416
<EOL>|2417,2418
Son|2418,2421
Died|2422,2426
_|2427,2428
_|2428,2429
_|2429,2430
SUBSTANCE|2431,2440
ABUSE|2441,2446
_|2447,2448
_|2448,2449
_|2449,2450
-|2451,2452
heroin|2453,2459
overdose|2460,2468
on|2469,2471
_|2472,2473
_|2473,2474
_|2474,2475
.|2475,2476
<EOL>|2476,2477
<EOL>|2478,2479
Physical|2479,2487
Exam|2488,2492
:|2492,2493
<EOL>|2493,2494
Physical|2494,2502
Exam|2503,2507
On|2508,2510
Admission|2511,2520
:|2520,2521
<EOL>|2521,2522
VITALS|2522,2528
:|2528,2529
_|2531,2532
_|2532,2533
_|2533,2534
1104|2535,2539
Temp|2540,2544
:|2544,2545
97.9|2546,2550
PO|2551,2553
BP|2554,2556
:|2556,2557
129|2558,2561
/|2561,2562
79|2562,2564
R|2565,2566
Lying|2567,2572
HR|2573,2575
:|2575,2576
82|2577,2579
<EOL>|2579,2580
RR|2580,2582
:|2582,2583
16|2584,2586
O2|2587,2589
sat|2590,2593
:|2593,2594
96|2595,2597
%|2597,2598
O2|2599,2601
delivery|2602,2610
:|2610,2611
Ra|2612,2614
<EOL>|2615,2616
<EOL>|2616,2617
General|2617,2624
:|2624,2625
Tearful|2626,2633
,|2633,2634
expressing|2635,2645
right|2646,2651
back|2652,2656
and|2657,2660
leg|2661,2664
pain|2665,2669
with|2670,2674
spasms|2675,2681
<EOL>|2682,2683
<EOL>|2683,2684
<EOL>|2684,2685
Chest|2685,2690
:|2690,2691
L|2692,2693
breast|2694,2700
incisions|2701,2710
well|2711,2715
healed|2716,2722
.|2722,2723
S|2724,2725
/|2725,2726
p|2726,2727
L|2728,2729
axilla|2730,2736
surgical|2737,2745
<EOL>|2745,2746
drain|2746,2751
removal|2752,2759
.|2759,2760
<EOL>|2760,2761
CV|2761,2763
:|2763,2764
Regular|2765,2772
rate|2773,2777
and|2778,2781
rhythm|2782,2788
,|2788,2789
normal|2790,2796
S1|2797,2799
+|2800,2801
S2|2802,2804
,|2804,2805
no|2806,2808
murmurs|2809,2816
<EOL>|2816,2817
Lungs|2817,2822
:|2822,2823
Clear|2824,2829
to|2830,2832
auscultation|2833,2845
bilaterally|2846,2857
,|2857,2858
no|2859,2861
wheezes|2862,2869
or|2870,2872
crackles|2873,2881
<EOL>|2881,2882
Abdomen|2882,2889
:|2889,2890
Soft|2891,2895
,|2895,2896
non-tender|2897,2907
,|2907,2908
non-distended|2909,2922
,|2922,2923
bowel|2924,2929
sounds|2930,2936
present|2937,2944
<EOL>|2944,2945
Ext|2945,2948
:|2948,2949
Warm|2950,2954
,|2954,2955
well|2956,2960
perfused|2961,2969
,|2969,2970
right|2971,2976
lower|2977,2982
extremity|2983,2992
is|2993,2995
tender|2996,3002
to|3003,3005
<EOL>|3005,3006
palpation|3006,3015
and|3016,3019
movement|3020,3028
limited|3029,3036
by|3037,3039
pain|3040,3044
.|3044,3045
Swelling|3046,3054
of|3055,3057
RLE|3058,3061
>|3062,3063
LLE|3064,3067
.|3067,3068
<EOL>|3068,3069
Palpable|3069,3077
2|3078,3079
+|3079,3080
_|3081,3082
_|3082,3083
_|3083,3084
pulses|3085,3091
bilaterally|3092,3103
.|3103,3104
<EOL>|3104,3105
Skin|3105,3109
:|3109,3110
Warm|3111,3115
,|3115,3116
dry|3117,3120
,|3120,3121
varicose|3122,3130
veins|3131,3136
noted|3137,3142
in|3143,3145
lower|3146,3151
extremities|3152,3163
.|3163,3164
<EOL>|3165,3166
Neuro|3166,3171
:|3171,3172
Grossly|3173,3180
oriented|3181,3189
<EOL>|3189,3190
MSK|3190,3193
exam|3194,3198
:|3198,3199
Right|3200,3205
SI|3206,3208
Joint|3209,3214
tenderness|3215,3225
.|3225,3226
Radicular|3227,3236
pain|3237,3241
worsened|3242,3250
<EOL>|3251,3252
with|3252,3256
<EOL>|3256,3257
back|3257,3261
flexion|3262,3269
and|3270,3273
relieved|3274,3282
with|3283,3287
extension|3288,3297
.|3297,3298
_|3299,3300
_|3300,3301
_|3301,3302
strength|3303,3311
<EOL>|3311,3312
bilaterally|3312,3323
w|3324,3325
/|3325,3326
hip|3327,3330
flexion|3331,3338
and|3339,3342
extension|3343,3352
,|3352,3353
knee|3354,3358
flexion|3359,3366
and|3367,3370
<EOL>|3370,3371
extension|3371,3380
,|3380,3381
foot|3382,3386
plantar|3387,3394
and|3395,3398
dorsiflexion|3399,3411
,|3411,3412
sensation|3413,3422
in|3423,3425
tact|3426,3430
<EOL>|3430,3431
bilaterally|3431,3442
<EOL>|3443,3444
<EOL>|3444,3445
_|3445,3446
_|3446,3447
_|3447,3448
Ortho|3449,3454
Spine|3455,3460
Exam|3461,3465
<EOL>|3465,3466
<EOL>|3466,3467
PE|3467,3469
:|3469,3470
<EOL>|3471,3472
VS|3472,3474
<EOL>|3474,3475
_|3475,3476
_|3476,3477
_|3477,3478
_|3479,3480
_|3480,3481
_|3481,3482
Temp|3483,3487
:|3487,3488
98.7|3489,3493
PO|3494,3496
BP|3497,3499
:|3499,3500
135|3501,3504
/|3504,3505
66|3505,3507
R|3508,3509
Lying|3510,3515
HR|3516,3518
:|3518,3519
99|3520,3522
RR|3523,3525
:|3525,3526
18|3527,3529
O2|3530,3532
<EOL>|3532,3533
sat|3533,3536
:|3536,3537
94|3538,3540
%|3540,3541
O2|3542,3544
delivery|3545,3553
:|3553,3554
Ra|3555,3557
<EOL>|3558,3559
_|3559,3560
_|3560,3561
_|3561,3562
_|3563,3564
_|3564,3565
_|3565,3566
Temp|3567,3571
:|3571,3572
98.7|3573,3577
PO|3578,3580
BP|3581,3583
:|3583,3584
135|3585,3588
/|3588,3589
66|3589,3591
R|3592,3593
Lying|3594,3599
HR|3600,3602
:|3602,3603
99|3604,3606
RR|3607,3609
:|3609,3610
18|3611,3613
O2|3614,3616
<EOL>|3616,3617
sat|3617,3620
:|3620,3621
94|3622,3624
%|3624,3625
O2|3626,3628
delivery|3629,3637
:|3637,3638
Ra|3639,3641
<EOL>|3642,3643
<EOL>|3643,3644
NAD|3644,3647
,|3647,3648
A|3649,3650
&|3650,3651
Ox4|3651,3654
<EOL>|3654,3655
nl|3655,3657
resp|3658,3662
effort|3663,3669
<EOL>|3669,3670
RRR|3670,3673
<EOL>|3673,3674
<EOL>|3676,3677
Sensory|3677,3684
:|3684,3685
<EOL>|3685,3686
UE|3686,3688
<EOL>|3689,3690
C5|3697,3699
C6|3708,3710
C7|3721,3723
C8|3731,3733
T1|3744,3746
<EOL>|3746,3747
(|3752,3753
lat|3753,3756
arm|3757,3760
)|3760,3761
(|3763,3764
thumb|3764,3769
)|3769,3770
(|3775,3776
mid|3776,3779
fing|3780,3784
)|3784,3785
(|3786,3787
sm|3787,3789
finger|3790,3796
)|3796,3797
(|3799,3800
med|3800,3803
arm|3804,3807
)|3807,3808
<EOL>|3808,3809
R|3809,3810
SILT|3815,3819
SILT|3826,3830
SILT|3838,3842
SILT|3850,3854
SILT|3863,3867
<EOL>|3867,3868
L|3868,3869
SILT|3874,3878
SILT|3885,3889
SILT|3897,3901
SILT|3909,3913
SILT|3922,3926
<EOL>|3926,3927
<EOL>|3927,3928
T2|3928,3930
-|3930,3931
L1|3931,3933
(|3934,3935
Trunk|3935,3940
)|3940,3941
<EOL>|3942,3943
SILT|3950,3954
<EOL>|3954,3955
<EOL>|3955,3956
_|3956,3957
_|3957,3958
_|3958,3959
<EOL>|3963,3964
L2|3969,3971
L3|3976,3978
L4|3984,3986
L5|3995,3997
S1|4005,4007
S2|4017,4019
<EOL>|4019,4020
(|4023,4024
Groin|4024,4029
)|4029,4030
(|4031,4032
Knee|4032,4036
)|4036,4037
(|4038,4039
Med|4039,4042
Calf|4043,4047
)|4047,4048
(|4049,4050
Grt|4050,4053
Toe|4054,4057
)|4057,4058
(|4059,4060
Sm|4060,4062
Toe|4063,4066
)|4066,4067
(|4068,4069
Post|4069,4073
Thigh|4074,4079
)|4079,4080
<EOL>|4080,4081
R|4081,4082
SILT|4086,4090
SILT|4093,4097
SILT|4101,4105
SILT|4112,4116
SILT|4121,4125
SILT|4132,4136
<EOL>|4137,4138
L|4138,4139
SILT|4143,4147
SILT|4150,4154
SILT|4158,4162
SILT|4169,4173
SILT|4178,4182
SILT|4189,4193
<EOL>|4194,4195
<EOL>|4195,4196
Motor|4196,4201
:|4201,4202
<EOL>|4202,4203
UE|4203,4205
Dlt|4208,4211
(|4211,4212
C5|4212,4214
)|4214,4215
Bic|4216,4219
(|4219,4220
C6|4220,4222
)|4222,4223
WE|4224,4226
(|4226,4227
C6|4227,4229
)|4229,4230
Tri|4231,4234
(|4234,4235
C7|4235,4237
)|4237,4238
WF|4239,4241
(|4241,4242
C7|4242,4244
)|4244,4245
FF|4246,4248
(|4248,4249
C8|4249,4251
)|4251,4252
FinAbd|4252,4258
(|4258,4259
T1|4259,4261
)|4261,4262
<EOL>|4262,4263
R|4263,4264
5|4270,4271
5|4278,4279
5|4286,4287
5|4293,4294
5|4301,4302
5|4308,4309
5|4314,4315
<EOL>|4315,4316
L|4316,4317
5|4323,4324
5|4331,4332
5|4339,4340
5|4346,4347
5|4354,4355
5|4361,4362
5|4367,4368
<EOL>|4368,4369
<EOL>|4369,4370
_|4370,4371
_|4371,4372
_|4372,4373
Flex|4375,4379
(|4379,4380
L1|4380,4382
)|4382,4383
Add|4384,4387
(|4387,4388
L2|4388,4390
)|4390,4391
Quad|4392,4396
(|4396,4397
L3|4397,4399
)|4399,4400
TA|4402,4404
(|4404,4405
L4|4405,4407
)|4407,4408
_|4409,4410
_|4410,4411
_|4411,4412
_|4413,4414
_|4414,4415
_|4415,4416
<EOL>|4416,4417
R|4417,4418
5|4424,4425
5|4432,4433
5|4440,4441
5|4450,4451
5|4457,4458
5|4464,4465
5|4474,4475
<EOL>|4481,4482
L|4482,4483
5|4489,4490
5|4497,4498
5|4505,4506
5|4515,4516
5|4522,4523
5|4529,4530
5|4539,4540
<EOL>|4540,4541
<EOL>|4541,4542
Reflexes|4542,4550
<EOL>|4551,4552
Bic|4556,4559
(|4559,4560
C4|4560,4562
-|4562,4563
5|4563,4564
)|4564,4565
BR|4567,4569
(|4569,4570
C5|4570,4572
-|4572,4573
6|4573,4574
)|4574,4575
Tri|4577,4580
(|4580,4581
C6|4581,4583
-|4583,4584
7|4584,4585
)|4585,4586
Pat|4588,4591
(|4591,4592
L3|4592,4594
-|4594,4595
4|4595,4596
)|4596,4597
Ach|4599,4602
(|4602,4603
L5|4603,4605
-|4605,4606
S1|4606,4608
)|4608,4609
<EOL>|4609,4610
R|4610,4611
2|4617,4618
2|4628,4629
2|4638,4639
2|4649,4650
2|4661,4662
<EOL>|4662,4663
L|4663,4664
2|4670,4671
2|4681,4682
2|4691,4692
2|4702,4703
2|4714,4715
<EOL>|4715,4716
<EOL>|4730,4731
_|4731,4732
_|4732,4733
_|4733,4734
:|4734,4735
Negative|4736,4744
<EOL>|4744,4745
Babinski|4745,4753
:|4753,4754
Downgoing|4756,4765
<EOL>|4765,4766
Clonus|4766,4772
:|4772,4773
No|4774,4776
beats|4777,4782
<EOL>|4782,4783
<EOL>|4783,4784
<EOL>|4785,4786
Pertinent|4786,4795
Results|4796,4803
:|4803,4804
<EOL>|4804,4805
IMAGING|4805,4812
:|4812,4813
<EOL>|4813,4814
MR|4814,4816
THORACIC|4817,4825
SPINE|4826,4831
W|4832,4833
/|4833,4834
O|4834,4835
CONTRAST|4836,4844
;|4844,4845
MR|4846,4848
_|4849,4850
_|4850,4851
_|4851,4852
SPINE|4853,4858
W|4859,4860
/|4860,4861
O|4861,4862
CONTRAST|4863,4871
_|4872,4873
_|4873,4874
_|4874,4875
<EOL>|4875,4876
IMPRESSION|4876,4886
:|4886,4887
<EOL>|4887,4888
1.|4888,4890
Severe|4891,4897
central|4898,4905
canal|4906,4911
narrowing|4912,4921
at|4922,4924
L4|4925,4927
-|4927,4928
5|4928,4929
level|4930,4935
from|4936,4940
<EOL>|4941,4942
degenerative|4942,4954
changes|4955,4962
.|4962,4963
<EOL>|4963,4964
2.|4964,4966
Large|4967,4972
right|4973,4978
paramedian|4979,4989
,|4989,4990
superior|4991,4999
disc|5000,5004
extrusion|5005,5014
L4|5015,5017
-|5017,5018
5|5018,5019
level|5020,5025
,|5025,5026
<EOL>|5027,5028
extends|5028,5035
into|5036,5040
<EOL>|5040,5041
right|5041,5046
L4|5047,5049
lateral|5050,5057
recess|5058,5064
,|5064,5065
mass|5066,5070
effect|5071,5077
on|5078,5080
exiting|5081,5088
right|5089,5094
L4|5095,5097
,|5097,5098
<EOL>|5099,5100
traversing|5100,5110
L5|5111,5113
<EOL>|5113,5114
nerves|5114,5120
,|5120,5121
severe|5122,5128
right|5129,5134
L4|5135,5137
-|5137,5138
5|5138,5139
foraminal|5140,5149
narrowing|5150,5159
.|5159,5160
.|5160,5161
<EOL>|5161,5162
3|5162,5163
.|5163,5164
Advanced|5165,5173
degenerative|5174,5186
changes|5187,5194
lumbar|5195,5201
spine|5202,5207
.|5207,5208
<EOL>|5208,5209
4.|5209,5211
Moderate|5212,5220
central|5221,5228
canal|5229,5234
narrowing|5235,5244
L2|5245,5247
-|5247,5248
L3|5248,5250
,|5250,5251
moderate|5252,5260
to|5261,5263
severe|5264,5270
at|5271,5273
<EOL>|5274,5275
L3|5275,5277
-|5277,5278
L4|5278,5280
levels|5281,5287
.|5287,5288
<EOL>|5288,5289
5.|5289,5291
Multilevel|5292,5302
significant|5303,5314
foraminal|5315,5324
narrowing|5325,5334
lumbar|5335,5341
spine|5342,5347
,|5347,5348
as|5349,5351
<EOL>|5352,5353
above|5353,5358
.|5358,5359
<EOL>|5359,5360
6.|5360,5362
Degenerative|5363,5375
changes|5376,5383
thoracic|5384,5392
spine|5393,5398
,|5398,5399
mild|5400,5404
-|5404,5405
to|5405,5407
-|5407,5408
moderate|5408,5416
central|5417,5424
<EOL>|5425,5426
canal|5426,5431
<EOL>|5431,5432
narrowing|5432,5441
,|5441,5442
foraminal|5443,5452
narrowing|5453,5462
.|5462,5463
<EOL>|5463,5464
<EOL>|5464,5465
CT|5465,5467
ABD|5468,5471
&|5472,5473
PELVIS|5474,5480
WITH|5481,5485
CONTRAST|5486,5494
_|5495,5496
_|5496,5497
_|5497,5498
<EOL>|5498,5499
IMPRESSION|5499,5509
:|5509,5510
<EOL>|5510,5511
<EOL>|5512,5513
1|5513,5514
.|5514,5515
No|5516,5518
acute|5519,5524
CT|5525,5527
findings|5528,5536
in|5537,5539
the|5540,5543
abdomen|5544,5551
or|5552,5554
pelvis|5555,5561
to|5562,5564
correlate|5565,5574
<EOL>|5575,5576
with|5576,5580
patient|5581,5588
's|5588,5590
<EOL>|5590,5591
reported|5591,5599
symptoms|5600,5608
.|5608,5609
Specifically|5611,5623
,|5623,5624
no|5625,5627
evidence|5628,5636
of|5637,5639
obstructive|5640,5651
<EOL>|5652,5653
renal|5653,5658
stone|5659,5664
or|5665,5667
<EOL>|5667,5668
pyelonephritis|5668,5682
.|5682,5683
<EOL>|5683,5684
2.|5684,5686
Sigmoid|5687,5694
diverticulosis|5695,5709
without|5712,5719
evidence|5720,5728
of|5729,5731
acute|5732,5737
<EOL>|5738,5739
diverticulitis|5739,5753
.|5753,5754
<EOL>|5754,5755
<EOL>|5755,5756
Admission|5756,5765
Labs|5766,5770
:|5770,5771
<EOL>|5771,5772
_|5772,5773
_|5773,5774
_|5774,5775
12|5776,5778
:|5778,5779
49PM|5779,5783
BLOOD|5784,5789
WBC|5790,5793
-|5793,5794
6.3|5794,5797
RBC|5798,5801
-|5801,5802
3|5802,5803
.|5803,5804
97|5804,5806
Hgb|5807,5810
-|5810,5811
11.9|5811,5815
Hct|5816,5819
-|5819,5820
37.2|5820,5824
MCV|5825,5828
-|5828,5829
94|5829,5831
<EOL>|5832,5833
MCH|5833,5836
-|5836,5837
30.0|5837,5841
MCHC|5842,5846
-|5846,5847
32.0|5847,5851
RDW|5852,5855
-|5855,5856
14.3|5856,5860
RDWSD|5861,5866
-|5866,5867
49|5867,5869
.|5869,5870
1|5870,5871
*|5871,5872
Plt|5873,5876
_|5877,5878
_|5878,5879
_|5879,5880
<EOL>|5880,5881
_|5881,5882
_|5882,5883
_|5883,5884
12|5885,5887
:|5887,5888
49PM|5888,5892
BLOOD|5893,5898
_|5899,5900
_|5900,5901
_|5901,5902
PTT|5903,5906
-|5906,5907
34.3|5907,5911
_|5912,5913
_|5913,5914
_|5914,5915
<EOL>|5915,5916
_|5916,5917
_|5917,5918
_|5918,5919
12|5920,5922
:|5922,5923
49PM|5923,5927
BLOOD|5928,5933
Glucose|5934,5941
-|5941,5942
117|5942,5945
*|5945,5946
UreaN|5947,5952
-|5952,5953
11|5953,5955
Creat|5956,5961
-|5961,5962
0.8|5962,5965
Na|5966,5968
-|5968,5969
143|5969,5972
<EOL>|5973,5974
K|5974,5975
-|5975,5976
4.3|5976,5979
Cl|5980,5982
-|5982,5983
106|5983,5986
HCO3|5987,5991
-|5991,5992
26|5992,5994
AnGap|5995,6000
-|6000,6001
11|6001,6003
<EOL>|6003,6004
<EOL>|6004,6005
_|6005,6006
_|6006,6007
_|6007,6008
10|6009,6011
:|6011,6012
06AM|6012,6016
BLOOD|6017,6022
WBC|6023,6026
-|6026,6027
5.8|6027,6030
RBC|6031,6034
-|6034,6035
2|6035,6036
.|6036,6037
81|6037,6039
*|6039,6040
Hgb|6041,6044
-|6044,6045
8|6045,6046
.|6046,6047
5|6047,6048
*|6048,6049
Hct|6050,6053
-|6053,6054
26|6054,6056
.|6056,6057
1|6057,6058
*|6058,6059
<EOL>|6060,6061
MCV|6061,6064
-|6064,6065
93|6065,6067
MCH|6068,6071
-|6071,6072
30.2|6072,6076
MCHC|6077,6081
-|6081,6082
32.6|6082,6086
RDW|6087,6090
-|6090,6091
14.0|6091,6095
RDWSD|6096,6101
-|6101,6102
47|6102,6104
.|6104,6105
6|6105,6106
*|6106,6107
Plt|6108,6111
_|6112,6113
_|6113,6114
_|6114,6115
<EOL>|6115,6116
_|6116,6117
_|6117,6118
_|6118,6119
05|6120,6122
:|6122,6123
53AM|6123,6127
BLOOD|6128,6133
WBC|6134,6137
-|6137,6138
6.6|6138,6141
RBC|6142,6145
-|6145,6146
2|6146,6147
.|6147,6148
88|6148,6150
*|6150,6151
Hgb|6152,6155
-|6155,6156
8|6156,6157
.|6157,6158
9|6158,6159
*|6159,6160
Hct|6161,6164
-|6164,6165
27|6165,6167
.|6167,6168
6|6168,6169
*|6169,6170
<EOL>|6171,6172
MCV|6172,6175
-|6175,6176
96|6176,6178
MCH|6179,6182
-|6182,6183
30.9|6183,6187
MCHC|6188,6192
-|6192,6193
32.2|6193,6197
RDW|6198,6201
-|6201,6202
14.4|6202,6206
RDWSD|6207,6212
-|6212,6213
50|6213,6215
.|6215,6216
4|6216,6217
*|6217,6218
Plt|6219,6222
_|6223,6224
_|6224,6225
_|6225,6226
<EOL>|6226,6227
_|6227,6228
_|6228,6229
_|6229,6230
04|6231,6233
:|6233,6234
30AM|6234,6238
BLOOD|6239,6244
WBC|6245,6248
-|6248,6249
6.9|6249,6252
RBC|6253,6256
-|6256,6257
3|6257,6258
.|6258,6259
40|6259,6261
*|6261,6262
Hgb|6263,6266
-|6266,6267
10|6267,6269
.|6269,6270
2|6270,6271
*|6271,6272
Hct|6273,6276
-|6276,6277
32|6277,6279
.|6279,6280
6|6280,6281
*|6281,6282
<EOL>|6283,6284
MCV|6284,6287
-|6287,6288
96|6288,6290
MCH|6291,6294
-|6294,6295
30.0|6295,6299
MCHC|6300,6304
-|6304,6305
31|6305,6307
.|6307,6308
3|6308,6309
*|6309,6310
RDW|6311,6314
-|6314,6315
14.4|6315,6319
RDWSD|6320,6325
-|6325,6326
50|6326,6328
.|6328,6329
3|6329,6330
*|6330,6331
Plt|6332,6335
_|6336,6337
_|6337,6338
_|6338,6339
<EOL>|6339,6340
_|6340,6341
_|6341,6342
_|6342,6343
10|6344,6346
:|6346,6347
06AM|6347,6351
BLOOD|6352,6357
Plt|6358,6361
_|6362,6363
_|6363,6364
_|6364,6365
<EOL>|6365,6366
_|6366,6367
_|6367,6368
_|6368,6369
04|6370,6372
:|6372,6373
30AM|6373,6377
BLOOD|6378,6383
Glucose|6384,6391
-|6391,6392
107|6392,6395
*|6395,6396
UreaN|6397,6402
-|6402,6403
10|6403,6405
Creat|6406,6411
-|6411,6412
0.7|6412,6415
Na|6416,6418
-|6418,6419
142|6419,6422
<EOL>|6423,6424
K|6424,6425
-|6425,6426
4.8|6426,6429
Cl|6430,6432
-|6432,6433
105|6433,6436
HCO3|6437,6441
-|6441,6442
25|6442,6444
AnGap|6445,6450
-|6450,6451
12|6451,6453
<EOL>|6453,6454
_|6454,6455
_|6455,6456
_|6456,6457
04|6458,6460
:|6460,6461
30AM|6461,6465
BLOOD|6466,6471
Glucose|6472,6479
-|6479,6480
147|6480,6483
*|6483,6484
UreaN|6485,6490
-|6490,6491
12|6491,6493
Creat|6494,6499
-|6499,6500
0.9|6500,6503
Na|6504,6506
-|6506,6507
142|6507,6510
<EOL>|6511,6512
K|6512,6513
-|6513,6514
4.8|6514,6517
Cl|6518,6520
-|6520,6521
99|6521,6523
HCO3|6524,6528
-|6528,6529
28|6529,6531
AnGap|6532,6537
-|6537,6538
15|6538,6540
<EOL>|6540,6541
_|6541,6542
_|6542,6543
_|6543,6544
08|6545,6547
:|6547,6548
49AM|6548,6552
BLOOD|6553,6558
Glucose|6559,6566
-|6566,6567
128|6567,6570
*|6570,6571
UreaN|6572,6577
-|6577,6578
10|6578,6580
Creat|6581,6586
-|6586,6587
0.9|6587,6590
Na|6591,6593
-|6593,6594
141|6594,6597
<EOL>|6598,6599
K|6599,6600
-|6600,6601
4.3|6601,6604
Cl|6605,6607
-|6607,6608
102|6608,6611
HCO3|6612,6616
-|6616,6617
28|6617,6619
AnGap|6620,6625
-|6625,6626
11|6626,6628
<EOL>|6628,6629
_|6629,6630
_|6630,6631
_|6631,6632
04|6633,6635
:|6635,6636
30AM|6636,6640
BLOOD|6641,6646
Calcium|6647,6654
-|6654,6655
8|6655,6656
.|6656,6657
2|6657,6658
*|6658,6659
Phos|6660,6664
-|6664,6665
2.9|6665,6668
Mg|6669,6671
-|6671,6672
2.0|6672,6675
<EOL>|6675,6676
_|6676,6677
_|6677,6678
_|6678,6679
08|6680,6682
:|6682,6683
49AM|6683,6687
BLOOD|6688,6693
Calcium|6694,6701
-|6701,6702
9.5|6702,6705
Phos|6706,6710
-|6710,6711
4.3|6711,6714
Mg|6715,6717
-|6717,6718
2.1|6718,6721
<EOL>|6721,6722
_|6722,6723
_|6723,6724
_|6724,6725
04|6726,6728
:|6728,6729
30AM|6729,6733
BLOOD|6734,6739
Calcium|6740,6747
-|6747,6748
8.8|6748,6751
Phos|6752,6756
-|6756,6757
4|6757,6758
.|6758,6759
6|6759,6760
*|6760,6761
Mg|6762,6764
-|6764,6765
2.1|6765,6768
<EOL>|6768,6769
<EOL>|6770,6771
Brief|6771,6776
Hospital|6777,6785
Course|6786,6792
:|6792,6793
<EOL>|6793,6794
Initial|6794,6801
Admission|6802,6811
:|6811,6812
<EOL>|6813,6814
ACTIVE|6814,6820
ISSUES|6821,6827
:|6827,6828
<EOL>|6828,6829
=|6829,6830
=|6830,6831
=|6831,6832
=|6832,6833
=|6833,6834
=|6834,6835
=|6835,6836
=|6836,6837
=|6837,6838
=|6838,6839
=|6839,6840
=|6840,6841
=|6841,6842
=|6842,6843
=|6843,6844
=|6844,6845
=|6845,6846
=|6846,6847
<EOL>|6847,6848
#|6848,6849
R|6850,6851
Low|6852,6855
Back|6856,6860
pain|6861,6865
and|6866,6869
Leg|6870,6873
Pain|6874,6878
<EOL>|6878,6879
#|6879,6880
Radiculopathy|6881,6894
<EOL>|6894,6895
Patient|6895,6902
presents|6903,6911
with|6912,6916
severe|6917,6923
right|6924,6929
lower|6930,6935
back|6936,6940
pain|6941,6945
with|6946,6950
<EOL>|6951,6952
prominent|6952,6961
<EOL>|6961,6962
lancinating|6962,6973
component|6974,6983
.|6983,6984
CT|6985,6987
A|6988,6989
/|6989,6990
P|6990,6991
with|6992,6996
no|6997,6999
evidence|7000,7008
of|7009,7011
visceral|7012,7020
<EOL>|7020,7021
pathology|7021,7030
or|7031,7033
nephrolithiasis|7034,7049
.|7049,7050
MRI|7051,7054
L|7055,7056
spine|7057,7062
with|7063,7067
significant|7068,7079
disc|7080,7084
<EOL>|7084,7085
bulge|7085,7090
at|7091,7093
L2|7094,7096
-|7096,7097
L3|7097,7099
and|7100,7103
L3|7104,7106
-|7106,7107
4|7107,7108
cause|7109,7114
severe|7115,7121
narrowing|7122,7131
of|7132,7134
the|7135,7138
spinal|7139,7145
<EOL>|7145,7146
canal|7146,7151
and|7152,7155
extrusion|7156,7165
at|7166,7168
L4|7169,7171
-|7171,7172
5|7172,7173
with|7174,7178
significant|7179,7190
L4|7191,7193
nerve|7194,7199
root|7200,7204
<EOL>|7204,7205
compression|7205,7216
,|7216,7217
likely|7218,7224
the|7225,7228
cause|7229,7234
of|7235,7237
patient|7238,7245
's|7245,7247
pain|7248,7252
.|7252,7253
She|7254,7257
was|7258,7261
<EOL>|7262,7263
recently|7263,7271
<EOL>|7271,7272
admitted|7272,7280
with|7281,7285
right|7286,7291
leg|7292,7295
pain|7296,7300
,|7300,7301
with|7302,7306
exam|7307,7311
notable|7312,7319
for|7320,7323
trochanteric|7324,7336
<EOL>|7336,7337
bursitis|7337,7345
,|7345,7346
now|7347,7350
s|7351,7352
/|7352,7353
p|7353,7354
injection|7355,7364
of|7365,7367
corticosteroid|7368,7382
.|7382,7383
Currently|7384,7393
<EOL>|7393,7394
neruovascularly|7394,7409
intact|7410,7416
,|7416,7417
with|7418,7422
no|7423,7425
evidence|7426,7434
of|7435,7437
cord|7438,7442
compression|7443,7454
by|7455,7457
<EOL>|7457,7458
history|7458,7465
or|7466,7468
on|7469,7471
exam|7472,7476
.|7476,7477
Per|7478,7481
ortho|7482,7487
spine|7488,7493
,|7493,7494
would|7495,7500
benefit|7501,7508
from|7509,7513
<EOL>|7513,7514
decompression|7514,7527
.|7527,7528
She|7529,7532
had|7533,7536
a|7537,7538
DECOMPRESSION|7539,7552
L2|7553,7555
-|7555,7556
S1|7556,7558
,|7558,7559
FUSION|7560,7566
L4|7567,7569
-|7569,7570
L5|7570,7572
,|7572,7573
<EOL>|7574,7575
DURAPLASTY|7575,7585
on|7586,7588
_|7589,7590
_|7590,7591
_|7591,7592
w|7593,7594
/|7594,7595
ortho-spine|7596,7607
once|7608,7612
her|7613,7616
INR|7617,7620
was|7621,7624
1.2|7625,7628
.|7628,7629
She|7630,7633
<EOL>|7634,7635
was|7635,7638
started|7639,7646
on|7647,7649
a|7650,7651
heparin|7652,7659
bridge|7660,7666
on|7667,7669
_|7670,7671
_|7671,7672
_|7672,7673
when|7674,7678
her|7679,7682
INR|7683,7686
dropped|7687,7694
<EOL>|7695,7696
below|7696,7701
2.0|7702,7705
and|7706,7709
transitioned|7710,7722
to|7723,7725
lovenox|7726,7733
bridge|7734,7740
to|7741,7743
coumadin|7744,7752
on|7753,7755
<EOL>|7756,7757
_|7757,7758
_|7758,7759
_|7759,7760
<EOL>|7760,7761
<EOL>|7761,7762
#|7762,7763
Dysuria|7764,7771
(|7772,7773
resolved|7773,7781
)|7781,7782
<EOL>|7782,7783
#|7783,7784
UTI|7785,7788
<EOL>|7788,7789
States|7789,7795
she|7796,7799
has|7800,7803
been|7804,7808
having|7809,7815
burning|7816,7823
pain|7824,7828
with|7829,7833
urination|7834,7843
recently|7844,7852
.|7852,7853
<EOL>|7853,7854
She|7854,7857
also|7858,7862
feels|7863,7868
that|7869,7873
she|7874,7877
needs|7878,7883
to|7884,7886
push|7887,7891
on|7892,7894
her|7895,7898
abdomen|7899,7906
to|7907,7909
urinate|7910,7917
.|7917,7918
<EOL>|7918,7919
Most|7919,7923
concerning|7924,7934
for|7935,7938
UTI|7939,7942
.|7942,7943
UA|7944,7946
demonstrating|7947,7960
large|7961,7966
leukocytes|7967,7977
and|7978,7981
8|7982,7983
<EOL>|7983,7984
WBC|7984,7987
.|7987,7988
However|7989,7996
,|7996,7997
urine|7998,8003
culture|8004,8011
showing|8012,8019
mixed|8020,8025
bacterial|8026,8035
flora|8036,8041
<EOL>|8041,8042
consistent|8042,8052
with|8053,8057
contamination|8058,8071
.|8071,8072
Will|8073,8077
treat|8078,8083
given|8084,8089
symptoms|8090,8098
.|8098,8099
<EOL>|8099,8100
Abdominal|8100,8109
pain|8110,8114
could|8115,8120
also|8121,8125
be|8126,8128
from|8129,8133
constipation|8134,8146
in|8147,8149
the|8150,8153
setting|8154,8161
of|8162,8164
<EOL>|8164,8165
opioid|8165,8171
use|8172,8175
.|8175,8176
Reports|8177,8184
resolution|8185,8195
of|8196,8198
symptoms|8199,8207
on|8208,8210
_|8211,8212
_|8212,8213
_|8213,8214
.|8214,8215
Was|8216,8219
treated|8220,8227
<EOL>|8228,8229
with|8229,8233
bactrim|8234,8241
DS|8242,8244
BID|8245,8248
for|8249,8252
3|8253,8254
days|8255,8259
starting|8260,8268
_|8269,8270
_|8270,8271
_|8271,8272
and|8273,8276
ending|8277,8283
_|8284,8285
_|8285,8286
_|8286,8287
.|8287,8288
<EOL>|8289,8290
<EOL>|8290,8291
CHRONIC|8291,8298
ISSUES|8299,8305
:|8305,8306
<EOL>|8306,8307
=|8307,8308
=|8308,8309
=|8309,8310
=|8310,8311
=|8311,8312
=|8312,8313
=|8313,8314
=|8314,8315
=|8315,8316
=|8316,8317
=|8317,8318
=|8318,8319
=|8319,8320
=|8320,8321
=|8321,8322
=|8322,8323
=|8323,8324
=|8324,8325
=|8325,8326
<EOL>|8326,8327
#|8327,8328
History|8329,8336
of|8337,8339
DVT|8340,8343
/|8343,8344
PE|8344,8346
<EOL>|8346,8347
#|8347,8348
Antiphospholipid|8349,8365
antibody|8366,8374
syndrome|8375,8383
:|8383,8384
<EOL>|8384,8385
Lupus|8385,8390
anticoagulant|8391,8404
positive|8405,8413
in|8414,8416
_|8417,8418
_|8418,8419
_|8419,8420
.|8420,8421
Had|8422,8425
bilateral|8426,8435
PE|8436,8438
in|8439,8441
_|8442,8443
_|8443,8444
_|8444,8445
.|8445,8446
<EOL>|8446,8447
She|8447,8450
has|8451,8454
been|8455,8459
taking|8460,8466
her|8467,8470
home|8471,8475
dose|8476,8480
of|8481,8483
warfarin|8484,8492
(|8493,8494
7.5|8494,8497
mg|8498,8500
_|8501,8502
_|8502,8503
_|8503,8504
and|8505,8508
<EOL>|8509,8510
5|8510,8511
<EOL>|8511,8512
mg|8512,8514
other|8515,8520
days|8521,8525
)|8525,8526
.|8526,8527
Warfarin|8528,8536
held|8537,8541
on|8542,8544
admission|8545,8554
for|8555,8558
procedure|8559,8568
with|8569,8573
<EOL>|8574,8575
heparin|8575,8582
drip|8583,8587
until|8588,8593
procedure|8594,8603
.|8603,8604
<EOL>|8605,8606
<EOL>|8606,8607
#|8607,8608
AAA|8609,8612
<EOL>|8612,8613
Has|8613,8616
a|8617,8618
reported|8619,8627
history|8628,8635
of|8636,8638
AAA|8639,8642
in|8643,8645
chart|8646,8651
,|8651,8652
but|8653,8656
does|8657,8661
not|8662,8665
follow|8666,8672
up|8673,8675
<EOL>|8675,8676
with|8676,8680
anyone|8681,8687
for|8688,8691
surveillance|8692,8704
and|8705,8708
CT|8709,8711
abd|8712,8715
/|8715,8716
pelvis|8716,8722
did|8723,8726
not|8727,8730
show|8731,8735
an|8736,8738
<EOL>|8738,8739
abdominal|8739,8748
aortic|8749,8755
aneurysm|8756,8764
.|8764,8765
<EOL>|8765,8766
<EOL>|8766,8767
#|8767,8768
Vitamin|8769,8776
D|8777,8778
deficiency|8779,8789
:|8789,8790
<EOL>|8790,8791
-|8791,8792
Continued|8793,8802
Vitamin|8803,8810
D|8811,8812
_|8813,8814
_|8814,8815
_|8815,8816
daily|8817,8822
<EOL>|8822,8823
<EOL>|8823,8824
#|8824,8825
OSA|8826,8829
<EOL>|8829,8830
-|8830,8831
Remained|8832,8840
on|8841,8843
CPAP|8844,8848
<EOL>|8849,8850
<EOL>|8850,8851
#|8851,8852
Other|8852,8857
Home|8858,8862
Meds|8863,8867
:|8867,8868
<EOL>|8868,8869
-|8869,8870
Continued|8871,8880
omeprazole|8881,8891
20mg|8892,8896
BID|8897,8900
for|8901,8904
GERD|8905,8909
<EOL>|8909,8910
-|8910,8911
Continued|8912,8921
sertraline|8922,8932
150mg|8933,8938
PO|8939,8941
daily|8942,8947
for|8948,8951
depression|8952,8962
<EOL>|8962,8963
-|8963,8964
Continued|8965,8974
Albuterol|8975,8984
0.083|8985,8990
%|8990,8991
Neb|8992,8995
Soln|8996,9000
1|9001,9002
NEB|9003,9006
IH|9007,9009
Q6H|9010,9013
:|9013,9014
PRN|9014,9017
cough|9018,9023
,|9023,9024
<EOL>|9024,9025
wheeze|9025,9031
<EOL>|9031,9032
-|9032,9033
Held|9034,9038
ProAir|9039,9045
<EOL>|9045,9046
-|9046,9047
Held|9048,9052
trazadone|9053,9062
while|9063,9068
getting|9069,9076
opioids|9077,9084
<EOL>|9084,9085
-|9085,9086
Held|9087,9091
furosemide|9092,9102
20mg|9103,9107
PO|9108,9110
daily|9111,9116
PRN|9117,9120
:|9120,9121
takes|9122,9127
rarely|9128,9134
<EOL>|9135,9136
-|9136,9137
d|9138,9139
/|9139,9140
c|9140,9141
gabapentin|9142,9152
:|9152,9153
not|9154,9157
helping|9158,9165
and|9166,9169
not|9170,9173
taking|9174,9180
<EOL>|9180,9181
-|9181,9182
d|9183,9184
/|9184,9185
c|9185,9186
erythromycin|9187,9199
-|9199,9200
no|9201,9203
longer|9204,9210
taking|9211,9217
<EOL>|9217,9218
<EOL>|9218,9219
Admission|9219,9228
to|9229,9231
Ortho|9232,9237
spine|9238,9243
:|9243,9244
<EOL>|9244,9245
<EOL>|9245,9246
Ms.|9246,9249
_|9250,9251
_|9251,9252
_|9252,9253
is|9254,9256
a|9257,9258
_|9259,9260
_|9260,9261
_|9261,9262
female|9263,9269
with|9270,9274
a|9275,9276
past|9277,9281
medical|9282,9289
<EOL>|9290,9291
history|9291,9298
significant|9299,9310
for|9311,9314
OSA|9315,9318
,|9318,9319
cerebral|9320,9328
aneurysm|9329,9337
,|9337,9338
abdominal|9339,9348
aortic|9349,9355
<EOL>|9356,9357
aneurysm|9357,9365
,|9365,9366
antiphospholipid|9367,9383
syndrome|9384,9392
w|9393,9394
/|9394,9395
multiple|9396,9404
DVTs|9405,9409
and|9410,9413
one|9414,9417
<EOL>|9418,9419
event|9419,9424
of|9425,9427
bilateral|9428,9437
large|9438,9443
PEs|9444,9447
on|9448,9450
warfarin|9451,9459
,|9459,9460
BRCA1|9461,9466
mutation|9467,9475
w|9476,9477
/|9477,9478
<EOL>|9478,9479
L|9479,9480
-|9480,9481
sided|9481,9486
breast|9487,9493
cancer|9494,9500
s|9501,9502
/|9502,9503
p|9503,9504
lumpectomy|9505,9515
,|9515,9516
who|9517,9520
presents|9521,9529
with|9530,9534
over|9535,9539
one|9540,9543
<EOL>|9544,9545
month|9545,9550
of|9551,9553
right|9554,9559
lower|9560,9565
back|9566,9570
pain|9571,9575
with|9576,9580
radicular|9581,9590
pain|9591,9595
down|9596,9600
the|9601,9604
<EOL>|9605,9606
right|9606,9611
leg|9612,9615
pain|9616,9620
found|9621,9626
to|9627,9629
have|9630,9634
significant|9635,9646
disc|9647,9651
herniations|9652,9663
at|9664,9666
<EOL>|9667,9668
L2|9668,9670
-|9670,9671
L5|9671,9673
.|9673,9674
She|9675,9678
is|9679,9681
now|9682,9685
s|9686,9687
/|9687,9688
p|9688,9689
L2|9691,9693
-|9693,9694
5|9694,9695
lami|9696,9700
,|9700,9701
L4|9702,9704
-|9704,9705
5|9705,9706
discectomy|9707,9717
,|9717,9718
and|9719,9722
<EOL>|9723,9724
non-instrumented|9724,9740
fusion|9741,9747
c|9748,9749
/|9749,9750
b|9750,9751
durotomy|9752,9760
s|9761,9762
/|9762,9763
p|9763,9764
_|9765,9766
_|9766,9767
_|9767,9768
,|9768,9769
_|9770,9771
_|9771,9772
_|9772,9773
<EOL>|9773,9774
<EOL>|9775,9776
<EOL>|9776,9777
Post|9777,9781
op|9782,9784
course|9785,9791
:|9791,9792
<EOL>|9793,9794
Patient|9794,9801
was|9802,9805
admitted|9806,9814
to|9815,9817
the|9818,9821
_|9822,9823
_|9823,9824
_|9824,9825
Spine|9826,9831
Surgery|9832,9839
Service|9840,9847
and|9848,9851
<EOL>|9852,9853
taken|9853,9858
to|9859,9861
the|9862,9865
Operating|9866,9875
Room|9876,9880
for|9881,9884
the|9885,9888
above|9889,9894
procedure|9895,9904
.|9904,9905
Refer|9905,9910
to|9911,9913
the|9914,9917
<EOL>|9918,9919
dictated|9919,9927
operative|9928,9937
note|9938,9942
for|9943,9946
further|9947,9954
details|9955,9962
.|9962,9963
The|9963,9966
surgery|9967,9974
was|9975,9978
<EOL>|9979,9980
without|9980,9987
complication|9988,10000
and|10001,10004
the|10005,10008
patient|10009,10016
was|10017,10020
transferred|10021,10032
to|10033,10035
the|10036,10039
PACU|10040,10044
<EOL>|10045,10046
in|10046,10048
a|10049,10050
stable|10051,10057
condition|10058,10067
.|10067,10068
<EOL>|10068,10069
<EOL>|10069,10070
Postoperative|10070,10083
DVT|10084,10087
_|10088,10089
_|10089,10090
_|10090,10091
drip|10092,10096
post|10097,10101
<EOL>|10102,10103
op|10103,10105
with|10106,10110
trasition|10111,10120
back|10121,10125
to|10126,10128
lovenox|10129,10136
bridge|10137,10143
to|10144,10146
coumadin|10147,10155
on|10156,10158
_|10159,10160
_|10160,10161
_|10161,10162
.|10162,10163
<EOL>|10164,10165
Activity|10165,10173
remained|10174,10182
flat|10183,10187
/|10187,10188
bedrest|10188,10195
for|10196,10199
dural|10200,10205
tear|10206,10210
precautions|10211,10222
for|10223,10226
48|10227,10229
<EOL>|10230,10231
hours|10231,10236
.|10236,10237
<EOL>|10238,10239
<EOL>|10239,10240
Activity|10240,10248
was|10249,10252
advanced|10253,10261
after|10262,10267
48|10268,10270
hours|10271,10276
.|10276,10277
Intravenous|10278,10289
antibiotics|10290,10301
<EOL>|10302,10303
were|10303,10307
continued|10308,10317
for|10318,10321
24hrs|10322,10327
postop|10328,10334
per|10335,10338
standard|10339,10347
protocol|10348,10356
.|10356,10357
<EOL>|10357,10358
<EOL>|10358,10359
Initial|10359,10366
postop|10367,10373
pain|10374,10378
was|10379,10382
controlled|10383,10393
with|10394,10398
oral|10399,10403
and|10404,10407
IV|10408,10410
pain|10411,10415
<EOL>|10416,10417
medication|10417,10427
.|10427,10428
Diet|10428,10432
was|10433,10436
advanced|10437,10445
as|10446,10448
tolerated|10449,10458
.|10458,10459
Foley|10459,10464
was|10465,10468
removed|10469,10476
on|10477,10479
<EOL>|10480,10481
POD|10481,10484
#|10484,10485
3|10485,10486
.|10486,10487
Physical|10488,10496
therapy|10497,10504
and|10505,10508
Occupational|10509,10521
therapy|10522,10529
were|10530,10534
consulted|10535,10544
<EOL>|10545,10546
for|10546,10549
mobilization|10550,10562
OOB|10563,10566
to|10567,10569
ambulate|10570,10578
and|10579,10582
ADL|10583,10586
's|10586,10588
.|10588,10589
<EOL>|10589,10590
<EOL>|10590,10591
Post|10591,10595
op|10596,10598
course|10599,10605
was|10606,10609
notable|10610,10617
for|10618,10621
acute|10622,10627
blood|10628,10633
loss|10634,10638
anemia|10639,10645
,|10645,10646
<EOL>|10647,10648
constipation|10648,10660
,|10660,10661
pain|10662,10666
and|10667,10670
hypokalemia|10671,10682
.|10682,10683
Acute|10684,10689
blood|10690,10695
loss|10696,10700
anemia|10701,10707
is|10708,10710
<EOL>|10711,10712
stable|10712,10718
and|10719,10722
did|10723,10726
not|10727,10730
require|10731,10738
intervention|10739,10751
.|10751,10752
She|10753,10756
was|10757,10760
treated|10761,10768
with|10769,10773
<EOL>|10774,10775
Immediate|10775,10784
release|10785,10792
morphine|10793,10801
,|10801,10802
Valium|10803,10809
and|10810,10813
Tylenol|10814,10821
for|10822,10825
pain|10826,10830
control|10831,10838
.|10838,10839
<EOL>|10840,10841
Oral|10841,10845
Potassium|10846,10855
was|10856,10859
given|10860,10865
for|10866,10869
hypokalemia|10870,10881
of|10882,10884
3.3|10885,10888
on|10889,10891
_|10892,10893
_|10893,10894
_|10894,10895
.|10895,10896
Vitals|10897,10903
<EOL>|10904,10905
and|10905,10908
labs|10909,10913
are|10914,10917
otherwise|10918,10927
stable|10928,10934
.|10934,10935
<EOL>|10936,10937
<EOL>|10937,10938
Hospital|10938,10946
course|10947,10953
was|10954,10957
otherwise|10958,10967
unremarkable|10968,10980
.|10980,10981
On|10981,10983
the|10984,10987
day|10988,10991
of|10992,10994
<EOL>|10995,10996
discharge|10996,11005
the|11006,11009
patient|11010,11017
was|11018,11021
afebrile|11022,11030
with|11031,11035
stable|11036,11042
vital|11043,11048
signs|11049,11054
,|11054,11055
<EOL>|11056,11057
comfortable|11057,11068
on|11069,11071
oral|11072,11076
pain|11077,11081
control|11082,11089
and|11090,11093
tolerating|11094,11104
a|11105,11106
regular|11107,11114
diet|11115,11119
.|11119,11120
<EOL>|11120,11121
<EOL>|11121,11122
<EOL>|11123,11124
Medications|11124,11135
on|11136,11138
Admission|11139,11148
:|11148,11149
<EOL>|11149,11150
The|11150,11153
Preadmission|11154,11166
Medication|11167,11177
list|11178,11182
is|11183,11185
accurate|11186,11194
and|11195,11198
complete|11199,11207
.|11207,11208
<EOL>|11208,11209
1.|11209,11211
Acetaminophen|11212,11225
1000|11226,11230
mg|11231,11233
PO|11234,11236
Q8H|11237,11240
:|11240,11241
PRN|11241,11244
Pain|11245,11249
-|11250,11251
Mild|11252,11256
/|11256,11257
Fever|11257,11262
<EOL>|11263,11264
2.|11264,11266
Albuterol|11267,11276
0.083|11277,11282
%|11282,11283
Neb|11284,11287
Soln|11288,11292
1|11293,11294
NEB|11295,11298
IH|11299,11301
Q6H|11302,11305
:|11305,11306
PRN|11306,11309
cough|11310,11315
,|11315,11316
wheeze|11317,11323
<EOL>|11324,11325
3.|11325,11327
Atorvastatin|11328,11340
40|11341,11343
mg|11344,11346
PO|11347,11349
QPM|11350,11353
<EOL>|11354,11355
4.|11355,11357
Docusate|11358,11366
Sodium|11367,11373
100|11374,11377
mg|11378,11380
PO|11381,11383
BID|11384,11387
<EOL>|11388,11389
5.|11389,11391
Omeprazole|11392,11402
20|11403,11405
mg|11406,11408
PO|11409,11411
BID|11412,11415
<EOL>|11416,11417
6.|11417,11419
Polyethylene|11420,11432
Glycol|11433,11439
17|11440,11442
g|11443,11444
PO|11445,11447
DAILY|11448,11453
:|11453,11454
PRN|11454,11457
Constipation|11458,11470
-|11471,11472
First|11473,11478
<EOL>|11479,11480
Line|11480,11484
<EOL>|11485,11486
7.|11486,11488
Senna|11489,11494
8.6|11495,11498
mg|11499,11501
PO|11502,11504
HS|11505,11507
<EOL>|11508,11509
8.|11509,11511
Sertraline|11512,11522
150|11523,11526
mg|11527,11529
PO|11530,11532
DAILY|11533,11538
<EOL>|11539,11540
9.|11540,11542
TraZODone|11543,11552
50|11553,11555
mg|11556,11558
PO|11559,11561
QHS|11562,11565
:|11565,11566
PRN|11566,11569
sleep|11570,11575
<EOL>|11576,11577
10|11577,11579
.|11579,11580
Vitamin|11581,11588
D|11589,11590
_|11591,11592
_|11592,11593
_|11593,11594
UNIT|11595,11599
PO|11600,11602
DAILY|11603,11608
<EOL>|11609,11610
11.|11610,11613
Warfarin|11614,11622
7.5|11623,11626
mg|11627,11629
PO|11630,11632
2X|11633,11635
/|11635,11636
WEEK|11636,11640
(|11641,11642
_|11642,11643
_|11643,11644
_|11644,11645
)|11645,11646
<EOL>|11647,11648
12.|11648,11651
Lidocaine|11652,11661
5|11662,11663
%|11663,11664
Patch|11665,11670
1|11671,11672
PTCH|11673,11677
TD|11678,11680
QAM|11681,11684
right|11685,11690
hip|11691,11694
<EOL>|11695,11696
13.|11696,11699
Furosemide|11700,11710
20|11711,11713
mg|11714,11716
PO|11717,11719
DAILY|11720,11725
:|11725,11726
PRN|11726,11729
Leg|11730,11733
swelling|11734,11742
<EOL>|11743,11744
14.|11744,11747
ProAir|11748,11754
HFA|11755,11758
(|11759,11760
albuterol|11760,11769
sulfate|11770,11777
)|11777,11778
90|11779,11781
mcg|11782,11785
/|11785,11786
actuation|11786,11795
inhalation|11796,11806
<EOL>|11807,11808
Q4H|11808,11811
:|11811,11812
PRN|11812,11815
<EOL>|11816,11817
15.|11817,11820
Warfarin|11821,11829
5|11830,11831
mg|11832,11834
PO|11835,11837
5X|11838,11840
/|11840,11841
WEEK|11841,11845
(|11846,11847
_|11847,11848
_|11848,11849
_|11849,11850
)|11850,11851
<EOL>|11852,11853
16|11853,11855
.|11855,11856
Gabapentin|11857,11867
600|11868,11871
mg|11872,11874
PO|11875,11877
TID|11878,11881
<EOL>|11882,11883
17.|11883,11886
TraMADol|11887,11895
50|11896,11898
mg|11899,11901
PO|11902,11904
Q6H|11905,11908
:|11908,11909
PRN|11909,11912
Pain|11913,11917
-|11918,11919
Moderate|11920,11928
<EOL>|11929,11930
<EOL>|11930,11931
<EOL>|11932,11933
Discharge|11933,11942
Medications|11943,11954
:|11954,11955
<EOL>|11955,11956
1.|11956,11958
Diazepam|11960,11968
5|11969,11970
mg|11971,11973
PO|11974,11976
Q8H|11977,11980
:|11980,11981
PRN|11981,11984
pain|11985,11989
/|11989,11990
spasm|11990,11995
<EOL>|11996,11997
may|11997,12000
cause|12001,12006
drowsiness|12007,12017
<EOL>|12018,12019
RX|12019,12021
*|12022,12023
diazepam|12023,12031
5|12032,12033
mg|12034,12036
1|12037,12038
tablet|12039,12045
by|12046,12048
mouth|12049,12054
every|12055,12060
eight|12061,12066
(|12067,12068
8|12068,12069
)|12069,12070
hours|12071,12076
Disp|12077,12081
<EOL>|12082,12083
#|12083,12084
*|12084,12085
25|12085,12087
Tablet|12088,12094
Refills|12095,12102
:|12102,12103
*|12103,12104
0|12104,12105
<EOL>|12106,12107
2.|12107,12109
Enoxaparin|12111,12121
Sodium|12122,12128
110|12129,12132
mg|12133,12135
SC|12136,12138
Q12H|12139,12143
Antiphospholipid|12144,12160
Syndrome|12161,12169
<EOL>|12170,12171
Treatment|12171,12180
Bridge|12181,12187
Dosing|12188,12194
<EOL>|12196,12197
3.|12197,12199
Morphine|12201,12209
Sulfate|12210,12217
_|12218,12219
_|12219,12220
_|12220,12221
15|12222,12224
mg|12225,12227
PO|12228,12230
Q6H|12231,12234
:|12234,12235
PRN|12235,12238
Pain|12239,12243
-|12244,12245
Severe|12246,12252
<EOL>|12253,12254
please|12254,12260
do|12261,12263
not|12264,12267
operate|12268,12275
heavy|12276,12281
machinery|12282,12291
,|12291,12292
drink|12293,12298
alcohol|12299,12306
or|12307,12309
drive|12310,12315
<EOL>|12316,12317
RX|12317,12319
*|12320,12321
morphine|12321,12329
15|12330,12332
mg|12333,12335
1|12336,12337
tablet|12338,12344
(|12344,12345
s|12345,12346
)|12346,12347
by|12348,12350
mouth|12351,12356
every|12357,12362
six|12363,12366
(|12367,12368
6|12368,12369
)|12369,12370
hours|12371,12376
Disp|12377,12381
<EOL>|12382,12383
#|12383,12384
*|12384,12385
30|12385,12387
Tablet|12388,12394
Refills|12395,12402
:|12402,12403
*|12403,12404
0|12404,12405
<EOL>|12406,12407
4.|12407,12409
Furosemide|12411,12421
10|12422,12424
mg|12425,12427
PO|12428,12430
DAILY|12431,12436
:|12436,12437
PRN|12437,12440
Leg|12441,12444
swelling|12445,12453
<EOL>|12455,12456
5.|12456,12458
Acetaminophen|12460,12473
1000|12474,12478
mg|12479,12481
PO|12482,12484
Q8H|12485,12488
:|12488,12489
PRN|12489,12492
Pain|12493,12497
-|12498,12499
Mild|12500,12504
/|12504,12505
Fever|12505,12510
<EOL>|12512,12513
6.|12513,12515
Albuterol|12517,12526
0.083|12527,12532
%|12532,12533
Neb|12534,12537
Soln|12538,12542
1|12543,12544
NEB|12545,12548
IH|12549,12551
Q6H|12552,12555
:|12555,12556
PRN|12556,12559
cough|12560,12565
,|12565,12566
wheeze|12567,12573
<EOL>|12575,12576
7.|12576,12578
Atorvastatin|12580,12592
40|12593,12595
mg|12596,12598
PO|12599,12601
QPM|12602,12605
<EOL>|12607,12608
8.|12608,12610
Docusate|12612,12620
Sodium|12621,12627
100|12628,12631
mg|12632,12634
PO|12635,12637
BID|12638,12641
<EOL>|12643,12644
9.|12644,12646
Lidocaine|12648,12657
5|12658,12659
%|12659,12660
Patch|12661,12666
1|12667,12668
PTCH|12669,12673
TD|12674,12676
QAM|12677,12680
right|12681,12686
hip|12687,12690
<EOL>|12692,12693
10.|12693,12696
Omeprazole|12698,12708
20|12709,12711
mg|12712,12714
PO|12715,12717
BID|12718,12721
<EOL>|12723,12724
11.|12724,12727
Polyethylene|12729,12741
Glycol|12742,12748
17|12749,12751
g|12752,12753
PO|12754,12756
DAILY|12757,12762
:|12762,12763
PRN|12763,12766
Constipation|12767,12779
-|12780,12781
First|12782,12787
<EOL>|12788,12789
Line|12789,12793
<EOL>|12795,12796
12.|12796,12799
ProAir|12801,12807
HFA|12808,12811
(|12812,12813
albuterol|12813,12822
sulfate|12823,12830
)|12830,12831
90|12832,12834
mcg|12835,12838
/|12838,12839
actuation|12839,12848
inhalation|12849,12859
<EOL>|12860,12861
Q4H|12861,12864
:|12864,12865
PRN|12865,12868
<EOL>|12870,12871
13.|12871,12874
Senna|12876,12881
8.6|12882,12885
mg|12886,12888
PO|12889,12891
HS|12892,12894
<EOL>|12896,12897
14.|12897,12900
Sertraline|12902,12912
150|12913,12916
mg|12917,12919
PO|12920,12922
DAILY|12923,12928
<EOL>|12930,12931
15.|12931,12934
TraZODone|12936,12945
50|12946,12948
mg|12949,12951
PO|12952,12954
QHS|12955,12958
:|12958,12959
PRN|12959,12962
sleep|12963,12968
<EOL>|12970,12971
16|12971,12973
.|12973,12974
Vitamin|12976,12983
D|12984,12985
_|12986,12987
_|12987,12988
_|12988,12989
UNIT|12990,12994
PO|12995,12997
DAILY|12998,13003
<EOL>|13005,13006
17.|13006,13009
Warfarin|13011,13019
5|13020,13021
mg|13022,13024
PO|13025,13027
5X|13028,13030
/|13030,13031
WEEK|13031,13035
(|13036,13037
_|13037,13038
_|13038,13039
_|13039,13040
)|13040,13041
<EOL>|13043,13044
18.|13044,13047
Warfarin|13049,13057
7.5|13058,13061
mg|13062,13064
PO|13065,13067
2X|13068,13070
/|13070,13071
WEEK|13071,13075
(|13076,13077
_|13077,13078
_|13078,13079
_|13079,13080
)|13080,13081
<EOL>|13083,13084
<EOL>|13084,13085
<EOL>|13086,13087
Discharge|13087,13096
Disposition|13097,13108
:|13108,13109
<EOL>|13109,13110
Extended|13110,13118
Care|13119,13123
<EOL>|13123,13124
<EOL>|13125,13126
Facility|13126,13134
:|13134,13135
<EOL>|13135,13136
_|13136,13137
_|13137,13138
_|13138,13139
<EOL>|13139,13140
<EOL>|13141,13142
Discharge|13142,13151
Diagnosis|13152,13161
:|13161,13162
<EOL>|13162,13163
-|13163,13164
Lumbar|13164,13170
spinal|13171,13177
stenosis|13178,13186
.|13186,13187
<EOL>|13187,13188
-|13188,13189
Spondylolisthesis|13189,13206
,|13206,13207
L4|13208,13210
-|13210,13211
L5|13211,13213
.|13213,13214
<EOL>|13214,13215
-|13215,13216
UTI|13216,13219
<EOL>|13219,13220
-|13220,13221
Constipation|13221,13233
<EOL>|13233,13234
<EOL>|13234,13235
Secondary|13235,13244
Diagnoses|13245,13254
:|13254,13255
<EOL>|13255,13256
-|13256,13257
History|13258,13265
of|13266,13268
DVT|13269,13272
/|13272,13273
PE|13273,13275
<EOL>|13275,13276
-|13276,13277
Antiphospholipid|13278,13294
antibody|13295,13303
syndrome|13304,13312
<EOL>|13312,13313
-|13313,13314
AAA|13315,13318
<EOL>|13318,13319
-|13319,13320
OSA|13321,13324
on|13325,13327
CPAP|13328,13332
<EOL>|13333,13334
<EOL>|13334,13335
<EOL>|13336,13337
Discharge|13337,13346
Condition|13347,13356
:|13356,13357
<EOL>|13357,13358
Mental|13358,13364
Status|13365,13371
:|13371,13372
Clear|13373,13378
and|13379,13382
coherent|13383,13391
.|13391,13392
<EOL>|13392,13393
Level|13393,13398
of|13399,13401
Consciousness|13402,13415
:|13415,13416
Alert|13417,13422
and|13423,13426
interactive|13427,13438
.|13438,13439
<EOL>|13439,13440
Activity|13440,13448
Status|13449,13455
:|13455,13456
Ambulatory|13457,13467
-|13468,13469
requires|13470,13478
assistance|13479,13489
or|13490,13492
aid|13493,13496
(|13497,13498
walker|13498,13504
<EOL>|13505,13506
or|13506,13508
cane|13509,13513
)|13513,13514
.|13514,13515
<EOL>|13515,13516
<EOL>|13516,13517
<EOL>|13518,13519
Discharge|13519,13528
Instructions|13529,13541
:|13541,13542
<EOL>|13542,13543
It|13543,13545
was|13546,13549
a|13550,13551
pleasure|13552,13560
to|13561,13563
care|13564,13568
for|13569,13572
you|13573,13576
at|13577,13579
the|13580,13583
_|13584,13585
_|13585,13586
_|13586,13587
<EOL>|13588,13589
_|13589,13590
_|13590,13591
_|13591,13592
.|13592,13593
<EOL>|13595,13596
<EOL>|13596,13597
Why|13597,13600
did|13601,13604
you|13605,13608
come|13609,13613
to|13614,13616
the|13617,13620
hospital|13621,13629
?|13629,13630
<EOL>|13632,13633
-|13633,13634
You|13636,13639
came|13640,13644
to|13645,13647
the|13648,13651
hospital|13652,13660
because|13661,13668
you|13669,13672
were|13673,13677
having|13678,13684
worsening|13685,13694
<EOL>|13695,13696
back|13696,13700
pain|13701,13705
with|13706,13710
pain|13711,13715
radiating|13716,13725
down|13726,13730
your|13731,13735
right|13736,13741
leg|13742,13745
.|13745,13746
This|13747,13751
pain|13752,13756
<EOL>|13757,13758
started|13758,13765
about|13766,13771
a|13772,13773
month|13774,13779
ago|13780,13783
and|13784,13787
progressively|13788,13801
got|13802,13805
worse|13806,13811
,|13811,13812
making|13813,13819
it|13820,13822
<EOL>|13823,13824
difficult|13824,13833
to|13834,13836
walk|13837,13841
.|13841,13842
You|13843,13846
also|13847,13851
had|13852,13855
burning|13856,13863
pain|13864,13868
with|13869,13873
urination|13874,13883
.|13883,13884
<EOL>|13884,13885
<EOL>|13885,13886
What|13886,13890
did|13891,13894
you|13895,13898
receive|13899,13906
in|13907,13909
the|13910,13913
hospital|13914,13922
?|13922,13923
<EOL>|13925,13926
-|13926,13927
You|13928,13931
had|13932,13935
an|13936,13938
MRI|13939,13942
that|13943,13947
showed|13948,13954
significant|13955,13966
disc|13967,13971
herniation|13972,13982
in|13983,13985
your|13986,13990
<EOL>|13991,13992
lower|13992,13997
back|13998,14002
,|14002,14003
which|14004,14009
was|14010,14013
the|14014,14017
cause|14018,14023
of|14024,14026
your|14027,14031
pain|14032,14036
.|14036,14037
The|14038,14041
spine|14042,14047
surgeons|14048,14056
<EOL>|14057,14058
felt|14058,14062
that|14063,14067
you|14068,14071
would|14072,14077
benefit|14078,14085
from|14086,14090
surgery|14091,14098
given|14099,14104
that|14105,14109
your|14110,14114
pain|14115,14119
<EOL>|14120,14121
was|14121,14124
constant|14125,14133
and|14134,14137
worsening|14138,14147
over|14148,14152
the|14153,14156
past|14157,14161
month|14162,14167
.|14167,14168
We|14169,14171
gave|14172,14176
you|14177,14180
pain|14181,14185
<EOL>|14186,14187
medications|14187,14198
and|14199,14202
stopped|14203,14210
your|14211,14215
warfarin|14216,14224
until|14225,14230
it|14231,14233
was|14234,14237
safe|14238,14242
for|14243,14246
you|14247,14250
<EOL>|14251,14252
to|14252,14254
have|14255,14259
surgery|14260,14267
.|14267,14268
You|14269,14272
had|14273,14276
a|14277,14278
spinal|14279,14285
decompression|14286,14299
on|14300,14302
_|14303,14304
_|14304,14305
_|14305,14306
.|14306,14307
We|14308,14310
<EOL>|14311,14312
also|14312,14316
gave|14317,14321
you|14322,14325
antibiotics|14326,14337
for|14338,14341
your|14342,14346
burning|14347,14354
pain|14355,14359
with|14360,14364
urination|14365,14374
,|14374,14375
<EOL>|14376,14377
which|14377,14382
we|14383,14385
believe|14386,14393
was|14394,14397
caused|14398,14404
by|14405,14407
a|14408,14409
urinary|14410,14417
tract|14418,14423
infection|14424,14433
.|14433,14434
<EOL>|14435,14436
<EOL>|14436,14437
What|14437,14441
should|14442,14448
you|14449,14452
do|14453,14455
once|14456,14460
you|14461,14464
leave|14465,14470
the|14471,14474
hospital|14475,14483
?|14483,14484
<EOL>|14486,14487
<EOL>|14487,14488
Lumbar|14488,14494
Decompression|14495,14508
With|14509,14513
Fusion|14514,14520
:|14520,14521
<EOL>|14521,14522
<EOL>|14522,14523
You|14523,14526
have|14527,14531
undergone|14532,14541
the|14542,14545
following|14546,14555
operation|14556,14565
:|14565,14566
Lumbar|14567,14573
Decompression|14574,14587
<EOL>|14588,14589
With|14589,14593
Fusion|14594,14600
<EOL>|14600,14601
<EOL>|14601,14602
Immediately|14602,14613
after|14614,14619
the|14620,14623
operation|14624,14633
:|14633,14634
<EOL>|14634,14635
<EOL>|14635,14636
|14636,14637
Activity|14653,14661
:|14661,14662
You|14662,14665
should|14666,14672
not|14673,14676
lift|14677,14681
anything|14682,14690
greater|14691,14698
<EOL>|14699,14700
than|14700,14704
10|14705,14707
lbs|14708,14711
for|14712,14715
2|14716,14717
weeks|14718,14723
.|14723,14724
You|14724,14727
will|14728,14732
be|14733,14735
more|14736,14740
comfortable|14741,14752
if|14753,14755
you|14756,14759
do|14760,14762
<EOL>|14763,14764
not|14764,14767
sit|14768,14771
or|14772,14774
stand|14775,14780
more|14781,14785
than|14786,14790
~|14790,14791
45|14791,14793
minutes|14794,14801
without|14802,14809
getting|14810,14817
up|14818,14820
and|14821,14824
<EOL>|14825,14826
walking|14826,14833
around|14834,14840
.|14840,14841
<EOL>|14841,14842
<EOL>|14842,14843
|14843,14844
Rehabilitation|14860,14874
/|14874,14875
Physical|14876,14884
_|14885,14886
_|14886,14887
_|14887,14888
times|14889,14894
a|14895,14896
<EOL>|14897,14898
day|14898,14901
you|14902,14905
should|14906,14912
go|14913,14915
for|14916,14919
a|14920,14921
walk|14922,14926
for|14927,14930
_|14931,14932
_|14932,14933
_|14933,14934
minutes|14935,14942
as|14943,14945
part|14946,14950
of|14951,14953
your|14954,14958
<EOL>|14959,14960
recovery|14960,14968
.|14968,14969
You|14969,14972
can|14973,14976
walk|14977,14981
as|14982,14984
much|14985,14989
as|14990,14992
you|14993,14996
can|14997,15000
tolerate|15001,15009
.|15009,15010
Limit|15010,15015
any|15016,15019
kind|15020,15024
<EOL>|15025,15026
of|15026,15028
lifting|15029,15036
.|15036,15037
<EOL>|15037,15038
<EOL>|15038,15039
|15039,15040
Diet|15056,15060
:|15060,15061
Eat|15062,15065
a|15066,15067
normal|15068,15074
healthy|15075,15082
diet|15083,15087
.|15087,15088
You|15088,15091
may|15092,15095
have|15096,15100
<EOL>|15101,15102
some|15102,15106
constipation|15107,15119
after|15120,15125
surgery|15126,15133
.|15133,15134
You|15134,15137
have|15138,15142
been|15143,15147
given|15148,15153
medication|15154,15164
<EOL>|15165,15166
to|15166,15168
help|15169,15173
with|15174,15178
this|15179,15183
issue|15184,15189
.|15189,15190
<EOL>|15190,15191
<EOL>|15191,15192
|15192,15193
Brace|15209,15214
:|15214,15215
You|15215,15218
may|15219,15222
have|15223,15227
been|15228,15232
given|15233,15238
a|15239,15240
brace|15241,15246
.|15246,15247
If|15247,15249
you|15250,15253
<EOL>|15254,15255
have|15255,15259
been|15260,15264
given|15265,15270
a|15271,15272
brace|15273,15278
,|15278,15279
this|15279,15283
brace|15284,15289
is|15290,15292
to|15293,15295
be|15296,15298
worn|15299,15303
when|15304,15308
you|15309,15312
are|15313,15316
<EOL>|15317,15318
walking|15318,15325
.|15325,15326
You|15326,15329
may|15330,15333
take|15334,15338
it|15339,15341
off|15342,15345
when|15346,15350
sitting|15351,15358
in|15359,15361
a|15362,15363
chair|15364,15369
or|15370,15372
while|15373,15378
<EOL>|15379,15380
lying|15380,15385
in|15386,15388
bed|15389,15392
.|15392,15393
<EOL>|15393,15394
<EOL>|15394,15395
|15395,15396
Wound|15412,15417
Care|15418,15422
:|15422,15423
Please|15423,15429
keep|15430,15434
the|15435,15438
incision|15439,15447
covered|15448,15455
<EOL>|15456,15457
with|15457,15461
a|15462,15463
dry|15464,15467
dressing|15468,15476
on|15477,15479
until|15480,15485
your|15486,15490
follow|15491,15497
up|15498,15500
appointment|15501,15512
.|15512,15513
Do|15514,15516
not|15517,15520
<EOL>|15521,15522
soak|15522,15526
the|15527,15530
incision|15531,15539
in|15540,15542
a|15543,15544
bath|15545,15549
or|15550,15552
pool|15553,15557
.|15557,15558
If|15558,15560
the|15561,15564
incision|15565,15573
starts|15574,15580
<EOL>|15581,15582
draining|15582,15590
at|15591,15593
anytime|15594,15601
after|15602,15607
surgery|15608,15615
,|15615,15616
do|15616,15618
not|15619,15622
get|15623,15626
the|15627,15630
incision|15631,15639
<EOL>|15640,15641
wet|15641,15644
.|15644,15645
Call|15645,15649
the|15650,15653
office|15654,15660
at|15661,15663
that|15664,15668
time|15669,15673
.|15673,15674
<EOL>|15674,15675
<EOL>|15675,15676
|15676,15677
You|15693,15696
should|15697,15703
resume|15704,15710
taking|15711,15717
your|15718,15722
normal|15723,15729
home|15730,15734
<EOL>|15735,15736
medications|15736,15747
.|15747,15748
<EOL>|15748,15749
<EOL>|15749,15750
|15750,15751
You|15767,15770
have|15771,15775
also|15776,15780
been|15781,15785
given|15786,15791
Additional|15792,15802
Medications|15803,15814
<EOL>|15815,15816
to|15816,15818
control|15819,15826
your|15827,15831
pain|15832,15836
.|15836,15837
Please|15837,15843
allow|15844,15849
72|15850,15852
hours|15853,15858
for|15859,15862
refill|15863,15869
of|15870,15872
<EOL>|15873,15874
narcotic|15874,15882
prescriptions|15883,15896
,|15896,15897
so|15897,15899
please|15900,15906
plan|15907,15911
ahead|15912,15917
.|15917,15918
You|15918,15921
can|15922,15925
either|15926,15932
have|15933,15937
<EOL>|15938,15939
them|15939,15943
mailed|15944,15950
to|15951,15953
your|15954,15958
home|15959,15963
or|15964,15966
pick|15967,15971
them|15972,15976
up|15977,15979
at|15980,15982
the|15983,15986
clinic|15987,15993
located|15994,16001
<EOL>|16002,16003
on|16003,16005
_|16006,16007
_|16007,16008
_|16008,16009
.|16009,16010
We|16010,16012
are|16013,16016
not|16017,16020
allowed|16021,16028
to|16029,16031
call|16032,16036
in|16037,16039
or|16040,16042
fax|16043,16046
narcotic|16047,16055
<EOL>|16056,16057
prescriptions|16057,16070
(|16070,16071
oxycontin|16071,16080
,|16080,16081
oxycodone|16081,16090
,|16090,16091
percocet|16091,16099
)|16099,16100
to|16101,16103
your|16104,16108
pharmacy|16109,16117
.|16117,16118
In|16118,16120
<EOL>|16121,16122
addition|16122,16130
,|16130,16131
we|16131,16133
are|16134,16137
only|16138,16142
allowed|16143,16150
to|16151,16153
write|16154,16159
for|16160,16163
pain|16164,16168
medications|16169,16180
for|16181,16184
<EOL>|16185,16186
90|16186,16188
days|16189,16193
from|16194,16198
the|16199,16202
date|16203,16207
of|16208,16210
surgery|16211,16218
.|16218,16219
<EOL>|16219,16220
<EOL>|16220,16221
|16221,16222
Follow|16238,16244
up|16245,16247
:|16247,16248
<EOL>|16248,16249
<EOL>|16249,16250
Please|16265,16271
Call|16272,16276
the|16277,16280
office|16281,16287
and|16288,16291
make|16292,16296
an|16297,16299
appointment|16300,16311
<EOL>|16312,16313
for|16313,16316
2|16317,16318
weeks|16319,16324
after|16325,16330
the|16331,16334
day|16335,16338
of|16339,16341
your|16342,16346
operation|16347,16356
if|16357,16359
this|16360,16364
has|16365,16368
not|16369,16372
been|16373,16377
<EOL>|16378,16379
done|16379,16383
already|16384,16391
.|16391,16392
<EOL>|16392,16393
<EOL>|16393,16394
At|16409,16411
the|16412,16415
2|16416,16417
-|16417,16418
week|16418,16422
visit|16423,16428
we|16429,16431
will|16432,16436
check|16437,16442
your|16443,16447
<EOL>|16448,16449
incision|16449,16457
,|16457,16458
take|16458,16462
baseline|16463,16471
X-rays|16472,16478
and|16479,16482
answer|16483,16489
any|16490,16493
questions|16494,16503
.|16503,16504
We|16504,16506
may|16507,16510
at|16511,16513
<EOL>|16514,16515
that|16515,16519
time|16520,16524
start|16525,16530
physical|16531,16539
therapy|16540,16547
<EOL>|16547,16548
<EOL>|16548,16549
We|16565,16567
will|16568,16572
then|16573,16577
see|16578,16581
you|16582,16585
at|16586,16588
6|16589,16590
weeks|16591,16596
from|16597,16601
the|16602,16605
day|16606,16609
of|16610,16612
<EOL>|16613,16614
the|16614,16617
operation|16618,16627
and|16628,16631
at|16632,16634
that|16635,16639
time|16640,16644
release|16645,16652
you|16653,16656
to|16657,16659
full|16660,16664
activity|16665,16673
.|16673,16674
<EOL>|16674,16675
<EOL>|16675,16676
Please|16676,16682
call|16683,16687
the|16688,16691
office|16692,16698
if|16699,16701
you|16702,16705
have|16706,16710
a|16711,16712
fever|16713,16718
>|16718,16719
101.5|16719,16724
degrees|16725,16732
<EOL>|16733,16734
Fahrenheit|16734,16744
and|16745,16748
/|16748,16749
or|16749,16751
drainage|16752,16760
from|16761,16765
your|16766,16770
wound|16771,16776
.|16776,16777
<EOL>|16777,16778
<EOL>|16778,16779
Physical|16779,16787
Therapy|16788,16795
:|16795,16796
<EOL>|16796,16797
1|16797,16798
)|16798,16799
Weight|16799,16805
bearing|16806,16813
as|16814,16816
tolerated|16817,16826
.2|16826,16828
)|16828,16829
Gait|16829,16833
,|16833,16834
balance|16834,16841
training|16842,16850
.3|16850,16852
)|16852,16853
No|16853,16855
<EOL>|16856,16857
lifting|16857,16864
>|16865,16866
10|16866,16868
lbs|16869,16872
.4|16872,16874
)|16874,16875
No|16875,16877
significant|16878,16889
bending|16890,16897
/|16897,16898
twisting|16898,16906
.|16906,16907
<EOL>|16908,16909
Treatments|16909,16919
Frequency|16920,16929
:|16929,16930
<EOL>|16930,16931
Please|16931,16937
keep|16938,16942
the|16943,16946
incision|16947,16955
covered|16956,16963
with|16964,16968
a|16969,16970
dry|16971,16974
dressing|16975,16983
on|16984,16986
until|16987,16992
<EOL>|16993,16994
your|16994,16998
follow|16999,17005
up|17006,17008
appointment|17009,17020
.|17020,17021
Do|17022,17024
not|17025,17028
soak|17029,17033
the|17034,17037
incision|17038,17046
in|17047,17049
a|17050,17051
bath|17052,17056
<EOL>|17057,17058
or|17058,17060
pool|17061,17065
.|17065,17066
If|17066,17068
the|17069,17072
incision|17073,17081
starts|17082,17088
draining|17089,17097
at|17098,17100
anytime|17101,17108
after|17109,17114
<EOL>|17115,17116
surgery|17116,17123
,|17123,17124
do|17124,17126
not|17127,17130
get|17131,17134
the|17135,17138
incision|17139,17147
wet|17148,17151
.|17151,17152
Call|17152,17156
the|17157,17160
office|17161,17167
at|17168,17170
that|17171,17175
<EOL>|17176,17177
time|17177,17181
.|17181,17182
<EOL>|17182,17183
<EOL>|17184,17185
Followup|17185,17193
Instructions|17194,17206
:|17206,17207
<EOL>|17207,17208
_|17208,17209
_|17209,17210
_|17210,17211
<EOL>|17211,17212

