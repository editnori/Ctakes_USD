 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Procedure|Health Care Activity|SIMPLE_SEGMENT|48,57|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|48,62|false|false|false|C2598112||Admission Date
Finding|Body Substance|SIMPLE_SEGMENT|82,91|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|82,91|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|82,91|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|82,91|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|82,96|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|114,119|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|114,119|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|114,119|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|138,141|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|138,141|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|138,141|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|138,141|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|138,141|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|149,156|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|149,156|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Finding|Finding|SIMPLE_SEGMENT|158,165|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|SURGERY
Finding|Functional Concept|SIMPLE_SEGMENT|158,165|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|SURGERY
Finding|Idea or Concept|SIMPLE_SEGMENT|158,165|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|SURGERY
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|158,165|false|false|false|C0543467|Operative Surgical Procedures|SURGERY
Disorder|Injury or Poisoning|Allergies|180,192|false|false|false|C0161497;C2876788|Poisoning by sulfonamide;Poisoning by, adverse effect of and underdosing of sulfonamides|Sulfonamides
Drug|Antibiotic|Allergies|180,192|false|false|false|C0038760;C0599503;C3539179;C3539184;C3541962;C3541963|Sulfonamide Anti-Infective Agents;Sulfonamides;Sulfonamides, Gynecological;Sulfonamides, intestinal antiinfectives;Sulfonamides, ophthalmologic antiinfectives;Sulfonamides, topical|Sulfonamides
Drug|Organic Chemical|Allergies|180,192|false|false|false|C0038760;C0599503;C3539179;C3539184;C3541962;C3541963|Sulfonamide Anti-Infective Agents;Sulfonamides;Sulfonamides, Gynecological;Sulfonamides, intestinal antiinfectives;Sulfonamides, ophthalmologic antiinfectives;Sulfonamides, topical|Sulfonamides
Drug|Pharmacologic Substance|Allergies|180,192|false|false|false|C0038760;C0599503;C3539179;C3539184;C3541962;C3541963|Sulfonamide Anti-Infective Agents;Sulfonamides;Sulfonamides, Gynecological;Sulfonamides, intestinal antiinfectives;Sulfonamides, ophthalmologic antiinfectives;Sulfonamides, topical|Sulfonamides
Finding|Pathologic Function|Allergies|180,192|false|false|false|C0261773|Adverse reaction to sulfonamides|Sulfonamides
Drug|Organic Chemical|Allergies|195,202|false|false|false|C0009214|codeine|Codeine
Drug|Pharmacologic Substance|Allergies|195,202|false|false|false|C0009214|codeine|Codeine
Drug|Organic Chemical|Allergies|205,212|false|false|false|C0591139|Bactrim|Bactrim
Drug|Pharmacologic Substance|Allergies|205,212|false|false|false|C0591139|Bactrim|Bactrim
Finding|Functional Concept|Allergies|215,224|false|false|false|C1999232|Attending (action)|Attending
Anatomy|Body Location or Region|Chief Complaint|250,259|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|Chief Complaint|250,264|false|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|Chief Complaint|260,264|false|false|false|C2598155||pain
Finding|Functional Concept|Chief Complaint|260,264|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Chief Complaint|260,264|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Chief Complaint|269,277|false|false|false|C0042963|Vomiting|vomiting
Finding|Classification|Chief Complaint|280,285|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|286,294|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|286,294|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|298,316|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|307,316|false|false|false|C0945766||Procedure
Event|Occupational Activity|Chief Complaint|307,316|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|307,316|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|307,316|false|false|false|C0184661|Interventional procedure|Procedure
Procedure|Diagnostic Procedure|Chief Complaint|322,344|false|false|false|C0085704|Exploratory laparotomy|Exploratory laparotomy
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|334,344|false|false|false|C0023038|Laparotomy|laparotomy
Finding|Cell Function|Chief Complaint|346,351|false|false|false|C0024348;C1536403|Lysis;pathologic cytolysis|lysis
Finding|Pathologic Function|Chief Complaint|346,351|false|false|false|C0024348;C1536403|Lysis;pathologic cytolysis|lysis
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|346,364|false|false|false|C0012826|Lysis of adhesions|lysis of adhesions
Finding|Pathologic Function|Chief Complaint|355,364|false|false|false|C0001511|Tissue Adhesions|adhesions
Anatomy|Body Part, Organ, or Organ Component|Chief Complaint|372,377|false|false|false|C0021853|Intestines|bowel
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|372,387|false|false|false|C0741614|Bowel resection|bowel resection
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|378,387|false|false|false|C0015252;C0728940|Excision;removal technique|resection
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|393,410|false|false|false|C0192711;C0192741|Anastomosis of intestine;Anastomosis of small intestine to small intestine|enteroenterostomy
Finding|Body Substance|History of Present Illness|447,454|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|447,454|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|447,454|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|464,468|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|History of Present Illness|464,468|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Finding|History of Present Illness|483,495|false|false|false|C1548863|Consent Type - Hysterectomy|hysterectomy
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|483,495|false|false|false|C0020699|Hysterectomy|hysterectomy
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|500,507|false|false|false|C0042149|Uterus|uterine
Disorder|Neoplastic Process|History of Present Illness|509,517|false|false|false|C0023267;C0042133|Fibroid Tumor;Uterine Fibroids|fibroids
Anatomy|Body Location or Region|History of Present Illness|528,532|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|528,532|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|History of Present Illness|528,532|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|History of Present Illness|528,532|false|false|false|C0740941|Lung Problem|lung
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|528,542|false|false|false|C0396565|Lung excision|lung resection
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|533,542|false|false|false|C0015252;C0728940|Excision;removal technique|resection
Disorder|Neoplastic Process|History of Present Illness|547,556|false|false|false|C0007095|Carcinoid Tumor|carcinoid
Disorder|Neoplastic Process|History of Present Illness|547,562|false|false|false|C0007095|Carcinoid Tumor|carcinoid tumor
Disorder|Neoplastic Process|History of Present Illness|557,562|false|true|false|C0027651|Neoplasms|tumor
Finding|Finding|History of Present Illness|557,562|false|true|false|C1578706;C3273930|Tumor Mass|tumor
Finding|Intellectual Product|History of Present Illness|557,562|false|true|false|C1578706;C3273930|Tumor Mass|tumor
Procedure|Health Care Activity|History of Present Illness|579,587|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|579,587|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Procedure|Health Care Activity|History of Present Illness|579,600|false|false|false|C5442589|Surgical consultation|surgical consultation
Finding|Classification|History of Present Illness|588,600|false|false|false|C1546898;C1548374|Diagnosis Classification - Consultation;Document Type - Consultation|consultation
Finding|Intellectual Product|History of Present Illness|588,600|false|false|false|C1546898;C1548374|Diagnosis Classification - Consultation;Document Type - Consultation|consultation
Procedure|Health Care Activity|History of Present Illness|588,600|false|false|false|C0009818|Consultation|consultation
Anatomy|Body Location or Region|History of Present Illness|605,614|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|History of Present Illness|605,619|false|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|History of Present Illness|615,619|false|false|true|C2598155||pain
Finding|Functional Concept|History of Present Illness|615,619|false|false|true|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|615,619|false|false|true|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|History of Present Illness|621,627|false|false|false|C4255480||nausea
Finding|Sign or Symptom|History of Present Illness|621,627|false|false|false|C0027497|Nausea|nausea
Finding|Sign or Symptom|History of Present Illness|634,642|false|false|false|C0042963|Vomiting|vomiting
Finding|Body Substance|History of Present Illness|648,655|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|648,655|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|648,655|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Finding|History of Present Illness|668,672|false|false|false|C5575035|Well (answer to question)|well
Finding|Sign or Symptom|History of Present Illness|743,751|false|false|false|C0026821|Muscle Cramp|cramping
Anatomy|Body Location or Region|History of Present Illness|752,761|false|false|false|C0000726|Abdomen|abdominal
Attribute|Clinical Attribute|History of Present Illness|763,767|false|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|763,767|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|763,767|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|History of Present Illness|784,790|false|false|false|C4255480||nausea
Finding|Sign or Symptom|History of Present Illness|784,790|false|false|false|C0027497|Nausea|nausea
Finding|Finding|History of Present Illness|795,809|false|false|false|C0232599|Vomiting bile|bilious emesis
Finding|Body Substance|History of Present Illness|803,809|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Finding|Physiologic Function|History of Present Illness|803,809|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Finding|Sign or Symptom|History of Present Illness|803,809|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Disorder|Disease or Syndrome|History of Present Illness|818,823|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|History of Present Illness|818,823|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Disorder|Disease or Syndrome|History of Present Illness|857,862|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|History of Present Illness|882,894|false|false|false|C0449450|Presentation|presentation
Finding|Finding|History of Present Illness|915,919|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|History of Present Illness|915,919|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|History of Present Illness|915,919|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Body Substance|History of Present Illness|927,933|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Finding|Physiologic Function|History of Present Illness|927,933|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Finding|Sign or Symptom|History of Present Illness|927,933|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Finding|Finding|History of Present Illness|943,951|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|History of Present Illness|943,951|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|967,973|false|false|false|C0021853|Intestines|bowels
Finding|Finding|History of Present Illness|976,983|false|false|false|C4035626|3 times|3 times
Disorder|Disease or Syndrome|History of Present Illness|978,983|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Attribute|Clinical Attribute|History of Present Illness|1021,1025|false|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|1021,1025|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1021,1025|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Anatomy|Body Location or Region|History of Present Illness|1087,1098|false|false|false|C0021852;C4319010|Abdomen>Small bowel;Intestines, Small|small bowel
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1087,1098|false|false|false|C0021852;C4319010|Abdomen>Small bowel;Intestines, Small|small bowel
Disorder|Disease or Syndrome|History of Present Illness|1087,1110|false|false|false|C0235329|Small bowel obstruction|small bowel obstruction
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1093,1098|false|false|false|C0021853|Intestines|bowel
Disorder|Disease or Syndrome|History of Present Illness|1093,1110|false|false|false|C0021843|Intestinal Obstruction|bowel obstruction
Finding|Finding|History of Present Illness|1099,1110|false|false|false|C0028778|Obstruction|obstruction
Procedure|Diagnostic Procedure|History of Present Illness|1133,1144|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Procedure|Health Care Activity|History of Present Illness|1133,1144|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Disorder|Neoplastic Process|Past Medical History|1184,1193|false|false|false|C0007095|Carcinoid Tumor|carcinoid
Disorder|Neoplastic Process|Past Medical History|1184,1199|false|false|false|C0007095|Carcinoid Tumor|carcinoid tumor
Disorder|Neoplastic Process|Past Medical History|1194,1199|false|false|false|C0027651|Neoplasms|tumor
Finding|Finding|Past Medical History|1194,1199|false|false|false|C1578706;C3273930|Tumor Mass|tumor
Finding|Intellectual Product|Past Medical History|1194,1199|false|false|false|C1578706;C3273930|Tumor Mass|tumor
Finding|Idea or Concept|Past Medical History|1203,1208|false|false|false|C1552828|Table Frame - above|above
Drug|Organic Chemical|Past Medical History|1209,1216|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|Past Medical History|1209,1216|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|Past Medical History|1209,1216|false|false|false|C0042890|Vitamins|Vitamin
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Past Medical History|1209,1220|false|false|false|C0042845;C0086024;C2936883|Vitamin B12 [EPC];cobalamins;vitamin B12|Vitamin B12
Drug|Organic Chemical|Past Medical History|1209,1220|false|false|false|C0042845;C0086024;C2936883|Vitamin B12 [EPC];cobalamins;vitamin B12|Vitamin B12
Drug|Pharmacologic Substance|Past Medical History|1209,1220|false|false|false|C0042845;C0086024;C2936883|Vitamin B12 [EPC];cobalamins;vitamin B12|Vitamin B12
Drug|Vitamin|Past Medical History|1209,1220|false|false|false|C0042845;C0086024;C2936883|Vitamin B12 [EPC];cobalamins;vitamin B12|Vitamin B12
Procedure|Laboratory Procedure|Past Medical History|1209,1220|false|false|false|C0202252|VITAMIN B12 MEASUREMENT|Vitamin B12
Disorder|Disease or Syndrome|Past Medical History|1209,1231|false|false|false|C0042847|Vitamin B 12 Deficiency|Vitamin B12 deficiency
Finding|Finding|Past Medical History|1209,1231|false|false|false|C5886863|Decreased circulating vitamin B12 concentration|Vitamin B12 deficiency
Finding|Gene or Genome|Past Medical History|1217,1220|false|false|false|C1417635;C1420797;C3538796|NDUFB3 gene;TNFAIP1 gene;TNFAIP1 wt Allele|B12
Disorder|Disease or Syndrome|Past Medical History|1221,1231|false|false|false|C0162429|Malnutrition|deficiency
Finding|Functional Concept|Past Medical History|1221,1231|false|false|false|C0011155|Deficiency|deficiency
Disorder|Mental or Behavioral Dysfunction|Past Medical History|1232,1242|false|false|false|C0011570;C0011581;C0344315;C0812393|Cancer patients and suicide and depression;Depressed mood;Depressive disorder;Mental Depression|depression
Finding|Functional Concept|Past Medical History|1232,1242|false|false|false|C0460137;C1579931|Depression - motion|depression
Finding|Sign or Symptom|Past Medical History|1232,1242|false|false|false|C0460137;C1579931|Depression - motion|depression
Disorder|Disease or Syndrome|Past Medical History|1243,1257|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|hyperlipidemia
Finding|Finding|Past Medical History|1243,1257|false|false|false|C0428465|Serum lipids high (finding)|hyperlipidemia
Anatomy|Body Location or Region|Past Medical History|1271,1275|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1271,1275|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Past Medical History|1271,1275|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Past Medical History|1271,1275|false|false|false|C0740941|Lung Problem|lung
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1271,1285|false|false|false|C0396565|Lung excision|lung resection
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1276,1285|false|false|false|C0015252;C0728940|Excision;removal technique|resection
Finding|Finding|Past Medical History|1304,1316|false|false|false|C1548863|Consent Type - Hysterectomy|hysterectomy
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1304,1316|false|false|false|C0020699|Hysterectomy|hysterectomy
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1328,1333|false|false|false|C4048756|Right arm|R arm
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1330,1333|false|false|false|C0446516;C1140618;C1269078|Upper Extremity;Upper arm|arm
Disorder|Anatomical Abnormality|Past Medical History|1330,1333|false|false|false|C3495676|Anorectal Malformations|arm
Finding|Gene or Genome|Past Medical History|1330,1333|false|false|false|C1824218;C3715044|AKR1A1 wt Allele;ARMC9 gene|arm
Procedure|Diagnostic Procedure|Past Medical History|1330,1333|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Research Activity|Past Medical History|1330,1333|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1330,1333|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Finding|Finding|Past Medical History|1334,1341|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|Past Medical History|1334,1341|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|Past Medical History|1334,1341|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1334,1341|false|false|false|C0543467|Operative Surgical Procedures|surgery
Event|Activity|Family Medical History|1385,1397|false|false|false|C1880177|Contribution|contributory
Finding|Gene or Genome|General Exam|1415,1419|false|false|false|C1823816|C1orf210 gene|Temp
Procedure|Therapeutic or Preventive Procedure|General Exam|1415,1419|false|false|false|C0279848|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Temp
Disorder|Disease or Syndrome|General Exam|1451,1454|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|General Exam|1451,1454|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|General Exam|1451,1454|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|1451,1454|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|General Exam|1451,1454|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Finding|Finding|General Exam|1451,1454|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Part, Organ, or Organ Component|General Exam|1492,1497|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|General Exam|1492,1497|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|General Exam|1492,1497|false|false|false|C0795691|HEART PROBLEM|heart
Finding|Finding|General Exam|1526,1533|true|false|false|C0018808|Heart murmur|murmurs
Anatomy|Body Part, Organ, or Organ Component|General Exam|1546,1551|false|false|false|C0024109|Lung|lungs
Finding|Idea or Concept|General Exam|1552,1557|false|false|false|C1550016|Remote control command - Clear|clear
Procedure|Diagnostic Procedure|General Exam|1561,1573|false|false|false|C0004339|Auscultation|auscultation
Finding|Finding|General Exam|1575,1598|false|false|false|C0238844|Decreased breath sounds|decreased breath sounds
Finding|Body Substance|General Exam|1585,1591|false|false|false|C0225386|Breath|breath
Attribute|Clinical Attribute|General Exam|1585,1598|false|false|false|C0035234;C3484186|Respiratory Sounds|breath sounds
Phenomenon|Natural Phenomenon or Process|General Exam|1592,1598|false|true|false|C0037709||sounds
Finding|Finding|General Exam|1605,1609|false|false|false|C5575035|Well (answer to question)|well
Procedure|Therapeutic or Preventive Procedure|General Exam|1619,1630|false|false|false|C0039991|Thoracotomy|thoracotomy
Finding|Finding|General Exam|1619,1635|false|false|false|C5238882|Thoracotomy Scar|thoracotomy scar
Finding|Finding|General Exam|1631,1635|false|false|false|C0241158;C1419736;C2004491|Cicatrix;RPS4X gene;Scar Tissue|scar
Finding|Gene or Genome|General Exam|1631,1635|false|false|false|C0241158;C1419736;C2004491|Cicatrix;RPS4X gene;Scar Tissue|scar
Finding|Pathologic Function|General Exam|1631,1635|false|false|false|C0241158;C1419736;C2004491|Cicatrix;RPS4X gene;Scar Tissue|scar
Finding|Finding|General Exam|1636,1643|false|true|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|General Exam|1636,1643|false|true|false|C0150312;C0449450|Present;Presentation|present
Anatomy|Body Location or Region|General Exam|1644,1651|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|abdomen
Disorder|Neoplastic Process|General Exam|1644,1651|false|false|false|C0153662|Malignant neoplasm of abdomen|abdomen
Finding|Finding|General Exam|1644,1651|false|false|false|C0941288|Abdomen problem|abdomen
Finding|Finding|General Exam|1644,1656|false|false|false|C0426663|Abdomen soft|abdomen soft
Disorder|Disease or Syndrome|General Exam|1652,1656|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Disorder|Disease or Syndrome|General Exam|1663,1668|false|false|false|C0028754|Obesity|obese
Finding|Finding|General Exam|1680,1689|false|false|false|C0700124|Dilated|distended
Finding|Finding|General Exam|1691,1699|false|false|false|C2984079|Somewhat|somewhat
Procedure|Diagnostic Procedure|General Exam|1711,1720|false|false|false|C0030247|Palpation|palpation
Anatomy|Body Location or Region|General Exam|1738,1745|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|abdomen
Disorder|Neoplastic Process|General Exam|1738,1745|false|false|false|C0153662|Malignant neoplasm of abdomen|abdomen
Finding|Finding|General Exam|1738,1745|false|false|false|C0941288|Abdomen problem|abdomen
Finding|Finding|General Exam|1750,1758|true|false|false|C0427198|Protective muscle spasm|guarding
Finding|Mental Process|General Exam|1771,1781|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|General Exam|1771,1781|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Finding|General Exam|1783,1786|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|General Exam|1783,1786|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Anatomy|Cell Component|General Exam|1787,1794|false|false|false|C1660780|midline cell component|midline
Anatomy|Body Location or Region|General Exam|1795,1804|false|false|false|C0000726|Abdomen|abdominal
Disorder|Injury or Poisoning|General Exam|1795,1810|false|false|false|C4510895|Wound of abdomen|abdominal wound
Disorder|Injury or Poisoning|General Exam|1805,1810|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|wound
Finding|Body Substance|General Exam|1805,1810|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Functional Concept|General Exam|1805,1810|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Intellectual Product|General Exam|1805,1810|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Body Substance|General Exam|1821,1829|true|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Finding|Sign or Symptom|General Exam|1821,1829|true|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Procedure|Therapeutic or Preventive Procedure|General Exam|1821,1829|true|false|false|C0013103|Drainage procedure|drainage
Disorder|Disease or Syndrome|General Exam|1835,1843|false|false|false|C0041834|Erythema|erythema
Anatomy|Cell|General Exam|1880,1883|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|1891,1894|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|1891,1894|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|1891,1894|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|1900,1903|false|false|false|C0019046|Hemoglobin|HGB
Drug|Biologically Active Substance|General Exam|1900,1903|false|false|false|C0019046|Hemoglobin|HGB
Finding|Gene or Genome|General Exam|1900,1903|false|false|false|C1424337|CYGB gene|HGB
Lab|Laboratory or Test Result|General Exam|1900,1903|false|false|false|C0019029|Hemoglobin concentration|HGB
Procedure|Laboratory Procedure|General Exam|1909,1912|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Procedure|Therapeutic or Preventive Procedure|General Exam|1909,1912|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Disorder|Virus|General Exam|1918,1921|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|General Exam|1918,1921|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|1918,1921|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|1918,1921|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|1926,1929|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|1926,1929|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|General Exam|1926,1929|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|1926,1929|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|1926,1929|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|General Exam|1935,1939|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Finding|Body Substance|General Exam|1980,1986|false|false|false|C0024202|Lymph|LYMPHS
Drug|Antibiotic|General Exam|1992,1997|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Biomedical or Dental Material|General Exam|1992,1997|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Organic Chemical|General Exam|1992,1997|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Disorder|Disease or Syndrome|General Exam|2003,2006|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|EOS
Finding|Gene or Genome|General Exam|2003,2006|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|EOS
Procedure|Laboratory Procedure|General Exam|2036,2039|false|false|false|C0201617|Primed lymphocyte test|PLT
Drug|Biologically Active Substance|General Exam|2064,2071|false|false|false|C0017725|glucose|GLUCOSE
Drug|Organic Chemical|General Exam|2064,2071|false|false|false|C0017725|glucose|GLUCOSE
Drug|Pharmacologic Substance|General Exam|2064,2071|false|false|false|C0017725|glucose|GLUCOSE
Lab|Laboratory or Test Result|General Exam|2064,2071|false|false|false|C5781949|Glucose^1.5H post dose glucagon|GLUCOSE
Procedure|Laboratory Procedure|General Exam|2064,2071|false|false|false|C0337438|Glucose measurement|GLUCOSE
Drug|Biologically Active Substance|General Exam|2077,2081|false|false|false|C0041942|urea|UREA
Drug|Organic Chemical|General Exam|2077,2081|false|false|false|C0041942|urea|UREA
Drug|Pharmacologic Substance|General Exam|2077,2081|false|false|false|C0041942|urea|UREA
Procedure|Laboratory Procedure|General Exam|2077,2081|false|false|false|C0523961|Urea measurement|UREA
Drug|Biologically Active Substance|General Exam|2097,2103|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Element, Ion, or Isotope|General Exam|2097,2103|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Pharmacologic Substance|General Exam|2097,2103|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Finding|Physiologic Function|General Exam|2097,2103|false|false|false|C4553025|Sodium metabolic function|SODIUM
Procedure|Laboratory Procedure|General Exam|2097,2103|false|false|false|C0337443|Sodium measurement|SODIUM
Drug|Biologically Active Substance|General Exam|2109,2118|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Element, Ion, or Isotope|General Exam|2109,2118|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Food|General Exam|2109,2118|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Inorganic Chemical|General Exam|2109,2118|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Pharmacologic Substance|General Exam|2109,2118|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Finding|Physiologic Function|General Exam|2109,2118|false|false|false|C4553027|Potassium metabolic function|POTASSIUM
Procedure|Laboratory Procedure|General Exam|2109,2118|false|false|false|C0202194|Potassium measurement|POTASSIUM
Drug|Element, Ion, or Isotope|General Exam|2123,2131|false|false|false|C0008203;C0596019|Chlorides;chloride ion|CHLORIDE
Finding|Physiologic Function|General Exam|2123,2131|false|false|false|C4553021|Chloride metabolic function|CHLORIDE
Procedure|Laboratory Procedure|General Exam|2123,2131|false|false|false|C0201952|Chloride measurement|CHLORIDE
Drug|Biologically Active Substance|General Exam|2142,2145|false|false|false|C0007012|carbon dioxide|CO2
Drug|Inorganic Chemical|General Exam|2142,2145|false|false|false|C0007012|carbon dioxide|CO2
Finding|Finding|General Exam|2142,2145|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Finding|Gene or Genome|General Exam|2142,2145|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Drug|Element, Ion, or Isotope|General Exam|2149,2154|false|false|false|C0003075|Anions|ANION
Attribute|Clinical Attribute|General Exam|2149,2158|false|false|false|C0003074|Anion Gap|ANION GAP
Lab|Laboratory or Test Result|General Exam|2149,2158|false|false|false|C1509129|Anion gap result|ANION GAP
Procedure|Laboratory Procedure|General Exam|2149,2158|false|false|false|C0201889;C2189246|Anion gap measurement;blood anion gap (lab test)|ANION GAP
Drug|Amino Acid, Peptide, or Protein|General Exam|2155,2158|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Drug|Biologically Active Substance|General Exam|2155,2158|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Finding|Gene or Genome|General Exam|2155,2158|false|false|false|C1419277;C2984552|RASA1 gene;RASA1 wt Allele|GAP
Disorder|Neoplastic Process|General Exam|2176,2179|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|General Exam|2176,2179|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|General Exam|2176,2179|false|false|false|C0001899|Alanine Transaminase|ALT
Finding|Gene or Genome|General Exam|2176,2179|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|General Exam|2176,2179|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|General Exam|2176,2179|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|General Exam|2176,2179|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Drug|Amino Acid, Peptide, or Protein|General Exam|2180,2184|false|false|false|C0376147|SGPT - Glutamate pyruvate transaminase|SGPT
Drug|Enzyme|General Exam|2180,2184|false|false|false|C0376147|SGPT - Glutamate pyruvate transaminase|SGPT
Finding|Gene or Genome|General Exam|2180,2184|false|false|false|C1415274|GPT gene|SGPT
Procedure|Laboratory Procedure|General Exam|2180,2184|false|false|false|C0036828|Serum Alanine Transaminase Test|SGPT
Anatomy|Body Space or Junction|General Exam|2189,2192|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|General Exam|2189,2192|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|2189,2192|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|General Exam|2189,2192|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|General Exam|2189,2192|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Finding|Gene or Genome|General Exam|2189,2192|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|2193,2197|false|false|false|C0242192|SGOT - Glutamate oxaloacetate transaminase|SGOT
Drug|Enzyme|General Exam|2193,2197|false|false|false|C0242192|SGOT - Glutamate oxaloacetate transaminase|SGOT
Finding|Gene or Genome|General Exam|2193,2197|false|false|false|C1415181|GOT1 gene|SGOT
Procedure|Laboratory Procedure|General Exam|2193,2197|false|false|false|C0201899|Aspartate aminotransferase measurement|SGOT
Drug|Amino Acid, Peptide, or Protein|General Exam|2205,2208|false|false|false|C0022917|Lactate Dehydrogenase|LDH
Drug|Enzyme|General Exam|2205,2208|false|false|false|C0022917|Lactate Dehydrogenase|LDH
Finding|Finding|General Exam|2205,2208|false|false|false|C0851148|Lifetime Drinking History|LDH
Procedure|Laboratory Procedure|General Exam|2205,2208|false|false|false|C0202113|Lactate dehydrogenase measurement|LDH
Drug|Amino Acid, Peptide, or Protein|General Exam|2214,2217|false|false|false|C1663627|ALK protein, human|ALK
Drug|Enzyme|General Exam|2214,2217|false|false|false|C1663627|ALK protein, human|ALK
Finding|Gene or Genome|General Exam|2214,2217|false|false|false|C1332080;C1663627;C1704943|ALK gene;ALK protein, human;ALK wt Allele|ALK
Finding|Receptor|General Exam|2214,2217|false|false|false|C1332080;C1663627;C1704943|ALK gene;ALK protein, human;ALK wt Allele|ALK
Procedure|Diagnostic Procedure|General Exam|2233,2246|false|false|false|C0412620|CT of abdomen|CT of abdomen
Procedure|Diagnostic Procedure|General Exam|2233,2257|false|false|false|C1641132|CT of abdomen and pelvis|CT of abdomen and pelvis
Anatomy|Body Location or Region|General Exam|2239,2246|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|abdomen
Disorder|Neoplastic Process|General Exam|2239,2246|false|false|false|C0153662|Malignant neoplasm of abdomen|abdomen
Finding|Finding|General Exam|2239,2246|false|false|false|C0941288|Abdomen problem|abdomen
Anatomy|Body Location or Region|General Exam|2239,2250|false|false|false|C0000726|Abdomen|abdomen and
Anatomy|Body Location or Region|General Exam|2239,2257|false|false|false|C1508499|Abdominopelvic structure|abdomen and pelvis
Anatomy|Body Part, Organ, or Organ Component|General Exam|2251,2257|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Anatomy|Body Space or Junction|General Exam|2251,2257|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Disorder|Neoplastic Process|General Exam|2251,2257|false|false|false|C0153663|Malignant neoplasm of pelvis|pelvis
Finding|Finding|General Exam|2251,2257|false|false|false|C0812455|Pelvis problem|pelvis
Finding|Finding|General Exam|2271,2278|false|false|false|C0700124|Dilated|dilated
Finding|Finding|General Exam|2271,2284|false|false|false|C4697734|Dilated loops|dilated loops
Anatomy|Body Location or Region|General Exam|2289,2300|false|false|false|C0021852;C4319010|Abdomen>Small bowel;Intestines, Small|small bowel
Anatomy|Body Part, Organ, or Organ Component|General Exam|2289,2300|false|false|false|C0021852;C4319010|Abdomen>Small bowel;Intestines, Small|small bowel
Anatomy|Body Part, Organ, or Organ Component|General Exam|2295,2300|false|false|false|C0021853|Intestines|bowel
Anatomy|Body Location or Region|General Exam|2322,2333|false|false|false|C0021852;C4319010|Abdomen>Small bowel;Intestines, Small|small bowel
Anatomy|Body Part, Organ, or Organ Component|General Exam|2322,2333|false|false|false|C0021852;C4319010|Abdomen>Small bowel;Intestines, Small|small bowel
Anatomy|Body Part, Organ, or Organ Component|General Exam|2328,2333|false|false|false|C0021853|Intestines|bowel
Finding|Intellectual Product|General Exam|2328,2342|false|false|false|C1546561|Bowel contents|bowel contents
Finding|Conceptual Entity|General Exam|2334,2342|false|false|false|C0456205;C1552853|Contents;contents - HtmlLinkType|contents
Finding|Intellectual Product|General Exam|2334,2342|false|false|false|C0456205;C1552853|Contents;contents - HtmlLinkType|contents
Attribute|Clinical Attribute|General Exam|2347,2353|false|false|false|C4522154|Distal Resection Margin|distal
Finding|Finding|General Exam|2355,2364|false|false|false|C0344329;C0392748|Collapse (finding);Collapsed|collapsed
Finding|Functional Concept|General Exam|2355,2364|false|false|false|C0344329;C0392748|Collapse (finding);Collapsed|collapsed
Drug|Organic Chemical|General Exam|2398,2406|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|General Exam|2398,2406|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|General Exam|2398,2406|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Finding|Functional Concept|General Exam|2398,2406|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|General Exam|2398,2406|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|General Exam|2410,2417|false|false|false|C1550516|Target Awareness - partial|partial
Anatomy|Body Part, Organ, or Organ Component|General Exam|2425,2430|false|false|false|C0021853|Intestines|bowel
Disorder|Disease or Syndrome|General Exam|2425,2442|false|false|false|C0021843|Intestinal Obstruction|bowel obstruction
Finding|Finding|General Exam|2431,2442|false|false|false|C0028778|Obstruction|obstruction
Finding|Functional Concept|General Exam|2462,2469|false|false|false|C0392747|Changing|changes
Finding|Functional Concept|General Exam|2483,2488|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|General Exam|2489,2493|false|false|false|C0035561|Bone structure of rib|ribs
Finding|Idea or Concept|General Exam|2507,2512|false|false|false|C1552828|Table Frame - above|above
Drug|Organic Chemical|General Exam|2525,2532|false|false|false|C0607422|Abdoman (drug)|abdoman
Drug|Pharmacologic Substance|General Exam|2525,2532|false|false|false|C0607422|Abdoman (drug)|abdoman
Anatomy|Body Part, Organ, or Organ Component|General Exam|2537,2543|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Anatomy|Body Space or Junction|General Exam|2537,2543|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Disorder|Neoplastic Process|General Exam|2537,2543|false|false|false|C0153663|Malignant neoplasm of pelvis|pelvis
Finding|Finding|General Exam|2537,2543|false|false|false|C0812455|Pelvis problem|pelvis
Finding|Intellectual Product|General Exam|2551,2559|false|false|false|C1552654|Parameterized Data Type - Interval|Interval
Finding|Idea or Concept|General Exam|2560,2569|false|false|false|C1546960|Patient Outcome - Worsening|worsening
Anatomy|Body Location or Region|General Exam|2573,2584|false|false|false|C0021852;C4319010|Abdomen>Small bowel;Intestines, Small|small bowel
Anatomy|Body Part, Organ, or Organ Component|General Exam|2573,2584|false|false|false|C0021852;C4319010|Abdomen>Small bowel;Intestines, Small|small bowel
Disorder|Disease or Syndrome|General Exam|2573,2596|false|false|false|C0235329|Small bowel obstruction|small bowel obstruction
Anatomy|Body Part, Organ, or Organ Component|General Exam|2579,2584|false|false|false|C0021853|Intestines|bowel
Disorder|Disease or Syndrome|General Exam|2579,2596|false|false|false|C0021843|Intestinal Obstruction|bowel obstruction
Finding|Finding|General Exam|2585,2596|false|false|false|C0028778|Obstruction|obstruction
Disorder|Cell or Molecular Dysfunction|General Exam|2598,2608|false|false|false|C0599156|Transition Mutation|Transition
Event|Activity|General Exam|2598,2608|false|false|false|C2700061|Transition (action)|Transition
Finding|Functional Concept|General Exam|2624,2628|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Finding|Body Substance|General Exam|2647,2654|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|General Exam|2647,2654|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|General Exam|2647,2654|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|General Exam|2693,2698|false|false|false|C1705923|Study Object|study
Procedure|Research Activity|General Exam|2693,2698|false|false|false|C0008972;C0947630;C2603343|Clinical Research;Scientific Study;Study|study
Finding|Functional Concept|General Exam|2705,2710|false|false|false|C1883002|Sequence Chromatogram|Trace
Finding|Functional Concept|General Exam|2711,2715|false|false|false|C0332296|Free of (attribute)|free
Finding|Pathologic Function|General Exam|2711,2721|false|false|false|C0013687|effusion|free fluid
Drug|Substance|General Exam|2716,2721|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|General Exam|2716,2721|false|false|false|C1546638|Fluid Specimen Code|fluid
Anatomy|Body Part, Organ, or Organ Component|General Exam|2729,2735|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Anatomy|Body Space or Junction|General Exam|2729,2735|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Disorder|Neoplastic Process|General Exam|2729,2735|false|false|false|C0153663|Malignant neoplasm of pelvis|pelvis
Finding|Finding|General Exam|2729,2735|false|false|false|C0812455|Pelvis problem|pelvis
Finding|Finding|General Exam|2739,2745|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|General Exam|2739,2745|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Functional Concept|General Exam|2746,2757|false|false|false|C0205463|Physiological|physiologic
Finding|Body Substance|General Exam|2778,2783|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|2778,2783|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|2778,2783|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Finding|General Exam|2778,2790|false|false|false|C0278030|Color of urine|URINE  COLOR
Drug|Biomedical or Dental Material|General Exam|2785,2790|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|COLOR
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|2785,2790|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|COLOR
Finding|Body Substance|General Exam|2829,2834|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|2829,2834|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|2829,2834|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Disorder|Disease or Syndrome|General Exam|2829,2841|false|false|false|C0018965|Hematuria|URINE  BLOOD
Disorder|Disease or Syndrome|General Exam|2836,2841|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|2836,2841|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Biologically Active Substance|General Exam|2845,2852|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|NITRITE
Drug|Inorganic Chemical|General Exam|2845,2852|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|NITRITE
Drug|Pharmacologic Substance|General Exam|2845,2852|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|NITRITE
Finding|Finding|General Exam|2853,2856|false|false|false|C5848551|Neg - answer|NEG
Drug|Amino Acid, Peptide, or Protein|General Exam|2857,2864|false|false|false|C0033684|Proteins|PROTEIN
Drug|Biologically Active Substance|General Exam|2857,2864|false|false|false|C0033684|Proteins|PROTEIN
Finding|Conceptual Entity|General Exam|2857,2864|false|false|false|C1521746|Protein Info|PROTEIN
Procedure|Laboratory Procedure|General Exam|2857,2864|false|false|false|C0202202|Protein measurement|PROTEIN
Drug|Biologically Active Substance|General Exam|2869,2876|false|false|false|C0017725|glucose|GLUCOSE
Drug|Organic Chemical|General Exam|2869,2876|false|false|false|C0017725|glucose|GLUCOSE
Drug|Pharmacologic Substance|General Exam|2869,2876|false|false|false|C0017725|glucose|GLUCOSE
Lab|Laboratory or Test Result|General Exam|2869,2876|false|false|false|C5781949|Glucose^1.5H post dose glucagon|GLUCOSE
Procedure|Laboratory Procedure|General Exam|2869,2876|false|false|false|C0337438|Glucose measurement|GLUCOSE
Finding|Finding|General Exam|2877,2880|false|false|false|C5848551|Neg - answer|NEG
Drug|Organic Chemical|General Exam|2881,2887|false|false|false|C0022634|Ketones|KETONE
Drug|Biologically Active Substance|General Exam|2891,2900|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|BILIRUBIN
Drug|Organic Chemical|General Exam|2891,2900|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|BILIRUBIN
Drug|Pharmacologic Substance|General Exam|2891,2900|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|BILIRUBIN
Procedure|Laboratory Procedure|General Exam|2891,2900|false|false|false|C0201913;C0863174|Bilirubin, total measurement;blood bilirubin level test|BILIRUBIN
Finding|Finding|General Exam|2901,2904|false|false|false|C5848551|Neg - answer|NEG
Finding|Finding|General Exam|2915,2918|false|false|false|C5848551|Neg - answer|NEG
Finding|Finding|General Exam|2932,2935|false|false|false|C5848551|Neg - answer|NEG
Finding|Body Substance|General Exam|2948,2953|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|2948,2953|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|2948,2953|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Lab|Laboratory or Test Result|General Exam|2948,2958|false|false|false|C0221752;C2188659|Red blood cells urine positive|URINE  RBC
Anatomy|Cell|General Exam|2955,2958|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|2955,2958|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|2955,2958|false|false|false|C0014792|Erythrocytes|RBC
Finding|Functional Concept|General Exam|2967,2975|false|false|false|C1510439|bacteria aspects|BACTERIA
Disorder|Disease or Syndrome|General Exam|2976,2979|false|false|false|C0011860|Diabetes Mellitus, Non-Insulin-Dependent|MOD
Drug|Food|General Exam|2980,2985|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Drug|Immunologic Factor|General Exam|2980,2985|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|2980,2985|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Drug|Pharmacologic Substance|General Exam|2980,2985|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Disorder|Disease or Syndrome|General Exam|2992,2995|false|false|false|C0267963|Exocrine pancreatic insufficiency|EPI
Drug|Amino Acid, Peptide, or Protein|General Exam|2992,2995|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Drug|Biologically Active Substance|General Exam|2992,2995|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Drug|Hormone|General Exam|2992,2995|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Drug|Organic Chemical|General Exam|2992,2995|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Drug|Pharmacologic Substance|General Exam|2992,2995|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Finding|Gene or Genome|General Exam|2992,2995|false|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|EPI
Finding|Intellectual Product|General Exam|2992,2995|false|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|EPI
Procedure|Diagnostic Procedure|General Exam|2992,2995|false|false|false|C0162734;C3641909|Echo-Planar Imaging;Electronic Portal Imaging|EPI
Finding|Body Substance|General Exam|3010,3015|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|3010,3015|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|3010,3015|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Finding|General Exam|3010,3023|false|false|false|C0455910|Mucus in urine (finding)|URINE  MUCOUS
Finding|Body Substance|General Exam|3017,3023|false|false|false|C0026727;C2753459|Mucus (substance);mucus layer|MUCOUS
Drug|Biologically Active Substance|General Exam|3042,3049|false|false|false|C0017725|glucose|GLUCOSE
Drug|Organic Chemical|General Exam|3042,3049|false|false|false|C0017725|glucose|GLUCOSE
Drug|Pharmacologic Substance|General Exam|3042,3049|false|false|false|C0017725|glucose|GLUCOSE
Lab|Laboratory or Test Result|General Exam|3042,3049|false|false|false|C5781949|Glucose^1.5H post dose glucagon|GLUCOSE
Procedure|Laboratory Procedure|General Exam|3042,3049|false|false|false|C0337438|Glucose measurement|GLUCOSE
Drug|Biologically Active Substance|General Exam|3055,3059|false|false|false|C0041942|urea|UREA
Drug|Organic Chemical|General Exam|3055,3059|false|false|false|C0041942|urea|UREA
Drug|Pharmacologic Substance|General Exam|3055,3059|false|false|false|C0041942|urea|UREA
Procedure|Laboratory Procedure|General Exam|3055,3059|false|false|false|C0523961|Urea measurement|UREA
Drug|Biologically Active Substance|General Exam|3075,3081|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Element, Ion, or Isotope|General Exam|3075,3081|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Pharmacologic Substance|General Exam|3075,3081|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Finding|Physiologic Function|General Exam|3075,3081|false|false|false|C4553025|Sodium metabolic function|SODIUM
Procedure|Laboratory Procedure|General Exam|3075,3081|false|false|false|C0337443|Sodium measurement|SODIUM
Drug|Biologically Active Substance|General Exam|3087,3096|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Element, Ion, or Isotope|General Exam|3087,3096|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Food|General Exam|3087,3096|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Inorganic Chemical|General Exam|3087,3096|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Pharmacologic Substance|General Exam|3087,3096|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Finding|Physiologic Function|General Exam|3087,3096|false|false|false|C4553027|Potassium metabolic function|POTASSIUM
Procedure|Laboratory Procedure|General Exam|3087,3096|false|false|false|C0202194|Potassium measurement|POTASSIUM
Drug|Element, Ion, or Isotope|General Exam|3101,3109|false|false|false|C0008203;C0596019|Chlorides;chloride ion|CHLORIDE
Finding|Physiologic Function|General Exam|3101,3109|false|false|false|C4553021|Chloride metabolic function|CHLORIDE
Procedure|Laboratory Procedure|General Exam|3101,3109|false|false|false|C0201952|Chloride measurement|CHLORIDE
Drug|Biologically Active Substance|General Exam|3120,3123|false|false|false|C0007012|carbon dioxide|CO2
Drug|Inorganic Chemical|General Exam|3120,3123|false|false|false|C0007012|carbon dioxide|CO2
Finding|Finding|General Exam|3120,3123|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Finding|Gene or Genome|General Exam|3120,3123|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Drug|Element, Ion, or Isotope|General Exam|3127,3132|false|false|false|C0003075|Anions|ANION
Attribute|Clinical Attribute|General Exam|3127,3136|false|false|false|C0003074|Anion Gap|ANION GAP
Lab|Laboratory or Test Result|General Exam|3127,3136|false|false|false|C1509129|Anion gap result|ANION GAP
Procedure|Laboratory Procedure|General Exam|3127,3136|false|false|false|C0201889;C2189246|Anion gap measurement;blood anion gap (lab test)|ANION GAP
Drug|Amino Acid, Peptide, or Protein|General Exam|3133,3136|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Drug|Biologically Active Substance|General Exam|3133,3136|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Finding|Gene or Genome|General Exam|3133,3136|false|false|false|C1419277;C2984552|RASA1 gene;RASA1 wt Allele|GAP
Disorder|Neoplastic Process|General Exam|3186,3189|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|General Exam|3186,3189|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|General Exam|3186,3189|false|false|false|C0001899|Alanine Transaminase|ALT
Finding|Gene or Genome|General Exam|3186,3189|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|General Exam|3186,3189|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|General Exam|3186,3189|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|General Exam|3186,3189|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Drug|Amino Acid, Peptide, or Protein|General Exam|3190,3194|false|false|false|C0376147|SGPT - Glutamate pyruvate transaminase|SGPT
Drug|Enzyme|General Exam|3190,3194|false|false|false|C0376147|SGPT - Glutamate pyruvate transaminase|SGPT
Finding|Gene or Genome|General Exam|3190,3194|false|false|false|C1415274|GPT gene|SGPT
Procedure|Laboratory Procedure|General Exam|3190,3194|false|false|false|C0036828|Serum Alanine Transaminase Test|SGPT
Anatomy|Body Space or Junction|General Exam|3199,3202|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|General Exam|3199,3202|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|3199,3202|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|General Exam|3199,3202|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|General Exam|3199,3202|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Finding|Gene or Genome|General Exam|3199,3202|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|3203,3207|false|false|false|C0242192|SGOT - Glutamate oxaloacetate transaminase|SGOT
Drug|Enzyme|General Exam|3203,3207|false|false|false|C0242192|SGOT - Glutamate oxaloacetate transaminase|SGOT
Finding|Gene or Genome|General Exam|3203,3207|false|false|false|C1415181|GOT1 gene|SGOT
Procedure|Laboratory Procedure|General Exam|3203,3207|false|false|false|C0201899|Aspartate aminotransferase measurement|SGOT
Drug|Amino Acid, Peptide, or Protein|General Exam|3215,3218|false|false|false|C0022917|Lactate Dehydrogenase|LDH
Drug|Enzyme|General Exam|3215,3218|false|false|false|C0022917|Lactate Dehydrogenase|LDH
Finding|Finding|General Exam|3215,3218|false|false|false|C0851148|Lifetime Drinking History|LDH
Procedure|Laboratory Procedure|General Exam|3215,3218|false|false|false|C0202113|Lactate dehydrogenase measurement|LDH
Drug|Amino Acid, Peptide, or Protein|General Exam|3224,3227|false|false|false|C1663627|ALK protein, human|ALK
Drug|Enzyme|General Exam|3224,3227|false|false|false|C1663627|ALK protein, human|ALK
Finding|Gene or Genome|General Exam|3224,3227|false|false|false|C1332080;C1663627;C1704943|ALK gene;ALK protein, human;ALK wt Allele|ALK
Finding|Receptor|General Exam|3224,3227|false|false|false|C1332080;C1663627;C1704943|ALK gene;ALK protein, human;ALK wt Allele|ALK
Drug|Amino Acid, Peptide, or Protein|General Exam|3264,3270|false|false|false|C0023764|lipase|LIPASE
Drug|Enzyme|General Exam|3264,3270|false|false|false|C0023764|lipase|LIPASE
Drug|Pharmacologic Substance|General Exam|3264,3270|false|false|false|C0023764|lipase|LIPASE
Procedure|Laboratory Procedure|General Exam|3264,3270|false|false|false|C0373670|Lipase measurement|LIPASE
Anatomy|Cell|General Exam|3288,3291|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|3299,3302|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|3299,3302|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|3299,3302|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|3308,3311|false|false|false|C0019046|Hemoglobin|HGB
Drug|Biologically Active Substance|General Exam|3308,3311|false|false|false|C0019046|Hemoglobin|HGB
Finding|Gene or Genome|General Exam|3308,3311|false|false|false|C1424337|CYGB gene|HGB
Lab|Laboratory or Test Result|General Exam|3308,3311|false|false|false|C0019029|Hemoglobin concentration|HGB
Procedure|Laboratory Procedure|General Exam|3317,3320|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Procedure|Therapeutic or Preventive Procedure|General Exam|3317,3320|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Disorder|Virus|General Exam|3326,3329|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|General Exam|3326,3329|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|3326,3329|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|3326,3329|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|3334,3337|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|3334,3337|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|General Exam|3334,3337|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|3334,3337|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|3334,3337|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|General Exam|3343,3347|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Finding|Body Substance|General Exam|3388,3394|false|false|false|C0024202|Lymph|LYMPHS
Drug|Antibiotic|General Exam|3400,3405|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Biomedical or Dental Material|General Exam|3400,3405|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Organic Chemical|General Exam|3400,3405|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Disorder|Disease or Syndrome|General Exam|3411,3414|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|EOS
Finding|Gene or Genome|General Exam|3411,3414|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|EOS
Procedure|Laboratory Procedure|General Exam|3444,3447|false|false|false|C0201617|Primed lymphocyte test|PLT
Finding|Idea or Concept|Hospital Course|3492,3496|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|Hospital Course|3492,3496|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Idea or Concept|Hospital Course|3528,3536|false|false|false|C1547192|Organization unit type - Hospital|hospital
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3551,3554|false|false|false|C0419179|NPO - Nothing by mouth|NPO
Drug|Substance|Hospital Course|3559,3565|false|false|false|C0302908|Liquid substance|fluids
Finding|Body Substance|Hospital Course|3559,3565|false|false|false|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3559,3565|false|false|false|C0016286|Fluid Therapy|fluids
Anatomy|Body Location or Region|Hospital Course|3593,3604|false|false|false|C3282907|Nasogastric|nasogastric
Finding|Functional Concept|Hospital Course|3593,3604|false|false|false|C0694637|Nasogastric Route of Administration|nasogastric
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3593,3609|false|false|false|C0812428|Nasogastric tube procedures|nasogastric tube
Finding|Functional Concept|Hospital Course|3605,3609|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|tube
Finding|Gene or Genome|Hospital Course|3605,3609|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|tube
Anatomy|Cell Component|Hospital Course|3628,3631|false|false|false|C2244316|proteasome-activating nucleotidase complex|pan
Disorder|Disease or Syndrome|Hospital Course|3628,3631|false|false|false|C0031036|Polyarteritis Nodosa|pan
Finding|Gene or Genome|Hospital Course|3628,3631|false|false|false|C5401218|ADA2 wt Allele|pan
Procedure|Health Care Activity|Hospital Course|3647,3658|false|false|false|C0886414|Body temperature measurement|temperature
Finding|Intellectual Product|Hospital Course|3689,3695|false|false|false|C0031082|Periodicals|serial
Finding|Finding|Hospital Course|3706,3714|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Finding|Functional Concept|Hospital Course|3706,3714|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Procedure|Health Care Activity|Hospital Course|3706,3714|false|false|false|C0031809|Physical Examination|physical
Finding|Finding|Hospital Course|3706,3719|false|false|false|C1509143|physical examination (physical finding)|physical exam
Procedure|Health Care Activity|Hospital Course|3706,3719|false|false|false|C0031809|Physical Examination|physical exam
Finding|Functional Concept|Hospital Course|3715,3719|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|Hospital Course|3715,3719|false|false|false|C0582103|Medical Examination|exam
Anatomy|Body Location or Region|Hospital Course|3725,3736|false|false|false|C3282907|Nasogastric|nasogastric
Finding|Functional Concept|Hospital Course|3725,3736|false|false|false|C0694637|Nasogastric Route of Administration|nasogastric
Finding|Functional Concept|Hospital Course|3738,3742|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|tube
Finding|Gene or Genome|Hospital Course|3738,3742|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|tube
Finding|Idea or Concept|Hospital Course|3758,3766|false|false|false|C1547192|Organization unit type - Hospital|hospital
Finding|Idea or Concept|Hospital Course|3767,3770|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|3767,3770|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Finding|Hospital Course|3767,3772|false|false|false|C3842676|Day 2|day 2
Anatomy|Body Location or Region|Hospital Course|3807,3816|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|Hospital Course|3807,3821|false|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|Hospital Course|3817,3821|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|3817,3821|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|3817,3821|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Procedure|Diagnostic Procedure|Hospital Course|3839,3852|false|false|false|C0412620|CT of abdomen|CT of abdomen
Anatomy|Body Location or Region|Hospital Course|3845,3852|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|abdomen
Disorder|Neoplastic Process|Hospital Course|3845,3852|false|false|false|C0153662|Malignant neoplasm of abdomen|abdomen
Finding|Finding|Hospital Course|3845,3852|false|false|false|C0941288|Abdomen problem|abdomen
Anatomy|Body Location or Region|Hospital Course|3845,3856|false|false|false|C0000726|Abdomen|abdomen and
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|3858,3864|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Anatomy|Body Space or Junction|Hospital Course|3858,3864|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Disorder|Neoplastic Process|Hospital Course|3858,3864|false|false|false|C0153663|Malignant neoplasm of pelvis|pelvis
Finding|Finding|Hospital Course|3858,3864|false|false|false|C0812455|Pelvis problem|pelvis
Finding|Functional Concept|Hospital Course|3888,3896|false|false|false|C0442805|Increase|increase
Finding|Intellectual Product|Hospital Course|3904,3910|false|false|false|C0542560|Academic degree|degree
Finding|Finding|Hospital Course|3915,3926|false|false|false|C0028778|Obstruction|obstruction
Finding|Finding|Hospital Course|3965,3974|false|false|false|C4738506|Operating|operating
Attribute|Clinical Attribute|Hospital Course|4004,4013|false|false|false|C0945766||procedure
Event|Occupational Activity|Hospital Course|4004,4013|false|false|false|C1546467|Act Class - procedure|procedure
Finding|Functional Concept|Hospital Course|4004,4013|false|false|false|C2700391|Procedure (set of actions)|procedure
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4004,4013|false|false|false|C0184661|Interventional procedure|procedure
Attribute|Clinical Attribute|Hospital Course|4034,4043|false|false|false|C0945766||procedure
Event|Occupational Activity|Hospital Course|4034,4043|false|false|false|C1546467|Act Class - procedure|procedure
Finding|Functional Concept|Hospital Course|4034,4043|false|false|false|C2700391|Procedure (set of actions)|procedure
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4034,4043|false|false|false|C0184661|Interventional procedure|procedure
Finding|Finding|Hospital Course|4044,4048|false|false|false|C5575035|Well (answer to question)|well
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4059,4062|false|false|false|C0419179|NPO - Nothing by mouth|NPO
Anatomy|Body Location or Region|Hospital Course|4069,4080|false|false|false|C3282907|Nasogastric|nasogastric
Finding|Functional Concept|Hospital Course|4069,4080|false|false|false|C0694637|Nasogastric Route of Administration|nasogastric
Finding|Functional Concept|Hospital Course|4082,4086|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|tube
Finding|Gene or Genome|Hospital Course|4082,4086|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|tube
Event|Activity|Hospital Course|4090,4095|false|false|false|C1882509|put - instruction imperative|place
Finding|Functional Concept|Hospital Course|4090,4095|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|Hospital Course|4090,4095|false|false|false|C1533810||place
Drug|Substance|Hospital Course|4116,4122|false|false|false|C0302908|Liquid substance|fluids
Finding|Body Substance|Hospital Course|4116,4122|false|false|false|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4116,4122|false|false|false|C0016286|Fluid Therapy|fluids
Attribute|Clinical Attribute|Hospital Course|4129,4133|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|4129,4133|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|4129,4133|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|Hospital Course|4167,4175|false|false|false|C0026549|morphine|morphine
Drug|Pharmacologic Substance|Hospital Course|4167,4175|false|false|false|C0026549|morphine|morphine
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4176,4179|false|false|false|C0149576|Structure of posterior cerebral artery|PCA
Disorder|Disease or Syndrome|Hospital Course|4176,4179|false|false|false|C0268398;C4275079|Familial lichen amyloidosis;Posterior cortical atrophy syndrome|PCA
Drug|Amino Acid, Peptide, or Protein|Hospital Course|4176,4179|false|false|false|C0030131;C0034330|p-Chloroamphetamine;pyrrolidonecarboxylic acid|PCA
Drug|Biologically Active Substance|Hospital Course|4176,4179|false|false|false|C0030131;C0034330|p-Chloroamphetamine;pyrrolidonecarboxylic acid|PCA
Drug|Indicator, Reagent, or Diagnostic Aid|Hospital Course|4176,4179|false|false|false|C0030131;C0034330|p-Chloroamphetamine;pyrrolidonecarboxylic acid|PCA
Drug|Organic Chemical|Hospital Course|4176,4179|false|false|false|C0030131;C0034330|p-Chloroamphetamine;pyrrolidonecarboxylic acid|PCA
Drug|Pharmacologic Substance|Hospital Course|4176,4179|false|false|false|C0030131;C0034330|p-Chloroamphetamine;pyrrolidonecarboxylic acid|PCA
Finding|Finding|Hospital Course|4176,4179|false|false|false|C0220723;C1549860;C1836722|CHOANAL ATRESIA, POSTERIOR;FLVCR1 gene;PCA Message Structure|PCA
Finding|Gene or Genome|Hospital Course|4176,4179|false|false|false|C0220723;C1549860;C1836722|CHOANAL ATRESIA, POSTERIOR;FLVCR1 gene;PCA Message Structure|PCA
Finding|Intellectual Product|Hospital Course|4176,4179|false|false|false|C0220723;C1549860;C1836722|CHOANAL ATRESIA, POSTERIOR;FLVCR1 gene;PCA Message Structure|PCA
Procedure|Laboratory Procedure|Hospital Course|4176,4179|false|false|false|C0030625;C0078944;C5968782|Passive Cutaneous Anaphylaxis;Patient controlled intravenous analgesia;Patient-Controlled Analgesia|PCA
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4176,4179|false|false|false|C0030625;C0078944;C5968782|Passive Cutaneous Anaphylaxis;Patient controlled intravenous analgesia;Patient-Controlled Analgesia|PCA
Anatomy|Body Location or Region|Hospital Course|4187,4198|false|false|false|C3282907|Nasogastric|nasogastric
Finding|Functional Concept|Hospital Course|4187,4198|false|false|false|C0694637|Nasogastric Route of Administration|nasogastric
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4187,4203|false|false|false|C0812428|Nasogastric tube procedures|nasogastric tube
Finding|Functional Concept|Hospital Course|4199,4203|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|tube
Finding|Gene or Genome|Hospital Course|4199,4203|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|tube
Finding|Gene or Genome|Hospital Course|4220,4224|false|false|false|C3469826;C3470073|DESI1 gene;SLC35G1 gene|post
Finding|Idea or Concept|Hospital Course|4228,4231|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|4228,4231|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Idea or Concept|Hospital Course|4251,4256|false|false|false|C1550016|Remote control command - Clear|clear
Finding|Finding|Hospital Course|4251,4263|false|false|false|C4264429|Clear liquid|clear liquid
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4251,4268|false|false|false|C2184084|Clear liquid diet|clear liquid diet
Drug|Biomedical or Dental Material|Hospital Course|4257,4263|false|false|false|C0302908;C1697794|Liquid Dosage Form;Liquid substance|liquid
Drug|Substance|Hospital Course|4257,4263|false|false|false|C0302908;C1697794|Liquid Dosage Form;Liquid substance|liquid
Finding|Finding|Hospital Course|4257,4263|false|false|false|C1304698|Liquid (finding)|liquid
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4257,4263|false|false|false|C0301571|Liquid diet|liquid
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4257,4268|false|false|false|C0301571|Liquid diet|liquid diet
Drug|Food|Hospital Course|4264,4268|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Finding|Functional Concept|Hospital Course|4264,4268|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|Hospital Course|4264,4268|false|false|false|C0012159|Diet therapy|diet
Finding|Finding|Hospital Course|4290,4294|false|false|false|C5575035|Well (answer to question)|well
Finding|Daily or Recreational Activity|Hospital Course|4345,4357|false|false|false|C0184625||regular diet
Drug|Food|Hospital Course|4353,4357|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Finding|Functional Concept|Hospital Course|4353,4357|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|Hospital Course|4353,4357|false|false|false|C0012159|Diet therapy|diet
Finding|Finding|Hospital Course|4376,4380|false|false|false|C5575035|Well (answer to question)|well
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4399,4404|false|false|false|C0021853|Intestines|bowel
Finding|Organism Function|Hospital Course|4399,4414|false|false|false|C0011135|Defecation|bowel movements
Finding|Organism Function|Hospital Course|4405,4414|false|false|false|C0026649|Movement|movements
Anatomy|Body Space or Junction|Hospital Course|4429,4433|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|4429,4433|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|4429,4433|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|4429,4433|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Sign or Symptom|Hospital Course|4429,4438|false|false|false|C0221776|Oral pain|oral pain
Attribute|Clinical Attribute|Hospital Course|4434,4438|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|4434,4438|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|4434,4438|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Pharmacologic Substance|Hospital Course|4439,4449|false|false|false|C0013227|Pharmaceutical Preparations|medication
Finding|Intellectual Product|Hospital Course|4439,4449|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Anatomy|Body Location or Region|Hospital Course|4457,4465|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|Hospital Course|4457,4465|false|false|false|C0332803|Surgical wound|incision
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4457,4465|false|false|false|C0184898|Surgical incisions|incision
Finding|Finding|Hospital Course|4478,4482|false|false|false|C5575035|Well (answer to question)|well
Finding|Finding|Hospital Course|4500,4506|false|false|false|C1554187|Gender Status - Intact|intact
Finding|Idea or Concept|Hospital Course|4559,4563|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|4559,4563|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|4559,4563|false|false|false|C1553498|home health encounter|home
Attribute|Clinical Attribute|Hospital Course|4573,4584|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|4573,4584|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|Hospital Course|4573,4584|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|4573,4597|false|false|false|C1627937|Medications on admission|Medications on Admission
Procedure|Health Care Activity|Hospital Course|4588,4597|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Disorder|Mental or Behavioral Dysfunction|Hospital Course|4609,4612|false|false|false|C1839839|MAJOR AFFECTIVE DISORDER 2|MDI
Finding|Intellectual Product|Hospital Course|4609,4612|false|false|false|C4049613|Myositis Damage Index|MDI
Finding|Gene or Genome|Hospital Course|4613,4616|false|false|false|C1422467|CIAO3 gene|prn
Finding|Sign or Symptom|Hospital Course|4617,4624|false|false|false|C0043144|Wheezing|wheezes
Drug|Organic Chemical|Hospital Course|4625,4632|false|false|false|C0720466|Flovent|Flovent
Drug|Pharmacologic Substance|Hospital Course|4625,4632|false|false|false|C0720466|Flovent|Flovent
Finding|Functional Concept|Hospital Course|4633,4640|false|false|false|C4319647|Inhaler (unit of presentation)|inhaler
Finding|Gene or Genome|Hospital Course|4641,4644|false|false|false|C1422467|CIAO3 gene|prn
Finding|Sign or Symptom|Hospital Course|4645,4652|false|false|false|C0043144|Wheezing|wheezes
Anatomy|Body Space or Junction|Hospital Course|4670,4674|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|4670,4674|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|4670,4674|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|4670,4674|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Drug|Organic Chemical|Hospital Course|4681,4692|false|false|false|C0074554|simvastatin|Simvastatin
Drug|Pharmacologic Substance|Hospital Course|4681,4692|false|false|false|C0074554|simvastatin|Simvastatin
Anatomy|Body Space or Junction|Hospital Course|4699,4703|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|4699,4703|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|4699,4703|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|4699,4703|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Anatomy|Body Space or Junction|Hospital Course|4727,4731|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|4727,4731|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|4727,4731|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|4727,4731|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Drug|Organic Chemical|Hospital Course|4749,4759|false|false|false|C0085934|Wellbutrin|Wellbutrin
Drug|Pharmacologic Substance|Hospital Course|4749,4759|false|false|false|C0085934|Wellbutrin|Wellbutrin
Anatomy|Body Space or Junction|Hospital Course|4766,4770|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|4766,4770|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|4766,4770|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|4766,4770|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Idea or Concept|Hospital Course|4779,4782|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|4779,4782|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Body Substance|Hospital Course|4785,4794|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|4785,4794|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|4785,4794|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|4785,4794|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|4785,4806|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|4795,4806|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|4795,4806|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|Hospital Course|4795,4806|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Hospital Course|4811,4820|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|Hospital Course|4811,4820|false|false|false|C0001927|albuterol|Albuterol
Drug|Organic Chemical|Hospital Course|4811,4828|false|false|false|C0543495|albuterol sulfate|Albuterol Sulfate
Drug|Pharmacologic Substance|Hospital Course|4811,4828|false|false|false|C0543495|albuterol sulfate|Albuterol Sulfate
Drug|Element, Ion, or Isotope|Hospital Course|4821,4828|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Inorganic Chemical|Hospital Course|4821,4828|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Pharmacologic Substance|Hospital Course|4821,4828|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Disorder|Disease or Syndrome|Hospital Course|4846,4849|false|false|false|C0015458|Facial Hemiatrophy|HFA
Procedure|Diagnostic Procedure|Hospital Course|4846,4849|false|false|false|C0430649|High frequency audiometry|HFA
Drug|Biomedical or Dental Material|Hospital Course|4850,4857|false|false|false|C1112870|Aerosol Dose Form|Aerosol
Finding|Functional Concept|Hospital Course|4858,4865|false|false|false|C4319647|Inhaler (unit of presentation)|Inhaler
Finding|Functional Concept|Hospital Course|4885,4895|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Finding|Organism Function|Hospital Course|4885,4895|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Finding|Sign or Symptom|Hospital Course|4931,4939|false|false|false|C0043144|Wheezing|wheezing
Attribute|Clinical Attribute|Hospital Course|4941,4960|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|Hospital Course|4941,4960|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|Hospital Course|4954,4960|false|false|false|C0225386|Breath|breath
Drug|Organic Chemical|Hospital Course|4967,4978|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Hospital Course|4967,4978|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Biomedical or Dental Material|Hospital Course|4997,5004|false|false|false|C1112870|Aerosol Dose Form|Aerosol
Finding|Functional Concept|Hospital Course|5024,5034|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Finding|Organism Function|Hospital Course|5024,5034|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Disorder|Mental or Behavioral Dysfunction|Hospital Course|5035,5038|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5035,5038|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|5035,5038|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|5035,5038|false|false|false|C1332410|BID gene|BID
Finding|Finding|Hospital Course|5040,5047|false|false|false|C4035627|2 times|2 times
Disorder|Disease or Syndrome|Hospital Course|5042,5047|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|Hospital Course|5050,5053|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|5050,5053|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|Hospital Course|5061,5070|false|false|false|C0030049|oxycodone|Oxycodone
Drug|Pharmacologic Substance|Hospital Course|5061,5070|false|false|false|C0030049|oxycodone|Oxycodone
Procedure|Laboratory Procedure|Hospital Course|5061,5070|false|false|false|C0524222|Oxycodone measurement|Oxycodone
Drug|Pharmacologic Substance|Hospital Course|5061,5084|false|false|false|C0717368|acetaminophen / oxycodone|Oxycodone-Acetaminophen
Drug|Organic Chemical|Hospital Course|5071,5084|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Hospital Course|5071,5084|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Procedure|Laboratory Procedure|Hospital Course|5071,5084|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Drug|Biomedical or Dental Material|Hospital Course|5092,5098|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|5108,5115|false|false|false|C0039225|Tablet Dosage Form|Tablets
Attribute|Clinical Attribute|Hospital Course|5154,5158|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|5154,5158|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|5154,5158|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Biomedical or Dental Material|Hospital Course|5169,5175|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|Hospital Course|5180,5187|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|5195,5203|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|Hospital Course|5195,5203|false|false|false|C1692318|docusate|Docusate
Drug|Organic Chemical|Hospital Course|5195,5210|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|Hospital Course|5195,5210|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|Hospital Course|5204,5210|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|5204,5210|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|5204,5210|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Finding|Physiologic Function|Hospital Course|5204,5210|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|5204,5210|false|false|false|C0337443|Sodium measurement|Sodium
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5218,5225|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|5218,5225|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|5218,5225|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5239,5246|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|5239,5246|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|5239,5246|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Disorder|Mental or Behavioral Dysfunction|Hospital Course|5250,5253|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5250,5253|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|5250,5253|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|5250,5253|false|false|false|C1332410|BID gene|BID
Disorder|Disease or Syndrome|Hospital Course|5258,5263|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|Hospital Course|5266,5269|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|5266,5269|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5281,5288|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|5281,5288|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|5281,5288|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Finding|Idea or Concept|Hospital Course|5293,5300|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|5308,5319|false|false|false|C0074554|simvastatin|Simvastatin
Drug|Pharmacologic Substance|Hospital Course|5308,5319|false|false|false|C0074554|simvastatin|Simvastatin
Drug|Biomedical or Dental Material|Hospital Course|5326,5332|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|5346,5352|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Intellectual Product|Hospital Course|5356,5360|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|Hospital Course|5356,5366|false|false|false|C3537736|Once A Day|once a day
Finding|Idea or Concept|Hospital Course|5363,5366|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|5363,5366|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Biomedical or Dental Material|Hospital Course|5377,5383|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|Hospital Course|5388,5395|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|5403,5412|false|false|false|C0040805|trazodone|Trazodone
Drug|Pharmacologic Substance|Hospital Course|5403,5412|false|false|false|C0040805|trazodone|Trazodone
Drug|Biomedical or Dental Material|Hospital Course|5420,5426|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|5440,5446|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Organic Chemical|Hospital Course|5467,5477|false|false|false|C0085934|Wellbutrin|Wellbutrin
Drug|Pharmacologic Substance|Hospital Course|5467,5477|false|false|false|C0085934|Wellbutrin|Wellbutrin
Drug|Biomedical or Dental Material|Hospital Course|5484,5490|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|5504,5510|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|Hospital Course|5522,5525|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|5522,5525|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Body Substance|Hospital Course|5532,5541|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|5532,5541|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|5532,5541|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|5532,5541|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|5532,5553|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|5532,5553|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|5542,5553|false|false|false|C2926604||Disposition
Procedure|Health Care Activity|Hospital Course|5542,5553|false|false|false|C0184758|Patient disposition|Disposition
Finding|Idea or Concept|Hospital Course|5555,5559|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|5555,5559|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|5555,5559|false|false|false|C1553498|home health encounter|Home
Finding|Body Substance|Hospital Course|5562,5571|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|5562,5571|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|5562,5571|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|5562,5571|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|5562,5581|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|5572,5581|false|false|false|C0945731||Diagnosis
Finding|Classification|Hospital Course|5572,5581|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|5572,5581|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|5572,5581|false|false|false|C0011900|Diagnosis|Diagnosis
Finding|Finding|Hospital Course|5583,5587|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|High
Finding|Idea or Concept|Hospital Course|5583,5587|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|High
Finding|Intellectual Product|Hospital Course|5583,5587|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|High
Finding|Finding|Hospital Course|5583,5593|false|false|false|C0205082;C4554016|Enneking High Surgical Grade;Severe (severity modifier)|High grade
Finding|Intellectual Product|Hospital Course|5583,5593|false|false|false|C0205082;C4554016|Enneking High Surgical Grade;Severe (severity modifier)|High grade
Finding|Classification|Hospital Course|5588,5593|false|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|grade
Finding|Finding|Hospital Course|5588,5593|false|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|grade
Anatomy|Body Location or Region|Hospital Course|5594,5605|false|false|false|C0021852;C4319010|Abdomen>Small bowel;Intestines, Small|small bowel
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5594,5605|false|false|false|C0021852;C4319010|Abdomen>Small bowel;Intestines, Small|small bowel
Disorder|Disease or Syndrome|Hospital Course|5594,5617|false|false|false|C0235329|Small bowel obstruction|small bowel obstruction
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5600,5605|false|false|false|C0021853|Intestines|bowel
Disorder|Disease or Syndrome|Hospital Course|5600,5617|false|false|false|C0021843|Intestinal Obstruction|bowel obstruction
Finding|Finding|Hospital Course|5606,5617|false|false|false|C0028778|Obstruction|obstruction
Finding|Intellectual Product|Discharge Condition|5658,5664|false|false|false|C1547311|Patient Condition Code - Stable|stable
Finding|Daily or Recreational Activity|Discharge Condition|5679,5691|false|false|false|C0184625||regular diet
Drug|Food|Discharge Condition|5687,5691|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Finding|Functional Concept|Discharge Condition|5687,5691|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|Discharge Condition|5687,5691|false|false|false|C0012159|Diet therapy|diet
Anatomy|Body Part, Organ, or Organ Component|Discharge Condition|5700,5705|false|false|false|C0021853|Intestines|bowel
Finding|Organism Function|Discharge Condition|5707,5716|false|false|false|C0026649|Movement|movements
Attribute|Clinical Attribute|Discharge Condition|5727,5731|false|false|false|C2598155||pain
Finding|Functional Concept|Discharge Condition|5727,5731|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Condition|5727,5731|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|Discharge Condition|5727,5739|false|false|false|C5548091|Demonstrates adequate pain control|pain control
Procedure|Therapeutic or Preventive Procedure|Discharge Condition|5727,5739|false|false|false|C0002766;C1304888|Pain control;Pain management (procedure)|pain control
Drug|Organic Chemical|Discharge Condition|5732,5739|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Pharmacologic Substance|Discharge Condition|5732,5739|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Substance|Discharge Condition|5732,5739|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Finding|Conceptual Entity|Discharge Condition|5732,5739|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Functional Concept|Discharge Condition|5732,5739|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Idea or Concept|Discharge Condition|5732,5739|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Intellectual Product|Discharge Instructions|5784,5790|false|false|false|C2348314|Doctor - Title|doctor
Finding|Intellectual Product|Discharge Instructions|5794,5812|false|false|false|C1549435;C1549986|Nurse Practitioner - Procedure Practitioner Identifier Code Type;nurse practitioner Degree/license/certificate|nurse practitioner
Finding|Finding|Discharge Instructions|5831,5840|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Finding|Idea or Concept|Discharge Instructions|5831,5840|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Finding|Intellectual Product|Discharge Instructions|5831,5840|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Finding|Pathologic Function|Discharge Instructions|5831,5840|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Phenomenon|Phenomenon or Process|Discharge Instructions|5831,5840|false|false|false|C0013956|Emergency Situation|Emergency
Procedure|Health Care Activity|Discharge Instructions|5831,5840|false|false|false|C1553500|emergency encounter|Emergency
Finding|Idea or Concept|Discharge Instructions|5841,5851|false|false|false|C1547537;C1548283;C1549615|Department - Charge type;Department - No suggested values defined;Organization Unit Type - Department|Department
Finding|Finding|Discharge Instructions|5895,5898|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Discharge Instructions|5895,5898|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Anatomy|Body Location or Region|Discharge Instructions|5899,5904|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Discharge Instructions|5899,5904|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Discharge Instructions|5899,5909|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|Discharge Instructions|5899,5909|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Discharge Instructions|5905,5909|false|false|false|C2598155||pain
Finding|Functional Concept|Discharge Instructions|5905,5909|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|5905,5909|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|Discharge Instructions|5911,5919|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|Discharge Instructions|5911,5919|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|Discharge Instructions|5911,5919|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|Discharge Instructions|5911,5919|false|false|false|C0033095||pressure
Finding|Finding|Discharge Instructions|5948,5951|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|New
Finding|Idea or Concept|Discharge Instructions|5948,5951|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|New
Finding|Idea or Concept|Discharge Instructions|5955,5964|false|false|false|C1546960|Patient Outcome - Worsening|worsening
Drug|Organic Chemical|Discharge Instructions|5965,5970|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|Discharge Instructions|5965,5970|false|false|false|C3815497|Cough (guaifenesin)|cough
Finding|Sign or Symptom|Discharge Instructions|5965,5970|false|false|false|C0010200|Coughing|cough
Attribute|Clinical Attribute|Discharge Instructions|5972,5991|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|Discharge Instructions|5972,5991|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|Discharge Instructions|5985,5991|false|false|false|C0225386|Breath|breath
Finding|Sign or Symptom|Discharge Instructions|5996,6002|false|false|false|C0043144|Wheezing|wheeze
Finding|Sign or Symptom|Discharge Instructions|6017,6025|false|false|false|C0042963|Vomiting|vomiting
Drug|Substance|Discharge Instructions|6047,6053|true|false|true|C0302908|Liquid substance|fluids
Finding|Body Substance|Discharge Instructions|6047,6053|true|false|true|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|6047,6053|true|false|true|C0016286|Fluid Therapy|fluids
Attribute|Clinical Attribute|Discharge Instructions|6063,6074|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|6063,6074|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|Discharge Instructions|6063,6074|false|false|false|C4284232|Medications|medications
Disorder|Disease or Syndrome|Discharge Instructions|6094,6104|false|false|false|C0011175|Dehydration|dehydrated
Finding|Sign or Symptom|Discharge Instructions|6122,6130|false|false|false|C0042963|Vomiting|vomiting
Finding|Finding|Discharge Instructions|6132,6140|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|Discharge Instructions|6132,6140|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Idea or Concept|Discharge Instructions|6152,6159|false|false|false|C0392360|Indication of (contextual qualifier)|reasons
Finding|Finding|Discharge Instructions|6161,6166|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|Signs
Finding|Functional Concept|Discharge Instructions|6161,6166|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|Signs
Finding|Finding|Discharge Instructions|6161,6181|false|false|false|C5924540|Signs of dehydration|Signs of dehydration
Disorder|Disease or Syndrome|Discharge Instructions|6170,6181|false|false|false|C0011175;C2062903|Dehydration;dehydration (Na, H2O)|dehydration
Disorder|Injury or Poisoning|Discharge Instructions|6170,6181|false|false|false|C0011175;C2062903|Dehydration;dehydration (Na, H2O)|dehydration
Procedure|Laboratory Procedure|Discharge Instructions|6170,6181|false|false|false|C4284399|Dehydration procedure|dehydration
Disorder|Disease or Syndrome|Discharge Instructions|6190,6199|false|false|false|C0043352|Xerostomia|dry mouth
Anatomy|Body Location or Region|Discharge Instructions|6194,6199|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Discharge Instructions|6194,6199|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Attribute|Clinical Attribute|Discharge Instructions|6208,6217|false|false|false|C0232117|Pulse Rate|heartbeat
Finding|Organ or Tissue Function|Discharge Instructions|6208,6217|false|false|false|C0425583|Heart beat|heartbeat
Finding|Mental Process|Discharge Instructions|6222,6229|false|false|false|C1527305|Feelings|feeling
Finding|Sign or Symptom|Discharge Instructions|6222,6235|false|false|false|C0849959|feeling dizzy|feeling dizzy
Finding|Sign or Symptom|Discharge Instructions|6230,6235|false|false|false|C0012833|Dizziness|dizzy
Finding|Finding|Discharge Instructions|6239,6244|false|false|false|C0039070;C4554554|Faint - appearance;Syncope|faint
Finding|Sign or Symptom|Discharge Instructions|6239,6244|false|false|false|C0039070;C4554554|Faint - appearance;Syncope|faint
Disorder|Disease or Syndrome|Discharge Instructions|6270,6275|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|Discharge Instructions|6270,6275|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Drug|Substance|Discharge Instructions|6290,6298|false|false|false|C0520510|Materials|material
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|6325,6330|false|false|false|C0021853|Intestines|bowel
Finding|Organism Function|Discharge Instructions|6325,6339|false|false|false|C0011135|Defecation|bowel movement
Finding|Organism Function|Discharge Instructions|6331,6339|false|false|false|C0026649|Movement|movement
Finding|Sign or Symptom|Discharge Instructions|6358,6365|false|false|false|C0085624|Burning sensation|burning
Disorder|Disease or Syndrome|Discharge Instructions|6389,6394|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|Discharge Instructions|6389,6394|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Body Substance|Discharge Instructions|6404,6409|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Functional Concept|Discharge Instructions|6404,6409|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Intellectual Product|Discharge Instructions|6404,6409|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Body Substance|Discharge Instructions|6427,6436|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Discharge Instructions|6427,6436|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Discharge Instructions|6427,6436|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Discharge Instructions|6427,6436|false|false|false|C0030685|Patient Discharge|discharge
Attribute|Clinical Attribute|Discharge Instructions|6445,6449|false|false|false|C2598155||pain
Finding|Functional Concept|Discharge Instructions|6445,6449|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|6445,6449|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Functional Concept|Discharge Instructions|6517,6521|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|Call
Finding|Gene or Genome|Discharge Instructions|6517,6521|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|Call
Finding|Intellectual Product|Discharge Instructions|6517,6521|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|Call
Finding|Mental Process|Discharge Instructions|6517,6521|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|Call
Attribute|Clinical Attribute|Discharge Instructions|6552,6556|false|false|false|C2598155||pain
Finding|Functional Concept|Discharge Instructions|6552,6556|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|6552,6556|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|Discharge Instructions|6569,6574|false|false|false|C1457868;C1550463|Observation Interpretation - worse;Worse|worse
Finding|Idea or Concept|Discharge Instructions|6569,6574|false|false|false|C1457868;C1550463|Observation Interpretation - worse;Worse|worse
Finding|Functional Concept|Discharge Instructions|6578,6585|false|false|false|C0392747|Changing|changes
Anatomy|Body Location or Region|Discharge Instructions|6586,6594|false|false|false|C1515974|Anatomic Site|location
Finding|Intellectual Product|Discharge Instructions|6586,6594|false|false|false|C1555588|Transaction counts and value totals - location|location
Anatomy|Body Location or Region|Discharge Instructions|6613,6618|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Discharge Instructions|6613,6618|false|false|false|C0741025|Chest problem|chest
Finding|Sign or Symptom|Discharge Instructions|6648,6654|false|false|false|C0085593|Chills|chills
Finding|Finding|Discharge Instructions|6659,6664|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|Discharge Instructions|6659,6664|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Intellectual Product|Discharge Instructions|6684,6691|false|false|false|C0542560|Academic degree|degrees
Finding|Intellectual Product|Discharge Instructions|6710,6717|false|false|false|C0542560|Academic degree|degrees
Finding|Functional Concept|Discharge Instructions|6733,6739|false|false|false|C0392747|Changing|change
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|6733,6739|false|false|false|C4319952|Change - procedure|change
Finding|Functional Concept|Discharge Instructions|6733,6742|false|false|false|C0392747|Changing|change in
Finding|Functional Concept|Discharge Instructions|6748,6756|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Discharge Instructions|6748,6756|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Finding|Discharge Instructions|6765,6768|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Discharge Instructions|6765,6768|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Functional Concept|Discharge Instructions|6769,6777|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Discharge Instructions|6769,6777|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Idea or Concept|Discharge Instructions|6783,6790|false|false|false|C2699424|Concern|concern
Finding|Idea or Concept|Discharge Instructions|6824,6828|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Discharge Instructions|6824,6828|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Discharge Instructions|6824,6828|false|false|false|C1553498|home health encounter|home
Attribute|Clinical Attribute|Discharge Instructions|6829,6840|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|6829,6840|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|Discharge Instructions|6829,6840|false|false|false|C4284232|Medications|medications
Drug|Pharmacologic Substance|Discharge Instructions|6897,6907|false|false|false|C0013227|Pharmaceutical Preparations|medication
Finding|Intellectual Product|Discharge Instructions|6897,6907|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Procedure|Health Care Activity|Discharge Instructions|6922,6926|false|false|false|C1515187|Take|take
Finding|Finding|Discharge Instructions|6932,6935|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Discharge Instructions|6932,6935|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Drug|Pharmacologic Substance|Discharge Instructions|6932,6947|false|false|false|C1718097|New medications|new medications
Attribute|Clinical Attribute|Discharge Instructions|6936,6947|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|6936,6947|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|Discharge Instructions|6936,6947|false|false|false|C4284232|Medications|medications
Drug|Amino Acid, Peptide, or Protein|Discharge Instructions|6985,6989|false|false|false|C1742913|REST protein, human|rest
Drug|Biologically Active Substance|Discharge Instructions|6985,6989|false|false|false|C1742913|REST protein, human|rest
Finding|Daily or Recreational Activity|Discharge Instructions|6985,6989|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Gene or Genome|Discharge Instructions|6985,6989|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Molecular Function|Discharge Instructions|6985,6989|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Disorder|Disease or Syndrome|Discharge Instructions|7020,7025|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|Discharge Instructions|7031,7034|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Discharge Instructions|7031,7034|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Substance|Discharge Instructions|7066,7072|false|false|false|C0302908|Liquid substance|fluids
Finding|Body Substance|Discharge Instructions|7066,7072|false|false|false|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|7066,7072|false|false|false|C0016286|Fluid Therapy|fluids
Event|Activity|Discharge Instructions|7080,7087|false|false|false|C0206244|Lifting|lifting
Finding|Daily or Recreational Activity|Discharge Instructions|7089,7096|false|false|false|C3812400|Weights - exercise activity|weights
Procedure|Laboratory Procedure|Discharge Instructions|7114,7117|false|false|false|C3161851|liquid-based cytology (procedure)|lbs
Attribute|Clinical Attribute|Discharge Instructions|7149,7156|false|false|false|C5444295||surgeon
Finding|Daily or Recreational Activity|Discharge Instructions|7165,7172|false|false|false|C0004379|Automobile Driving|driving
Disorder|Injury or Poisoning|Discharge Instructions|7192,7201|false|false|false|C0337246|Contact with machinery|machinery
Attribute|Clinical Attribute|Discharge Instructions|7215,7219|false|false|false|C2598155||pain
Finding|Functional Concept|Discharge Instructions|7215,7219|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|7215,7219|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|Discharge Instructions|7221,7232|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|7221,7232|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|Discharge Instructions|7221,7232|false|false|false|C4284232|Medications|medications
Anatomy|Body Location or Region|Discharge Instructions|7235,7243|false|false|false|C2338258|Cranial incision point|Incision
Disorder|Injury or Poisoning|Discharge Instructions|7235,7243|false|false|false|C0332803|Surgical wound|Incision
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|7235,7243|false|false|false|C0184898|Surgical incisions|Incision
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|7235,7248|false|false|false|C0150258|Incision care|Incision Care
Event|Activity|Discharge Instructions|7244,7248|false|false|false|C1947933|care activity|Care
Finding|Finding|Discharge Instructions|7244,7248|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|Discharge Instructions|7244,7248|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|Discharge Instructions|7269,7275|false|false|false|C2348314|Doctor - Title|doctor
Finding|Intellectual Product|Discharge Instructions|7279,7297|false|false|false|C1549435;C1549986|Nurse Practitioner - Procedure Practitioner Identifier Code Type;nurse practitioner Degree/license/certificate|nurse practitioner
Attribute|Clinical Attribute|Discharge Instructions|7321,7325|false|false|false|C2598155||pain
Finding|Functional Concept|Discharge Instructions|7321,7325|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|7321,7325|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|Discharge Instructions|7327,7335|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|Discharge Instructions|7327,7335|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Disorder|Disease or Syndrome|Discharge Instructions|7337,7344|false|false|false|C0041834|Erythema|redness
Finding|Finding|Discharge Instructions|7337,7344|false|false|false|C0332575|Redness|redness
Finding|Body Substance|Discharge Instructions|7349,7357|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Finding|Sign or Symptom|Discharge Instructions|7349,7357|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|7349,7357|false|false|false|C0013103|Drainage procedure|drainage
Anatomy|Body Location or Region|Discharge Instructions|7367,7375|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|Discharge Instructions|7367,7375|false|false|false|C0332803|Surgical wound|incision
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|7367,7375|false|false|false|C0184898|Surgical incisions|incision
Anatomy|Body Location or Region|Discharge Instructions|7377,7381|false|false|false|C1515974|Anatomic Site|site
Finding|Intellectual Product|Discharge Instructions|7377,7381|false|false|false|C1546778||site
Procedure|Health Care Activity|Discharge Instructions|7404,7409|false|false|false|C0150141|Bathing|baths
Finding|Functional Concept|Discharge Instructions|7421,7427|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|Discharge Instructions|7421,7427|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|Discharge Instructions|7421,7430|false|false|false|C0589120|Follow-up status|follow-up
Procedure|Health Care Activity|Discharge Instructions|7421,7430|false|false|false|C1522577|follow-up|follow-up
Event|Activity|Discharge Instructions|7431,7442|false|false|false|C0003629|Appointments|appointment
Procedure|Health Care Activity|Discharge Instructions|7471,7479|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|7471,7479|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Disorder|Injury or Poisoning|Discharge Instructions|7471,7489|false|false|false|C0332803|Surgical wound|surgical incisions
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|7471,7489|false|false|false|C0184898|Surgical incisions|surgical incisions
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|7480,7489|false|false|false|C0184898|Surgical incisions|incisions
Finding|Intellectual Product|Discharge Instructions|7497,7501|false|false|false|C1547225|Mild Severity of Illness Code|mild
Drug|Biomedical or Dental Material|Discharge Instructions|7502,7506|false|false|false|C1705308|Soap Dosage Form|soap
Finding|Finding|Discharge Instructions|7512,7516|false|false|false|C0582051|Feels warm|warm
Phenomenon|Natural Phenomenon or Process|Discharge Instructions|7512,7516|false|false|false|C0687712|warming process|warm
Drug|Inorganic Chemical|Discharge Instructions|7517,7522|false|false|false|C0043047;C1550678|Water Specimen;water|water
Drug|Pharmacologic Substance|Discharge Instructions|7517,7522|false|false|false|C0043047;C1550678|Water Specimen;water|water
Finding|Intellectual Product|Discharge Instructions|7517,7522|false|false|false|C1547961|Water - Specimen Source Codes|water
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|7517,7522|false|false|false|C0020311|Hydrotherapy|water
Disorder|Disease or Syndrome|Discharge Instructions|7531,7534|false|false|false|C0030587|Paroxysmal atrial tachycardia|pat
Drug|Organic Chemical|Discharge Instructions|7531,7534|false|false|false|C2825250|Fenamole|pat
Drug|Pharmacologic Substance|Discharge Instructions|7531,7534|false|false|false|C2825250|Fenamole|pat
Finding|Molecular Function|Discharge Instructions|7531,7534|false|false|false|C2247344;C2247346;C2248827|aspartate-prephenate aminotransferase activity;glutamate-prephenate aminotransferase activity;protein acetyltransferase activity|pat
Procedure|Diagnostic Procedure|Discharge Instructions|7531,7534|false|false|false|C3897364|Thermoacoustic Computed Tomography|pat
Event|Governmental or Regulatory Activity|Discharge Instructions|7539,7543|false|false|false|C1510751|Academic Research Enhancement Awards|area
Finding|Functional Concept|Discharge Instructions|7601,7607|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|Discharge Instructions|7601,7607|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|Discharge Instructions|7601,7610|false|false|false|C0589120|Follow-up status|follow-up
Procedure|Health Care Activity|Discharge Instructions|7601,7610|false|false|false|C1522577|follow-up|follow-up
Event|Activity|Discharge Instructions|7612,7623|false|false|false|C0003629|Appointments|appointment
Finding|Finding|Discharge Instructions|7681,7684|false|false|false|C5939094|Own|own
Finding|Finding|Discharge Instructions|7731,7744|false|false|false|C0241311|post operative (finding)|after surgery
Finding|Finding|Discharge Instructions|7737,7744|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|Discharge Instructions|7737,7744|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|Discharge Instructions|7737,7744|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|7737,7744|false|false|false|C0543467|Operative Surgical Procedures|surgery
Anatomy|Body Location or Region|Discharge Instructions|7767,7771|false|false|false|C1515974|Anatomic Site|site
Finding|Intellectual Product|Discharge Instructions|7767,7771|false|false|false|C1546778||site
Finding|Idea or Concept|Discharge Instructions|7778,7781|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Discharge Instructions|7778,7781|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Finding|Discharge Instructions|7786,7791|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|Discharge Instructions|7786,7791|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Disorder|Disease or Syndrome|Discharge Instructions|7795,7804|false|false|false|C0009450|Communicable Diseases|infection
Finding|Pathologic Function|Discharge Instructions|7795,7804|false|false|false|C3714514|Infection|infection
Disorder|Disease or Syndrome|Discharge Instructions|7817,7824|false|false|false|C0041834|Erythema|redness
Finding|Finding|Discharge Instructions|7817,7824|false|false|false|C0332575|Redness|redness
Attribute|Clinical Attribute|Discharge Instructions|7828,7832|false|false|false|C2598155||pain
Finding|Functional Concept|Discharge Instructions|7828,7832|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|7828,7832|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|Discharge Instructions|7834,7842|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|Discharge Instructions|7834,7842|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Phenomenon|Natural Phenomenon or Process|Discharge Instructions|7844,7848|false|false|false|C0028884|Odors|odor
Finding|Finding|Discharge Instructions|7860,7866|false|false|false|C4554530|Bloody|bloody
Procedure|Health Care Activity|Discharge Instructions|7871,7879|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|7880,7892|false|false|false|C3263700||Instructions
Finding|Intellectual Product|Discharge Instructions|7880,7892|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

