 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Procedure|Health Care Activity|SIMPLE_SEGMENT|45,54|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|45,59|false|false|false|C2598112||Admission Date
Finding|Body Substance|SIMPLE_SEGMENT|79,88|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|79,88|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|79,88|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|79,88|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|79,93|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|111,116|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|111,116|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|111,116|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|135,138|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|135,138|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|135,138|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|135,138|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|135,138|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|146,153|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|146,153|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Attribute|Clinical Attribute|SIMPLE_SEGMENT|167,176|false|false|false|C1717415||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|167,176|false|false|false|C0020517|Hypersensitivity|Allergies
Attribute|Clinical Attribute|SIMPLE_SEGMENT|188,197|false|false|false|C1717415||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|188,197|false|false|false|C0020517|Hypersensitivity|Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|200,222|true|false|false|C0041755|Adverse reaction to drug|Adverse Drug Reactions
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|208,212|false|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|Drug
Finding|Finding|SIMPLE_SEGMENT|208,212|false|false|false|C0740721|Drug problem|Drug
Finding|Pathologic Function|SIMPLE_SEGMENT|208,222|true|false|false|C0041755|Adverse reaction to drug|Drug Reactions
Finding|Functional Concept|SIMPLE_SEGMENT|225,234|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|SIMPLE_SEGMENT|243,258|false|false|false|C0277786|Chief complaint (finding)|Chief Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|249,258|false|false|false|C3864418||Complaint
Finding|Finding|SIMPLE_SEGMENT|249,258|false|false|false|C5441521|Complaint (finding)|Complaint
Finding|Organism Function|SIMPLE_SEGMENT|268,274|false|false|false|C0037817|Speech|speech
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|268,274|false|false|false|C0846595|Speech assessment|speech
Finding|Classification|SIMPLE_SEGMENT|277,282|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|SIMPLE_SEGMENT|283,291|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|283,291|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|295,313|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|304,313|false|false|false|C0945766||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|304,313|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|304,313|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|304,313|false|false|false|C0184661|Interventional procedure|Procedure
Finding|Conceptual Entity|SIMPLE_SEGMENT|322,329|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|322,329|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|322,329|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|322,332|false|false|false|C0262926|Medical History|History of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|322,348|false|false|false|C0488508||History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|322,348|false|false|false|C0262512|History of present illness (finding)|History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|333,340|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Idea or Concept|SIMPLE_SEGMENT|333,340|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Finding|SIMPLE_SEGMENT|333,348|false|false|false|C4264312|Present illness|Present Illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|341,348|false|false|false|C0221423|Illness (finding)|Illness
Finding|Idea or Concept|SIMPLE_SEGMENT|354,358|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|SIMPLE_SEGMENT|354,358|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Functional Concept|SIMPLE_SEGMENT|363,368|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|393,399|false|false|false|C0018792|Heart Atrium|Atrial
Attribute|Clinical Attribute|SIMPLE_SEGMENT|393,412|false|false|false|C2926591||Atrial fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|393,412|false|false|false|C0004238|Atrial Fibrillation|Atrial fibrillation
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|393,412|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Atrial fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|400,412|false|false|false|C0232197|Fibrillation|fibrillation
Drug|Organic Chemical|SIMPLE_SEGMENT|417,424|false|false|false|C3530466|Eliquis|Eliquis
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|417,424|false|false|false|C3530466|Eliquis|Eliquis
Finding|Intellectual Product|SIMPLE_SEGMENT|431,435|false|false|false|C1720092|Once - dosing instruction fragment|once
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|444,456|false|false|false|C0020538|Hypertensive disease|hypertension
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|458,472|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|hyperlipidemia
Finding|Finding|SIMPLE_SEGMENT|458,472|false|false|false|C0428465|Serum lipids high (finding)|hyperlipidemia
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|474,477|false|false|false|C0262212|Choroidal fissure|CHF
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|474,477|false|false|false|C0018802|Congestive heart failure|CHF
Finding|Functional Concept|SIMPLE_SEGMENT|490,498|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|SIMPLE_SEGMENT|490,498|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|SIMPLE_SEGMENT|490,498|false|false|false|C4706767|Transfer (immobility management)|transfer
Finding|Intellectual Product|SIMPLE_SEGMENT|522,527|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Intellectual Product|SIMPLE_SEGMENT|522,533|false|false|false|C1272517|Sudden onset (contextual qualifier) (qualifier value)|acute onset
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|535,545|false|false|false|C0013362|Dysarthria|dysarthria
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|550,553|false|false|false|C3813556|Cancer/Testis Antigen|CTA
Finding|Gene or Genome|SIMPLE_SEGMENT|550,553|false|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|550,553|false|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Finding|Finding|SIMPLE_SEGMENT|561,569|false|false|false|C0332149|Possible|possible
Finding|Idea or Concept|SIMPLE_SEGMENT|570,577|false|true|false|C1550516|Target Awareness - partial|partial
Finding|Pathologic Function|SIMPLE_SEGMENT|578,586|false|true|false|C0087086;C0302148|Blood Clot;Thrombus|thrombus
Finding|Pathologic Function|SIMPLE_SEGMENT|590,598|false|false|false|C1261287|Stenosis|stenosis
Event|Activity|SIMPLE_SEGMENT|612,620|false|false|false|C2919031|Division (action)|division
Finding|Idea or Concept|SIMPLE_SEGMENT|612,620|false|false|false|C1547541|Organization Unit Type - Division|division
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|612,620|false|false|false|C0152060;C1293097|Division (surgical procedure);Transection (procedure)|division
Event|Activity|SIMPLE_SEGMENT|660,670|false|false|false|C1283169||monitoring
Procedure|Health Care Activity|SIMPLE_SEGMENT|660,670|false|false|false|C0150369|Preventive monitoring|monitoring
Finding|Finding|SIMPLE_SEGMENT|675,683|false|false|false|C0332149|Possible|possible
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|684,696|false|false|false|C0162578|Thrombectomy|thrombectomy
Finding|Functional Concept|SIMPLE_SEGMENT|704,708|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|704,708|false|false|false|C0582103|Medical Examination|exam
Finding|Conceptual Entity|SIMPLE_SEGMENT|728,735|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|728,735|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|728,735|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Body Substance|SIMPLE_SEGMENT|750,757|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|750,757|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|750,757|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Body Substance|SIMPLE_SEGMENT|783,790|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|783,790|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|783,790|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|837,843|false|false|false|C4048877|Dinner|dinner
Finding|Intellectual Product|SIMPLE_SEGMENT|861,865|false|false|false|C1720594|Then - dosing instruction fragment|then
Finding|Finding|SIMPLE_SEGMENT|945,949|false|false|false|C5575035|Well (answer to question)|well
Finding|Intellectual Product|SIMPLE_SEGMENT|971,975|false|false|false|C1720594|Then - dosing instruction fragment|Then
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|988,991|false|false|false|C0029121|Oppositional Defiant Disorder|odd
Finding|Gene or Genome|SIMPLE_SEGMENT|988,991|false|false|false|C1415068;C1418191|GJA1 gene;OSR1 gene|odd
Finding|Finding|SIMPLE_SEGMENT|992,1001|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|992,1001|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|SIMPLE_SEGMENT|992,1001|false|false|false|C2229507|sensory exam|sensation
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1028,1032|false|false|false|C0446516|Upper arm|arms
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1028,1032|false|false|false|C5782111||arms
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1028,1032|false|false|false|C0206655|Alveolar rhabdomyosarcoma|arms
Finding|Gene or Genome|SIMPLE_SEGMENT|1028,1032|false|false|false|C2681631;C5575339|Adherence to Refills and Medications Scale;KIDINS220 gene|arms
Finding|Intellectual Product|SIMPLE_SEGMENT|1028,1032|false|false|false|C2681631;C5575339|Adherence to Refills and Medications Scale;KIDINS220 gene|arms
Finding|Intellectual Product|SIMPLE_SEGMENT|1138,1142|false|false|false|C1720594|Then - dosing instruction fragment|Then
Finding|Classification|SIMPLE_SEGMENT|1149,1155|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|1149,1155|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|1149,1155|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|1149,1155|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Finding|SIMPLE_SEGMENT|1211,1215|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|1211,1215|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|1211,1215|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Finding|SIMPLE_SEGMENT|1250,1254|false|false|false|C1299581|Able (qualifier value)|able
Finding|Gene or Genome|SIMPLE_SEGMENT|1284,1289|false|false|false|C1424898|RXFP2 gene|great
Finding|Finding|SIMPLE_SEGMENT|1290,1300|false|false|false|C1299586|Has difficulty doing (qualifier value)|difficulty
Finding|Finding|SIMPLE_SEGMENT|1333,1340|false|false|false|C3888388|Usually|usually
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1373,1377|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1373,1377|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|1373,1377|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1373,1377|false|false|false|C0562271|Examination of knee joint|knee
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1373,1389|false|false|false|C5575606||knee replacement
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1373,1389|false|false|false|C0086511|Knee Replacement Arthroplasty|knee replacement
Finding|Functional Concept|SIMPLE_SEGMENT|1378,1389|false|false|false|C0559956|Replacement|replacement
Procedure|Health Care Activity|SIMPLE_SEGMENT|1378,1389|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|replacement
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1378,1389|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|replacement
Finding|Idea or Concept|SIMPLE_SEGMENT|1459,1465|false|false|false|C1550031|Unlock|unlock
Finding|Idea or Concept|SIMPLE_SEGMENT|1480,1488|false|false|false|C1546466|Problems - What subject filter|problems
Finding|Classification|SIMPLE_SEGMENT|1500,1506|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|1500,1506|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|1500,1506|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|1500,1506|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Finding|SIMPLE_SEGMENT|1524,1534|false|false|false|C1299586|Has difficulty doing (qualifier value)|difficulty
Finding|Idea or Concept|SIMPLE_SEGMENT|1580,1584|false|false|false|C1705313|Term (lexical)|word
Finding|Finding|SIMPLE_SEGMENT|1585,1592|true|false|false|C0037088;C0243095;C2825141|Experimental Finding;Finding;Signs and Symptoms|finding
Finding|Sign or Symptom|SIMPLE_SEGMENT|1585,1592|true|false|false|C0037088;C0243095;C2825141|Experimental Finding;Finding;Signs and Symptoms|finding
Finding|Finding|SIMPLE_SEGMENT|1594,1604|false|false|false|C1299586|Has difficulty doing (qualifier value)|difficulty
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1643,1649|false|false|true|C5890614||person
Finding|Intellectual Product|SIMPLE_SEGMENT|1643,1649|false|false|true|C1522390|Person Info|person
Finding|Finding|SIMPLE_SEGMENT|1659,1667|false|false|false|C3843660|Too much|too much
Finding|Finding|SIMPLE_SEGMENT|1663,1667|false|false|false|C4281574|Much|much
Finding|Mental Process|SIMPLE_SEGMENT|1743,1748|false|false|false|C0004448|Awareness|aware
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|1756,1766|false|false|false|C0013362|Dysarthria|dysarthria
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1822,1828|false|false|false|C0038454|Cerebrovascular accident|stroke
Finding|Finding|SIMPLE_SEGMENT|1822,1828|false|false|false|C5977286|Stroke (heart beat)|stroke
Finding|Intellectual Product|SIMPLE_SEGMENT|1830,1834|false|false|false|C1720594|Then - dosing instruction fragment|Then
Finding|Finding|SIMPLE_SEGMENT|1945,1949|false|false|false|C1299581|Able (qualifier value)|able
Finding|Functional Concept|SIMPLE_SEGMENT|2013,2019|false|false|false|C0234621|Visual|visual
Finding|Finding|SIMPLE_SEGMENT|2013,2027|true|false|false|C0750280|Visual changes|visual changes
Finding|Functional Concept|SIMPLE_SEGMENT|2020,2027|true|false|false|C0392747|Changing|changes
Finding|Finding|SIMPLE_SEGMENT|2032,2040|true|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Sign or Symptom|SIMPLE_SEGMENT|2032,2040|true|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2045,2053|false|false|false|C0030554|Paresthesia|tingling
Finding|Sign or Symptom|SIMPLE_SEGMENT|2045,2053|false|false|false|C2242996|Has tingling sensation|tingling
Finding|Sign or Symptom|SIMPLE_SEGMENT|2068,2076|true|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Finding|Finding|SIMPLE_SEGMENT|2121,2125|false|false|false|C1299581|Able (qualifier value)|able
Event|Activity|SIMPLE_SEGMENT|2153,2158|true|false|false|C5966184|Issue (action)|issue
Finding|Finding|SIMPLE_SEGMENT|2153,2158|true|false|false|C0033213;C1706387|Issue (document);Problem|issue
Finding|Intellectual Product|SIMPLE_SEGMENT|2153,2158|true|false|false|C0033213;C1706387|Issue (document);Problem|issue
Finding|Finding|SIMPLE_SEGMENT|2173,2178|false|false|false|C0392703|Shakes|shaky
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|2201,2204|false|false|false|C0015063|Ethyl Methanesulfonate|EMS
Drug|Organic Chemical|SIMPLE_SEGMENT|2201,2204|false|false|false|C0015063|Ethyl Methanesulfonate|EMS
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2201,2204|false|false|false|C0015063|Ethyl Methanesulfonate|EMS
Finding|Gene or Genome|SIMPLE_SEGMENT|2201,2204|false|false|false|C5203240|EMSLR gene|EMS
Procedure|Health Care Activity|SIMPLE_SEGMENT|2201,2204|false|false|false|C0013961|Emergency Medical Services|EMS
Finding|Intellectual Product|SIMPLE_SEGMENT|2218,2223|false|false|false|C1697238|NIH stroke scale|NIHSS
Finding|Organism Function|SIMPLE_SEGMENT|2243,2249|false|false|false|C0037817|Speech|speech
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2243,2249|false|false|false|C0846595|Speech assessment|speech
Finding|Functional Concept|SIMPLE_SEGMENT|2284,2292|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|2284,2292|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Organism Function|SIMPLE_SEGMENT|2370,2376|false|false|false|C0037817|Speech|speech
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2370,2376|false|false|false|C0846595|Speech assessment|speech
Finding|Idea or Concept|SIMPLE_SEGMENT|2417,2422|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Intellectual Product|SIMPLE_SEGMENT|2417,2422|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Drug|Organic Chemical|SIMPLE_SEGMENT|2440,2444|false|false|false|C0067518|N-(4-aminophenethyl)spiroperidol|naps
Finding|Finding|SIMPLE_SEGMENT|2450,2457|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|hearing
Finding|Physiologic Function|SIMPLE_SEGMENT|2450,2457|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|hearing
Finding|Intellectual Product|SIMPLE_SEGMENT|2461,2465|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|poor
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|2470,2478|false|false|false|C0168634|BaseLine dental cement|baseline
Finding|Idea or Concept|SIMPLE_SEGMENT|2470,2478|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Finding|Finding|SIMPLE_SEGMENT|2501,2508|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|hearing
Finding|Physiologic Function|SIMPLE_SEGMENT|2501,2508|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|hearing
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2509,2513|false|false|false|C0001175|Acquired Immunodeficiency Syndrome|aids
Finding|Sign or Symptom|SIMPLE_SEGMENT|2580,2587|false|false|false|C0013428|Dysuria|dysuria
Finding|Sign or Symptom|SIMPLE_SEGMENT|2612,2630|false|false|false|C0948396|Frequent headache|frequent headaches
Finding|Sign or Symptom|SIMPLE_SEGMENT|2621,2630|false|false|false|C0018681|Headache|headaches
Finding|Sign or Symptom|SIMPLE_SEGMENT|2668,2676|false|false|false|C0018681|Headache|headache
Drug|Organic Chemical|SIMPLE_SEGMENT|2702,2710|false|false|false|C0040610|tramadol|tramadol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2702,2710|false|false|false|C0040610|tramadol|tramadol
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2702,2710|false|false|false|C1266765|Tramadol measurement (procedure)|tramadol
Drug|Organic Chemical|SIMPLE_SEGMENT|2716,2729|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2716,2729|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2716,2729|false|false|false|C0373527|Acetaminophen measurement|acetaminophen
Finding|Functional Concept|SIMPLE_SEGMENT|2738,2744|false|false|false|C1948027|Couple (action)|couple
Finding|Sign or Symptom|SIMPLE_SEGMENT|2773,2782|false|false|false|C0018681|Headache|headaches
Finding|Sign or Symptom|SIMPLE_SEGMENT|2832,2840|false|false|false|C0018681|Headache|headache
Finding|Finding|SIMPLE_SEGMENT|2844,2854|false|false|false|C0240795|positional|positional
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2923,2929|false|false|false|C0944911||weight
Finding|Finding|SIMPLE_SEGMENT|2923,2929|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|SIMPLE_SEGMENT|2923,2929|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|SIMPLE_SEGMENT|2923,2929|false|false|false|C1305866|Weighing patient|weight
Finding|Finding|SIMPLE_SEGMENT|2923,2934|false|false|false|C1262477;C3540682|Losing Weight (question);Weight Loss|weight loss
Finding|Intellectual Product|SIMPLE_SEGMENT|2923,2934|false|false|false|C1262477;C3540682|Losing Weight (question);Weight Loss|weight loss
Finding|Finding|SIMPLE_SEGMENT|2930,2934|false|false|false|C5890125|Loss (adaptation)|loss
Finding|Idea or Concept|SIMPLE_SEGMENT|2965,2969|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|SIMPLE_SEGMENT|2965,2969|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Gene or Genome|SIMPLE_SEGMENT|2970,2973|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2994,2997|false|false|false|C3161851|liquid-based cytology (procedure)|lbs
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3018,3021|false|false|false|C3161851|liquid-based cytology (procedure)|lbs
Finding|Organism Function|SIMPLE_SEGMENT|3027,3035|false|false|false|C0003618|Desire for food|appetite
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3040,3045|false|false|false|C1410088|Still|still
Finding|Idea or Concept|SIMPLE_SEGMENT|3046,3050|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Finding|Sign or Symptom|SIMPLE_SEGMENT|3089,3095|false|false|false|C0020175|Hunger|hungry
Finding|Finding|SIMPLE_SEGMENT|3170,3176|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Finding|Intellectual Product|SIMPLE_SEGMENT|3170,3176|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Finding|Mental Process|SIMPLE_SEGMENT|3170,3176|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3250,3255|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|3273,3279|false|false|false|C4048877|Dinner|dinner
Finding|Classification|SIMPLE_SEGMENT|3338,3344|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|3338,3344|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|3338,3344|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|3338,3344|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Social Behavior|SIMPLE_SEGMENT|3430,3435|false|false|false|C0545082|Visit|visit
Finding|Gene or Genome|SIMPLE_SEGMENT|3457,3462|false|false|false|C4321205|MELTF-AS1 gene|plane
Finding|Finding|SIMPLE_SEGMENT|3503,3512|false|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|3503,3512|false|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Finding|Finding|SIMPLE_SEGMENT|3517,3537|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Finding|Functional Concept|SIMPLE_SEGMENT|3522,3529|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|3522,3529|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|3522,3529|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|3522,3529|false|false|false|C0199168|Medical service|Medical
Finding|Finding|SIMPLE_SEGMENT|3522,3537|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|3530,3537|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|3530,3537|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|3530,3537|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3554,3560|false|false|false|C0018792|Heart Atrium|Atrial
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3554,3573|false|false|false|C2926591||Atrial fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3554,3573|false|false|false|C0004238|Atrial Fibrillation|Atrial fibrillation
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3554,3573|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Atrial fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3561,3573|false|false|false|C0232197|Fibrillation|fibrillation
Drug|Organic Chemical|SIMPLE_SEGMENT|3577,3584|false|false|false|C3530466|Eliquis|Eliquis
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3577,3584|false|false|false|C3530466|Eliquis|Eliquis
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|3585,3588|false|false|false|C0262212|Choroidal fissure|CHF
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3585,3588|false|false|false|C0018802|Congestive heart failure|CHF
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3589,3609|false|false|false|C0020443|Hypercholesterolemia|Hypercholesterolemia
Finding|Finding|SIMPLE_SEGMENT|3589,3609|false|false|false|C1522133|Hypercholesterolemia result|Hypercholesterolemia
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3610,3622|false|false|false|C0020538|Hypertensive disease|Hypertension
Finding|Functional Concept|SIMPLE_SEGMENT|3625,3631|false|false|false|C0728831|Social|Social
Finding|Finding|SIMPLE_SEGMENT|3625,3639|false|false|false|C0424945;C3714536|Social History;Social and personal history|Social History
Finding|Conceptual Entity|SIMPLE_SEGMENT|3632,3639|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|3632,3639|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|3632,3639|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Classification|SIMPLE_SEGMENT|3645,3651|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|SIMPLE_SEGMENT|3645,3651|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|SIMPLE_SEGMENT|3645,3651|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|SIMPLE_SEGMENT|3645,3651|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Finding|SIMPLE_SEGMENT|3645,3659|false|false|false|C0241889|Family Medical History|Family History
Finding|Conceptual Entity|SIMPLE_SEGMENT|3652,3659|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|3652,3659|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|3652,3659|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Conceptual Entity|SIMPLE_SEGMENT|3661,3667|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Idea or Concept|SIMPLE_SEGMENT|3661,3667|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Finding|SIMPLE_SEGMENT|3670,3676|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|SIMPLE_SEGMENT|3670,3676|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|3688,3701|false|false|false|C0036341|Schizophrenia|schizophrenia
Finding|Idea or Concept|SIMPLE_SEGMENT|3702,3708|false|false|false|C1546508|Relationship - Mother|Mother
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|3711,3714|false|false|false|C0262212|Choroidal fissure|CHF
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3711,3714|false|false|false|C0018802|Congestive heart failure|CHF
Finding|Conceptual Entity|SIMPLE_SEGMENT|3715,3722|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Finding|Idea or Concept|SIMPLE_SEGMENT|3715,3722|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3725,3731|false|false|false|C0038454|Cerebrovascular accident|stroke
Finding|Finding|SIMPLE_SEGMENT|3725,3731|false|false|false|C5977286|Stroke (heart beat)|stroke
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3733,3740|false|false|false|C0007272|Carotid Arteries|carotid
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3733,3749|false|false|false|C0007282|Carotid Stenosis|carotid stenosis
Finding|Pathologic Function|SIMPLE_SEGMENT|3741,3749|false|false|false|C1261287|Stenosis|stenosis
Finding|Finding|SIMPLE_SEGMENT|3752,3760|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|3752,3760|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|3752,3760|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|3752,3765|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|3752,3765|false|false|false|C0031809|Physical Examination|Physical Exam
Finding|Functional Concept|SIMPLE_SEGMENT|3761,3765|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|3761,3765|false|false|false|C0582103|Medical Examination|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|3767,3776|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Finding|Functional Concept|SIMPLE_SEGMENT|3777,3781|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|SIMPLE_SEGMENT|3777,3781|false|false|false|C0582103|Medical Examination|EXAM
Finding|Classification|SIMPLE_SEGMENT|3849,3856|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|SIMPLE_SEGMENT|3849,3856|false|false|false|C3812897|General medical service|General
Finding|Finding|SIMPLE_SEGMENT|3858,3863|false|false|false|C0234422|Awake (finding)|Awake
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3892,3895|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3892,3895|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3892,3895|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|3892,3895|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3892,3895|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Finding|Finding|SIMPLE_SEGMENT|3892,3895|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3897,3902|false|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3914,3921|false|false|false|C0036410|Sclera|scleral
Finding|Finding|SIMPLE_SEGMENT|3914,3929|true|false|false|C0240962|Scleral icterus|scleral icterus
Finding|Sign or Symptom|SIMPLE_SEGMENT|3922,3929|true|false|false|C0022346|Icterus|icterus
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3937,3940|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3937,3940|false|false|false|C0026987|Myelofibrosis|MMM
Finding|Finding|SIMPLE_SEGMENT|3945,3952|true|false|false|C0221198|Lesion|lesions
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3962,3972|false|false|false|C0521367|Oropharyngeal|oropharynx
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3974,3978|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Anatomy|Cell Component|SIMPLE_SEGMENT|3974,3978|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Finding|Finding|SIMPLE_SEGMENT|3974,3978|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|Neck
Finding|Functional Concept|SIMPLE_SEGMENT|3980,3986|false|false|false|C0332254|Supple|Supple
Finding|Finding|SIMPLE_SEGMENT|3991,4006|true|false|false|C1320474|Nuchal Rigidity|nuchal rigidity
Finding|Sign or Symptom|SIMPLE_SEGMENT|3998,4006|true|false|false|C0026837|Muscle Rigidity|rigidity
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3998,4006|true|false|false|C0700109|plastic property - rigidity|rigidity
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4008,4017|false|false|false|C0024109|Lung|Pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4008,4017|false|false|false|C2707265||Pulmonary
Finding|Finding|SIMPLE_SEGMENT|4008,4017|false|false|false|C4522268|Pulmonary (intended site)|Pulmonary
Event|Occupational Activity|SIMPLE_SEGMENT|4026,4030|false|false|false|C0043227|Work|work
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|4026,4043|false|false|false|C0043229|Work of Breathing|work of breathing
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4034,4043|false|false|false|C5885990||breathing
Finding|Finding|SIMPLE_SEGMENT|4034,4043|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|SIMPLE_SEGMENT|4034,4043|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|SIMPLE_SEGMENT|4034,4043|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|SIMPLE_SEGMENT|4034,4043|false|false|false|C1160636|respiratory system process|breathing
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4045,4052|false|false|false|C0018787|Heart|Cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|4045,4052|false|false|false|C1314974|Cardiac attachment|Cardiac
Finding|Finding|SIMPLE_SEGMENT|4059,4063|false|false|false|C0582051|Feels warm|warm
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|4059,4063|false|false|false|C0687712|warming process|warm
Finding|Finding|SIMPLE_SEGMENT|4065,4069|false|false|false|C5575035|Well (answer to question)|well
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4080,4087|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4080,4087|false|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Finding|Finding|SIMPLE_SEGMENT|4080,4087|false|false|false|C0941288|Abdomen problem|Abdomen
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4089,4093|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4110,4121|false|false|false|C0015385;C0278454|All extremities;Limb structure|Extremities
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4130,4135|false|false|false|C1717255||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|4130,4135|false|false|false|C0013604|Edema|edema
Anatomy|Body System|SIMPLE_SEGMENT|4137,4141|false|false|false|C1123023;C4520765|Skin;Skin, Human|Skin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4137,4141|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|Skin
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4137,4141|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|Skin
Finding|Body Substance|SIMPLE_SEGMENT|4137,4141|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|Skin
Finding|Intellectual Product|SIMPLE_SEGMENT|4137,4141|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|Skin
Finding|Pathologic Function|SIMPLE_SEGMENT|4143,4153|false|false|false|C0013491|Ecchymosis|ecchymoses
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4159,4163|false|false|false|C0230444|Shin|shin
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4185,4189|false|false|false|C0230444|Shin|shin
Finding|Mental Process|SIMPLE_SEGMENT|4207,4213|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4207,4220|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|SIMPLE_SEGMENT|4207,4220|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4214,4220|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|4214,4220|false|false|false|C1546481|What subject filter - Status|Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4222,4227|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|4222,4227|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4222,4227|false|false|false|C0718338|Alert brand of caffeine|Alert
Finding|Finding|SIMPLE_SEGMENT|4222,4227|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|4222,4227|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|4222,4227|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Finding|SIMPLE_SEGMENT|4243,4247|false|false|false|C1299581|Able (qualifier value)|Able
Finding|Conceptual Entity|SIMPLE_SEGMENT|4258,4265|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|4258,4265|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|4258,4265|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|4297,4301|false|false|false|C1299581|Able (qualifier value)|able
Finding|Intellectual Product|SIMPLE_SEGMENT|4305,4309|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|name
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4343,4351|true|false|false|C2706915||Language
Finding|Intellectual Product|SIMPLE_SEGMENT|4343,4351|true|false|false|C0033348|Programming Languages|Language
Finding|Finding|SIMPLE_SEGMENT|4367,4373|false|false|false|C1554187|Gender Status - Intact|intact
Finding|Finding|SIMPLE_SEGMENT|4374,4384|false|false|false|C0205341;C2018025|Repeat;speech fluency repetition (physical finding)|repetition
Finding|Functional Concept|SIMPLE_SEGMENT|4374,4384|false|false|false|C0205341;C2018025|Repeat;speech fluency repetition (physical finding)|repetition
Finding|Mental Process|SIMPLE_SEGMENT|4389,4402|false|false|false|C0162340|Comprehension|comprehension
Finding|Finding|SIMPLE_SEGMENT|4411,4418|false|false|false|C0233743|Prosody|prosody
Finding|Finding|SIMPLE_SEGMENT|4453,4457|false|false|false|C1299581|Able (qualifier value)|Able
Finding|Intellectual Product|SIMPLE_SEGMENT|4461,4465|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|name
Finding|Finding|SIMPLE_SEGMENT|4471,4475|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|SIMPLE_SEGMENT|4471,4475|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|SIMPLE_SEGMENT|4471,4475|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Finding|SIMPLE_SEGMENT|4480,4483|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|SIMPLE_SEGMENT|4480,4483|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|SIMPLE_SEGMENT|4484,4493|false|false|false|C3898838;C4321352|Frequency;How Often|frequency
Finding|Finding|SIMPLE_SEGMENT|4504,4508|false|false|false|C1299581|Able (qualifier value)|Able
Finding|Finding|SIMPLE_SEGMENT|4525,4535|false|false|false|C1299586|Has difficulty doing (qualifier value)|difficulty
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|4540,4550|true|false|false|C0013362|Dysarthria|dysarthria
Finding|Finding|SIMPLE_SEGMENT|4552,4556|false|false|false|C1299581|Able (qualifier value)|Able
Anatomy|Cell Component|SIMPLE_SEGMENT|4573,4580|false|false|false|C1660780|midline cell component|midline
Finding|Idea or Concept|SIMPLE_SEGMENT|4621,4629|false|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|4621,4632|false|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|4633,4640|true|false|false|C0003635|Apraxias|apraxia
Event|Event|SIMPLE_SEGMENT|4644,4651|false|false|false|C5969868|Neglect (event)|neglect
Finding|Finding|SIMPLE_SEGMENT|4644,4651|false|false|false|C0521874|Victim of neglect (finding)|neglect
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4655,4662|false|false|false|C0037303|Bone structure of cranium|Cranial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4655,4669|false|false|false|C0010268|Cranial Nerves|Cranial Nerves
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4655,4669|false|false|false|C0004992;C0496937|Benign neoplasm of cranial nerves;Neoplasm of uncertain or unknown behavior of cranial nerves|Cranial Nerves
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4663,4669|false|false|false|C0027740|Nerve|Nerves
Finding|Finding|SIMPLE_SEGMENT|4689,4694|false|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4728,4737|false|false|false|C0028738|Nystagmus|nystagmus
Finding|Finding|SIMPLE_SEGMENT|4746,4754|false|false|false|C0036019|Saccades|saccades
Finding|Finding|SIMPLE_SEGMENT|4763,4776|false|false|false|C0518608|Social confrontation skill|confrontation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4763,4776|false|false|false|C0700282;C1444674|Confrontation;Confrontation visual field test|confrontation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4763,4776|false|false|false|C0700282;C1444674|Confrontation;Confrontation visual field test|confrontation
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4782,4788|false|false|false|C0015450|Face|Facial
Finding|Finding|SIMPLE_SEGMENT|4782,4798|false|false|false|C0517999|facial sensation|Facial sensation
Finding|Finding|SIMPLE_SEGMENT|4789,4798|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|4789,4798|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|SIMPLE_SEGMENT|4789,4798|false|false|false|C2229507|sensory exam|sensation
Finding|Finding|SIMPLE_SEGMENT|4799,4805|false|false|false|C1554187|Gender Status - Intact|intact
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4809,4814|false|false|false|C1570446|TNFSF14 protein, human|light
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4809,4814|false|false|false|C1570446|TNFSF14 protein, human|light
Finding|Finding|SIMPLE_SEGMENT|4809,4814|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Functional Concept|SIMPLE_SEGMENT|4809,4814|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Gene or Genome|SIMPLE_SEGMENT|4809,4814|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|4809,4814|false|false|false|C0023693|Light|light
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4809,4814|false|false|false|C0031765|Phototherapy|light
Finding|Physiologic Function|SIMPLE_SEGMENT|4809,4820|false|false|false|C0423553|Light touch|light touch
Finding|Mental Process|SIMPLE_SEGMENT|4815,4820|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|4815,4820|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4815,4820|false|false|false|C0152054|Therapeutic Touch|touch
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4835,4838|false|false|false|C2338708;C3496273;C3496274|Lamina VII of gray matter of spinal cord;layer VII (Cajal);lobule VII|VII
Finding|Intellectual Product|SIMPLE_SEGMENT|4835,4838|false|false|false|C0445385|Roman numeral VII|VII
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4843,4849|false|false|false|C0015450|Face|facial
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4843,4855|true|false|false|C0427055|Facial Paresis|facial droop
Finding|Finding|SIMPLE_SEGMENT|4843,4855|true|false|false|C4022719|Unilateral facial palsy|facial droop
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4857,4863|false|false|false|C0015450|Face|facial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4864,4875|false|false|false|C1995013|Set of muscles|musculature
Finding|Conceptual Entity|SIMPLE_SEGMENT|4876,4885|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Finding|SIMPLE_SEGMENT|4876,4885|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4887,4891|false|false|false|C0228488;C2327388|Cerebellar pyramis;Lamina VIII of gray matter of spinal cord|VIII
Finding|Gene or Genome|SIMPLE_SEGMENT|4887,4891|false|false|false|C0445599;C1413661|COX8A gene;Roman numeral VIII|VIII
Finding|Intellectual Product|SIMPLE_SEGMENT|4887,4891|false|false|false|C0445599;C1413661|COX8A gene;Roman numeral VIII|VIII
Finding|Finding|SIMPLE_SEGMENT|4893,4900|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|Hearing
Finding|Physiologic Function|SIMPLE_SEGMENT|4893,4900|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|Hearing
Finding|Finding|SIMPLE_SEGMENT|4901,4907|false|false|false|C1554187|Gender Status - Intact|intact
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4911,4917|false|false|false|C0016129;C0851278;C4299059|Fingers;Fingers not including thumb;Upper extremity>Finger|finger
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4918,4926|false|false|false|C1177045|Snap brand of resin|snapping
Finding|Finding|SIMPLE_SEGMENT|4950,4957|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|hearing
Finding|Physiologic Function|SIMPLE_SEGMENT|4950,4957|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|hearing
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4958,4962|false|false|false|C0001175|Acquired Immunodeficiency Syndrome|aids
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4972,4978|false|false|false|C0700374|Palate|Palate
Finding|Idea or Concept|SIMPLE_SEGMENT|5011,5019|false|false|false|C0808080|Strength (attribute)|strength
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5050,5056|false|false|false|C0040408|Tongue|Tongue
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5050,5056|false|false|false|C0153933|Benign neoplasm of tongue|Tongue
Procedure|Health Care Activity|SIMPLE_SEGMENT|5050,5056|false|false|false|C0872394|Procedure on tongue|Tongue
Anatomy|Cell Component|SIMPLE_SEGMENT|5070,5077|false|false|false|C1660780|midline cell component|midline
Finding|Idea or Concept|SIMPLE_SEGMENT|5083,5087|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Finding|Idea or Concept|SIMPLE_SEGMENT|5100,5108|false|false|false|C0808080|Strength (attribute)|Strength
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5119,5125|false|false|false|C0040408|Tongue|tongue
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5119,5125|false|false|false|C0153933|Benign neoplasm of tongue|tongue
Procedure|Health Care Activity|SIMPLE_SEGMENT|5119,5125|false|false|false|C0872394|Procedure on tongue|tongue
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5129,5134|false|false|false|C0007966|Cheek structure|cheek
Finding|Functional Concept|SIMPLE_SEGMENT|5135,5142|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|testing
Finding|Intellectual Product|SIMPLE_SEGMENT|5135,5142|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|testing
Finding|Functional Concept|SIMPLE_SEGMENT|5146,5151|false|false|false|C1513492|motor movement|Motor
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5160,5164|false|false|false|C0012173;C1337615|Bulk (conceptual);Dietary Fiber|bulk
Drug|Food|SIMPLE_SEGMENT|5160,5164|false|false|false|C0012173;C1337615|Bulk (conceptual);Dietary Fiber|bulk
Finding|Pathologic Function|SIMPLE_SEGMENT|5189,5203|true|false|false|C1504476|Pronator drift|pronator drift
Finding|Organism Function|SIMPLE_SEGMENT|5221,5230|false|false|false|C0026649|Movement|movements
Finding|Sign or Symptom|SIMPLE_SEGMENT|5240,5246|false|false|false|C0040822|Tremor|tremor
Finding|Sign or Symptom|SIMPLE_SEGMENT|5250,5259|false|false|false|C0232766|Asterixis|asterixis
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5421,5426|false|false|false|C1570446|TNFSF14 protein, human|light
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5421,5426|false|false|false|C1570446|TNFSF14 protein, human|light
Finding|Finding|SIMPLE_SEGMENT|5421,5426|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Functional Concept|SIMPLE_SEGMENT|5421,5426|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Gene or Genome|SIMPLE_SEGMENT|5421,5426|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|5421,5426|false|false|false|C0023693|Light|light
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5421,5426|false|false|false|C0031765|Phototherapy|light
Finding|Physiologic Function|SIMPLE_SEGMENT|5421,5432|false|false|false|C0423553|Light touch|light touch
Finding|Mental Process|SIMPLE_SEGMENT|5427,5432|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|5427,5432|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5427,5432|false|false|false|C0152054|Therapeutic Touch|touch
Procedure|Health Care Activity|SIMPLE_SEGMENT|5444,5455|false|false|false|C0886414|Body temperature measurement|temperature
Finding|Finding|SIMPLE_SEGMENT|5468,5477|false|false|false|C0392756;C0442797|Decreasing;Reduced|Decreased
Finding|Finding|SIMPLE_SEGMENT|5468,5493|false|false|false|C1295585|Decreased vibratory sense|Decreased vibratory sense
Finding|Organism Function|SIMPLE_SEGMENT|5478,5493|false|false|false|C0234198||vibratory sense
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|5488,5493|false|false|false|C0036658|Sensory perception|sense
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5501,5505|false|false|false|C0016504|Foot|feet
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5512,5518|false|false|false|C0003086|Ankle|ankles
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5520,5525|false|false|false|C0022417;C0392905;C1269611|Articular system;Joints|Joint
Anatomy|Body System|SIMPLE_SEGMENT|5520,5525|false|false|false|C0022417;C0392905;C1269611|Articular system;Joints|Joint
Finding|Finding|SIMPLE_SEGMENT|5520,5525|false|false|false|C0575044|Joint problem|Joint
Finding|Physiologic Function|SIMPLE_SEGMENT|5520,5540|false|false|false|C0423561|Joint position sense|Joint position sense
Finding|Organism Function|SIMPLE_SEGMENT|5526,5540|false|false|false|C0234219|Position Sense|position sense
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|5535,5540|false|false|false|C0036658|Sensory perception|sense
Finding|Finding|SIMPLE_SEGMENT|5541,5547|false|false|false|C1554187|Gender Status - Intact|intact
Finding|Gene or Genome|SIMPLE_SEGMENT|5555,5560|false|false|false|C1424898|RXFP2 gene|great
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5555,5565|false|false|false|C0018534|Hallux structure|great toes
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5561,5565|false|false|false|C0040357;C4299090|Lower extremity>Toes;Toes|toes
Finding|Mental Process|SIMPLE_SEGMENT|5570,5580|true|false|false|C0015347|Extinction, Psychological|extinction
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5584,5587|false|false|false|C0011195;C1848296|DOSAGE-SENSITIVE SEX REVERSAL;Dejerine-Sottas Disease|DSS
Drug|Organic Chemical|SIMPLE_SEGMENT|5584,5587|false|false|false|C0719637|DSS brand of docusate sodium|DSS
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5584,5587|false|false|false|C0719637|DSS brand of docusate sodium|DSS
Finding|Gene or Genome|SIMPLE_SEGMENT|5584,5587|false|false|false|C1417820;C2698419;C2698698;C5890838|MPZ wt Allele;NR0B1 gene;NR0B1 wt Allele;PMP22 wt Allele|DSS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5589,5596|false|false|false|C0015458|Facial Hemiatrophy|Romberg
Finding|Functional Concept|SIMPLE_SEGMENT|5597,5603|false|false|false|C0332197|Absent|absent
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5597,5603|false|false|false|C5237010|Expression Negative|absent
Finding|Finding|SIMPLE_SEGMENT|5607,5615|false|false|false|C0034929;C0596002|Observation of reflex;Reflex action|Reflexes
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|5607,5615|false|false|false|C0034929;C0596002|Observation of reflex;Reflex action|Reflexes
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5607,5615|false|false|false|C0436145|Examination of reflexes|Reflexes
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5620,5623|false|false|false|C0175372;C3495985|Structure of inferior brachium of corpora quadrigemina;nucleus of the brachium of the inferior colliculus|Bic
Drug|Organic Chemical|SIMPLE_SEGMENT|5620,5623|false|false|false|C0063382|imidazole mustard|Bic
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5620,5623|false|false|false|C0063382|imidazole mustard|Bic
Finding|Gene or Genome|SIMPLE_SEGMENT|5620,5623|false|false|false|C1537811;C2681931|MIR155 gene;MIR155HG gene|Bic
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5620,5623|false|false|false|C5202575|BIC Regimen|Bic
Finding|Gene or Genome|SIMPLE_SEGMENT|5626,5629|false|false|false|C0814229;C3891460|TRI-AAT9-1 gene;Temptation and Restraint Inventory|Tri
Finding|Intellectual Product|SIMPLE_SEGMENT|5626,5629|false|false|false|C0814229;C3891460|TRI-AAT9-1 gene;Temptation and Restraint Inventory|Tri
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5638,5641|false|false|false|C0030587|Paroxysmal atrial tachycardia|Pat
Drug|Organic Chemical|SIMPLE_SEGMENT|5638,5641|false|false|false|C2825250|Fenamole|Pat
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5638,5641|false|false|false|C2825250|Fenamole|Pat
Finding|Molecular Function|SIMPLE_SEGMENT|5638,5641|false|false|false|C2247344;C2247346;C2248827|aspartate-prephenate aminotransferase activity;glutamate-prephenate aminotransferase activity;protein acetyltransferase activity|Pat
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5638,5641|false|false|false|C3897364|Thermoacoustic Computed Tomography|Pat
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|5644,5647|false|false|false|C0001080|Achondroplasia|Ach
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5644,5647|false|false|false|C0001041|acetylcholine|Ach
Drug|Organic Chemical|SIMPLE_SEGMENT|5644,5647|false|false|false|C0001041|acetylcholine|Ach
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5644,5647|false|false|false|C0001041|acetylcholine|Ach
Finding|Gene or Genome|SIMPLE_SEGMENT|5644,5647|false|false|false|C0234238;C1333543;C1705145|Ache;FGFR3 gene;FGFR3 wt Allele|Ach
Finding|Sign or Symptom|SIMPLE_SEGMENT|5644,5647|false|false|false|C0234238;C1333543;C1705145|Ache;FGFR3 gene;FGFR3 wt Allele|Ach
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5714,5721|false|false|false|C0230463;C0442036|Plantar (qualifier value);Sole of Foot|Plantar
Finding|Finding|SIMPLE_SEGMENT|5722,5730|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Intellectual Product|SIMPLE_SEGMENT|5722,5730|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Mental Process|SIMPLE_SEGMENT|5722,5730|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5735,5741|false|false|false|C1879367|Flexor (Anatomical coordinate)|flexor
Finding|Functional Concept|SIMPLE_SEGMENT|5757,5769|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|Coordination
Finding|Idea or Concept|SIMPLE_SEGMENT|5757,5769|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|Coordination
Finding|Physiologic Function|SIMPLE_SEGMENT|5757,5769|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|Coordination
Finding|Mental Process|SIMPLE_SEGMENT|5774,5783|false|false|false|C0162425||intention
Finding|Sign or Symptom|SIMPLE_SEGMENT|5774,5790|true|false|false|C0234376;C4551520|Action Tremor;Intention tremor|intention tremor
Finding|Sign or Symptom|SIMPLE_SEGMENT|5784,5790|true|false|false|C0040822|Tremor|tremor
Finding|Finding|SIMPLE_SEGMENT|5796,5805|true|false|false|C0234162|Cerebellar Dysmetria|dysmetria
Drug|Organic Chemical|SIMPLE_SEGMENT|5809,5812|false|false|false|C0033228|fenofibrate|FNF
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5809,5812|false|false|false|C0033228|fenofibrate|FNF
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5837,5841|false|false|false|C0018870|Heel|heel
Finding|Finding|SIMPLE_SEGMENT|5850,5859|true|false|false|C0234162|Cerebellar Dysmetria|dysmetria
Finding|Finding|SIMPLE_SEGMENT|5861,5867|false|false|false|C1299582|Unable|Unable
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5878,5882|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5878,5882|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5878,5882|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5878,5882|false|false|false|C0562271|Examination of knee joint|knee
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5890,5894|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5890,5894|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5890,5894|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5890,5894|false|false|false|C0562271|Examination of knee joint|knee
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5890,5902|false|false|false|C0187769|Operative procedure on knee|knee surgery
Finding|Finding|SIMPLE_SEGMENT|5895,5902|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|SIMPLE_SEGMENT|5895,5902|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|SIMPLE_SEGMENT|5895,5902|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5895,5902|false|false|false|C0543467|Operative Surgical Procedures|surgery
Finding|Finding|SIMPLE_SEGMENT|5907,5911|false|false|false|C0016928|Gait|Gait
Finding|Finding|SIMPLE_SEGMENT|5913,5919|false|false|false|C1299582|Unable|unable
Finding|Body Substance|SIMPLE_SEGMENT|5933,5940|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|5933,5940|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|5933,5940|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5959,5967|false|false|false|C0168634|BaseLine dental cement|baseline
Finding|Idea or Concept|SIMPLE_SEGMENT|5959,5967|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Finding|Body Substance|SIMPLE_SEGMENT|5969,5978|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|5969,5978|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|5969,5978|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|5969,5978|false|false|false|C0030685|Patient Discharge|DISCHARGE
Finding|Functional Concept|SIMPLE_SEGMENT|5979,5983|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|SIMPLE_SEGMENT|5979,5983|false|false|false|C0582103|Medical Examination|EXAM
Finding|Idea or Concept|SIMPLE_SEGMENT|5991,5995|false|false|false|C1511726|Data|Data
Finding|Gene or Genome|SIMPLE_SEGMENT|6021,6025|false|false|false|C1823816|C1orf210 gene|Temp
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6021,6025|false|false|false|C0279848|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Temp
Finding|Finding|SIMPLE_SEGMENT|6126,6134|false|false|false|C1314680;C1705822;C2053584|Transfer Technique;delivery (history)|delivery
Finding|Functional Concept|SIMPLE_SEGMENT|6126,6134|false|false|false|C1314680;C1705822;C2053584|Transfer Technique;delivery (history)|delivery
Finding|Organism Function|SIMPLE_SEGMENT|6126,6134|false|false|false|C1314680;C1705822;C2053584|Transfer Technique;delivery (history)|delivery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6126,6134|false|false|false|C0011209|Obstetric Delivery|delivery
Finding|Classification|SIMPLE_SEGMENT|6140,6147|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|SIMPLE_SEGMENT|6140,6147|false|false|false|C3812897|General medical service|General
Finding|Finding|SIMPLE_SEGMENT|6149,6154|false|false|false|C0234422|Awake (finding)|Awake
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6183,6186|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6183,6186|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6183,6186|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|6183,6186|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6183,6186|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Finding|Finding|SIMPLE_SEGMENT|6183,6186|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6188,6193|false|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6205,6212|false|false|false|C0036410|Sclera|scleral
Finding|Finding|SIMPLE_SEGMENT|6205,6220|true|false|false|C0240962|Scleral icterus|scleral icterus
Finding|Sign or Symptom|SIMPLE_SEGMENT|6213,6220|true|false|false|C0022346|Icterus|icterus
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6228,6231|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6228,6231|false|false|false|C0026987|Myelofibrosis|MMM
Finding|Finding|SIMPLE_SEGMENT|6236,6243|true|false|false|C0221198|Lesion|lesions
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6253,6263|false|false|false|C0521367|Oropharyngeal|oropharynx
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6265,6269|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Anatomy|Cell Component|SIMPLE_SEGMENT|6265,6269|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Finding|Finding|SIMPLE_SEGMENT|6265,6269|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|Neck
Finding|Functional Concept|SIMPLE_SEGMENT|6271,6277|false|false|false|C0332254|Supple|Supple
Finding|Finding|SIMPLE_SEGMENT|6282,6297|true|false|false|C1320474|Nuchal Rigidity|nuchal rigidity
Finding|Sign or Symptom|SIMPLE_SEGMENT|6289,6297|true|false|false|C0026837|Muscle Rigidity|rigidity
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|6289,6297|true|false|false|C0700109|plastic property - rigidity|rigidity
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6299,6308|false|false|false|C0024109|Lung|Pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6299,6308|false|false|false|C2707265||Pulmonary
Finding|Finding|SIMPLE_SEGMENT|6299,6308|false|false|false|C4522268|Pulmonary (intended site)|Pulmonary
Event|Occupational Activity|SIMPLE_SEGMENT|6317,6321|false|false|false|C0043227|Work|work
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|6317,6334|false|false|false|C0043229|Work of Breathing|work of breathing
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6325,6334|false|false|false|C5885990||breathing
Finding|Finding|SIMPLE_SEGMENT|6325,6334|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|SIMPLE_SEGMENT|6325,6334|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|SIMPLE_SEGMENT|6325,6334|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|SIMPLE_SEGMENT|6325,6334|false|false|false|C1160636|respiratory system process|breathing
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6336,6343|false|false|false|C0018787|Heart|Cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|6336,6343|false|false|false|C1314974|Cardiac attachment|Cardiac
Finding|Finding|SIMPLE_SEGMENT|6353,6357|false|false|false|C0582051|Feels warm|warm
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|6353,6357|false|false|false|C0687712|warming process|warm
Finding|Finding|SIMPLE_SEGMENT|6359,6363|false|false|false|C5575035|Well (answer to question)|well
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6374,6381|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6374,6381|false|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Finding|Finding|SIMPLE_SEGMENT|6374,6381|false|false|false|C0941288|Abdomen problem|Abdomen
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6383,6387|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6404,6415|false|false|false|C0015385;C0278454|All extremities;Limb structure|Extremities
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6424,6429|false|false|false|C1717255||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|6424,6429|false|false|false|C0013604|Edema|edema
Anatomy|Body System|SIMPLE_SEGMENT|6431,6435|false|false|false|C1123023;C4520765|Skin;Skin, Human|Skin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6431,6435|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|Skin
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6431,6435|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|Skin
Finding|Body Substance|SIMPLE_SEGMENT|6431,6435|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|Skin
Finding|Intellectual Product|SIMPLE_SEGMENT|6431,6435|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|Skin
Finding|Pathologic Function|SIMPLE_SEGMENT|6437,6447|false|false|false|C0013491|Ecchymosis|ecchymoses
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6453,6457|false|false|false|C0230444|Shin|shin
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6479,6483|false|false|false|C0230444|Shin|shin
Finding|Mental Process|SIMPLE_SEGMENT|6501,6507|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6501,6514|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|SIMPLE_SEGMENT|6501,6514|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6508,6514|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|6508,6514|false|false|false|C1546481|What subject filter - Status|Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6516,6521|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|6516,6521|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6516,6521|false|false|false|C0718338|Alert brand of caffeine|Alert
Finding|Finding|SIMPLE_SEGMENT|6516,6521|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|6516,6521|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|6516,6521|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6535,6541|false|false|false|C5890614||person
Finding|Intellectual Product|SIMPLE_SEGMENT|6535,6541|false|false|false|C1522390|Person Info|person
Finding|Finding|SIMPLE_SEGMENT|6557,6561|false|false|false|C1299581|Able (qualifier value)|Able
Drug|Organic Chemical|SIMPLE_SEGMENT|6565,6571|false|false|false|C0163712|Relate - vinyl resin|relate
Finding|Conceptual Entity|SIMPLE_SEGMENT|6572,6579|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|6572,6579|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|6572,6579|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6623,6631|false|false|false|C2706915||Language
Finding|Intellectual Product|SIMPLE_SEGMENT|6623,6631|false|false|false|C0033348|Programming Languages|Language
Finding|Finding|SIMPLE_SEGMENT|6647,6653|false|false|false|C1554187|Gender Status - Intact|intact
Finding|Mental Process|SIMPLE_SEGMENT|6654,6667|false|false|false|C0162340|Comprehension|comprehension
Finding|Finding|SIMPLE_SEGMENT|6676,6683|false|false|false|C0233743|Prosody|prosody
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|6721,6731|true|false|false|C0013362|Dysarthria|dysarthria
Finding|Finding|SIMPLE_SEGMENT|6733,6737|false|false|false|C1299581|Able (qualifier value)|Able
Finding|Functional Concept|SIMPLE_SEGMENT|6741,6747|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|SIMPLE_SEGMENT|6741,6747|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Anatomy|Cell Component|SIMPLE_SEGMENT|6753,6760|false|false|false|C1660780|midline cell component|midline
Finding|Idea or Concept|SIMPLE_SEGMENT|6801,6809|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|6801,6812|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|6813,6820|false|false|false|C0003635|Apraxias|apraxia
Event|Event|SIMPLE_SEGMENT|6824,6831|false|false|false|C5969868|Neglect (event)|neglect
Finding|Finding|SIMPLE_SEGMENT|6824,6831|false|false|false|C0521874|Victim of neglect (finding)|neglect
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6835,6842|false|false|false|C0037303|Bone structure of cranium|Cranial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6835,6849|false|false|false|C0010268|Cranial Nerves|Cranial Nerves
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6835,6849|false|false|false|C0004992;C0496937|Benign neoplasm of cranial nerves;Neoplasm of uncertain or unknown behavior of cranial nerves|Cranial Nerves
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6843,6849|false|false|false|C0027740|Nerve|Nerves
Finding|Finding|SIMPLE_SEGMENT|6869,6874|false|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6908,6917|false|false|false|C0028738|Nystagmus|nystagmus
Finding|Finding|SIMPLE_SEGMENT|6926,6934|false|false|false|C0036019|Saccades|saccades
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6939,6945|false|false|false|C0015450|Face|Facial
Finding|Finding|SIMPLE_SEGMENT|6939,6955|false|false|false|C0517999|facial sensation|Facial sensation
Finding|Finding|SIMPLE_SEGMENT|6946,6955|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|6946,6955|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|SIMPLE_SEGMENT|6946,6955|false|false|false|C2229507|sensory exam|sensation
Finding|Finding|SIMPLE_SEGMENT|6956,6962|false|false|false|C1554187|Gender Status - Intact|intact
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6966,6971|false|false|false|C1570446|TNFSF14 protein, human|light
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6966,6971|false|false|false|C1570446|TNFSF14 protein, human|light
Finding|Finding|SIMPLE_SEGMENT|6966,6971|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Functional Concept|SIMPLE_SEGMENT|6966,6971|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Gene or Genome|SIMPLE_SEGMENT|6966,6971|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|6966,6971|false|false|false|C0023693|Light|light
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6966,6971|false|false|false|C0031765|Phototherapy|light
Finding|Physiologic Function|SIMPLE_SEGMENT|6966,6977|false|false|false|C0423553|Light touch|light touch
Finding|Mental Process|SIMPLE_SEGMENT|6972,6977|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|6972,6977|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6972,6977|false|false|false|C0152054|Therapeutic Touch|touch
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6979,6982|false|false|false|C2338708;C3496273;C3496274|Lamina VII of gray matter of spinal cord;layer VII (Cajal);lobule VII|VII
Finding|Intellectual Product|SIMPLE_SEGMENT|6979,6982|false|false|false|C0445385|Roman numeral VII|VII
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6987,6993|false|false|false|C0015450|Face|facial
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6987,6999|true|false|false|C0427055|Facial Paresis|facial droop
Finding|Finding|SIMPLE_SEGMENT|6987,6999|true|false|false|C4022719|Unilateral facial palsy|facial droop
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7001,7007|false|false|false|C0015450|Face|facial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7008,7019|false|false|false|C1995013|Set of muscles|musculature
Finding|Conceptual Entity|SIMPLE_SEGMENT|7020,7029|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Finding|SIMPLE_SEGMENT|7020,7029|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7031,7035|false|false|false|C0228488;C2327388|Cerebellar pyramis;Lamina VIII of gray matter of spinal cord|VIII
Finding|Gene or Genome|SIMPLE_SEGMENT|7031,7035|false|false|false|C0445599;C1413661|COX8A gene;Roman numeral VIII|VIII
Finding|Intellectual Product|SIMPLE_SEGMENT|7031,7035|false|false|false|C0445599;C1413661|COX8A gene;Roman numeral VIII|VIII
Finding|Finding|SIMPLE_SEGMENT|7037,7044|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|Hearing
Finding|Physiologic Function|SIMPLE_SEGMENT|7037,7044|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|Hearing
Finding|Finding|SIMPLE_SEGMENT|7045,7051|false|false|false|C1554187|Gender Status - Intact|intact
Finding|Social Behavior|SIMPLE_SEGMENT|7055,7067|false|false|false|C0871703|conversation|conversation
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7076,7082|false|false|false|C0700374|Palate|Palate
Finding|Idea or Concept|SIMPLE_SEGMENT|7115,7123|false|false|false|C0808080|Strength (attribute)|strength
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7154,7160|false|false|false|C0040408|Tongue|Tongue
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7154,7160|false|false|false|C0153933|Benign neoplasm of tongue|Tongue
Procedure|Health Care Activity|SIMPLE_SEGMENT|7154,7160|false|false|false|C0872394|Procedure on tongue|Tongue
Anatomy|Cell Component|SIMPLE_SEGMENT|7174,7181|false|false|false|C1660780|midline cell component|midline
Finding|Idea or Concept|SIMPLE_SEGMENT|7187,7191|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Finding|Functional Concept|SIMPLE_SEGMENT|7206,7211|false|false|false|C1513492|motor movement|Motor
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7220,7224|false|false|false|C0012173;C1337615|Bulk (conceptual);Dietary Fiber|bulk
Drug|Food|SIMPLE_SEGMENT|7220,7224|false|false|false|C0012173;C1337615|Bulk (conceptual);Dietary Fiber|bulk
Finding|Pathologic Function|SIMPLE_SEGMENT|7249,7263|true|false|false|C1504476|Pronator drift|pronator drift
Finding|Organism Function|SIMPLE_SEGMENT|7281,7290|false|false|false|C0026649|Movement|movements
Finding|Sign or Symptom|SIMPLE_SEGMENT|7300,7306|false|false|false|C0040822|Tremor|tremor
Finding|Sign or Symptom|SIMPLE_SEGMENT|7310,7319|false|false|false|C0232766|Asterixis|asterixis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7330,7334|false|false|false|C0224234|Structure of deltoid muscle|Delt
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7336,7339|false|false|false|C0175372;C3495985|Structure of inferior brachium of corpora quadrigemina;nucleus of the brachium of the inferior colliculus|Bic
Drug|Organic Chemical|SIMPLE_SEGMENT|7336,7339|false|false|false|C0063382|imidazole mustard|Bic
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7336,7339|false|false|false|C0063382|imidazole mustard|Bic
Finding|Gene or Genome|SIMPLE_SEGMENT|7336,7339|false|false|false|C1537811;C2681931|MIR155 gene;MIR155HG gene|Bic
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7336,7339|false|false|false|C5202575|BIC Regimen|Bic
Finding|Gene or Genome|SIMPLE_SEGMENT|7341,7344|false|false|false|C0814229;C3891460|TRI-AAT9-1 gene;Temptation and Restraint Inventory|Tri
Finding|Intellectual Product|SIMPLE_SEGMENT|7341,7344|false|false|false|C0814229;C3891460|TRI-AAT9-1 gene;Temptation and Restraint Inventory|Tri
Finding|Gene or Genome|SIMPLE_SEGMENT|7351,7354|false|false|false|C1537570;C3539626|LGR5 gene;LGR5 wt Allele|FEx
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7370,7373|false|false|false|C0030481|Tropical Spastic Paraparesis|Ham
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7370,7373|false|false|false|C1570167;C3853311|ATF7IP protein, human;Ham|Ham
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7370,7373|false|false|false|C1570167;C3853311|ATF7IP protein, human;Ham|Ham
Drug|Food|SIMPLE_SEGMENT|7370,7373|false|false|false|C1570167;C3853311|ATF7IP protein, human;Ham|Ham
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7370,7373|false|false|false|C0279477|altretamine/doxorubicin/melphalan protocol|Ham
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7379,7382|false|false|false|C0017110;C1550641;C1704673|Gas - SpecimenType;Gas Dosage Form;Gases|Gas
Drug|Chemical Viewed Structurally|SIMPLE_SEGMENT|7379,7382|false|false|false|C0017110;C1550641;C1704673|Gas - SpecimenType;Gas Dosage Form;Gases|Gas
Drug|Substance|SIMPLE_SEGMENT|7379,7382|false|false|false|C0017110;C1550641;C1704673|Gas - SpecimenType;Gas Dosage Form;Gases|Gas
Finding|Gene or Genome|SIMPLE_SEGMENT|7379,7382|false|false|false|C0596601;C1414950;C1439341;C1540252;C1546643;C2266618;C2986619;C3812826;C5890923|GALNS gene;GALNS wt Allele;GAST gene;GAST wt Allele;Gas - Specimen Source Codes;PAGR1 gene;PAGR1 wt Allele;gastrointestinal gas;germacrene-A synthase activity|Gas
Finding|Intellectual Product|SIMPLE_SEGMENT|7379,7382|false|false|false|C0596601;C1414950;C1439341;C1540252;C1546643;C2266618;C2986619;C3812826;C5890923|GALNS gene;GALNS wt Allele;GAST gene;GAST wt Allele;Gas - Specimen Source Codes;PAGR1 gene;PAGR1 wt Allele;gastrointestinal gas;germacrene-A synthase activity|Gas
Finding|Molecular Function|SIMPLE_SEGMENT|7379,7382|false|false|false|C0596601;C1414950;C1439341;C1540252;C1546643;C2266618;C2986619;C3812826;C5890923|GALNS gene;GALNS wt Allele;GAST gene;GAST wt Allele;Gas - Specimen Source Codes;PAGR1 gene;PAGR1 wt Allele;gastrointestinal gas;germacrene-A synthase activity|Gas
Finding|Sign or Symptom|SIMPLE_SEGMENT|7379,7382|false|false|false|C0596601;C1414950;C1439341;C1540252;C1546643;C2266618;C2986619;C3812826;C5890923|GALNS gene;GALNS wt Allele;GAST gene;GAST wt Allele;Gas - Specimen Source Codes;PAGR1 gene;PAGR1 wt Allele;gastrointestinal gas;germacrene-A synthase activity|Gas
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7503,7507|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|Knee
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7503,7507|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|Knee
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|7503,7507|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|Knee
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7503,7507|false|false|false|C0562271|Examination of knee joint|Knee
Finding|Finding|SIMPLE_SEGMENT|7526,7539|false|true|false|C0455610|History of surgery|prior surgery
Finding|Finding|SIMPLE_SEGMENT|7532,7539|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|SIMPLE_SEGMENT|7532,7539|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|SIMPLE_SEGMENT|7532,7539|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7532,7539|false|false|false|C0543467|Operative Surgical Procedures|surgery
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7566,7571|false|false|false|C1570446|TNFSF14 protein, human|light
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7566,7571|false|false|false|C1570446|TNFSF14 protein, human|light
Finding|Finding|SIMPLE_SEGMENT|7566,7571|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Functional Concept|SIMPLE_SEGMENT|7566,7571|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Gene or Genome|SIMPLE_SEGMENT|7566,7571|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|7566,7571|false|false|false|C0023693|Light|light
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7566,7571|false|false|false|C0031765|Phototherapy|light
Finding|Physiologic Function|SIMPLE_SEGMENT|7566,7577|false|false|false|C0423553|Light touch|light touch
Finding|Mental Process|SIMPLE_SEGMENT|7572,7577|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|7572,7577|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7572,7577|false|false|false|C0152054|Therapeutic Touch|touch
Finding|Functional Concept|SIMPLE_SEGMENT|7592,7604|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|Coordination
Finding|Idea or Concept|SIMPLE_SEGMENT|7592,7604|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|Coordination
Finding|Physiologic Function|SIMPLE_SEGMENT|7592,7604|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|Coordination
Finding|Mental Process|SIMPLE_SEGMENT|7609,7618|false|false|false|C0162425||intention
Finding|Sign or Symptom|SIMPLE_SEGMENT|7609,7625|true|false|false|C0234376;C4551520|Action Tremor;Intention tremor|intention tremor
Finding|Sign or Symptom|SIMPLE_SEGMENT|7619,7625|true|false|false|C0040822|Tremor|tremor
Finding|Finding|SIMPLE_SEGMENT|7631,7640|true|false|false|C0234162|Cerebellar Dysmetria|dysmetria
Drug|Organic Chemical|SIMPLE_SEGMENT|7644,7647|false|false|false|C0033228|fenofibrate|FNF
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7644,7647|false|false|false|C0033228|fenofibrate|FNF
Finding|Finding|SIMPLE_SEGMENT|7664,7668|false|false|false|C0016928|Gait|Gait
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7688,7696|false|false|false|C0168634|BaseLine dental cement|baseline
Finding|Idea or Concept|SIMPLE_SEGMENT|7688,7696|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7730,7735|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|7730,7735|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|7736,7739|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|7744,7747|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7744,7747|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7744,7747|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7753,7756|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7753,7756|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|7753,7756|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|7753,7756|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7762,7765|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7762,7765|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|7773,7776|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|7773,7776|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7773,7776|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7773,7776|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|7780,7783|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7780,7783|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|7780,7783|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|7780,7783|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7780,7783|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7789,7793|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7820,7823|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7840,7845|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|7840,7845|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Antibiotic|SIMPLE_SEGMENT|7861,7866|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7861,7866|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|SIMPLE_SEGMENT|7861,7866|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7871,7874|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|Eos
Finding|Gene or Genome|SIMPLE_SEGMENT|7871,7874|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|Eos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7973,7978|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|7973,7978|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7983,7986|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7983,7986|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8008,8013|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|8008,8013|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|8008,8021|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|8008,8021|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8008,8021|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8014,8021|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|8014,8021|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8014,8021|false|false|false|C0017725|glucose|Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|8014,8021|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8014,8021|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|SIMPLE_SEGMENT|8065,8069|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8065,8069|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8065,8069|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8094,8099|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|8094,8099|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8100,8105|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|SIMPLE_SEGMENT|8100,8105|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|SIMPLE_SEGMENT|8100,8105|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8100,8105|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8134,8139|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|8134,8139|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8134,8147|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8140,8147|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|8140,8147|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|8140,8147|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8140,8147|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|8140,8147|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|8140,8147|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8140,8147|false|false|false|C0201925|Calcium measurement|Calcium
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8193,8198|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|8193,8198|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8210,8213|false|false|false|C0023821|High Density Lipoproteins|HDL
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8210,8213|false|false|false|C0023821|High Density Lipoproteins|HDL
Finding|Gene or Genome|SIMPLE_SEGMENT|8210,8213|false|false|false|C3715113|HSD11B1 wt Allele|HDL
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8210,8213|false|false|false|C0392885|High density lipoprotein measurement|HDL
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8253,8258|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|8253,8258|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8260,8265|false|false|false|C0019018|Glycosylated hemoglobin A|HbA1c
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8260,8265|false|false|false|C0019018|Glycosylated hemoglobin A|HbA1c
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8260,8265|false|false|false|C0202054|Glucohemoglobin measurement|HbA1c
Finding|Gene or Genome|SIMPLE_SEGMENT|8270,8273|false|false|false|C1416571|KCNH1 gene|eAG
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8290,8295|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|8290,8295|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8319,8324|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|8319,8324|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8325,8328|false|false|false|C2708739||TSH
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8325,8328|false|false|false|C0040160|thyrotropin|TSH
Drug|Hormone|SIMPLE_SEGMENT|8325,8328|false|false|false|C0040160|thyrotropin|TSH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8325,8328|false|false|false|C0040160|thyrotropin|TSH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8325,8328|false|false|false|C0202230|Thyroid stimulating hormone measurement|TSH
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8346,8351|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|8346,8351|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Finding|Finding|SIMPLE_SEGMENT|8360,8363|false|false|false|C5848551|Neg - answer|NEG
Finding|Body Substance|SIMPLE_SEGMENT|8376,8381|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|8376,8381|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|8376,8381|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Finding|SIMPLE_SEGMENT|8376,8387|false|false|false|C0278030|Color of urine|URINE Color
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8382,8387|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|Color
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|8382,8387|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|Color
Drug|Organic Chemical|SIMPLE_SEGMENT|8388,8393|false|false|false|C4047917|Cereal plant straw|Straw
Finding|Idea or Concept|SIMPLE_SEGMENT|8401,8406|false|false|false|C1550016|Remote control command - Clear|Clear
Finding|Body Substance|SIMPLE_SEGMENT|8426,8431|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|8426,8431|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|8426,8431|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8426,8437|false|false|false|C0018965|Hematuria|URINE Blood
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8432,8437|false|false|false|C0851353|Blood and lymphatic system disorders|Blood
Finding|Body Substance|SIMPLE_SEGMENT|8432,8437|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Finding|Finding|SIMPLE_SEGMENT|8438,8441|false|false|false|C5848551|Neg - answer|NEG
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8442,8449|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|Nitrite
Drug|Inorganic Chemical|SIMPLE_SEGMENT|8442,8449|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|Nitrite
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8442,8449|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|Nitrite
Finding|Finding|SIMPLE_SEGMENT|8450,8453|false|false|false|C5848551|Neg - answer|NEG
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8454,8461|false|false|false|C0033684|Proteins|Protein
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8454,8461|false|false|false|C0033684|Proteins|Protein
Finding|Conceptual Entity|SIMPLE_SEGMENT|8454,8461|false|false|false|C1521746|Protein Info|Protein
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8454,8461|false|false|false|C0202202|Protein measurement|Protein
Finding|Finding|SIMPLE_SEGMENT|8462,8465|false|false|false|C5848551|Neg - answer|NEG
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8467,8474|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|8467,8474|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8467,8474|false|false|false|C0017725|glucose|Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|8467,8474|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8467,8474|false|false|false|C0337438|Glucose measurement|Glucose
Finding|Finding|SIMPLE_SEGMENT|8475,8478|false|false|false|C5848551|Neg - answer|NEG
Drug|Organic Chemical|SIMPLE_SEGMENT|8479,8485|false|false|false|C0022634|Ketones|Ketone
Finding|Finding|SIMPLE_SEGMENT|8486,8489|false|false|false|C5848551|Neg - answer|NEG
Finding|Finding|SIMPLE_SEGMENT|8498,8501|false|false|false|C5848551|Neg - answer|NEG
Finding|Finding|SIMPLE_SEGMENT|8510,8513|false|false|false|C5848551|Neg - answer|NEG
Finding|Finding|SIMPLE_SEGMENT|8527,8530|false|false|false|C5848551|Neg - answer|NEG
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8540,8543|false|false|false|C3813556|Cancer/Testis Antigen|CTA
Finding|Gene or Genome|SIMPLE_SEGMENT|8540,8543|false|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8540,8543|false|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Anatomy|Body Location or Region|SIMPLE_SEGMENT|8544,8548|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8544,8548|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8544,8548|false|false|false|C0362076|Problems with head|head
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8544,8548|false|false|false|C0876917|Procedure on head|head
Anatomy|Body Location or Region|SIMPLE_SEGMENT|8549,8553|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|SIMPLE_SEGMENT|8549,8553|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|SIMPLE_SEGMENT|8549,8553|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Finding|Idea or Concept|SIMPLE_SEGMENT|8558,8565|false|false|false|C0871010|Opinions|opinion
Finding|Intellectual Product|SIMPLE_SEGMENT|8572,8582|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|8572,8582|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Functional Concept|SIMPLE_SEGMENT|8599,8603|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8599,8620|false|false|false|C0226231|Structure of left vertebral artery|left vertebral artery
Finding|Pathologic Function|SIMPLE_SEGMENT|8599,8630|false|false|false|C4536452|Occlusion of left vertebral artery (disorder)|left vertebral artery occlusion
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8604,8613|false|false|false|C0549207|Bone structure of spine|vertebral
Anatomy|Body Location or Region|SIMPLE_SEGMENT|8604,8620|false|false|false|C0042559;C4695118|Head+Neck>Vertebral artery;Structure of vertebral artery|vertebral artery
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8604,8620|false|false|false|C0042559;C4695118|Head+Neck>Vertebral artery;Structure of vertebral artery|vertebral artery
Finding|Pathologic Function|SIMPLE_SEGMENT|8604,8630|false|false|false|C0265104|Vertebral artery obstruction (disorder)|vertebral artery occlusion
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8614,8620|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|SIMPLE_SEGMENT|8614,8620|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Finding|Pathologic Function|SIMPLE_SEGMENT|8614,8630|false|false|false|C0264995|Occlusion of artery (disorder)|artery occlusion
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|8621,8630|false|false|false|C0001168|Complete obstruction|occlusion
Finding|Finding|SIMPLE_SEGMENT|8621,8630|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Functional Concept|SIMPLE_SEGMENT|8621,8630|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|8621,8630|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Pathologic Function|SIMPLE_SEGMENT|8621,8630|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Idea or Concept|SIMPLE_SEGMENT|8665,8673|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|8665,8676|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Finding|Pathologic Function|SIMPLE_SEGMENT|8677,8685|true|false|false|C0022116|Ischemia|ischemia
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8677,8685|true|false|false|C4321499|Ischemia Procedure|ischemia
Finding|Finding|SIMPLE_SEGMENT|8691,8699|false|false|false|C2984079|Somewhat|Somewhat
Event|Activity|SIMPLE_SEGMENT|8714,8724|false|false|false|C0599946|Attenuation|attenuated
Finding|Functional Concept|SIMPLE_SEGMENT|8725,8729|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Finding|Social Behavior|SIMPLE_SEGMENT|8733,8741|false|false|false|C0678975|inferiority|inferior
Drug|Chemical Viewed Structurally|SIMPLE_SEGMENT|8742,8748|false|false|false|C1881507|Macromolecular Branch|branch
Finding|Idea or Concept|SIMPLE_SEGMENT|8759,8767|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|8759,8770|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|8777,8786|true|false|false|C0001168|Complete obstruction|occlusion
Finding|Finding|SIMPLE_SEGMENT|8777,8786|true|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Functional Concept|SIMPLE_SEGMENT|8777,8786|true|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|8777,8786|true|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Pathologic Function|SIMPLE_SEGMENT|8777,8786|true|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Intellectual Product|SIMPLE_SEGMENT|8795,8800|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Anatomy|Body Location or Region|SIMPLE_SEGMENT|8801,8813|false|false|false|C0524466|Intracranial|intracranial
Finding|Functional Concept|SIMPLE_SEGMENT|8801,8813|false|false|false|C1522213|Intracranial Route of Administration|intracranial
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|8814,8825|false|false|false|C0000768|Congenital Abnormality|abnormality
Finding|Finding|SIMPLE_SEGMENT|8814,8825|false|false|false|C1704258|Abnormality|abnormality
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8841,8848|false|false|false|C0881943||CT head
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8841,8848|false|false|false|C0202691|CAT scan of head|CT head
Anatomy|Body Location or Region|SIMPLE_SEGMENT|8844,8848|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8844,8848|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8844,8848|false|false|false|C0362076|Problems with head|head
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8844,8848|false|false|false|C0876917|Procedure on head|head
Finding|Gene or Genome|SIMPLE_SEGMENT|8855,8858|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8855,8858|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|SIMPLE_SEGMENT|8855,8858|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8855,8863|false|false|false|C0412674|MRI of head|MRI head
Anatomy|Body Location or Region|SIMPLE_SEGMENT|8859,8863|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8859,8863|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8859,8863|false|false|false|C0362076|Problems with head|head
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8859,8863|false|false|false|C0876917|Procedure on head|head
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|8868,8876|false|false|false|C0009924|Contrast Media|contrast
Finding|Intellectual Product|SIMPLE_SEGMENT|8877,8887|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|8877,8887|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|8895,8900|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Anatomy|Body Location or Region|SIMPLE_SEGMENT|8901,8913|false|false|false|C0524466|Intracranial|intracranial
Finding|Functional Concept|SIMPLE_SEGMENT|8901,8913|false|false|false|C1522213|Intracranial Route of Administration|intracranial
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|8914,8925|true|false|false|C0000768|Congenital Abnormality|abnormality
Finding|Finding|SIMPLE_SEGMENT|8914,8925|true|false|false|C1704258|Abnormality|abnormality
Finding|Gene or Genome|SIMPLE_SEGMENT|8945,8950|true|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Finding|Pathologic Function|SIMPLE_SEGMENT|8962,8972|false|false|false|C0021308|Infarction|infarction
Finding|Pathologic Function|SIMPLE_SEGMENT|8976,8986|false|false|false|C0019080|Hemorrhage|hemorrhage
Finding|Finding|SIMPLE_SEGMENT|9001,9005|false|false|false|C4321394|Foci|foci
Finding|Finding|SIMPLE_SEGMENT|9012,9016|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|SIMPLE_SEGMENT|9012,9016|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|SIMPLE_SEGMENT|9012,9016|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|9017,9023|false|false|false|C1710082|Signal|signal
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9041,9052|false|false|false|C0815275|Subcortical|subcortical
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9058,9086|false|false|false|C0228157|Periventricular white matter|periventricular white matter
Anatomy|Tissue|SIMPLE_SEGMENT|9074,9086|false|false|false|C0682708|White matter|white matter
Finding|Functional Concept|SIMPLE_SEGMENT|9120,9127|false|false|false|C0392747|Changing|changes
Finding|Intellectual Product|SIMPLE_SEGMENT|9135,9142|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|9135,9142|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9143,9155|false|false|false|C0225988|Structure of small blood vessel (organ)|small vessel
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9149,9155|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9149,9155|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9156,9163|false|false|false|C0012634|Disease|disease
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|9170,9173|false|false|false|C0430462|Transthoracic echocardiography|TTE
Finding|Intellectual Product|SIMPLE_SEGMENT|9174,9184|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|9174,9184|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Finding|SIMPLE_SEGMENT|9200,9206|true|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Finding|Functional Concept|SIMPLE_SEGMENT|9200,9206|true|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Finding|Intellectual Product|SIMPLE_SEGMENT|9200,9206|true|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Finding|Pathologic Function|SIMPLE_SEGMENT|9210,9225|true|false|false|C0040038|Thromboembolism|thromboembolism
Finding|Finding|SIMPLE_SEGMENT|9250,9256|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|SIMPLE_SEGMENT|9250,9256|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Pathologic Function|SIMPLE_SEGMENT|9272,9280|false|false|false|C0087086;C0302148|Blood Clot;Thrombus|thrombus
Finding|Finding|SIMPLE_SEGMENT|9272,9290|false|false|false|C4717432|Thrombus formation|thrombus formation
Finding|Functional Concept|SIMPLE_SEGMENT|9281,9290|false|false|false|C1522492|Formation|formation
Phenomenon|Biologic Function|SIMPLE_SEGMENT|9281,9290|false|false|false|C0220781|Anabolism|formation
Finding|Functional Concept|SIMPLE_SEGMENT|9304,9308|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9309,9320|false|false|false|C0018827|Heart Ventricle|ventricular
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|9321,9329|false|false|false|C0039155|Systole|systolic
Finding|Finding|SIMPLE_SEGMENT|9330,9338|false|true|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|SIMPLE_SEGMENT|9330,9338|false|true|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|SIMPLE_SEGMENT|9330,9338|false|true|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|SIMPLE_SEGMENT|9330,9338|false|true|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Mental Process|SIMPLE_SEGMENT|9346,9353|false|false|false|C0542559|contextual factors|setting
Finding|Conceptual Entity|SIMPLE_SEGMENT|9371,9382|false|false|false|C2827666|Variability|variability
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9390,9400|false|false|false|C0003811|Cardiac Arrhythmia|arrhythmia
Finding|Intellectual Product|SIMPLE_SEGMENT|9402,9406|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Finding|Finding|SIMPLE_SEGMENT|9410,9418|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|SIMPLE_SEGMENT|9410,9418|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9431,9454|false|false|false|C0040961|Tricuspid Valve Insufficiency|tricuspid regurgitation
Finding|Finding|SIMPLE_SEGMENT|9441,9454|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|SIMPLE_SEGMENT|9441,9454|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|SIMPLE_SEGMENT|9441,9454|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9463,9472|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9463,9472|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|9463,9472|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Finding|SIMPLE_SEGMENT|9473,9481|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|SIMPLE_SEGMENT|9473,9481|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|9473,9481|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|9473,9481|false|false|false|C0033095||pressure
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9495,9506|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9495,9506|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9495,9515|false|false|false|C0031039|Pericardial effusion|pericardial effusion
Finding|Body Substance|SIMPLE_SEGMENT|9495,9515|false|false|false|C1253937|Pericardial effusion body substance|pericardial effusion
Finding|Body Substance|SIMPLE_SEGMENT|9507,9515|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|SIMPLE_SEGMENT|9507,9515|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|9507,9515|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|SIMPLE_SEGMENT|9518,9523|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|Brief
Finding|Idea or Concept|SIMPLE_SEGMENT|9524,9532|false|false|false|C1547192|Organization unit type - Hospital|Hospital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9524,9539|false|false|false|C0488549||Hospital Course
Finding|Finding|SIMPLE_SEGMENT|9524,9539|false|false|false|C0489547|Hospital course|Hospital Course
Finding|Idea or Concept|SIMPLE_SEGMENT|9558,9562|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|SIMPLE_SEGMENT|9558,9562|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9579,9583|false|false|false|C0004238|Atrial Fibrillation|AFib
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|9579,9583|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|AFib
Drug|Organic Chemical|SIMPLE_SEGMENT|9587,9594|false|false|false|C3530466|Eliquis|Eliquis
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9587,9594|false|false|false|C3530466|Eliquis|Eliquis
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|9596,9599|false|false|false|C0262212|Choroidal fissure|CHF
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9596,9599|false|false|false|C0018802|Congestive heart failure|CHF
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9607,9610|false|false|false|C0020538|Hypertensive disease|HTN
Finding|Intellectual Product|SIMPLE_SEGMENT|9628,9640|false|false|false|C1272517|Sudden onset (contextual qualifier) (qualifier value)|sudden onset
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|9641,9651|false|false|false|C0013362|Dysarthria|dysarthria
Finding|Finding|SIMPLE_SEGMENT|9653,9661|false|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Finding|Idea or Concept|SIMPLE_SEGMENT|9653,9661|false|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9662,9665|false|false|false|C0446516;C1140618;C1269078|Upper Extremity;Upper arm|arm
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|9662,9665|false|false|false|C3495676|Anorectal Malformations|arm
Finding|Gene or Genome|SIMPLE_SEGMENT|9662,9665|false|false|false|C1824218;C3715044|AKR1A1 wt Allele;ARMC9 gene|arm
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|9662,9665|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Research Activity|SIMPLE_SEGMENT|9662,9665|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9662,9665|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Finding|Organism Function|SIMPLE_SEGMENT|9667,9676|false|false|false|C0026649|Movement|movements
Finding|Intellectual Product|SIMPLE_SEGMENT|9682,9686|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|poor
Finding|Finding|SIMPLE_SEGMENT|9682,9694|false|false|false|C0234964|Poor balance (finding)|poor balance
Drug|Organic Chemical|SIMPLE_SEGMENT|9687,9694|false|false|false|C4319618|Balance (substance)|balance
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9687,9694|false|false|false|C4319618|Balance (substance)|balance
Finding|Finding|SIMPLE_SEGMENT|9687,9694|false|false|false|C0014653;C0560184|Ability to balance;Equilibrium|balance
Finding|Organism Function|SIMPLE_SEGMENT|9687,9694|false|false|false|C0014653;C0560184|Ability to balance;Equilibrium|balance
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|9687,9694|false|false|false|C2174421|examination of balance|balance
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9706,9714|false|false|false|C0168634|BaseLine dental cement|baseline
Finding|Idea or Concept|SIMPLE_SEGMENT|9706,9714|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Finding|Intellectual Product|SIMPLE_SEGMENT|9717,9722|false|false|false|C1697238|NIH stroke scale|NIHSS
Finding|Organism Function|SIMPLE_SEGMENT|9738,9744|false|false|false|C0037817|Speech|speech
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|9738,9744|false|false|false|C0846595|Speech assessment|speech
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9762,9765|false|false|false|C3813556|Cancer/Testis Antigen|CTA
Finding|Gene or Genome|SIMPLE_SEGMENT|9762,9765|false|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|9762,9765|false|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9766,9770|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9766,9770|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9766,9770|false|false|false|C0362076|Problems with head|head
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9766,9770|false|false|false|C0876917|Procedure on head|head
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9766,9779|false|false|false|C0460004|Head and neck structure|head and neck
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9775,9779|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|SIMPLE_SEGMENT|9775,9779|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|SIMPLE_SEGMENT|9775,9779|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Finding|Idea or Concept|SIMPLE_SEGMENT|9810,9817|false|false|false|C2699424|Concern|concern
Finding|Functional Concept|SIMPLE_SEGMENT|9822,9826|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Drug|Chemical Viewed Structurally|SIMPLE_SEGMENT|9830,9836|false|false|false|C1881507|Macromolecular Branch|branch
Event|Activity|SIMPLE_SEGMENT|9837,9848|false|false|false|C0599946|Attenuation|attenuation
Finding|Pathologic Function|SIMPLE_SEGMENT|9865,9873|false|false|false|C1261287|Stenosis|stenosis
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|9877,9886|false|false|false|C0001168|Complete obstruction|occlusion
Finding|Finding|SIMPLE_SEGMENT|9877,9886|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Functional Concept|SIMPLE_SEGMENT|9877,9886|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|9877,9886|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Pathologic Function|SIMPLE_SEGMENT|9877,9886|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Finding|SIMPLE_SEGMENT|9930,9943|false|false|false|C0518609|Consideration|consideration
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9947,9959|false|false|false|C0162578|Thrombectomy|thrombectomy
Finding|Intellectual Product|SIMPLE_SEGMENT|9964,9969|false|false|false|C1697238|NIH stroke scale|NIHSS
Event|Activity|SIMPLE_SEGMENT|9975,9982|false|false|false|C1706079||arrival
Finding|Functional Concept|SIMPLE_SEGMENT|9975,9982|false|false|false|C1555577|arrival - ActRelationshipType|arrival
Finding|Conceptual Entity|SIMPLE_SEGMENT|10008,10017|false|false|false|C4527371|Candidate|candidate
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10054,10060|false|false|false|C0038454|Cerebrovascular accident|stroke
Finding|Finding|SIMPLE_SEGMENT|10054,10060|false|false|false|C5977286|Stroke (heart beat)|stroke
Event|Occupational Activity|SIMPLE_SEGMENT|10061,10068|false|false|false|C0557854|Services|service
Finding|Idea or Concept|SIMPLE_SEGMENT|10061,10068|false|false|false|C3245478|ActInformationPrivacyReason - service|service
Finding|Idea or Concept|SIMPLE_SEGMENT|10081,10091|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|SIMPLE_SEGMENT|10081,10091|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Finding|Finding|SIMPLE_SEGMENT|10095,10103|false|false|false|C0332149|Possible|possible
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10104,10107|false|true|false|C0007787;C0917805|Transient Cerebral Ischemia;Transient Ischemic Attack|TIA
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10111,10117|false|false|false|C0038454|Cerebrovascular accident|stroke
Finding|Finding|SIMPLE_SEGMENT|10111,10117|false|false|false|C5977286|Stroke (heart beat)|stroke
Finding|Functional Concept|SIMPLE_SEGMENT|10131,10139|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|10131,10139|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Procedure|Health Care Activity|SIMPLE_SEGMENT|10153,10162|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Gene or Genome|SIMPLE_SEGMENT|10164,10167|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10164,10167|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|SIMPLE_SEGMENT|10164,10167|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10164,10172|false|false|false|C0412674|MRI of head|MRI head
Anatomy|Body Location or Region|SIMPLE_SEGMENT|10168,10172|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10168,10172|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10168,10172|false|false|false|C0362076|Problems with head|head
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10168,10172|false|false|false|C0876917|Procedure on head|head
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|10178,10186|false|false|false|C0009924|Contrast Media|contrast
Finding|Idea or Concept|SIMPLE_SEGMENT|10200,10208|false|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|10200,10211|false|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10212,10218|true|false|false|C0038454|Cerebrovascular accident|stroke
Finding|Finding|SIMPLE_SEGMENT|10212,10218|true|false|false|C5977286|Stroke (heart beat)|stroke
Finding|Intellectual Product|SIMPLE_SEGMENT|10220,10227|false|false|false|C0684224|Report (document)|Reports
Procedure|Health Care Activity|SIMPLE_SEGMENT|10220,10227|false|false|false|C0700287|Reporting|Reports
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10236,10250|false|false|false|C0013516|Echocardiography|echocardiogram
Finding|Classification|SIMPLE_SEGMENT|10255,10265|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|10255,10265|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10266,10269|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|10266,10269|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|10266,10269|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10266,10269|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|SIMPLE_SEGMENT|10266,10269|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|10266,10269|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|SIMPLE_SEGMENT|10266,10269|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10266,10269|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Finding|Gene or Genome|SIMPLE_SEGMENT|10266,10269|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|SIMPLE_SEGMENT|10266,10269|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Intellectual Product|SIMPLE_SEGMENT|10300,10305|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10306,10314|false|false|false|C2926606||findings
Finding|Functional Concept|SIMPLE_SEGMENT|10306,10314|false|false|false|C2607943|findings aspects|findings
Finding|Idea or Concept|SIMPLE_SEGMENT|10360,10367|false|false|false|C2699424|Concern|concern
Finding|Finding|SIMPLE_SEGMENT|10384,10390|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Finding|Intellectual Product|SIMPLE_SEGMENT|10384,10390|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Finding|Mental Process|SIMPLE_SEGMENT|10384,10390|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Finding|Finding|SIMPLE_SEGMENT|10396,10400|false|false|false|C1299581|Able (qualifier value)|able
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|10412,10416|false|false|false|C0001288|Activity of daily living (function)|ADLs
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|10421,10426|false|false|false|C1998602|Meal (occasion for eating)|meals
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10448,10451|false|false|false|C1431931|ALF protein, human|ALF
Drug|Biologically Active Substance|SIMPLE_SEGMENT|10448,10451|false|false|false|C1431931|ALF protein, human|ALF
Finding|Gene or Genome|SIMPLE_SEGMENT|10448,10451|false|false|false|C1332077;C1704942|GTF2A1L gene;GTF2A1L wt Allele|ALF
Finding|Gene or Genome|SIMPLE_SEGMENT|10469,10472|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Finding|Intellectual Product|SIMPLE_SEGMENT|10505,10510|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Functional Concept|SIMPLE_SEGMENT|10511,10517|true|false|false|C0392747|Changing|change
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10511,10517|true|false|false|C4319952|Change - procedure|change
Finding|Intellectual Product|SIMPLE_SEGMENT|10550,10554|false|false|false|C1720092|Once - dosing instruction fragment|once
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|10587,10590|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10587,10590|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|10587,10590|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|SIMPLE_SEGMENT|10587,10590|false|false|false|C1332410|BID gene|BID
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10591,10601|false|false|false|C0013227|Pharmaceutical Preparations|medication
Finding|Intellectual Product|SIMPLE_SEGMENT|10591,10601|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|10644,10647|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10644,10647|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|10644,10647|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|SIMPLE_SEGMENT|10644,10647|false|false|false|C1332410|BID gene|BID
Finding|Conceptual Entity|SIMPLE_SEGMENT|10663,10672|false|false|false|C4527371|Candidate|candidate
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|10682,10685|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10682,10685|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|10682,10685|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|SIMPLE_SEGMENT|10682,10685|false|false|false|C1332410|BID gene|BID
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10697,10700|false|false|false|C1114365||age
Drug|Biologically Active Substance|SIMPLE_SEGMENT|10697,10700|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|SIMPLE_SEGMENT|10697,10700|false|false|false|C0162574|Glycation End Products, Advanced|age
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10705,10711|false|false|false|C0944911||weight
Finding|Finding|SIMPLE_SEGMENT|10705,10711|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|SIMPLE_SEGMENT|10705,10711|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|SIMPLE_SEGMENT|10705,10711|false|false|false|C1305866|Weighing patient|weight
Drug|Organic Chemical|SIMPLE_SEGMENT|10733,10745|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10733,10745|false|false|false|C0286651|atorvastatin|atorvastatin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10755,10769|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|hyperlipidemia
Finding|Finding|SIMPLE_SEGMENT|10755,10769|false|false|false|C0428465|Serum lipids high (finding)|hyperlipidemia
Drug|Biologically Active Substance|SIMPLE_SEGMENT|10771,10774|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Drug|Organic Chemical|SIMPLE_SEGMENT|10771,10774|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10771,10774|false|false|false|C0202117|Low density lipoprotein cholesterol measurement|LDL
Anatomy|Body System|SIMPLE_SEGMENT|10784,10794|false|false|false|C0007226|Cardiovascular system|cardiology
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|10823,10828|false|false|false|C0030471;C1305231|Nasal sinus;Sinus - general anatomical term|sinus
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|10823,10828|false|false|false|C0016169|pathologic fistula|sinus
Drug|Organic Chemical|SIMPLE_SEGMENT|10823,10828|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10823,10828|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10829,10835|false|false|false|C0488347||pauses
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10845,10854|false|false|false|C0039451|Telemetry|telemetry
Finding|Idea or Concept|SIMPLE_SEGMENT|10887,10891|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|10887,10891|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|10887,10891|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|10892,10900|false|false|false|C0004147|atenolol|atenolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10892,10900|false|false|false|C0004147|atenolol|atenolol
Finding|Idea or Concept|SIMPLE_SEGMENT|10929,10933|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|10929,10933|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|10929,10933|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|10935,10942|false|false|false|C0012265|digoxin|digoxin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10935,10942|false|false|false|C0012265|digoxin|digoxin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10935,10942|false|false|false|C0337449|Digoxin measurement|digoxin
Finding|Finding|SIMPLE_SEGMENT|10947,10952|false|false|false|C0587267;C3810854|Close;Closed|close
Finding|Functional Concept|SIMPLE_SEGMENT|10947,10952|false|false|false|C0587267;C3810854|Close;Closed|close
Anatomy|Body System|SIMPLE_SEGMENT|10953,10963|false|false|false|C0007226|Cardiovascular system|cardiology
Finding|Idea or Concept|SIMPLE_SEGMENT|10983,10987|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|10983,10987|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|10983,10987|false|false|false|C1553498|home health encounter|home
Finding|Finding|SIMPLE_SEGMENT|11006,11011|false|false|false|C0587267;C3810854|Close;Closed|close
Finding|Functional Concept|SIMPLE_SEGMENT|11006,11011|false|false|false|C0587267;C3810854|Close;Closed|close
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11012,11015|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|11012,11015|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|11012,11015|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|11012,11015|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|SIMPLE_SEGMENT|11012,11015|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|11012,11015|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|SIMPLE_SEGMENT|11012,11015|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11012,11015|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Finding|Gene or Genome|SIMPLE_SEGMENT|11012,11015|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|SIMPLE_SEGMENT|11012,11015|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Finding|SIMPLE_SEGMENT|11023,11032|false|false|false|C0687129;C1550450|Encounter due to vagabond status;Living Arrangement - Transient|Transient
Finding|Organism Function|SIMPLE_SEGMENT|11041,11047|false|false|false|C0037817|Speech|speech
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|11041,11047|false|false|false|C0846595|Speech assessment|speech
Finding|Finding|SIMPLE_SEGMENT|11052,11063|false|false|false|C1444783|Instability|instability
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11069,11072|false|false|false|C0007787;C0917805|Transient Cerebral Ischemia;Transient Ischemic Attack|TIA
Procedure|Health Care Activity|SIMPLE_SEGMENT|11079,11086|false|false|false|C0009818|Consultation|consult
Finding|Idea or Concept|SIMPLE_SEGMENT|11101,11105|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|11101,11105|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|11101,11105|false|false|false|C1553498|home health encounter|home
Finding|Idea or Concept|SIMPLE_SEGMENT|11111,11115|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|11111,11115|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|11111,11115|false|false|false|C1553498|home health encounter|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|11111,11124|false|false|false|C0020043|Home visit (procedure)|home services
Event|Occupational Activity|SIMPLE_SEGMENT|11116,11124|false|false|false|C0557854|Services|services
Procedure|Health Care Activity|SIMPLE_SEGMENT|11116,11124|false|false|false|C1704289|Clinical Service|services
Drug|Organic Chemical|SIMPLE_SEGMENT|11138,11150|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11138,11150|false|false|false|C0286651|atorvastatin|atorvastatin
Finding|Idea or Concept|SIMPLE_SEGMENT|11173,11177|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|11173,11177|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|11173,11177|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|11178,11186|false|false|false|C1831808|apixaban|apixaban
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11178,11186|false|false|false|C1831808|apixaban|apixaban
Drug|Organic Chemical|SIMPLE_SEGMENT|11191,11202|false|false|false|C0723712|Therapeutic brand of coal tar|therapeutic
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11191,11202|false|false|false|C0723712|Therapeutic brand of coal tar|therapeutic
Finding|Functional Concept|SIMPLE_SEGMENT|11191,11202|false|false|false|C0302350;C1547427|Therapeutic;Therapeutic - Location Service Code|therapeutic
Finding|Intellectual Product|SIMPLE_SEGMENT|11191,11202|false|false|false|C0302350;C1547427|Therapeutic;Therapeutic - Location Service Code|therapeutic
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11191,11202|false|false|false|C0087111|Therapeutic procedure|therapeutic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11220,11226|false|false|false|C0038454|Cerebrovascular accident|stroke
Finding|Finding|SIMPLE_SEGMENT|11220,11226|false|false|false|C5977286|Stroke (heart beat)|stroke
Finding|Body Substance|SIMPLE_SEGMENT|11243,11252|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|11243,11252|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|11243,11252|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|11243,11252|false|false|false|C0030685|Patient Discharge|discharge
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11258,11264|false|false|false|C0038454|Cerebrovascular accident|stroke
Finding|Finding|SIMPLE_SEGMENT|11258,11264|false|false|false|C5977286|Stroke (heart beat)|stroke
Finding|Intellectual Product|SIMPLE_SEGMENT|11258,11269|false|false|false|C1277291|Stroke risk|stroke risk
Finding|Idea or Concept|SIMPLE_SEGMENT|11265,11269|false|false|false|C0035647|Risk|risk
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11265,11277|false|false|false|C1830376||risk factors
Finding|Finding|SIMPLE_SEGMENT|11265,11277|false|false|false|C0035648;C0455624;C1553898|History of - risk factor;risk factors;risk factors - observation list|risk factors
Finding|Intellectual Product|SIMPLE_SEGMENT|11265,11277|false|false|false|C0035648;C0455624;C1553898|History of - risk factor;risk factors;risk factors - observation list|risk factors
Finding|Classification|SIMPLE_SEGMENT|11308,11311|false|false|false|C4521595|United States Military enlisted E3 (qualifier value)|A1c
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|11308,11311|false|false|false|C0474680|Hemoglobin A1c measurement|A1c
Finding|Finding|SIMPLE_SEGMENT|11320,11326|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Finding|Idea or Concept|SIMPLE_SEGMENT|11320,11326|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Finding|Intellectual Product|SIMPLE_SEGMENT|11327,11334|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|11327,11334|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Finding|Functional Concept|SIMPLE_SEGMENT|11345,11349|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11345,11366|false|false|false|C0226231|Structure of left vertebral artery|left vertebral artery
Finding|Pathologic Function|SIMPLE_SEGMENT|11345,11376|false|false|false|C4536452|Occlusion of left vertebral artery (disorder)|left vertebral artery occlusion
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11350,11359|false|false|false|C0549207|Bone structure of spine|vertebral
Anatomy|Body Location or Region|SIMPLE_SEGMENT|11350,11366|false|false|false|C0042559;C4695118|Head+Neck>Vertebral artery;Structure of vertebral artery|vertebral artery
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11350,11366|false|false|false|C0042559;C4695118|Head+Neck>Vertebral artery;Structure of vertebral artery|vertebral artery
Finding|Pathologic Function|SIMPLE_SEGMENT|11350,11376|false|false|false|C0265104|Vertebral artery obstruction (disorder)|vertebral artery occlusion
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11360,11366|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|SIMPLE_SEGMENT|11360,11366|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Finding|Pathologic Function|SIMPLE_SEGMENT|11360,11376|false|false|false|C0264995|Occlusion of artery (disorder)|artery occlusion
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|11367,11376|false|false|false|C0001168|Complete obstruction|occlusion
Finding|Finding|SIMPLE_SEGMENT|11367,11376|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Functional Concept|SIMPLE_SEGMENT|11367,11376|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|11367,11376|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Pathologic Function|SIMPLE_SEGMENT|11367,11376|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Finding|SIMPLE_SEGMENT|11382,11390|false|false|false|C2984079|Somewhat|somewhat
Event|Activity|SIMPLE_SEGMENT|11405,11415|false|false|false|C0599946|Attenuation|attenuated
Finding|Functional Concept|SIMPLE_SEGMENT|11416,11420|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Finding|Social Behavior|SIMPLE_SEGMENT|11424,11432|false|false|false|C0678975|inferiority|inferior
Drug|Chemical Viewed Structurally|SIMPLE_SEGMENT|11433,11439|false|false|false|C1881507|Macromolecular Branch|branch
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11443,11457|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|Hyperlipidemia
Finding|Finding|SIMPLE_SEGMENT|11443,11457|false|false|false|C0428465|Serum lipids high (finding)|Hyperlipidemia
Drug|Biologically Active Substance|SIMPLE_SEGMENT|11459,11462|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Drug|Organic Chemical|SIMPLE_SEGMENT|11459,11462|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|11459,11462|false|false|false|C0202117|Low density lipoprotein cholesterol measurement|LDL
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11470,11477|false|false|false|C0028754|Obesity|Obesity
Finding|Finding|SIMPLE_SEGMENT|11470,11477|false|false|false|C4759928|BODY MASS INDEX QUANTITATIVE TRAIT LOCUS 20|Obesity
Finding|Idea or Concept|SIMPLE_SEGMENT|11484,11491|true|false|false|C2699424|Concern|concern
Drug|Organic Chemical|SIMPLE_SEGMENT|11502,11507|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11502,11507|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Finding|Organism Function|SIMPLE_SEGMENT|11502,11507|false|false|false|C0037313|Sleep|sleep
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11502,11513|false|false|false|C0037315|Sleep Apnea Syndromes|sleep apnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|11508,11513|false|false|false|C0003578|Apnea|apnea
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11540,11549|false|false|false|C0945731||diagnosis
Finding|Classification|SIMPLE_SEGMENT|11540,11549|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|11540,11549|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|11540,11549|false|false|false|C0011900|Diagnosis|diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|11553,11567|false|false|false|C0013516|Echocardiography|echocardiogram
Finding|Intellectual Product|SIMPLE_SEGMENT|11597,11602|false|false|false|C1705923|Study Object|study
Procedure|Research Activity|SIMPLE_SEGMENT|11597,11602|false|false|false|C0008972;C0947630;C2603343|Clinical Research;Scientific Study;Study|study
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11605,11608|false|false|false|C0002880;C0272325|Autoimmune hemolytic anemia;Factor 8 deficiency, acquired|AHA
Drug|Organic Chemical|SIMPLE_SEGMENT|11605,11608|false|false|false|C0050451|acetohydroxamic acid|AHA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11605,11608|false|false|false|C0050451|acetohydroxamic acid|AHA
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|11609,11612|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Enzyme|SIMPLE_SEGMENT|11609,11612|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Organic Chemical|SIMPLE_SEGMENT|11609,11612|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11609,11612|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Finding|Gene or Genome|SIMPLE_SEGMENT|11609,11612|false|false|false|C1412553|ARSA gene|ASA
Anatomy|Cell Component|SIMPLE_SEGMENT|11613,11617|false|false|false|C1167518|viral nucleocapsid location|Core
Finding|Body Substance|SIMPLE_SEGMENT|11613,11617|false|false|false|C3274653|Core Specimen|Core
Finding|Functional Concept|SIMPLE_SEGMENT|11618,11626|false|false|false|C1879489|Measures (attribute)|Measures
Finding|Functional Concept|SIMPLE_SEGMENT|11631,11639|false|false|false|C0475224|Ischemic|Ischemic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11631,11646|false|false|false|C0948008|Ischemic stroke|Ischemic Stroke
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11640,11646|false|false|false|C0038454|Cerebrovascular accident|Stroke
Finding|Finding|SIMPLE_SEGMENT|11640,11646|false|false|false|C5977286|Stroke (heart beat)|Stroke
Finding|Finding|SIMPLE_SEGMENT|11651,11660|false|false|false|C0687129;C1550450|Encounter due to vagabond status;Living Arrangement - Transient|Transient
Finding|Functional Concept|SIMPLE_SEGMENT|11661,11669|false|true|false|C0475224|Ischemic|Ischemic
Finding|Finding|SIMPLE_SEGMENT|11671,11677|false|false|false|C1261512;C1304680|Attack (finding);Attack behavior|Attack
Finding|Social Behavior|SIMPLE_SEGMENT|11671,11677|false|false|false|C1261512;C1304680|Attack (finding);Attack behavior|Attack
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11681,11690|false|false|false|C0011168|Deglutition Disorders|Dysphagia
Procedure|Health Care Activity|SIMPLE_SEGMENT|11681,11700|false|false|false|C0500456|Screening for dysphagia|Dysphagia screening
Finding|Finding|SIMPLE_SEGMENT|11691,11700|false|false|false|C0220909;C1305399;C1409616|Aspects of disease screening;Screening - procedure intent;Special screening finding|screening
Finding|Functional Concept|SIMPLE_SEGMENT|11691,11700|false|false|false|C0220909;C1305399;C1409616|Aspects of disease screening;Screening - procedure intent;Special screening finding|screening
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|11691,11700|false|false|false|C0199230;C0220908;C1698960;C1710031;C1710032|Disease Screening;Screening;Screening for cancer;Screening procedure;research subject screening|screening
Procedure|Health Care Activity|SIMPLE_SEGMENT|11691,11700|false|false|false|C0199230;C0220908;C1698960;C1710031;C1710032|Disease Screening;Screening;Screening for cancer;Screening procedure;research subject screening|screening
Procedure|Research Activity|SIMPLE_SEGMENT|11691,11700|false|false|false|C0199230;C0220908;C1698960;C1710031;C1710032|Disease Screening;Screening;Screening for cancer;Screening procedure;research subject screening|screening
Finding|Functional Concept|SIMPLE_SEGMENT|11715,11721|false|false|false|C1512806|Intake|intake
Procedure|Health Care Activity|SIMPLE_SEGMENT|11715,11721|false|false|false|C3251814;C4521161|Intake (treatment);Measurement of fluid intake|intake
Finding|Finding|SIMPLE_SEGMENT|11727,11730|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Gene or Genome|SIMPLE_SEGMENT|11727,11730|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Idea or Concept|SIMPLE_SEGMENT|11727,11730|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Intellectual Product|SIMPLE_SEGMENT|11727,11730|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Anatomy|Body Location or Region|SIMPLE_SEGMENT|11776,11779|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11776,11779|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11776,11779|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11776,11791|false|false|false|C0853245|DVT prophylaxis|DVT Prophylaxis
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11780,11791|false|false|false|C0199176|Prophylactic treatment|Prophylaxis
Finding|Finding|SIMPLE_SEGMENT|11810,11813|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Gene or Genome|SIMPLE_SEGMENT|11810,11813|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Idea or Concept|SIMPLE_SEGMENT|11810,11813|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Intellectual Product|SIMPLE_SEGMENT|11810,11813|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Finding|SIMPLE_SEGMENT|11840,11847|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|SIMPLE_SEGMENT|11840,11847|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11840,11847|false|false|false|C0087111|Therapeutic procedure|therapy
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|11864,11867|false|false|false|C0082420|Endoglin, human|end
Drug|Immunologic Factor|SIMPLE_SEGMENT|11864,11867|false|false|false|C0082420|Endoglin, human|end
Finding|Functional Concept|SIMPLE_SEGMENT|11864,11867|false|false|false|C1366583;C1561490;C1704837|ENG gene;ENG wt Allele;end - ActRelationshipCheckpoint|end
Finding|Gene or Genome|SIMPLE_SEGMENT|11864,11867|false|false|false|C1366583;C1561490;C1704837|ENG gene;ENG wt Allele;end - ActRelationshipCheckpoint|end
Finding|Idea or Concept|SIMPLE_SEGMENT|11871,11879|false|false|false|C1547192|Organization unit type - Hospital|hospital
Finding|Idea or Concept|SIMPLE_SEGMENT|11880,11883|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|11880,11883|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Finding|SIMPLE_SEGMENT|11880,11885|false|false|false|C3842676|Day 2|day 2
Finding|Finding|SIMPLE_SEGMENT|11892,11895|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Gene or Genome|SIMPLE_SEGMENT|11892,11895|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Idea or Concept|SIMPLE_SEGMENT|11892,11895|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Intellectual Product|SIMPLE_SEGMENT|11892,11895|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Drug|Biologically Active Substance|SIMPLE_SEGMENT|11907,11910|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Drug|Organic Chemical|SIMPLE_SEGMENT|11907,11910|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|11907,11910|false|false|false|C0202117|Low density lipoprotein cholesterol measurement|LDL
Finding|Finding|SIMPLE_SEGMENT|11927,11930|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Gene or Genome|SIMPLE_SEGMENT|11927,11930|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Idea or Concept|SIMPLE_SEGMENT|11927,11930|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Intellectual Product|SIMPLE_SEGMENT|11927,11930|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Drug|Biologically Active Substance|SIMPLE_SEGMENT|11932,11935|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Drug|Organic Chemical|SIMPLE_SEGMENT|11932,11935|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|11932,11935|false|false|false|C0202117|Low density lipoprotein cholesterol measurement|LDL
Drug|Organic Chemical|SIMPLE_SEGMENT|11964,11970|false|false|false|C0360714|Hydroxymethylglutaryl-CoA Reductase Inhibitors|statin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11964,11970|false|false|false|C0360714|Hydroxymethylglutaryl-CoA Reductase Inhibitors|statin
Finding|Gene or Genome|SIMPLE_SEGMENT|11964,11970|false|false|false|C1414273|EEF1A2 gene|statin
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11964,11978|false|false|false|C1278454|Administration of prophylactic statin|statin therapy
Finding|Finding|SIMPLE_SEGMENT|11971,11978|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|SIMPLE_SEGMENT|11971,11978|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11971,11978|false|false|false|C0087111|Therapeutic procedure|therapy
Drug|Organic Chemical|SIMPLE_SEGMENT|11994,12005|false|false|false|C0074554|simvastatin|simvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11994,12005|false|false|false|C0074554|simvastatin|simvastatin
Drug|Organic Chemical|SIMPLE_SEGMENT|12013,12024|false|false|false|C0074554|simvastatin|simvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12013,12024|false|false|false|C0074554|simvastatin|simvastatin
Drug|Organic Chemical|SIMPLE_SEGMENT|12046,12058|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12046,12058|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Organic Chemical|SIMPLE_SEGMENT|12075,12087|false|false|false|C0965129|rosuvastatin|rosuvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12075,12087|false|false|false|C0965129|rosuvastatin|rosuvastatin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|12106,12109|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Drug|Organic Chemical|SIMPLE_SEGMENT|12106,12109|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|12106,12109|false|false|false|C0202117|Low density lipoprotein cholesterol measurement|LDL
Finding|Finding|SIMPLE_SEGMENT|12121,12124|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Gene or Genome|SIMPLE_SEGMENT|12121,12124|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Idea or Concept|SIMPLE_SEGMENT|12121,12124|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Intellectual Product|SIMPLE_SEGMENT|12121,12124|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Drug|Biologically Active Substance|SIMPLE_SEGMENT|12138,12141|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Drug|Organic Chemical|SIMPLE_SEGMENT|12138,12141|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|12138,12141|false|false|false|C0202117|Low density lipoprotein cholesterol measurement|LDL
Drug|Biologically Active Substance|SIMPLE_SEGMENT|12145,12148|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Drug|Organic Chemical|SIMPLE_SEGMENT|12145,12148|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|12145,12148|false|false|false|C0202117|Low density lipoprotein cholesterol measurement|LDL
Finding|Idea or Concept|SIMPLE_SEGMENT|12154,12160|false|false|false|C0392360|Indication of (contextual qualifier)|reason
Drug|Organic Chemical|SIMPLE_SEGMENT|12176,12182|false|false|false|C0360714|Hydroxymethylglutaryl-CoA Reductase Inhibitors|Statin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12176,12182|false|false|false|C0360714|Hydroxymethylglutaryl-CoA Reductase Inhibitors|Statin
Finding|Gene or Genome|SIMPLE_SEGMENT|12176,12182|false|false|false|C1414273|EEF1A2 gene|Statin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12183,12193|false|false|false|C0013227|Pharmaceutical Preparations|medication
Finding|Intellectual Product|SIMPLE_SEGMENT|12183,12193|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Finding|Pathologic Function|SIMPLE_SEGMENT|12183,12201|false|false|false|C0013182|Drug Allergy|medication allergy
Finding|Finding|SIMPLE_SEGMENT|12194,12201|false|false|false|C0020517;C0489531;C1314973;C1527304;C1547542;C3539909|Allergic Reaction;Allergic disposition;Allergy - Charge Type Reason;History of allergies;Hypersensitivity;Response to antigens|allergy
Finding|Idea or Concept|SIMPLE_SEGMENT|12194,12201|false|false|false|C0020517;C0489531;C1314973;C1527304;C1547542;C3539909|Allergic Reaction;Allergic disposition;Allergy - Charge Type Reason;History of allergies;Hypersensitivity;Response to antigens|allergy
Finding|Pathologic Function|SIMPLE_SEGMENT|12194,12201|false|false|false|C0020517;C0489531;C1314973;C1527304;C1547542;C3539909|Allergic Reaction;Allergic disposition;Allergy - Charge Type Reason;History of allergies;Hypersensitivity;Response to antigens|allergy
Finding|Physiologic Function|SIMPLE_SEGMENT|12194,12201|false|false|false|C0020517;C0489531;C1314973;C1527304;C1547542;C3539909|Allergic Reaction;Allergic disposition;Allergy - Charge Type Reason;History of allergies;Hypersensitivity;Response to antigens|allergy
Finding|Idea or Concept|SIMPLE_SEGMENT|12212,12219|false|false|false|C0392360|Indication of (contextual qualifier)|reasons
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12234,12243|false|false|false|C0804815||physician
Finding|Intellectual Product|SIMPLE_SEGMENT|12253,12261|false|false|false|C0237607;C3245512|Experience (Practice);HL7PublishingSubSection - practice|practice
Finding|Mental Process|SIMPLE_SEGMENT|12253,12261|false|false|false|C0237607;C3245512|Experience (Practice);HL7PublishingSubSection - practice|practice
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12269,12278|false|false|false|C0804815||physician
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12284,12293|false|false|false|C0804815||physician
Finding|Gene or Genome|SIMPLE_SEGMENT|12294,12297|false|false|false|C2986617|ANPEP wt Allele|APN
Finding|Idea or Concept|SIMPLE_SEGMENT|12305,12315|false|false|false|C1546966|Primary Observer's Qualification - Pharmacist|pharmacist
Drug|Biologically Active Substance|SIMPLE_SEGMENT|12320,12323|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Drug|Organic Chemical|SIMPLE_SEGMENT|12320,12323|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|12320,12323|false|false|false|C0202117|Low density lipoprotein cholesterol measurement|LDL
Finding|Individual Behavior|SIMPLE_SEGMENT|12349,12356|false|false|false|C0037369;C0453996;C1548578|Location characteristic ID - Smoking;Smoking;Tobacco smoking behavior|Smoking
Finding|Intellectual Product|SIMPLE_SEGMENT|12349,12356|false|false|false|C0037369;C0453996;C1548578|Location characteristic ID - Smoking;Smoking;Tobacco smoking behavior|Smoking
Finding|Individual Behavior|SIMPLE_SEGMENT|12349,12366|false|false|false|C0085134|Cessation of smoking|Smoking cessation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|12349,12366|false|false|false|C1095963|Smoking cessation therapy|Smoking cessation
Event|Activity|SIMPLE_SEGMENT|12357,12366|false|false|false|C1880019|Cessation|cessation
Finding|Finding|SIMPLE_SEGMENT|12367,12377|false|false|false|C0740209;C2148587|Encounter due to counseling;duration of counseling|counseling
Procedure|Health Care Activity|SIMPLE_SEGMENT|12367,12377|false|false|false|C0010210;C0542296|Counseling;Counselling service|counseling
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|12367,12377|false|false|false|C0010210;C0542296|Counseling;Counselling service|counseling
Finding|Finding|SIMPLE_SEGMENT|12388,12391|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Gene or Genome|SIMPLE_SEGMENT|12388,12391|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Idea or Concept|SIMPLE_SEGMENT|12388,12391|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Intellectual Product|SIMPLE_SEGMENT|12388,12391|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Idea or Concept|SIMPLE_SEGMENT|12402,12408|true|false|false|C0392360|Indication of (contextual qualifier)|reason
Finding|Finding|SIMPLE_SEGMENT|12430,12436|false|false|false|C1299582|Unable|unable
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12456,12462|false|false|false|C0038454|Cerebrovascular accident|Stroke
Finding|Finding|SIMPLE_SEGMENT|12456,12462|false|false|false|C5977286|Stroke (heart beat)|Stroke
Procedure|Educational Activity|SIMPLE_SEGMENT|12456,12472|false|false|false|C4303794|Education about stroke|Stroke education
Finding|Classification|SIMPLE_SEGMENT|12463,12472|false|false|false|C0013622;C0013658;C0424927|Details of education;Educational Status;Educational aspects|education
Finding|Finding|SIMPLE_SEGMENT|12463,12472|false|false|false|C0013622;C0013658;C0424927|Details of education;Educational Status;Educational aspects|education
Procedure|Educational Activity|SIMPLE_SEGMENT|12463,12472|false|false|false|C0013621;C0039401|Education (procedure);Knowledge acquisition|education
Finding|Idea or Concept|SIMPLE_SEGMENT|12494,12498|false|false|false|C0035647|Risk|risk
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12494,12506|false|false|false|C1830376||risk factors
Finding|Finding|SIMPLE_SEGMENT|12494,12506|false|false|false|C0035648;C0455624;C1553898|History of - risk factor;risk factors;risk factors - observation list|risk factors
Finding|Intellectual Product|SIMPLE_SEGMENT|12494,12506|false|false|false|C0035648;C0455624;C1553898|History of - risk factor;risk factors;risk factors - observation list|risk factors
Event|Activity|SIMPLE_SEGMENT|12516,12524|false|false|false|C1879547|activation [action]|activate
Finding|Functional Concept|SIMPLE_SEGMENT|12516,12524|false|false|false|C1515877;C3853838|activate - Data Operation;activate biological process|activate
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|12525,12528|false|false|false|C0015063|Ethyl Methanesulfonate|EMS
Drug|Organic Chemical|SIMPLE_SEGMENT|12525,12528|false|false|false|C0015063|Ethyl Methanesulfonate|EMS
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12525,12528|false|false|false|C0015063|Ethyl Methanesulfonate|EMS
Finding|Gene or Genome|SIMPLE_SEGMENT|12525,12528|false|false|false|C5203240|EMSLR gene|EMS
Procedure|Health Care Activity|SIMPLE_SEGMENT|12525,12528|false|false|false|C0013961|Emergency Medical Services|EMS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12533,12539|false|false|false|C0038454|Cerebrovascular accident|stroke
Finding|Finding|SIMPLE_SEGMENT|12533,12539|false|false|false|C5977286|Stroke (heart beat)|stroke
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12541,12547|false|false|false|C0038454|Cerebrovascular accident|stroke
Finding|Finding|SIMPLE_SEGMENT|12541,12547|false|false|false|C5977286|Stroke (heart beat)|stroke
Finding|Conceptual Entity|SIMPLE_SEGMENT|12548,12555|false|false|false|C0871599;C1549021;C1578603;C1578605;C4553014|Cautionary Warning;System Alert;Warning - AcknowledgementDetailType;Warning - EquipmentAlertLevel;Warning - Error severity|warning
Finding|Idea or Concept|SIMPLE_SEGMENT|12548,12555|false|false|false|C0871599;C1549021;C1578603;C1578605;C4553014|Cautionary Warning;System Alert;Warning - AcknowledgementDetailType;Warning - EquipmentAlertLevel;Warning - Error severity|warning
Finding|Intellectual Product|SIMPLE_SEGMENT|12548,12555|false|false|false|C0871599;C1549021;C1578603;C1578605;C4553014|Cautionary Warning;System Alert;Warning - AcknowledgementDetailType;Warning - EquipmentAlertLevel;Warning - Error severity|warning
Event|Governmental or Regulatory Activity|SIMPLE_SEGMENT|12548,12561|false|false|false|C0871598|warning signs|warning signs
Finding|Finding|SIMPLE_SEGMENT|12556,12561|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|SIMPLE_SEGMENT|12556,12561|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Sign or Symptom|SIMPLE_SEGMENT|12556,12574|false|false|false|C0037088|Signs and Symptoms|signs and symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|12566,12574|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|12566,12574|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12588,12599|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12588,12599|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|SIMPLE_SEGMENT|12588,12599|false|false|false|C4284232|Medications|medications
Finding|Functional Concept|SIMPLE_SEGMENT|12601,12605|false|false|false|C0686904|Patient need for (contextual qualifier)|need
Finding|Functional Concept|SIMPLE_SEGMENT|12601,12609|false|false|false|C0686904|Patient need for (contextual qualifier)|need for
Procedure|Health Care Activity|SIMPLE_SEGMENT|12610,12618|false|false|false|C1522577|follow-up|followup
Finding|Finding|SIMPLE_SEGMENT|12654,12657|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Gene or Genome|SIMPLE_SEGMENT|12654,12657|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Idea or Concept|SIMPLE_SEGMENT|12654,12657|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Intellectual Product|SIMPLE_SEGMENT|12654,12657|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Event|Activity|SIMPLE_SEGMENT|12669,12679|false|false|false|C1516048|Assessed|Assessment
Finding|Intellectual Product|SIMPLE_SEGMENT|12669,12679|false|false|false|C0679207|Knowledge acquisition using a method of assessment|Assessment
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|12669,12679|false|false|false|C0028708;C0031809;C0220825;C0542573;C0549068;C0549070;C0549071;C0549072;C0549073;C0549074;C0549075;C0549076;C0549078;C0549079;C0549080;C1161151;C1261322;C2237115|Evaluation;Evaluation procedure;Nutrition Assessment;Personal care assessment;Physical Examination;assessment of cognitive functions|Assessment
Procedure|Health Care Activity|SIMPLE_SEGMENT|12669,12679|false|false|false|C0028708;C0031809;C0220825;C0542573;C0549068;C0549070;C0549071;C0549072;C0549073;C0549074;C0549075;C0549076;C0549078;C0549079;C0549080;C1161151;C1261322;C2237115|Evaluation;Evaluation procedure;Nutrition Assessment;Personal care assessment;Physical Examination;assessment of cognitive functions|Assessment
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|12669,12698|false|false|false|C0431070|Assessment for rehabilitation|Assessment for rehabilitation
Finding|Finding|SIMPLE_SEGMENT|12684,12698|false|false|false|C0007237;C0034992|Encounter due to care involving use of rehabilitation procedures;Rehabilitation aspects|rehabilitation
Finding|Functional Concept|SIMPLE_SEGMENT|12684,12698|false|false|false|C0007237;C0034992|Encounter due to care involving use of rehabilitation procedures;Rehabilitation aspects|rehabilitation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|12684,12698|false|false|false|C0034991|Rehabilitation therapy|rehabilitation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|12702,12707|false|false|false|C0034991|Rehabilitation therapy|rehab
Event|Occupational Activity|SIMPLE_SEGMENT|12708,12716|false|false|false|C0557854|Services|services
Procedure|Health Care Activity|SIMPLE_SEGMENT|12708,12716|false|false|false|C1704289|Clinical Service|services
Finding|Finding|SIMPLE_SEGMENT|12734,12737|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Gene or Genome|SIMPLE_SEGMENT|12734,12737|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Idea or Concept|SIMPLE_SEGMENT|12734,12737|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Intellectual Product|SIMPLE_SEGMENT|12734,12737|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Drug|Organic Chemical|SIMPLE_SEGMENT|12763,12769|false|false|false|C0360714|Hydroxymethylglutaryl-CoA Reductase Inhibitors|statin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12763,12769|false|false|false|C0360714|Hydroxymethylglutaryl-CoA Reductase Inhibitors|statin
Finding|Gene or Genome|SIMPLE_SEGMENT|12763,12769|false|false|false|C1414273|EEF1A2 gene|statin
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|12763,12777|false|false|false|C1278454|Administration of prophylactic statin|statin therapy
Finding|Finding|SIMPLE_SEGMENT|12770,12777|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|SIMPLE_SEGMENT|12770,12777|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|12770,12777|false|false|false|C0087111|Therapeutic procedure|therapy
Finding|Finding|SIMPLE_SEGMENT|12783,12786|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Gene or Genome|SIMPLE_SEGMENT|12783,12786|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Idea or Concept|SIMPLE_SEGMENT|12783,12786|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Intellectual Product|SIMPLE_SEGMENT|12783,12786|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Drug|Biologically Active Substance|SIMPLE_SEGMENT|12799,12802|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Drug|Organic Chemical|SIMPLE_SEGMENT|12799,12802|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|12799,12802|false|false|false|C0202117|Low density lipoprotein cholesterol measurement|LDL
Finding|Idea or Concept|SIMPLE_SEGMENT|12809,12815|false|false|false|C0392360|Indication of (contextual qualifier)|reason
Drug|Organic Chemical|SIMPLE_SEGMENT|12831,12837|false|false|false|C0360714|Hydroxymethylglutaryl-CoA Reductase Inhibitors|Statin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12831,12837|false|false|false|C0360714|Hydroxymethylglutaryl-CoA Reductase Inhibitors|Statin
Finding|Gene or Genome|SIMPLE_SEGMENT|12831,12837|false|false|false|C1414273|EEF1A2 gene|Statin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12838,12848|false|false|false|C0013227|Pharmaceutical Preparations|medication
Finding|Intellectual Product|SIMPLE_SEGMENT|12838,12848|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Finding|Pathologic Function|SIMPLE_SEGMENT|12838,12856|false|false|false|C0013182|Drug Allergy|medication allergy
Finding|Finding|SIMPLE_SEGMENT|12849,12856|false|false|false|C0020517;C0489531;C1314973;C1527304;C1547542;C3539909|Allergic Reaction;Allergic disposition;Allergy - Charge Type Reason;History of allergies;Hypersensitivity;Response to antigens|allergy
Finding|Idea or Concept|SIMPLE_SEGMENT|12849,12856|false|false|false|C0020517;C0489531;C1314973;C1527304;C1547542;C3539909|Allergic Reaction;Allergic disposition;Allergy - Charge Type Reason;History of allergies;Hypersensitivity;Response to antigens|allergy
Finding|Pathologic Function|SIMPLE_SEGMENT|12849,12856|false|false|false|C0020517;C0489531;C1314973;C1527304;C1547542;C3539909|Allergic Reaction;Allergic disposition;Allergy - Charge Type Reason;History of allergies;Hypersensitivity;Response to antigens|allergy
Finding|Physiologic Function|SIMPLE_SEGMENT|12849,12856|false|false|false|C0020517;C0489531;C1314973;C1527304;C1547542;C3539909|Allergic Reaction;Allergic disposition;Allergy - Charge Type Reason;History of allergies;Hypersensitivity;Response to antigens|allergy
Finding|Idea or Concept|SIMPLE_SEGMENT|12867,12874|false|false|false|C0392360|Indication of (contextual qualifier)|reasons
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12889,12898|false|false|false|C0804815||physician
Finding|Intellectual Product|SIMPLE_SEGMENT|12908,12916|false|false|false|C0237607;C3245512|Experience (Practice);HL7PublishingSubSection - practice|practice
Finding|Mental Process|SIMPLE_SEGMENT|12908,12916|false|false|false|C0237607;C3245512|Experience (Practice);HL7PublishingSubSection - practice|practice
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12924,12933|false|false|false|C0804815||physician
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12939,12948|false|false|false|C0804815||physician
Finding|Gene or Genome|SIMPLE_SEGMENT|12949,12952|false|false|false|C2986617|ANPEP wt Allele|APN
Finding|Idea or Concept|SIMPLE_SEGMENT|12960,12970|false|false|false|C1546966|Primary Observer's Qualification - Pharmacist|pharmacist
Drug|Biologically Active Substance|SIMPLE_SEGMENT|12975,12978|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Drug|Organic Chemical|SIMPLE_SEGMENT|12975,12978|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|12975,12978|false|false|false|C0202117|Low density lipoprotein cholesterol measurement|LDL
Finding|Finding|SIMPLE_SEGMENT|13033,13040|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|SIMPLE_SEGMENT|13033,13040|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|13033,13040|false|false|false|C0087111|Therapeutic procedure|therapy
Finding|Finding|SIMPLE_SEGMENT|13046,13049|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Gene or Genome|SIMPLE_SEGMENT|13046,13049|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Idea or Concept|SIMPLE_SEGMENT|13046,13049|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Intellectual Product|SIMPLE_SEGMENT|13046,13049|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Gene or Genome|SIMPLE_SEGMENT|13051,13055|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|Type
Finding|Intellectual Product|SIMPLE_SEGMENT|13051,13055|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|Type
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13061,13073|false|false|false|C5214487|Antiplatelet|Antiplatelet
Finding|Finding|SIMPLE_SEGMENT|13080,13095|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|Anticoagulation
Finding|Physiologic Function|SIMPLE_SEGMENT|13080,13095|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|Anticoagulation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|13080,13095|false|false|false|C0003281|Anticoagulation Therapy|Anticoagulation
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|13123,13127|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|13123,13127|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|13123,13127|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|13123,13127|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Finding|SIMPLE_SEGMENT|13128,13143|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Finding|Physiologic Function|SIMPLE_SEGMENT|13128,13143|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|13128,13143|false|false|false|C0003281|Anticoagulation Therapy|anticoagulation
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|13162,13168|false|false|false|C0018792|Heart Atrium|atrial
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13170,13182|false|false|false|C0232197|Fibrillation|fibrillation
Finding|Pathologic Function|SIMPLE_SEGMENT|13183,13190|false|false|false|C0016385|Cardiac Flutter|flutter
Finding|Finding|SIMPLE_SEGMENT|13196,13199|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Gene or Genome|SIMPLE_SEGMENT|13196,13199|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Idea or Concept|SIMPLE_SEGMENT|13196,13199|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Intellectual Product|SIMPLE_SEGMENT|13196,13199|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Functional Concept|SIMPLE_SEGMENT|13219,13228|false|false|false|C1516691|Cognitive|Cognitive
Finding|Finding|SIMPLE_SEGMENT|13229,13239|false|false|false|C5441521|Complaint (finding)|complaints
Finding|Gene or Genome|SIMPLE_SEGMENT|13242,13245|false|false|false|C1417635;C1420797;C3538796|NDUFB3 gene;TNFAIP1 gene;TNFAIP1 wt Allele|B12
Finding|Intellectual Product|SIMPLE_SEGMENT|13252,13260|false|false|false|C3241998|one time|one time
Finding|Finding|SIMPLE_SEGMENT|13256,13260|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|13256,13260|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|13256,13260|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|13264,13279|false|false|false|C0242297|Dietary Supplementation|supplementation
Finding|Intellectual Product|SIMPLE_SEGMENT|13281,13285|false|false|false|C1720594|Then - dosing instruction fragment|then
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|13292,13296|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|13292,13296|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|13292,13296|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|13292,13296|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Gene or Genome|SIMPLE_SEGMENT|13297,13300|false|false|false|C1417635;C1420797;C3538796|NDUFB3 gene;TNFAIP1 gene;TNFAIP1 wt Allele|B12
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|13302,13317|false|false|false|C0242297|Dietary Supplementation|supplementation
Finding|Functional Concept|SIMPLE_SEGMENT|13320,13330|false|false|false|C0521023|treponemal|Treponemal
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|13331,13341|false|false|false|C0003241;C3495458|Antibodies;antibodies (medication)|antibodies
Drug|Immunologic Factor|SIMPLE_SEGMENT|13331,13341|false|false|false|C0003241;C3495458|Antibodies;antibodies (medication)|antibodies
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13331,13341|false|false|false|C0003241;C3495458|Antibodies;antibodies (medication)|antibodies
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|13331,13350|false|false|false|C0855852|Antibody NOS negative|antibodies negative
Finding|Classification|SIMPLE_SEGMENT|13342,13350|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|13342,13350|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|13342,13350|false|false|false|C5237010|Expression Negative|negative
Finding|Idea or Concept|SIMPLE_SEGMENT|13353,13361|false|false|false|C0750591|consider|consider
Finding|Functional Concept|SIMPLE_SEGMENT|13362,13371|false|false|false|C1516691|Cognitive|cognitive
Procedure|Health Care Activity|SIMPLE_SEGMENT|13382,13390|false|false|false|C0034927|Patient referral|referral
Finding|Classification|SIMPLE_SEGMENT|13394,13404|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|13394,13404|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Finding|SIMPLE_SEGMENT|13409,13415|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Finding|Intellectual Product|SIMPLE_SEGMENT|13409,13415|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Finding|Mental Process|SIMPLE_SEGMENT|13409,13415|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Finding|Finding|SIMPLE_SEGMENT|13417,13429|true|false|false|C1299586|Has difficulty doing (qualifier value)|difficulties
Event|Activity|SIMPLE_SEGMENT|13453,13464|false|false|false|C4321457|Examination|examination
Procedure|Health Care Activity|SIMPLE_SEGMENT|13453,13464|false|false|false|C0031809;C0582103|Medical Examination;Physical Examination|examination
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13467,13471|false|false|false|C0004238|Atrial Fibrillation|Afib
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|13467,13471|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Afib
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|13482,13487|false|false|false|C0030471;C1305231|Nasal sinus;Sinus - general anatomical term|sinus
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|13482,13487|false|false|false|C0016169|pathologic fistula|sinus
Drug|Organic Chemical|SIMPLE_SEGMENT|13482,13487|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13482,13487|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13488,13494|false|false|false|C0488347||pauses
Drug|Organic Chemical|SIMPLE_SEGMENT|13505,13512|false|false|false|C0012265|digoxin|digoxin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13505,13512|false|false|false|C0012265|digoxin|digoxin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|13505,13512|false|false|false|C0337449|Digoxin measurement|digoxin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13559,13562|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|13559,13562|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|13559,13562|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|13559,13562|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|SIMPLE_SEGMENT|13559,13562|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|13559,13562|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|SIMPLE_SEGMENT|13559,13562|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13559,13562|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Finding|Gene or Genome|SIMPLE_SEGMENT|13559,13562|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|SIMPLE_SEGMENT|13559,13562|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Drug|Organic Chemical|SIMPLE_SEGMENT|13591,13602|false|false|false|C0723712|Therapeutic brand of coal tar|therapeutic
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13591,13602|false|false|false|C0723712|Therapeutic brand of coal tar|therapeutic
Finding|Functional Concept|SIMPLE_SEGMENT|13591,13602|false|false|false|C0302350;C1547427|Therapeutic;Therapeutic - Location Service Code|therapeutic
Finding|Intellectual Product|SIMPLE_SEGMENT|13591,13602|false|false|false|C0302350;C1547427|Therapeutic;Therapeutic - Location Service Code|therapeutic
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|13591,13602|false|false|false|C0087111|Therapeutic procedure|therapeutic
Drug|Organic Chemical|SIMPLE_SEGMENT|13613,13620|false|false|false|C3530466|Eliquis|Eliquis
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13613,13620|false|false|false|C3530466|Eliquis|Eliquis
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|13629,13632|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|13629,13632|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|13629,13632|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|SIMPLE_SEGMENT|13629,13632|false|false|false|C1332410|BID gene|BID
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13653,13656|false|false|false|C1114365||age
Drug|Biologically Active Substance|SIMPLE_SEGMENT|13653,13656|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|SIMPLE_SEGMENT|13653,13656|false|false|false|C0162574|Glycation End Products, Advanced|age
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13661,13667|false|false|false|C0944911||weight
Finding|Finding|SIMPLE_SEGMENT|13661,13667|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|SIMPLE_SEGMENT|13661,13667|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|SIMPLE_SEGMENT|13661,13667|false|false|false|C1305866|Weighing patient|weight
Drug|Organic Chemical|SIMPLE_SEGMENT|13692,13704|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13692,13704|false|false|false|C0286651|atorvastatin|atorvastatin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13707,13710|false|false|false|C0020538|Hypertensive disease|HTN
Finding|Idea or Concept|SIMPLE_SEGMENT|13713,13721|false|false|false|C0549178|Continuous|continue
Finding|Idea or Concept|SIMPLE_SEGMENT|13722,13726|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|13722,13726|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|13722,13726|false|false|false|C1553498|home health encounter|home
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13727,13744|false|false|false|C0003364|Antihypertensive Agents|antihypertensives
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|13756,13764|false|false|false|C0041199|Troponin|troponin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|13756,13764|false|false|false|C0041199|Troponin|troponin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|13756,13764|false|false|false|C0523952|Troponin measurement|troponin
Finding|Conceptual Entity|SIMPLE_SEGMENT|13766,13774|false|false|false|C1514893;C2699488|Resolution;physiologic resolution|RESOLVED
Finding|Pathologic Function|SIMPLE_SEGMENT|13766,13774|false|false|false|C1514893;C2699488|Resolution;physiologic resolution|RESOLVED
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|13778,13786|false|false|false|C0041199|Troponin|Troponin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|13778,13786|false|false|false|C0041199|Troponin|Troponin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|13778,13786|false|false|false|C0523952|Troponin measurement|Troponin
Finding|Classification|SIMPLE_SEGMENT|13804,13812|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|13804,13812|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|13804,13812|false|false|false|C5237010|Expression Negative|negative
Procedure|Health Care Activity|SIMPLE_SEGMENT|13816,13825|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Finding|SIMPLE_SEGMENT|13828,13840|false|false|false|C0586553|Raised TSH level|elevated TSH
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13837,13840|false|false|false|C2708739||TSH
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|13837,13840|false|false|false|C0040160|thyrotropin|TSH
Drug|Hormone|SIMPLE_SEGMENT|13837,13840|false|false|false|C0040160|thyrotropin|TSH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13837,13840|false|false|false|C0040160|thyrotropin|TSH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|13837,13840|false|false|false|C0202230|Thyroid stimulating hormone measurement|TSH
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13869,13872|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|13869,13872|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|13869,13872|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|13869,13872|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|SIMPLE_SEGMENT|13869,13872|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|13869,13872|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|SIMPLE_SEGMENT|13869,13872|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13869,13872|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Finding|Gene or Genome|SIMPLE_SEGMENT|13869,13872|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|SIMPLE_SEGMENT|13869,13872|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13879,13890|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13879,13890|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|13879,13890|false|false|false|C4284232|Medications|Medications
Finding|Finding|SIMPLE_SEGMENT|13879,13903|false|false|false|C1627937|Medications on admission|Medications on Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|13894,13903|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13922,13932|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|13922,13932|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|13922,13937|false|false|false|C0746470|MEDICATION LIST|Medication list
Finding|Intellectual Product|SIMPLE_SEGMENT|13933,13937|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Drug|Organic Chemical|SIMPLE_SEGMENT|13954,13962|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13954,13962|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|SIMPLE_SEGMENT|13954,13962|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Finding|Functional Concept|SIMPLE_SEGMENT|13954,13962|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|SIMPLE_SEGMENT|13954,13962|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Organic Chemical|SIMPLE_SEGMENT|13967,13975|false|false|false|C0004147|atenolol|Atenolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13967,13975|false|false|false|C0004147|atenolol|Atenolol
Drug|Organic Chemical|SIMPLE_SEGMENT|13995,14003|false|false|false|C1831808|apixaban|Apixaban
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13995,14003|false|false|false|C1831808|apixaban|Apixaban
Drug|Organic Chemical|SIMPLE_SEGMENT|14024,14032|false|false|false|C0126174|losartan|Losartan
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14024,14032|false|false|false|C0126174|losartan|Losartan
Drug|Organic Chemical|SIMPLE_SEGMENT|14024,14042|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14024,14042|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|14033,14042|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|14033,14042|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Food|SIMPLE_SEGMENT|14033,14042|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|14033,14042|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14033,14042|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Finding|Physiologic Function|SIMPLE_SEGMENT|14033,14042|false|false|false|C4553027|Potassium metabolic function|Potassium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|14033,14042|false|false|false|C0202194|Potassium measurement|Potassium
Drug|Organic Chemical|SIMPLE_SEGMENT|14062,14069|false|false|false|C0012265|digoxin|Digoxin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14062,14069|false|false|false|C0012265|digoxin|Digoxin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|14062,14069|false|false|false|C0337449|Digoxin measurement|Digoxin
Drug|Antibiotic|SIMPLE_SEGMENT|14092,14104|false|false|false|C0282386|levofloxacin|LevoFLOXacin
Drug|Organic Chemical|SIMPLE_SEGMENT|14092,14104|false|false|false|C0282386|levofloxacin|LevoFLOXacin
Finding|Body Substance|SIMPLE_SEGMENT|14124,14133|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|14124,14133|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|14124,14133|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|14124,14133|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|14124,14145|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14134,14145|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14134,14145|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|14134,14145|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|SIMPLE_SEGMENT|14151,14163|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14151,14163|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|SIMPLE_SEGMENT|14182,14194|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14182,14194|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|14203,14209|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|SIMPLE_SEGMENT|14213,14221|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|14216,14221|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|14216,14221|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Intellectual Product|SIMPLE_SEGMENT|14222,14226|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|14255,14261|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|SIMPLE_SEGMENT|14262,14269|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|14278,14292|false|false|false|C0042845;C3714801|Cyanocobalamin Drug Class;vitamin B12|Cyanocobalamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14278,14292|false|false|false|C0042845;C3714801|Cyanocobalamin Drug Class;vitamin B12|Cyanocobalamin
Drug|Vitamin|SIMPLE_SEGMENT|14278,14292|false|false|false|C0042845;C3714801|Cyanocobalamin Drug Class;vitamin B12|Cyanocobalamin
Drug|Organic Chemical|SIMPLE_SEGMENT|14315,14329|false|false|false|C0042845;C3714801|Cyanocobalamin Drug Class;vitamin B12|cyanocobalamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14315,14329|false|false|false|C0042845;C3714801|Cyanocobalamin Drug Class;vitamin B12|cyanocobalamin
Drug|Vitamin|SIMPLE_SEGMENT|14315,14329|false|false|false|C0042845;C3714801|Cyanocobalamin Drug Class;vitamin B12|cyanocobalamin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|14315,14344|false|false|false|C0202252|VITAMIN B12 MEASUREMENT|cyanocobalamin (vitamin B-12)
Drug|Organic Chemical|SIMPLE_SEGMENT|14331,14338|false|false|false|C0042890|Vitamins|vitamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14331,14338|false|false|false|C0042890|Vitamins|vitamin
Drug|Vitamin|SIMPLE_SEGMENT|14331,14338|false|false|false|C0042890|Vitamins|vitamin
Drug|Organic Chemical|SIMPLE_SEGMENT|14331,14340|false|false|false|C0042849;C1704763;C5442122|B Vitamin Family;VITAMIN B;vitamin B complex|vitamin B
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14331,14340|false|false|false|C0042849;C1704763;C5442122|B Vitamin Family;VITAMIN B;vitamin B complex|vitamin B
Drug|Vitamin|SIMPLE_SEGMENT|14331,14340|false|false|false|C0042849;C1704763;C5442122|B Vitamin Family;VITAMIN B;vitamin B complex|vitamin B
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|14331,14343|false|false|false|C0042845;C0086024|cobalamins;vitamin B12|vitamin B-12
Drug|Organic Chemical|SIMPLE_SEGMENT|14331,14343|false|false|false|C0042845;C0086024|cobalamins;vitamin B12|vitamin B-12
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14331,14343|false|false|false|C0042845;C0086024|cobalamins;vitamin B12|vitamin B-12
Drug|Vitamin|SIMPLE_SEGMENT|14331,14343|false|false|false|C0042845;C0086024|cobalamins;vitamin B12|vitamin B-12
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|14331,14343|false|false|false|C0202252|VITAMIN B12 MEASUREMENT|vitamin B-12
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|14355,14361|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|SIMPLE_SEGMENT|14365,14373|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|14368,14373|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|14368,14373|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Intellectual Product|SIMPLE_SEGMENT|14375,14379|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|14396,14402|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|SIMPLE_SEGMENT|14403,14410|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|14419,14427|false|false|false|C1831808|apixaban|Apixaban
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14419,14427|false|false|false|C1831808|apixaban|Apixaban
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|14438,14441|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|14438,14441|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|14438,14441|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|SIMPLE_SEGMENT|14438,14441|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|14448,14456|false|false|false|C0004147|atenolol|Atenolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14448,14456|false|false|false|C0004147|atenolol|Atenolol
Drug|Antibiotic|SIMPLE_SEGMENT|14478,14490|false|false|false|C0282386|levofloxacin|LevoFLOXacin
Drug|Organic Chemical|SIMPLE_SEGMENT|14478,14490|false|false|false|C0282386|levofloxacin|LevoFLOXacin
Drug|Organic Chemical|SIMPLE_SEGMENT|14512,14520|false|false|false|C0126174|losartan|Losartan
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14512,14520|false|false|false|C0126174|losartan|Losartan
Drug|Organic Chemical|SIMPLE_SEGMENT|14512,14530|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14512,14530|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|14521,14530|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|14521,14530|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Food|SIMPLE_SEGMENT|14521,14530|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|14521,14530|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14521,14530|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Finding|Physiologic Function|SIMPLE_SEGMENT|14521,14530|false|false|false|C4553027|Potassium metabolic function|Potassium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|14521,14530|false|false|false|C0202194|Potassium measurement|Potassium
Finding|Body Substance|SIMPLE_SEGMENT|14551,14560|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|14551,14560|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|14551,14560|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|14551,14560|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14551,14572|false|false|false|C4019243||Discharge Disposition
Finding|Finding|SIMPLE_SEGMENT|14551,14572|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14561,14572|false|false|false|C2926604||Disposition
Procedure|Health Care Activity|SIMPLE_SEGMENT|14561,14572|false|false|false|C0184758|Patient disposition|Disposition
Finding|Idea or Concept|SIMPLE_SEGMENT|14574,14578|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|SIMPLE_SEGMENT|14574,14578|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|SIMPLE_SEGMENT|14574,14578|false|false|false|C1553498|home health encounter|Home
Event|Occupational Activity|SIMPLE_SEGMENT|14584,14591|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|14584,14591|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Finding|Intellectual Product|SIMPLE_SEGMENT|14594,14602|false|false|false|C4695111|ADMIN.FACILITY|Facility
Finding|Body Substance|SIMPLE_SEGMENT|14610,14619|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|14610,14619|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|14610,14619|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|14610,14619|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|14610,14629|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14620,14629|false|false|false|C0945731||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|14620,14629|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|14620,14629|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|14620,14629|false|false|false|C0011900|Diagnosis|Diagnosis
Finding|Finding|SIMPLE_SEGMENT|14631,14640|false|false|false|C0687129;C1550450|Encounter due to vagabond status;Living Arrangement - Transient|transient
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|14641,14651|false|false|false|C0013362|Dysarthria|dysarthria
Disorder|Neoplastic Process|SIMPLE_SEGMENT|14656,14665|true|false|false|C0027627|Neoplasm Metastasis|secondary
Finding|Functional Concept|SIMPLE_SEGMENT|14656,14665|true|false|false|C1522484|metastatic qualifier|secondary
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14669,14672|false|false|false|C0007787;C0917805|Transient Cerebral Ischemia;Transient Ischemic Attack|TIA
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14676,14682|false|true|false|C0038454|Cerebrovascular accident|stroke
Finding|Finding|SIMPLE_SEGMENT|14676,14682|false|true|false|C5977286|Stroke (heart beat)|stroke
Finding|Intellectual Product|SIMPLE_SEGMENT|14683,14687|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Drug|Organic Chemical|SIMPLE_SEGMENT|14688,14695|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14688,14695|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|SIMPLE_SEGMENT|14688,14695|false|false|false|C0042890|Vitamins|Vitamin
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|14688,14699|false|false|false|C0042845;C0086024;C2936883|Vitamin B12 [EPC];cobalamins;vitamin B12|Vitamin B12
Drug|Organic Chemical|SIMPLE_SEGMENT|14688,14699|false|false|false|C0042845;C0086024;C2936883|Vitamin B12 [EPC];cobalamins;vitamin B12|Vitamin B12
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14688,14699|false|false|false|C0042845;C0086024;C2936883|Vitamin B12 [EPC];cobalamins;vitamin B12|Vitamin B12
Drug|Vitamin|SIMPLE_SEGMENT|14688,14699|false|false|false|C0042845;C0086024;C2936883|Vitamin B12 [EPC];cobalamins;vitamin B12|Vitamin B12
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|14688,14699|false|false|false|C0202252|VITAMIN B12 MEASUREMENT|Vitamin B12
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14688,14710|false|false|false|C0042847|Vitamin B 12 Deficiency|Vitamin B12 deficiency
Finding|Finding|SIMPLE_SEGMENT|14688,14710|false|false|false|C5886863|Decreased circulating vitamin B12 concentration|Vitamin B12 deficiency
Finding|Gene or Genome|SIMPLE_SEGMENT|14696,14699|false|false|false|C1417635;C1420797;C3538796|NDUFB3 gene;TNFAIP1 gene;TNFAIP1 wt Allele|B12
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14700,14710|false|false|false|C0162429|Malnutrition|deficiency
Finding|Functional Concept|SIMPLE_SEGMENT|14700,14710|false|false|false|C0011155|Deficiency|deficiency
Finding|Body Substance|SIMPLE_SEGMENT|14713,14722|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|14713,14722|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|14713,14722|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|14713,14722|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14723,14732|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14723,14732|false|false|false|C0012634|Disease|Condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|14723,14732|false|false|false|C1705253|Logical Condition|Condition
Finding|Mental Process|SIMPLE_SEGMENT|14734,14740|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14734,14747|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|SIMPLE_SEGMENT|14734,14747|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14741,14747|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|14741,14747|false|false|false|C1546481|What subject filter - Status|Status
Finding|Idea or Concept|SIMPLE_SEGMENT|14749,14754|false|false|false|C1550016|Remote control command - Clear|Clear
Finding|Finding|SIMPLE_SEGMENT|14759,14767|false|false|false|C4068804|Coherent|coherent
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14769,14791|false|false|false|C4050479||Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|14769,14791|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|14778,14791|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|SIMPLE_SEGMENT|14778,14791|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14793,14798|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|14793,14798|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14793,14798|false|false|false|C0718338|Alert brand of caffeine|Alert
Finding|Finding|SIMPLE_SEGMENT|14793,14798|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|14793,14798|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|14793,14798|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|14803,14814|false|false|false|C1704675|Interaction|interactive
Event|Activity|SIMPLE_SEGMENT|14816,14824|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|14816,14824|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|SIMPLE_SEGMENT|14816,14824|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14825,14831|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|14825,14831|false|false|false|C1546481|What subject filter - Status|Status
Finding|Functional Concept|SIMPLE_SEGMENT|14833,14843|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|SIMPLE_SEGMENT|14833,14843|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|SIMPLE_SEGMENT|14833,14843|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|SIMPLE_SEGMENT|14833,14843|false|false|false|C1561560|ambulatory encounter|Ambulatory
Finding|Social Behavior|SIMPLE_SEGMENT|14855,14865|false|false|false|C0018896|Helping Behavior|assistance
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|14869,14872|false|false|false|C1454018|AICDA protein, human|aid
Drug|Enzyme|SIMPLE_SEGMENT|14869,14872|false|false|false|C1454018|AICDA protein, human|aid
Finding|Gene or Genome|SIMPLE_SEGMENT|14869,14872|false|false|false|C1421876;C3540469|AICDA gene;AICDA wt Allele|aid
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|14869,14872|false|false|false|C0021588;C0280108|AID - Artificial insemination by donor;dacarbazine/doxorubicin/ifosfamide protocol|aid
Finding|Body Substance|SIMPLE_SEGMENT|14894,14903|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|14894,14903|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|14894,14903|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|14894,14903|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14894,14916|false|false|false|C3669312||Discharge Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|14894,14916|false|false|false|C4282220|Discharge instructions|Discharge Instructions
Procedure|Health Care Activity|SIMPLE_SEGMENT|14894,14916|false|false|false|C2266673|hospital discharge instructions (treatment)|Discharge Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14904,14916|false|false|false|C3263700||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|14904,14916|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Finding|Gene or Genome|SIMPLE_SEGMENT|14918,14922|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Finding|Functional Concept|SIMPLE_SEGMENT|14962,14970|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|14962,14970|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Organism Function|SIMPLE_SEGMENT|14982,14988|false|false|false|C0037817|Speech|speech
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|14982,14988|false|false|false|C0846595|Speech assessment|speech
Finding|Idea or Concept|SIMPLE_SEGMENT|14997,15004|false|false|false|C2699424|Concern|concern
Finding|Intellectual Product|SIMPLE_SEGMENT|15012,15017|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|ACUTE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15012,15033|false|false|false|C5392833|Acute Ischemic Stroke|ACUTE ISCHEMIC STROKE
Finding|Functional Concept|SIMPLE_SEGMENT|15018,15026|false|false|false|C0475224|Ischemic|ISCHEMIC
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15018,15033|false|false|false|C0948008|Ischemic stroke|ISCHEMIC STROKE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15027,15033|false|false|false|C0038454|Cerebrovascular accident|STROKE
Finding|Finding|SIMPLE_SEGMENT|15027,15033|false|false|false|C5977286|Stroke (heart beat)|STROKE
Attribute|Clinical Attribute|SIMPLE_SEGMENT|15037,15046|false|false|false|C3864998||condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15037,15046|false|false|false|C0012634|Disease|condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|15037,15046|false|false|false|C1705253|Logical Condition|condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15055,15060|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|SIMPLE_SEGMENT|15055,15060|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Anatomy|Body Location or Region|SIMPLE_SEGMENT|15062,15068|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|15062,15068|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Drug|Biologically Active Substance|SIMPLE_SEGMENT|15079,15085|false|false|false|C0030054|oxygen|oxygen
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|15079,15085|false|false|false|C0030054|oxygen|oxygen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|15079,15085|false|false|false|C0030054|oxygen|oxygen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|15079,15085|false|false|false|C0184633|Oxygen Therapy Care|oxygen
Drug|Food|SIMPLE_SEGMENT|15090,15099|false|false|false|C0678695|Nutrients|nutrients
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|15107,15112|false|false|false|C0006104;C4266577|Brain;Head>Brain|brain
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15107,15112|false|false|false|C0006111|Brain Diseases|brain
Drug|Organic Chemical|SIMPLE_SEGMENT|15130,15134|false|false|false|C0009074|clotrimazole|clot
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|15130,15134|false|false|false|C0009074|clotrimazole|clot
Finding|Pathologic Function|SIMPLE_SEGMENT|15130,15134|false|false|false|C0302148|Blood Clot|clot
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|15140,15145|false|false|false|C0006104;C4266577|Brain;Head>Brain|brain
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15140,15145|false|false|false|C0006111|Brain Diseases|brain
Finding|Idea or Concept|SIMPLE_SEGMENT|15153,15157|false|false|false|C1552020|Role Class - part|part
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|15166,15170|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|15166,15170|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Finding|Intellectual Product|SIMPLE_SEGMENT|15166,15170|false|false|false|C1551342|Document Body|body
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|15226,15230|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|15226,15230|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Finding|Intellectual Product|SIMPLE_SEGMENT|15226,15230|false|false|false|C1551342|Document Body|body
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|15235,15241|false|false|false|C0010957|Tissue damage|damage
Finding|Functional Concept|SIMPLE_SEGMENT|15235,15241|false|false|false|C1883709;C2681922|Damage;MAGEE1 gene|damage
Finding|Gene or Genome|SIMPLE_SEGMENT|15235,15241|false|false|false|C1883709;C2681922|Damage;MAGEE1 gene|damage
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|15249,15254|false|false|false|C0006104;C4266577|Brain;Head>Brain|brain
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15249,15254|false|false|false|C0006111|Brain Diseases|brain
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15283,15288|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|SIMPLE_SEGMENT|15283,15288|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|15283,15295|false|false|false|C0678861;C0920762|Arterial blood supply;Vascular blood supply|blood supply
Finding|Physiologic Function|SIMPLE_SEGMENT|15283,15295|false|false|false|C0678861;C0920762|Arterial blood supply;Vascular blood supply|blood supply
Event|Activity|SIMPLE_SEGMENT|15289,15295|false|false|false|C1999230|Providing (action)|supply
Finding|Functional Concept|SIMPLE_SEGMENT|15289,15295|false|false|false|C0243163;C1561604;C4760136|Supply (process);Supply (system);supply aspects|supply
Finding|Idea or Concept|SIMPLE_SEGMENT|15289,15295|false|false|false|C0243163;C1561604;C4760136|Supply (process);Supply (system);supply aspects|supply
Finding|Conceptual Entity|SIMPLE_SEGMENT|15312,15319|false|false|false|C1883525;C2346866|Assortment;Variety (taxon)|variety
Finding|Functional Concept|SIMPLE_SEGMENT|15324,15332|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|15324,15332|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Gene or Genome|SIMPLE_SEGMENT|15347,15350|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|15347,15350|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|SIMPLE_SEGMENT|15347,15350|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|15359,15364|false|false|false|C0006104;C4266577|Brain;Head>Brain|brain
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15359,15364|false|false|false|C0006111|Brain Diseases|brain
Finding|Idea or Concept|SIMPLE_SEGMENT|15379,15387|false|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|15379,15390|false|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15391,15397|false|false|false|C0038454|Cerebrovascular accident|stroke
Finding|Finding|SIMPLE_SEGMENT|15391,15397|false|false|false|C5977286|Stroke (heart beat)|stroke
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15401,15404|false|false|false|C0007787;C0917805|Transient Cerebral Ischemia;Transient Ischemic Attack|TIA
Finding|Functional Concept|SIMPLE_SEGMENT|15411,15419|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|15411,15419|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Drug|Organic Chemical|SIMPLE_SEGMENT|15436,15443|false|false|false|C0163712|Relate - vinyl resin|related
Finding|Finding|SIMPLE_SEGMENT|15436,15443|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Finding|Functional Concept|SIMPLE_SEGMENT|15436,15443|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15448,15453|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|SIMPLE_SEGMENT|15448,15453|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Finding|SIMPLE_SEGMENT|15448,15462|false|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|blood pressure
Finding|Organism Function|SIMPLE_SEGMENT|15448,15462|false|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|blood pressure
Procedure|Health Care Activity|SIMPLE_SEGMENT|15448,15462|false|false|false|C0005824|Blood pressure determination|blood pressure
Finding|Finding|SIMPLE_SEGMENT|15454,15462|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|SIMPLE_SEGMENT|15454,15462|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|15454,15462|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|15454,15462|false|false|false|C0033095||pressure
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15464,15475|false|false|false|C0011175;C2062903|Dehydration;dehydration (Na, H2O)|dehydration
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|15464,15475|false|false|false|C0011175;C2062903|Dehydration;dehydration (Na, H2O)|dehydration
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|15464,15475|false|false|false|C4284399|Dehydration procedure|dehydration
Drug|Organic Chemical|SIMPLE_SEGMENT|15477,15484|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|15477,15484|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Finding|Intellectual Product|SIMPLE_SEGMENT|15477,15484|false|false|false|C1547288|Alcohol - Recreational Drug Use Code|alcohol
Finding|Finding|SIMPLE_SEGMENT|15477,15488|false|false|false|C0001948;C0552479|Alcohol consumption;history of alcohol use|alcohol use
Finding|Individual Behavior|SIMPLE_SEGMENT|15477,15488|false|false|false|C0001948;C0552479|Alcohol consumption;history of alcohol use|alcohol use
Finding|Functional Concept|SIMPLE_SEGMENT|15485,15488|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|SIMPLE_SEGMENT|15485,15488|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Finding|SIMPLE_SEGMENT|15495,15506|false|false|false|C3811910|combination - answer to question|combination
Attribute|Clinical Attribute|SIMPLE_SEGMENT|15548,15559|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|15548,15559|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|SIMPLE_SEGMENT|15548,15559|false|false|false|C4284232|Medications|medications
Drug|Organic Chemical|SIMPLE_SEGMENT|15581,15589|false|false|false|C1831808|apixaban|apixaban
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|15581,15589|false|false|false|C1831808|apixaban|apixaban
Drug|Organic Chemical|SIMPLE_SEGMENT|15617,15624|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|15617,15624|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|SIMPLE_SEGMENT|15617,15624|false|false|false|C0042890|Vitamins|Vitamin
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|15617,15628|false|false|false|C0042845;C0086024;C2936883|Vitamin B12 [EPC];cobalamins;vitamin B12|Vitamin B12
Drug|Organic Chemical|SIMPLE_SEGMENT|15617,15628|false|false|false|C0042845;C0086024;C2936883|Vitamin B12 [EPC];cobalamins;vitamin B12|Vitamin B12
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|15617,15628|false|false|false|C0042845;C0086024;C2936883|Vitamin B12 [EPC];cobalamins;vitamin B12|Vitamin B12
Drug|Vitamin|SIMPLE_SEGMENT|15617,15628|false|false|false|C0042845;C0086024;C2936883|Vitamin B12 [EPC];cobalamins;vitamin B12|Vitamin B12
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|15617,15628|false|false|false|C0202252|VITAMIN B12 MEASUREMENT|Vitamin B12
Finding|Gene or Genome|SIMPLE_SEGMENT|15625,15628|false|false|false|C1417635;C1420797;C3538796|NDUFB3 gene;TNFAIP1 gene;TNFAIP1 wt Allele|B12
Drug|Food|SIMPLE_SEGMENT|15635,15645|false|false|false|C0242295|Dietary Supplements|supplement
Finding|Functional Concept|SIMPLE_SEGMENT|15635,15645|false|false|false|C1549514;C1947943;C2348609|Supplement;Supplement (document);Supplement - Diet Code Specification Type|supplement
Finding|Idea or Concept|SIMPLE_SEGMENT|15635,15645|false|false|false|C1549514;C1947943;C2348609|Supplement;Supplement (document);Supplement - Diet Code Specification Type|supplement
Finding|Intellectual Product|SIMPLE_SEGMENT|15635,15645|false|false|false|C1549514;C1947943;C2348609|Supplement;Supplement (document);Supplement - Diet Code Specification Type|supplement
Attribute|Clinical Attribute|SIMPLE_SEGMENT|15670,15681|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|15670,15681|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|SIMPLE_SEGMENT|15670,15681|false|false|false|C4284232|Medications|medications
Finding|Intellectual Product|SIMPLE_SEGMENT|15725,15737|false|false|false|C1547426|Location Service Code - Primary Care|primary care
Procedure|Health Care Activity|SIMPLE_SEGMENT|15725,15737|false|false|false|C0033137|Primary Health Care|primary care
Event|Activity|SIMPLE_SEGMENT|15733,15737|false|false|false|C1947933|care activity|care
Finding|Finding|SIMPLE_SEGMENT|15733,15737|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|15733,15737|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Attribute|Clinical Attribute|SIMPLE_SEGMENT|15738,15747|false|false|false|C0804815||physician
Attribute|Clinical Attribute|SIMPLE_SEGMENT|15853,15859|false|false|false|C0488347||pauses
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|15863,15870|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|15863,15870|false|false|false|C1314974|Cardiac attachment|cardiac
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|15863,15881|false|false|false|C0150496|Cardiac monitoring|cardiac monitoring
Event|Activity|SIMPLE_SEGMENT|15871,15881|false|false|false|C1283169||monitoring
Procedure|Health Care Activity|SIMPLE_SEGMENT|15871,15881|false|false|false|C0150369|Preventive monitoring|monitoring
Finding|Functional Concept|SIMPLE_SEGMENT|15913,15921|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|15913,15921|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Finding|SIMPLE_SEGMENT|15942,15951|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Idea or Concept|SIMPLE_SEGMENT|15942,15951|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Intellectual Product|SIMPLE_SEGMENT|15942,15951|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Pathologic Function|SIMPLE_SEGMENT|15942,15951|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|15942,15951|false|false|false|C0013956|Emergency Situation|emergency
Procedure|Health Care Activity|SIMPLE_SEGMENT|15942,15951|false|false|false|C1553500|emergency encounter|emergency
Finding|Functional Concept|SIMPLE_SEGMENT|15952,15959|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Idea or Concept|SIMPLE_SEGMENT|15952,15959|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Intellectual Product|SIMPLE_SEGMENT|15952,15959|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|15952,15959|false|false|false|C0199168|Medical service|medical
Finding|Intellectual Product|SIMPLE_SEGMENT|15960,15969|false|false|false|C0004268;C4281780|Attention;Attention - G-code|attention
Finding|Mental Process|SIMPLE_SEGMENT|15960,15969|false|false|false|C0004268;C4281780|Attention;Attention - G-code|attention
Finding|Finding|SIMPLE_SEGMENT|15981,15990|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Finding|Idea or Concept|SIMPLE_SEGMENT|15981,15990|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Finding|Intellectual Product|SIMPLE_SEGMENT|15981,15990|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Finding|Pathologic Function|SIMPLE_SEGMENT|15981,15990|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|15981,15990|false|false|false|C0013956|Emergency Situation|Emergency
Procedure|Health Care Activity|SIMPLE_SEGMENT|15981,15990|false|false|false|C1553500|emergency encounter|Emergency
Finding|Functional Concept|SIMPLE_SEGMENT|15991,15998|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|15991,15998|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|15991,15998|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|15991,15998|false|false|false|C0199168|Medical service|Medical
Event|Occupational Activity|SIMPLE_SEGMENT|16000,16008|false|false|false|C0557854|Services|Services
Procedure|Health Care Activity|SIMPLE_SEGMENT|16000,16008|false|false|false|C1704289|Clinical Service|Services
Finding|Intellectual Product|SIMPLE_SEGMENT|16050,16059|false|false|false|C0004268;C4281780|Attention;Attention - G-code|attention
Finding|Mental Process|SIMPLE_SEGMENT|16050,16059|false|false|false|C0004268;C4281780|Attention;Attention - G-code|attention
Finding|Intellectual Product|SIMPLE_SEGMENT|16068,16080|false|false|false|C1272517|Sudden onset (contextual qualifier) (qualifier value)|sudden onset
Finding|Mental Process|SIMPLE_SEGMENT|16085,16096|false|false|false|C0546816|Persistence|persistence
Finding|Functional Concept|SIMPLE_SEGMENT|16106,16114|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|16106,16114|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Idea or Concept|SIMPLE_SEGMENT|16125,16132|false|false|false|C1550516|Target Awareness - partial|partial
Drug|Organic Chemical|SIMPLE_SEGMENT|16136,16144|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|16136,16144|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|SIMPLE_SEGMENT|16136,16144|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Finding|Functional Concept|SIMPLE_SEGMENT|16136,16144|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|SIMPLE_SEGMENT|16136,16144|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Finding|SIMPLE_SEGMENT|16145,16149|false|false|false|C5890125|Loss (adaptation)|loss
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|16145,16159|false|false|false|C0042798;C0456909|Blindness;Low Vision|loss of vision
Finding|Finding|SIMPLE_SEGMENT|16145,16159|false|false|false|C3665346;C3665386|Abnormal vision;Unspecified visual loss|loss of vision
Finding|Sign or Symptom|SIMPLE_SEGMENT|16145,16159|false|false|false|C3665346;C3665386|Abnormal vision;Unspecified visual loss|loss of vision
Attribute|Clinical Attribute|SIMPLE_SEGMENT|16153,16159|false|false|false|C2707266||vision
Finding|Organism Function|SIMPLE_SEGMENT|16153,16159|false|false|false|C0042789|Vision|vision
Finding|Finding|SIMPLE_SEGMENT|16169,16173|false|false|false|C5890125|Loss (adaptation)|loss
Finding|Functional Concept|SIMPLE_SEGMENT|16181,16188|false|false|false|C5891046|Oral Intake Ability|ability
Finding|Intellectual Product|SIMPLE_SEGMENT|16181,16191|false|false|false|C5420000|Ability Question|ability to
Anatomy|Body Location or Region|SIMPLE_SEGMENT|16214,16219|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|16214,16219|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Finding|SIMPLE_SEGMENT|16229,16233|false|false|false|C5890125|Loss (adaptation)|loss
Finding|Functional Concept|SIMPLE_SEGMENT|16241,16248|false|false|false|C5891046|Oral Intake Ability|ability
Finding|Intellectual Product|SIMPLE_SEGMENT|16241,16251|false|false|false|C5420000|Ability Question|ability to
Finding|Sign or Symptom|SIMPLE_SEGMENT|16296,16304|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|16324,16328|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|16324,16328|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Finding|Intellectual Product|SIMPLE_SEGMENT|16324,16328|false|false|false|C1551342|Document Body|body
Anatomy|Body Location or Region|SIMPLE_SEGMENT|16366,16370|false|false|false|C0015450;C4266571|Face;Head>Face|face
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|16366,16370|false|false|false|C3160739|FANCONI ANEMIA, COMPLEMENTATION GROUP E|face
Finding|Gene or Genome|SIMPLE_SEGMENT|16366,16370|false|false|false|C1414531;C1423759;C2828055|ELOVL6 gene;FANCE gene;FANCE wt Allele|face
Finding|Finding|SIMPLE_SEGMENT|16380,16384|false|false|false|C5890125|Loss (adaptation)|loss
Finding|Sign or Symptom|SIMPLE_SEGMENT|16380,16397|false|false|false|C0028643|Numbness|loss of sensation
Finding|Finding|SIMPLE_SEGMENT|16388,16397|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|16388,16397|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|SIMPLE_SEGMENT|16388,16397|false|false|false|C2229507|sensory exam|sensation
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|16417,16421|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|16417,16421|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Finding|Intellectual Product|SIMPLE_SEGMENT|16417,16421|false|false|false|C1551342|Document Body|body
Procedure|Health Care Activity|SIMPLE_SEGMENT|16460,16468|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|16469,16481|false|false|false|C3263700||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|16469,16481|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

