 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|46,55|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|46,55|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|46,60|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|80,89|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|80,89|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|80,94|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|136,139|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|147,154|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|147,154|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|156,164|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|SIMPLE_SEGMENT|167,176|false|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|167,176|false|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|167,176|false|false|false|C0020517|Hypersensitivity|Allergies
Drug|Antibiotic|SIMPLE_SEGMENT|179,190|false|false|false|C0002645|amoxicillin|amoxicillin
Drug|Organic Chemical|SIMPLE_SEGMENT|179,190|false|false|false|C0002645|amoxicillin|amoxicillin
Event|Event|SIMPLE_SEGMENT|179,190|false|false|false|||amoxicillin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|193,197|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|193,197|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|193,197|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Event|Event|SIMPLE_SEGMENT|193,197|false|false|false|||iron
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|193,197|false|false|false|C0337439|Iron measurement|iron
Event|Event|SIMPLE_SEGMENT|200,209|false|false|false|||Attending
Finding|Functional Concept|SIMPLE_SEGMENT|200,209|false|false|false|C1999232|Attending (action)|Attending
Finding|Classification|SIMPLE_SEGMENT|218,223|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|SIMPLE_SEGMENT|224,232|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|224,232|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|236,254|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|245,254|false|false|false|C0945766||Procedure
Event|Event|SIMPLE_SEGMENT|245,254|false|false|false|||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|245,254|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|245,254|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|245,254|false|false|false|C0184661|Interventional procedure|Procedure
Event|Event|SIMPLE_SEGMENT|262,268|false|false|false|||attach
Finding|Intellectual Product|SIMPLE_SEGMENT|262,268|false|false|false|C1314972;C2598091|Claims attachment;HIPAA attachments|attach
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|262,268|false|false|false|C3714578|Fix|attach
Procedure|Health Care Activity|SIMPLE_SEGMENT|290,299|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|SIMPLE_SEGMENT|300,304|false|false|false|||LABS
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|300,304|false|false|false|C0587081|Laboratory test finding|LABS
Event|Event|SIMPLE_SEGMENT|336,339|false|false|false|||PLT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|336,339|false|false|false|C0201617|Primed lymphocyte test|PLT
Drug|Antibiotic|SIMPLE_SEGMENT|379,384|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|379,384|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Organic Chemical|SIMPLE_SEGMENT|379,384|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Event|Event|SIMPLE_SEGMENT|379,384|false|false|false|||MONOS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|390,393|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|EOS
Event|Event|SIMPLE_SEGMENT|390,393|false|false|false|||EOS
Finding|Gene or Genome|SIMPLE_SEGMENT|390,393|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|EOS
Anatomy|Cell|SIMPLE_SEGMENT|496,499|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|504,507|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|504,507|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|504,507|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|513,516|false|false|false|C0019046|Hemoglobin|HGB
Drug|Biologically Active Substance|SIMPLE_SEGMENT|513,516|false|false|false|C0019046|Hemoglobin|HGB
Event|Event|SIMPLE_SEGMENT|513,516|false|false|false|||HGB
Finding|Gene or Genome|SIMPLE_SEGMENT|513,516|false|false|false|C1424337|CYGB gene|HGB
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|513,516|false|false|false|C0019029|Hemoglobin concentration|HGB
Event|Event|SIMPLE_SEGMENT|522,525|false|false|false|||HCT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|522,525|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|522,525|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Disorder|Virus|SIMPLE_SEGMENT|531,534|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|531,534|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|531,534|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|531,534|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|531,534|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|539,542|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|539,542|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|539,542|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|539,542|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|539,542|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|539,542|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|SIMPLE_SEGMENT|548,552|false|false|false|||MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|548,552|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|592,595|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Enzyme|SIMPLE_SEGMENT|592,595|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Organic Chemical|SIMPLE_SEGMENT|592,595|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|592,595|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Event|Event|SIMPLE_SEGMENT|592,595|false|false|false|||ASA
Finding|Gene or Genome|SIMPLE_SEGMENT|592,595|false|false|false|C1412553|ARSA gene|ASA
Event|Event|SIMPLE_SEGMENT|596,599|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|596,599|false|false|false|C5848551|Neg - answer|NEG
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|600,607|false|false|false|C0161679|Toxic effect of ethyl alcohol|ETHANOL
Drug|Organic Chemical|SIMPLE_SEGMENT|600,607|false|false|false|C0001962;C3854029;C3854030|CNS depressants ethanol;antiseptics ethanol;ethanol|ETHANOL
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|600,607|false|false|false|C0001962;C3854029;C3854030|CNS depressants ethanol;antiseptics ethanol;ethanol|ETHANOL
Event|Event|SIMPLE_SEGMENT|600,607|false|false|false|||ETHANOL
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|600,607|false|false|false|C0202304|Ethanol measurement|ETHANOL
Event|Event|SIMPLE_SEGMENT|608,611|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|608,611|false|false|false|C5848551|Neg - answer|NEG
Event|Event|SIMPLE_SEGMENT|622,625|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|622,625|false|false|false|C5848551|Neg - answer|NEG
Event|Event|SIMPLE_SEGMENT|637,640|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|637,640|false|false|false|C5848551|Neg - answer|NEG
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|655,662|false|false|false|C0001924;C5966160|Albumin;Albumins|ALBUMIN
Drug|Biologically Active Substance|SIMPLE_SEGMENT|655,662|false|false|false|C0001924;C5966160|Albumin;Albumins|ALBUMIN
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|655,662|false|false|false|C0001924;C5966160|Albumin;Albumins|ALBUMIN
Event|Event|SIMPLE_SEGMENT|655,662|false|false|false|||ALBUMIN
Finding|Gene or Genome|SIMPLE_SEGMENT|655,662|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|ALBUMIN
Finding|Physiologic Function|SIMPLE_SEGMENT|655,662|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|ALBUMIN
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|655,662|false|false|false|C0201838|Albumin measurement|ALBUMIN
Drug|Biologically Active Substance|SIMPLE_SEGMENT|667,674|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|667,674|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Inorganic Chemical|SIMPLE_SEGMENT|667,674|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|667,674|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Vitamin|SIMPLE_SEGMENT|667,674|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Event|Event|SIMPLE_SEGMENT|667,674|false|false|false|||CALCIUM
Finding|Physiologic Function|SIMPLE_SEGMENT|667,674|false|false|false|C4553026|Calcium metabolic function|CALCIUM
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|667,674|false|false|false|C0201925|Calcium measurement|CALCIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|679,688|false|false|false|C0031603;C1601799|Phosphates;phosphate ion|PHOSPHATE
Drug|Inorganic Chemical|SIMPLE_SEGMENT|679,688|false|false|false|C0031603;C1601799|Phosphates;phosphate ion|PHOSPHATE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|679,688|false|false|false|C0031603;C1601799|Phosphates;phosphate ion|PHOSPHATE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|679,688|false|false|false|C0523826|Phosphate measurement|PHOSPHATE
Drug|Biologically Active Substance|SIMPLE_SEGMENT|694,703|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|694,703|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Drug|Inorganic Chemical|SIMPLE_SEGMENT|694,703|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|694,703|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|694,703|false|false|false|C0373675|Magnesium measurement|MAGNESIUM
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|722,728|false|false|false|C0023764|lipase|LIPASE
Drug|Enzyme|SIMPLE_SEGMENT|722,728|false|false|false|C0023764|lipase|LIPASE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|722,728|false|false|false|C0023764|lipase|LIPASE
Event|Event|SIMPLE_SEGMENT|722,728|false|false|false|||LIPASE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|722,728|false|false|false|C0373670|Lipase measurement|LIPASE
Disorder|Neoplastic Process|SIMPLE_SEGMENT|746,749|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|746,749|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|SIMPLE_SEGMENT|746,749|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|SIMPLE_SEGMENT|746,749|false|false|false|||ALT
Finding|Gene or Genome|SIMPLE_SEGMENT|746,749|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|SIMPLE_SEGMENT|746,749|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|SIMPLE_SEGMENT|746,749|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|746,749|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|750,754|false|false|false|C0376147|SGPT - Glutamate pyruvate transaminase|SGPT
Drug|Enzyme|SIMPLE_SEGMENT|750,754|false|false|false|C0376147|SGPT - Glutamate pyruvate transaminase|SGPT
Event|Event|SIMPLE_SEGMENT|750,754|false|false|false|||SGPT
Finding|Gene or Genome|SIMPLE_SEGMENT|750,754|false|false|false|C1415274|GPT gene|SGPT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|750,754|false|false|false|C0036828|Serum Alanine Transaminase Test|SGPT
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|759,762|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|SIMPLE_SEGMENT|759,762|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|759,762|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|SIMPLE_SEGMENT|759,762|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|SIMPLE_SEGMENT|759,762|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|SIMPLE_SEGMENT|759,762|false|false|false|||AST
Finding|Gene or Genome|SIMPLE_SEGMENT|759,762|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|763,767|false|false|false|C0242192|SGOT - Glutamate oxaloacetate transaminase|SGOT
Drug|Enzyme|SIMPLE_SEGMENT|763,767|false|false|false|C0242192|SGOT - Glutamate oxaloacetate transaminase|SGOT
Event|Event|SIMPLE_SEGMENT|763,767|false|false|false|||SGOT
Finding|Gene or Genome|SIMPLE_SEGMENT|763,767|false|false|false|C1415181|GOT1 gene|SGOT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|763,767|false|false|false|C0201899|Aspartate aminotransferase measurement|SGOT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|772,775|false|false|false|C1663627|ALK protein, human|ALK
Drug|Enzyme|SIMPLE_SEGMENT|772,775|false|false|false|C1663627|ALK protein, human|ALK
Event|Event|SIMPLE_SEGMENT|772,775|false|false|false|||ALK
Finding|Gene or Genome|SIMPLE_SEGMENT|772,775|false|false|false|C1332080;C1663627;C1704943|ALK gene;ALK protein, human;ALK wt Allele|ALK
Finding|Receptor|SIMPLE_SEGMENT|772,775|false|false|false|C1332080;C1663627;C1704943|ALK gene;ALK protein, human;ALK wt Allele|ALK
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|772,780|false|false|false|C0002059|Alkaline Phosphatase|ALK PHOS
Drug|Enzyme|SIMPLE_SEGMENT|772,780|false|false|false|C0002059|Alkaline Phosphatase|ALK PHOS
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|772,780|false|false|false|C0201850|Alkaline phosphatase measurement|ALK PHOS
Event|Event|SIMPLE_SEGMENT|776,780|false|false|false|||PHOS
Event|Event|SIMPLE_SEGMENT|784,787|false|false|false|||TOT
Drug|Biologically Active Substance|SIMPLE_SEGMENT|812,819|false|false|false|C0017725|glucose|GLUCOSE
Drug|Organic Chemical|SIMPLE_SEGMENT|812,819|false|false|false|C0017725|glucose|GLUCOSE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|812,819|false|false|false|C0017725|glucose|GLUCOSE
Event|Event|SIMPLE_SEGMENT|812,819|false|false|false|||GLUCOSE
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|812,819|false|false|false|C5781949|Glucose^1.5H post dose glucagon|GLUCOSE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|812,819|false|false|false|C0337438|Glucose measurement|GLUCOSE
Drug|Biologically Active Substance|SIMPLE_SEGMENT|825,829|false|false|false|C0041942|urea|UREA
Drug|Organic Chemical|SIMPLE_SEGMENT|825,829|false|false|false|C0041942|urea|UREA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|825,829|false|false|false|C0041942|urea|UREA
Event|Event|SIMPLE_SEGMENT|825,829|false|false|false|||UREA
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|825,829|false|false|false|C0523961|Urea measurement|UREA
Drug|Biologically Active Substance|SIMPLE_SEGMENT|845,851|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|845,851|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|845,851|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Event|Event|SIMPLE_SEGMENT|845,851|false|false|false|||SODIUM
Finding|Physiologic Function|SIMPLE_SEGMENT|845,851|false|false|false|C4553025|Sodium metabolic function|SODIUM
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|845,851|false|false|false|C0337443|Sodium measurement|SODIUM
Drug|Biologically Active Substance|SIMPLE_SEGMENT|857,866|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|857,866|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Food|SIMPLE_SEGMENT|857,866|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Inorganic Chemical|SIMPLE_SEGMENT|857,866|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|857,866|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Event|Event|SIMPLE_SEGMENT|857,866|false|false|false|||POTASSIUM
Finding|Physiologic Function|SIMPLE_SEGMENT|857,866|false|false|false|C4553027|Potassium metabolic function|POTASSIUM
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|857,866|false|false|false|C0202194|Potassium measurement|POTASSIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|871,879|false|false|false|C0008203;C0596019|Chlorides;chloride ion|CHLORIDE
Event|Event|SIMPLE_SEGMENT|871,879|false|false|false|||CHLORIDE
Finding|Physiologic Function|SIMPLE_SEGMENT|871,879|false|false|false|C4553021|Chloride metabolic function|CHLORIDE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|871,879|false|false|false|C0201952|Chloride measurement|CHLORIDE
Drug|Biologically Active Substance|SIMPLE_SEGMENT|890,893|false|false|false|C0007012|carbon dioxide|CO2
Drug|Inorganic Chemical|SIMPLE_SEGMENT|890,893|false|false|false|C0007012|carbon dioxide|CO2
Event|Event|SIMPLE_SEGMENT|890,893|false|false|false|||CO2
Finding|Finding|SIMPLE_SEGMENT|890,893|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Finding|Gene or Genome|SIMPLE_SEGMENT|890,893|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|897,902|false|false|false|C0003075|Anions|ANION
Attribute|Clinical Attribute|SIMPLE_SEGMENT|897,906|false|false|false|C0003074|Anion Gap|ANION GAP
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|897,906|false|false|false|C1509129|Anion gap result|ANION GAP
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|897,906|false|false|false|C0201889;C2189246|Anion gap measurement;blood anion gap (lab test)|ANION GAP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|903,906|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Drug|Biologically Active Substance|SIMPLE_SEGMENT|903,906|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Event|Event|SIMPLE_SEGMENT|903,906|false|false|false|||GAP
Finding|Gene or Genome|SIMPLE_SEGMENT|903,906|false|false|false|C1419277;C2984552|RASA1 gene;RASA1 wt Allele|GAP
Finding|Body Substance|SIMPLE_SEGMENT|922,927|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|922,927|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|922,927|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|922,934|false|false|false|C0018965|Hematuria|URINE  BLOOD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|929,934|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|929,934|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|929,934|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Event|Event|SIMPLE_SEGMENT|935,938|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|935,938|false|false|false|C5848551|Neg - answer|NEG
Drug|Biologically Active Substance|SIMPLE_SEGMENT|939,946|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|NITRITE
Drug|Inorganic Chemical|SIMPLE_SEGMENT|939,946|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|NITRITE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|939,946|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|NITRITE
Finding|Finding|SIMPLE_SEGMENT|947,950|false|false|false|C5848551|Neg - answer|NEG
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|951,958|false|false|false|C0033684|Proteins|PROTEIN
Drug|Biologically Active Substance|SIMPLE_SEGMENT|951,958|false|false|false|C0033684|Proteins|PROTEIN
Event|Event|SIMPLE_SEGMENT|951,958|false|false|false|||PROTEIN
Finding|Conceptual Entity|SIMPLE_SEGMENT|951,958|false|false|false|C1521746|Protein Info|PROTEIN
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|951,958|false|false|false|C0202202|Protein measurement|PROTEIN
Event|Event|SIMPLE_SEGMENT|959,962|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|959,962|false|false|false|C5848551|Neg - answer|NEG
Drug|Biologically Active Substance|SIMPLE_SEGMENT|964,971|false|false|false|C0017725|glucose|GLUCOSE
Drug|Organic Chemical|SIMPLE_SEGMENT|964,971|false|false|false|C0017725|glucose|GLUCOSE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|964,971|false|false|false|C0017725|glucose|GLUCOSE
Event|Event|SIMPLE_SEGMENT|964,971|false|false|false|||GLUCOSE
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|964,971|false|false|false|C5781949|Glucose^1.5H post dose glucagon|GLUCOSE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|964,971|false|false|false|C0337438|Glucose measurement|GLUCOSE
Event|Event|SIMPLE_SEGMENT|972,975|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|972,975|false|false|false|C5848551|Neg - answer|NEG
Drug|Organic Chemical|SIMPLE_SEGMENT|976,982|false|false|false|C0022634|Ketones|KETONE
Drug|Biologically Active Substance|SIMPLE_SEGMENT|987,996|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|BILIRUBIN
Drug|Organic Chemical|SIMPLE_SEGMENT|987,996|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|BILIRUBIN
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|987,996|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|BILIRUBIN
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|987,996|false|false|false|C0201913;C0863174|Bilirubin, total measurement;blood bilirubin level test|BILIRUBIN
Event|Event|SIMPLE_SEGMENT|997,1000|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|997,1000|false|false|false|C5848551|Neg - answer|NEG
Event|Event|SIMPLE_SEGMENT|1031,1034|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|1031,1034|false|false|false|C5848551|Neg - answer|NEG
Finding|Body Substance|SIMPLE_SEGMENT|1047,1052|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|1047,1052|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|1047,1052|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Finding|SIMPLE_SEGMENT|1047,1059|false|false|false|C0278030|Color of urine|URINE  COLOR
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|1054,1059|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|COLOR
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|1054,1059|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|COLOR
Event|Event|SIMPLE_SEGMENT|1054,1059|false|false|false|||COLOR
Drug|Organic Chemical|SIMPLE_SEGMENT|1060,1065|false|false|false|C4047917|Cereal plant straw|Straw
Event|Event|SIMPLE_SEGMENT|1066,1072|false|false|false|||APPEAR
Finding|Idea or Concept|SIMPLE_SEGMENT|1073,1078|false|false|false|C1550016|Remote control command - Clear|CLEAR
Finding|Body Substance|SIMPLE_SEGMENT|1098,1103|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|1098,1103|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|1098,1103|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Finding|SIMPLE_SEGMENT|1114,1117|false|false|false|C5848551|Neg - answer|NEG
Finding|Finding|SIMPLE_SEGMENT|1127,1130|false|false|false|C5848551|Neg - answer|NEG
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|1131,1138|false|false|false|C0221793;C0376196|Opiate Alkaloids;Opiates|opiates
Drug|Organic Chemical|SIMPLE_SEGMENT|1131,1138|false|false|false|C0221793;C0376196|Opiate Alkaloids;Opiates|opiates
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1131,1138|false|false|false|C0221793;C0376196|Opiate Alkaloids;Opiates|opiates
Event|Event|SIMPLE_SEGMENT|1131,1138|false|false|false|||opiates
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1131,1138|false|false|false|C0242401|Opiate Measurement|opiates
Event|Event|SIMPLE_SEGMENT|1139,1142|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|1139,1142|false|false|false|C5848551|Neg - answer|NEG
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|1144,1151|false|false|false|C0274659|Poisoning by cocaine|cocaine
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|1144,1151|false|false|false|C0009170|cocaine|cocaine
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|1144,1151|false|false|false|C0009170|cocaine|cocaine
Drug|Organic Chemical|SIMPLE_SEGMENT|1144,1151|false|false|false|C0009170|cocaine|cocaine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1144,1151|false|false|false|C0009170|cocaine|cocaine
Event|Event|SIMPLE_SEGMENT|1144,1151|false|false|false|||cocaine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1144,1151|false|false|false|C0202362|Cocaine measurement|cocaine
Event|Event|SIMPLE_SEGMENT|1152,1155|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|1152,1155|false|false|false|C5848551|Neg - answer|NEG
Finding|Finding|SIMPLE_SEGMENT|1165,1168|false|false|false|C5848551|Neg - answer|NEG
Finding|Finding|SIMPLE_SEGMENT|1177,1180|false|false|false|C5848551|Neg - answer|NEG
Event|Event|SIMPLE_SEGMENT|1189,1192|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|1189,1192|false|false|false|C5848551|Neg - answer|NEG
Finding|Body Substance|SIMPLE_SEGMENT|1205,1210|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|1205,1210|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|1205,1210|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Event|Event|SIMPLE_SEGMENT|1212,1215|false|false|false|||UCG
Event|Event|SIMPLE_SEGMENT|1216,1224|false|false|false|||NEGATIVE
Finding|Classification|SIMPLE_SEGMENT|1216,1224|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|NEGATIVE
Finding|Finding|SIMPLE_SEGMENT|1216,1224|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|NEGATIVE
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1216,1224|false|false|false|C5237010|Expression Negative|NEGATIVE
Finding|Body Substance|SIMPLE_SEGMENT|1237,1242|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|1237,1242|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|1237,1242|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Event|Event|SIMPLE_SEGMENT|1250,1256|false|false|false|||RANDOM
Event|Event|SIMPLE_SEGMENT|1268,1272|false|false|false|||LABS
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1268,1272|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1302,1307|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|1302,1307|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|1302,1307|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1332,1337|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|1332,1337|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|1332,1337|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1338,1341|false|false|false|C2708739||TSH
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1338,1341|false|false|false|C0040160|thyrotropin|TSH
Drug|Hormone|SIMPLE_SEGMENT|1338,1341|false|false|false|C0040160|thyrotropin|TSH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1338,1341|false|false|false|C0040160|thyrotropin|TSH
Event|Event|SIMPLE_SEGMENT|1338,1341|false|false|false|||TSH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1338,1341|false|false|false|C0202230|Thyroid stimulating hormone measurement|TSH
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1359,1364|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|1359,1364|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|1359,1364|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Finding|Functional Concept|SIMPLE_SEGMENT|1365,1369|false|false|false|C0332296|Free of (attribute)|Free
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1365,1372|false|false|false|C0202225|T4 free measurement|Free T4
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1389,1394|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|1389,1394|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|1389,1394|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|1395,1402|false|false|false|C0042890|Vitamins|VITAMIN
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1395,1402|false|false|false|C0042890|Vitamins|VITAMIN
Drug|Vitamin|SIMPLE_SEGMENT|1395,1402|false|false|false|C0042890|Vitamins|VITAMIN
Drug|Organic Chemical|SIMPLE_SEGMENT|1395,1405|false|false|false|C0039840|thiamine|VITAMIN B1
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1395,1405|false|false|false|C0039840|thiamine|VITAMIN B1
Drug|Vitamin|SIMPLE_SEGMENT|1395,1405|false|false|false|C0039840|thiamine|VITAMIN B1
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1395,1405|false|false|false|C0373727|Thiamine measurement|VITAMIN B1
Finding|Body Substance|SIMPLE_SEGMENT|1406,1417|false|false|false|C0370231;C1546552;C1608383|whole blood;whole blood specimen|WHOLE BLOOD
Finding|Intellectual Product|SIMPLE_SEGMENT|1406,1417|false|false|false|C0370231;C1546552;C1608383|whole blood;whole blood specimen|WHOLE BLOOD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1412,1417|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|1412,1417|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|1412,1417|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1418,1421|false|false|false|C1956415|Paroxysmal nocturnal dyspnea|PND
Event|Event|SIMPLE_SEGMENT|1418,1421|false|false|false|||PND
Finding|Gene or Genome|SIMPLE_SEGMENT|1418,1421|false|false|false|C1417807;C4552608|NPPA gene;NPPA wt Allele|PND
Event|Event|SIMPLE_SEGMENT|1423,1428|false|false|false|||MICRO
Finding|Conceptual Entity|SIMPLE_SEGMENT|1423,1428|false|false|false|C3811161;C4049106|Micro (prefix);Microbiology - Laboratory Class|MICRO
Finding|Intellectual Product|SIMPLE_SEGMENT|1423,1428|false|false|false|C3811161;C4049106|Micro (prefix);Microbiology - Laboratory Class|MICRO
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1423,1428|false|false|false|C0085672|Microbiology procedure|MICRO
Finding|Body Substance|SIMPLE_SEGMENT|1449,1454|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|1449,1454|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|1449,1454|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Idea or Concept|SIMPLE_SEGMENT|1486,1491|false|false|false|C1546485|Diagnosis Type - Final|FINAL
Finding|Intellectual Product|SIMPLE_SEGMENT|1486,1498|false|false|false|C0460114|Final report|FINAL REPORT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1492,1498|false|false|false|C4255046||REPORT
Event|Event|SIMPLE_SEGMENT|1492,1498|false|false|false|||REPORT
Finding|Intellectual Product|SIMPLE_SEGMENT|1492,1498|false|false|false|C0684224|Report (document)|REPORT
Procedure|Health Care Activity|SIMPLE_SEGMENT|1492,1498|false|false|false|C0700287|Reporting|REPORT
Finding|Body Substance|SIMPLE_SEGMENT|1507,1512|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|1507,1512|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|1507,1512|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1507,1520|false|false|false|C0430404|Urine culture|URINE CULTURE
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|1513,1520|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|SIMPLE_SEGMENT|1513,1520|false|false|false|||CULTURE
Finding|Functional Concept|SIMPLE_SEGMENT|1513,1520|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|SIMPLE_SEGMENT|1513,1520|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1513,1520|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Event|Event|SIMPLE_SEGMENT|1522,1527|false|false|false|||Final
Finding|Idea or Concept|SIMPLE_SEGMENT|1522,1527|false|false|false|C1546485|Diagnosis Type - Final|Final
Event|Event|SIMPLE_SEGMENT|1540,1545|false|false|false|||MIXED
Anatomy|Cell|SIMPLE_SEGMENT|1569,1575|false|false|false|C1947989|Colony (cells or organisms)|COLONY
Event|Event|SIMPLE_SEGMENT|1584,1594|false|false|false|||CONSISTENT
Finding|Idea or Concept|SIMPLE_SEGMENT|1584,1594|false|false|false|C0332290|Consistent with|CONSISTENT
Anatomy|Body System|SIMPLE_SEGMENT|1601,1605|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1601,1605|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1601,1605|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Event|Event|SIMPLE_SEGMENT|1601,1605|false|false|false|||SKIN
Finding|Body Substance|SIMPLE_SEGMENT|1601,1605|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|SIMPLE_SEGMENT|1601,1605|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Event|Event|SIMPLE_SEGMENT|1615,1616|false|false|false|||/
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1619,1626|false|false|false|C0017420;C0559522|Genital system;Genitalia|GENITAL
Anatomy|Body System|SIMPLE_SEGMENT|1619,1626|false|false|false|C0017420;C0559522|Genital system;Genitalia|GENITAL
Finding|Body Substance|SIMPLE_SEGMENT|1619,1626|false|false|false|C1546649;C1550642|Specimen Type - Genital|GENITAL
Finding|Intellectual Product|SIMPLE_SEGMENT|1619,1626|false|false|false|C1546649;C1550642|Specimen Type - Genital|GENITAL
Event|Event|SIMPLE_SEGMENT|1627,1640|false|false|false|||CONTAMINATION
Finding|Idea or Concept|SIMPLE_SEGMENT|1627,1640|false|false|false|C2349974|Contamination|CONTAMINATION
Phenomenon|Human-caused Phenomenon or Process|SIMPLE_SEGMENT|1627,1640|false|false|false|C0259846|adulteration|CONTAMINATION
Event|Event|SIMPLE_SEGMENT|1644,1651|false|false|false|||IMAGING
Finding|Finding|SIMPLE_SEGMENT|1644,1651|false|false|false|C0740845|Imaging problem|IMAGING
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1644,1651|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|IMAGING
Finding|Body Substance|SIMPLE_SEGMENT|1668,1677|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|1668,1677|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|1668,1677|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|1668,1677|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|SIMPLE_SEGMENT|1678,1682|false|false|false|||LABS
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1678,1682|false|false|false|C0587081|Laboratory test finding|LABS
Event|Event|SIMPLE_SEGMENT|1703,1707|false|false|false|||labs
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1703,1707|true|false|false|C0587081|Laboratory test finding|labs
Finding|Idea or Concept|SIMPLE_SEGMENT|1711,1714|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|1711,1714|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|1718,1727|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|1718,1727|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|1718,1727|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|1718,1727|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|1718,1727|false|false|false|C0030685|Patient Discharge|discharge
Finding|Body Substance|SIMPLE_SEGMENT|1729,1738|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|1729,1738|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|1729,1738|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|1729,1738|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|SIMPLE_SEGMENT|1739,1747|false|false|false|||PHYSICAL
Finding|Finding|SIMPLE_SEGMENT|1739,1747|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|SIMPLE_SEGMENT|1739,1747|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|1739,1747|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|SIMPLE_SEGMENT|1739,1752|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAM
Procedure|Health Care Activity|SIMPLE_SEGMENT|1739,1752|false|false|false|C0031809|Physical Examination|PHYSICAL EXAM
Event|Event|SIMPLE_SEGMENT|1748,1752|false|false|false|||EXAM
Finding|Functional Concept|SIMPLE_SEGMENT|1748,1752|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|SIMPLE_SEGMENT|1748,1752|false|false|false|C0582103|Medical Examination|EXAM
Event|Event|SIMPLE_SEGMENT|1779,1785|false|false|false|||VITALS
Event|Event|SIMPLE_SEGMENT|1796,1800|false|false|false|||Temp
Finding|Gene or Genome|SIMPLE_SEGMENT|1796,1800|false|false|false|C1823816|C1orf210 gene|Temp
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1796,1800|false|false|false|C0279848|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Temp
Event|Event|SIMPLE_SEGMENT|1829,1831|false|false|false|||HR
Event|Event|SIMPLE_SEGMENT|1860,1868|false|false|false|||delivery
Finding|Finding|SIMPLE_SEGMENT|1860,1868|false|false|false|C1314680;C1705822;C2053584|Transfer Technique;delivery (history)|delivery
Finding|Functional Concept|SIMPLE_SEGMENT|1860,1868|false|false|false|C1314680;C1705822;C2053584|Transfer Technique;delivery (history)|delivery
Finding|Organism Function|SIMPLE_SEGMENT|1860,1868|false|false|false|C1314680;C1705822;C2053584|Transfer Technique;delivery (history)|delivery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1860,1868|false|false|false|C0011209|Obstetric Delivery|delivery
Event|Event|SIMPLE_SEGMENT|1875,1882|false|false|false|||GENERAL
Finding|Classification|SIMPLE_SEGMENT|1875,1882|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|1875,1882|false|false|false|C3812897|General medical service|GENERAL
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1885,1888|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1885,1888|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1885,1888|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|1885,1888|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1885,1888|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|SIMPLE_SEGMENT|1885,1888|false|false|false|||NAD
Finding|Finding|SIMPLE_SEGMENT|1885,1888|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Event|Event|SIMPLE_SEGMENT|1890,1897|false|false|false|||sitting
Event|Event|SIMPLE_SEGMENT|1911,1918|false|false|false|||smiling
Finding|Social Behavior|SIMPLE_SEGMENT|1911,1918|false|false|false|C0037363|Smiling|smiling
Event|Event|SIMPLE_SEGMENT|1920,1926|false|false|false|||moving
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1927,1931|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1927,1931|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1927,1931|false|false|false|C0362076|Problems with head|head
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1927,1931|false|false|false|C0876917|Procedure on head|head
Event|Event|SIMPLE_SEGMENT|1932,1938|false|false|false|||around
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1939,1943|false|false|false|C0015392|Eye|EYES
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1939,1943|false|false|false|C5848506||EYES
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1945,1951|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1945,1951|false|false|false|C0036412|Scleral Diseases|Sclera
Event|Event|SIMPLE_SEGMENT|1945,1951|false|false|false|||Sclera
Procedure|Health Care Activity|SIMPLE_SEGMENT|1945,1951|false|false|false|C2228481|examination of sclera|Sclera
Event|Event|SIMPLE_SEGMENT|1952,1961|false|false|false|||anicteric
Finding|Finding|SIMPLE_SEGMENT|1952,1961|false|false|false|C0205180|Anicteric|anicteric
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|1974,1983|true|false|false|C1272883|Injection|injection
Event|Event|SIMPLE_SEGMENT|1974,1983|false|false|false|||injection
Finding|Functional Concept|SIMPLE_SEGMENT|1974,1983|true|false|false|C1828121|Injection Route of Administration|injection
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1974,1983|true|false|false|C0021485;C1533685|Injection of therapeutic agent;Injection procedure|injection
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1986,1993|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|SIMPLE_SEGMENT|1986,1993|false|false|false|C1314974|Cardiac attachment|CARDIAC
Event|Event|SIMPLE_SEGMENT|1995,1998|false|false|false|||RRR
Event|Event|SIMPLE_SEGMENT|2022,2029|false|false|false|||murmurs
Finding|Finding|SIMPLE_SEGMENT|2022,2029|true|false|false|C0018808|Heart murmur|murmurs
Finding|Finding|SIMPLE_SEGMENT|2030,2034|true|false|false|C0232267|Pericardial friction rub|rubs
Event|Event|SIMPLE_SEGMENT|2035,2042|false|false|false|||gallops
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2044,2048|false|false|false|C0231832|Respiratory rate|RESP
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2044,2048|false|false|false|C0851355|Respiratory, thoracic and mediastinal disorders|RESP
Event|Event|SIMPLE_SEGMENT|2044,2048|false|false|false|||RESP
Event|Event|SIMPLE_SEGMENT|2050,2055|false|false|false|||Clear
Finding|Idea or Concept|SIMPLE_SEGMENT|2050,2055|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|SIMPLE_SEGMENT|2059,2071|false|false|false|||auscultation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2059,2071|false|false|false|C0004339|Auscultation|auscultation
Event|Event|SIMPLE_SEGMENT|2088,2095|false|false|false|||wheezes
Finding|Sign or Symptom|SIMPLE_SEGMENT|2088,2095|true|false|false|C0043144|Wheezing|wheezes
Event|Event|SIMPLE_SEGMENT|2097,2104|false|false|false|||rhonchi
Finding|Finding|SIMPLE_SEGMENT|2097,2104|true|false|false|C0035508|Rhonchi|rhonchi
Event|Event|SIMPLE_SEGMENT|2108,2113|false|false|false|||rales
Finding|Finding|SIMPLE_SEGMENT|2108,2113|false|false|false|C0034642;C0240859|Basilar Rales;Rales|rales
Event|Event|SIMPLE_SEGMENT|2118,2127|false|false|false|||increased
Finding|Finding|SIMPLE_SEGMENT|2118,2127|true|false|false|C0442805;C5236002|Increase;Increased (finding)|increased
Finding|Functional Concept|SIMPLE_SEGMENT|2118,2127|true|false|false|C0442805;C5236002|Increase;Increased (finding)|increased
Finding|Sign or Symptom|SIMPLE_SEGMENT|2118,2145|true|false|false|C0859927|Increased work of breathing|increased work of breathing
Event|Event|SIMPLE_SEGMENT|2128,2132|false|false|false|||work
Event|Occupational Activity|SIMPLE_SEGMENT|2128,2132|true|false|false|C0043227|Work|work
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|2128,2145|true|false|false|C0043229|Work of Breathing|work of breathing
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2136,2145|false|false|false|C5885990||breathing
Event|Event|SIMPLE_SEGMENT|2136,2145|false|false|false|||breathing
Finding|Finding|SIMPLE_SEGMENT|2136,2145|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|SIMPLE_SEGMENT|2136,2145|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|SIMPLE_SEGMENT|2136,2145|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|SIMPLE_SEGMENT|2136,2145|false|false|false|C1160636|respiratory system process|breathing
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2147,2154|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2147,2154|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Event|Event|SIMPLE_SEGMENT|2147,2154|false|false|false|||ABDOMEN
Finding|Finding|SIMPLE_SEGMENT|2147,2154|false|false|false|C0941288|Abdomen problem|ABDOMEN
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2163,2169|false|false|false|C0021853|Intestines|bowels
Event|Event|SIMPLE_SEGMENT|2170,2176|false|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|2170,2176|false|false|false|C0037709||sounds
Event|Event|SIMPLE_SEGMENT|2182,2191|false|false|false|||distended
Finding|Finding|SIMPLE_SEGMENT|2182,2191|false|false|false|C0700124|Dilated|distended
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2205,2216|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Drug|Food|SIMPLE_SEGMENT|2218,2224|false|false|false|C5890763||Pulses
Event|Event|SIMPLE_SEGMENT|2218,2224|false|false|false|||Pulses
Finding|Physiologic Function|SIMPLE_SEGMENT|2218,2224|false|false|false|C0391850|Physiologic pulse|Pulses
Procedure|Health Care Activity|SIMPLE_SEGMENT|2218,2224|false|false|false|C0034107|Pulse taking|Pulses
Event|Event|SIMPLE_SEGMENT|2225,2227|false|false|false|||DP
Finding|Conceptual Entity|SIMPLE_SEGMENT|2228,2234|false|false|false|C0442038;C0920847|Circumpennate;Radial|Radial
Anatomy|Body System|SIMPLE_SEGMENT|2251,2255|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2251,2255|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2251,2255|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Event|Event|SIMPLE_SEGMENT|2251,2255|false|false|false|||SKIN
Finding|Body Substance|SIMPLE_SEGMENT|2251,2255|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|SIMPLE_SEGMENT|2251,2255|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Event|Event|SIMPLE_SEGMENT|2257,2261|false|false|false|||Warm
Finding|Finding|SIMPLE_SEGMENT|2257,2261|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|2257,2261|false|false|false|C0687712|warming process|Warm
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|2263,2266|false|false|false|C1855179|CATARACT, ANTERIOR POLAR|Cap
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|2263,2266|false|false|false|C0006935|capsule (pharmacologic)|Cap
Event|Event|SIMPLE_SEGMENT|2263,2266|false|false|false|||Cap
Finding|Gene or Genome|SIMPLE_SEGMENT|2263,2266|false|false|false|C1416891;C1418551;C1419093;C1422073;C1422760;C2985259;C4522312|BRD4 gene;BRD4 wt Allele;CAP1 gene;HACD1 gene;LNPEP gene;SERPINB6 gene;SORBS1 gene|Cap
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2263,2266|false|false|false|C0278651;C0280547;C1879916|CAP Regimen;cisplatin/cyclophosphamide/doxorubicin protocol;cyclophosphamide/doxorubicin/prednisone protocol|Cap
Event|Event|SIMPLE_SEGMENT|2267,2273|false|false|false|||refill
Finding|Idea or Concept|SIMPLE_SEGMENT|2267,2273|false|false|false|C0807726|refill|refill
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2282,2286|true|false|false|C5779629|Eruption of skin (disorder)|rash
Event|Event|SIMPLE_SEGMENT|2282,2286|false|false|false|||rash
Finding|Pathologic Function|SIMPLE_SEGMENT|2282,2286|true|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Sign or Symptom|SIMPLE_SEGMENT|2282,2286|true|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Event|Event|SIMPLE_SEGMENT|2288,2298|false|false|false|||NEUROLOGIC
Event|Event|SIMPLE_SEGMENT|2300,2306|false|false|false|||Speech
Finding|Organism Function|SIMPLE_SEGMENT|2300,2306|false|false|false|C0037817|Speech|Speech
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2300,2306|false|false|false|C0846595|Speech assessment|Speech
Event|Event|SIMPLE_SEGMENT|2325,2333|false|false|false|||improved
Finding|Finding|SIMPLE_SEGMENT|2325,2333|false|false|false|C0184511;C1561611;C4084203|Admission Level of Care Code - Improved;Improved;Improved - answer to question|improved
Finding|Intellectual Product|SIMPLE_SEGMENT|2325,2333|false|false|false|C0184511;C1561611;C4084203|Admission Level of Care Code - Improved;Improved;Improved - answer to question|improved
Event|Event|SIMPLE_SEGMENT|2344,2350|false|false|false|||speaks
Finding|Finding|SIMPLE_SEGMENT|2344,2350|false|false|true|C0600116|Does speak|speaks
Finding|Gene or Genome|SIMPLE_SEGMENT|2355,2361|false|false|false|C1424587|LITAF gene|simple
Event|Event|SIMPLE_SEGMENT|2362,2371|false|false|false|||sentences
Finding|Intellectual Product|SIMPLE_SEGMENT|2362,2371|false|false|false|C0876929|Sentence|sentences
Event|Event|SIMPLE_SEGMENT|2373,2380|false|false|false|||Sitting
Finding|Finding|SIMPLE_SEGMENT|2373,2380|false|false|false|C0277814;C2584297|Sitting Function;Sitting position|Sitting
Finding|Physiologic Function|SIMPLE_SEGMENT|2373,2380|false|false|false|C0277814;C2584297|Sitting Function;Sitting position|Sitting
Event|Event|SIMPLE_SEGMENT|2396,2400|false|false|false|||able
Finding|Finding|SIMPLE_SEGMENT|2396,2400|false|false|false|C1299581|Able (qualifier value)|able
Event|Event|SIMPLE_SEGMENT|2404,2408|false|false|false|||move
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2409,2424|false|false|false|C0278454|All extremities|all extremities
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2413,2424|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2458,2465|false|false|false|C0016129|Fingers|fingers
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2466,2470|false|false|false|C0040357;C4299090|Lower extremity>Toes;Toes|toes
Event|Event|SIMPLE_SEGMENT|2487,2495|false|false|false|||sticking
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2496,2501|false|false|false|C0040067|Thumb structure|thumb
Event|Event|SIMPLE_SEGMENT|2502,2504|false|false|false|||up
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|2506,2511|false|false|false|C0004936;C1306597|Mental disorders;Psychiatric problem|PSYCH
Event|Event|SIMPLE_SEGMENT|2506,2511|false|false|false|||PSYCH
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2513,2518|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|2513,2518|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2513,2518|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|SIMPLE_SEGMENT|2513,2518|false|false|false|||Alert
Finding|Finding|SIMPLE_SEGMENT|2513,2518|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|2513,2518|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|2513,2518|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|SIMPLE_SEGMENT|2523,2528|false|false|false|||awake
Finding|Finding|SIMPLE_SEGMENT|2523,2528|false|false|false|C0234422|Awake (finding)|awake
Event|Event|SIMPLE_SEGMENT|2530,2538|false|false|false|||pleasant
Finding|Mental Process|SIMPLE_SEGMENT|2530,2538|false|false|false|C2987187|Pleasant|pleasant
Event|Event|SIMPLE_SEGMENT|2540,2547|false|false|false|||smiling
Finding|Social Behavior|SIMPLE_SEGMENT|2540,2547|false|false|false|C0037363|Smiling|smiling
Finding|Intellectual Product|SIMPLE_SEGMENT|2552,2557|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|Brief
Finding|Idea or Concept|SIMPLE_SEGMENT|2558,2566|false|false|false|C1547192|Organization unit type - Hospital|Hospital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2558,2573|false|false|false|C0488549||Hospital Course
Finding|Finding|SIMPLE_SEGMENT|2558,2573|false|false|false|C0489547|Hospital course|Hospital Course
Finding|Intellectual Product|SIMPLE_SEGMENT|2575,2580|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|BRIEF
Finding|Idea or Concept|SIMPLE_SEGMENT|2581,2589|false|false|false|C1547192|Organization unit type - Hospital|HOSPITAL
Event|Event|SIMPLE_SEGMENT|2590,2597|false|false|false|||SUMMARY
Finding|Intellectual Product|SIMPLE_SEGMENT|2590,2597|false|false|false|C1552616;C1706244|Summary (document);summary - ActRelationshipSubset|SUMMARY
Event|Event|SIMPLE_SEGMENT|2639,2646|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|2639,2646|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|2639,2646|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|2639,2646|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|2639,2649|false|false|false|C0262926|Medical History|history of
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|2650,2667|false|false|false|C0855228|Eating disorder symptom|disordered eating
Event|Event|SIMPLE_SEGMENT|2661,2667|false|false|false|||eating
Finding|Organism Function|SIMPLE_SEGMENT|2661,2667|false|false|false|C0013470|Eating|eating
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2669,2673|false|false|false|C0038436;C0878676|6-pyruvoyl-tetrahydropterin synthase deficiency;Post-Traumatic Stress Disorder|PTSD
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|2669,2673|false|false|false|C0038436;C0878676|6-pyruvoyl-tetrahydropterin synthase deficiency;Post-Traumatic Stress Disorder|PTSD
Event|Event|SIMPLE_SEGMENT|2669,2673|false|false|false|||PTSD
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|2675,2678|false|false|false|C0270549|Generalized Anxiety Disorder|GAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2675,2678|false|false|false|C0017785|Glutamate Decarboxylase|GAD
Drug|Enzyme|SIMPLE_SEGMENT|2675,2678|false|false|false|C0017785|Glutamate Decarboxylase|GAD
Event|Event|SIMPLE_SEGMENT|2675,2678|false|false|false|||GAD
Finding|Gene or Genome|SIMPLE_SEGMENT|2675,2678|false|false|false|C1414925;C5575531|GAD1 gene;GAD1 wt Allele|GAD
Finding|Finding|SIMPLE_SEGMENT|2685,2690|false|false|false|C0030318|Panic|panic
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|2685,2699|false|false|false|C0030319|Panic Disorder|panic disorder
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2691,2699|false|false|false|C0012634|Disease|disorder
Event|Event|SIMPLE_SEGMENT|2691,2699|false|false|false|||disorder
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|2701,2711|false|false|false|C0011570;C0011581;C0344315;C0812393|Cancer patients and suicide and depression;Depressed mood;Depressive disorder;Mental Depression|depression
Event|Event|SIMPLE_SEGMENT|2701,2711|false|false|false|||depression
Finding|Functional Concept|SIMPLE_SEGMENT|2701,2711|false|false|false|C0460137;C1579931|Depression - motion|depression
Finding|Sign or Symptom|SIMPLE_SEGMENT|2701,2711|false|false|false|C0460137;C1579931|Depression - motion|depression
Finding|Conceptual Entity|SIMPLE_SEGMENT|2716,2726|false|false|false|C0205245;C0542341;C2700217|Function (attribute);Functional;Functional Relationship|functional
Finding|Functional Concept|SIMPLE_SEGMENT|2716,2726|false|false|false|C0205245;C0542341;C2700217|Function (attribute);Functional;Functional Relationship|functional
Event|Event|SIMPLE_SEGMENT|2727,2739|false|false|false|||neurological
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2741,2749|false|false|false|C0012634|Disease|disorder
Event|Event|SIMPLE_SEGMENT|2741,2749|false|false|false|||disorder
Event|Event|SIMPLE_SEGMENT|2750,2760|false|false|false|||presenting
Event|Event|SIMPLE_SEGMENT|2768,2775|false|false|false|||therapy
Finding|Finding|SIMPLE_SEGMENT|2768,2775|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|SIMPLE_SEGMENT|2768,2775|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2768,2775|false|false|false|C0087111|Therapeutic procedure|therapy
Event|Event|SIMPLE_SEGMENT|2776,2783|false|false|false|||session
Event|Event|SIMPLE_SEGMENT|2776,2783|false|false|false|C1883016|Activity Session|session
Finding|Conceptual Entity|SIMPLE_SEGMENT|2776,2783|false|false|false|C1883017|Session|session
Event|Event|SIMPLE_SEGMENT|2789,2797|false|false|false|||weakness
Finding|Sign or Symptom|SIMPLE_SEGMENT|2789,2797|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Finding|Finding|SIMPLE_SEGMENT|2800,2808|false|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Finding|Idea or Concept|SIMPLE_SEGMENT|2800,2808|false|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2800,2817|false|false|false|C0013384|Dyskinetic syndrome|abnormal movement
Finding|Finding|SIMPLE_SEGMENT|2800,2817|false|false|false|C0558189|Abnormal movement|abnormal movement
Event|Event|SIMPLE_SEGMENT|2809,2817|false|false|false|||movement
Finding|Organism Function|SIMPLE_SEGMENT|2809,2817|false|false|false|C0026649|Movement|movement
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|2823,2830|false|false|false|C0003537|Aphasia|aphasia
Event|Event|SIMPLE_SEGMENT|2823,2830|false|false|false|||aphasia
Event|Event|SIMPLE_SEGMENT|2849,2854|false|false|false|||acute
Finding|Intellectual Product|SIMPLE_SEGMENT|2849,2854|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Conceptual Entity|SIMPLE_SEGMENT|2856,2866|false|false|false|C0205245;C0542341;C2700217|Function (attribute);Functional;Functional Relationship|functional
Finding|Functional Concept|SIMPLE_SEGMENT|2856,2866|false|false|false|C0205245;C0542341;C2700217|Function (attribute);Functional;Functional Relationship|functional
Event|Event|SIMPLE_SEGMENT|2880,2887|false|false|false|||episode
Event|Event|SIMPLE_SEGMENT|2897,2906|false|false|false|||evaluated
Event|Event|SIMPLE_SEGMENT|2925,2935|false|false|false|||psychology
Finding|Functional Concept|SIMPLE_SEGMENT|2925,2935|false|false|false|C1524060|psychology qualifier|psychology
Event|Event|SIMPLE_SEGMENT|2940,2944|false|false|false|||felt
Event|Event|SIMPLE_SEGMENT|2954,2964|false|false|false|||consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|2954,2964|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|2954,2969|false|false|false|C0332290|Consistent with|consistent with
Event|Event|SIMPLE_SEGMENT|2970,2980|false|false|false|||functional
Finding|Conceptual Entity|SIMPLE_SEGMENT|2970,2980|false|false|false|C0205245;C0542341;C2700217|Function (attribute);Functional;Functional Relationship|functional
Finding|Functional Concept|SIMPLE_SEGMENT|2970,2980|false|false|false|C0205245;C0542341;C2700217|Function (attribute);Functional;Functional Relationship|functional
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2982,3003|false|false|false|C0027765|nervous system disorder|neurological disorder
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2995,3003|false|false|false|C0012634|Disease|disorder
Event|Event|SIMPLE_SEGMENT|2995,3003|false|false|false|||disorder
Event|Event|SIMPLE_SEGMENT|3005,3012|false|false|false|||similar
Event|Event|SIMPLE_SEGMENT|3026,3038|false|false|false|||presentation
Finding|Idea or Concept|SIMPLE_SEGMENT|3026,3038|false|false|false|C0449450|Presentation|presentation
Event|Event|SIMPLE_SEGMENT|3045,3050|false|false|false|||began
Event|Event|SIMPLE_SEGMENT|3051,3058|false|false|false|||working
Finding|Gene or Genome|SIMPLE_SEGMENT|3088,3093|false|false|false|C1424898|RXFP2 gene|great
Event|Event|SIMPLE_SEGMENT|3094,3105|false|false|false|||improvement
Finding|Conceptual Entity|SIMPLE_SEGMENT|3094,3105|false|false|false|C2986411|Improvement|improvement
Finding|Finding|SIMPLE_SEGMENT|3110,3114|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|3110,3114|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|3110,3114|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|SIMPLE_SEGMENT|3118,3127|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|3118,3127|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|3118,3127|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|3118,3127|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|3118,3127|false|false|false|C0030685|Patient Discharge|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|3131,3136|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|SIMPLE_SEGMENT|3137,3142|false|false|false|||rehab
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3137,3142|false|false|false|C0034991|Rehabilitation therapy|rehab
Finding|Idea or Concept|SIMPLE_SEGMENT|3146,3158|false|false|false|C1548597|Marketing basis - Transitional|TRANSITIONAL
Event|Event|SIMPLE_SEGMENT|3159,3165|false|false|false|||ISSUES
Event|Event|SIMPLE_SEGMENT|3192,3197|false|false|false|||rehab
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3192,3197|false|false|false|C0034991|Rehabilitation therapy|rehab
Event|Event|SIMPLE_SEGMENT|3209,3217|false|false|false|||continue
Event|Event|SIMPLE_SEGMENT|3218,3228|false|false|false|||aggressive
Finding|Individual Behavior|SIMPLE_SEGMENT|3218,3228|false|false|false|C0001807;C1547300;C1548760|Aggressive behavior;Precaution Code - Aggressive;Risk Codes - Aggressive|aggressive
Finding|Intellectual Product|SIMPLE_SEGMENT|3218,3228|false|false|false|C0001807;C1547300;C1548760|Aggressive behavior;Precaution Code - Aggressive;Risk Codes - Aggressive|aggressive
Event|Event|SIMPLE_SEGMENT|3252,3263|false|false|false|||improvement
Finding|Conceptual Entity|SIMPLE_SEGMENT|3252,3263|false|true|false|C2986411|Improvement|improvement
Finding|Conceptual Entity|SIMPLE_SEGMENT|3268,3278|false|false|false|C0205245;C0542341;C2700217|Function (attribute);Functional;Functional Relationship|functional
Finding|Functional Concept|SIMPLE_SEGMENT|3268,3278|false|false|false|C0205245;C0542341;C2700217|Function (attribute);Functional;Functional Relationship|functional
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3268,3285|false|false|false|C2707028||functional status
Finding|Finding|SIMPLE_SEGMENT|3268,3285|false|false|false|C0489534;C0598463|Functional Status;functional status (history)|functional status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3279,3285|false|false|false|C5889824||status
Event|Event|SIMPLE_SEGMENT|3279,3285|false|false|false|||status
Finding|Idea or Concept|SIMPLE_SEGMENT|3279,3285|false|false|false|C1546481|What subject filter - Status|status
Event|Event|SIMPLE_SEGMENT|3294,3303|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|3294,3303|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|3294,3303|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|3294,3303|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|3294,3303|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|SIMPLE_SEGMENT|3312,3318|false|false|false|||ensure
Finding|Body Substance|SIMPLE_SEGMENT|3319,3326|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|3319,3326|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|3319,3326|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|SIMPLE_SEGMENT|3319,3330|false|false|false|C0332310|Has patient|patient has
Event|Event|SIMPLE_SEGMENT|3331,3337|false|false|false|||follow
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3351,3354|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|3351,3354|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3351,3354|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3351,3354|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|SIMPLE_SEGMENT|3351,3354|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|3351,3354|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|SIMPLE_SEGMENT|3351,3354|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3351,3354|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|SIMPLE_SEGMENT|3351,3354|false|false|false|||PCP
Finding|Gene or Genome|SIMPLE_SEGMENT|3351,3354|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|SIMPLE_SEGMENT|3351,3354|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Event|SIMPLE_SEGMENT|3363,3372|false|false|false|||therapist
Finding|Body Substance|SIMPLE_SEGMENT|3378,3385|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|3378,3385|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|3378,3385|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3415,3421|false|false|false|C4255480||nausea
Event|Event|SIMPLE_SEGMENT|3415,3421|false|false|false|||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|3415,3421|false|false|false|C0027497|Nausea|nausea
Event|Event|SIMPLE_SEGMENT|3425,3433|false|false|false|||appetite
Finding|Organism Function|SIMPLE_SEGMENT|3425,3433|false|false|false|C0003618|Desire for food|appetite
Event|Event|SIMPLE_SEGMENT|3435,3443|false|false|false|||improved
Event|Event|SIMPLE_SEGMENT|3452,3460|false|false|false|||continue
Drug|Organic Chemical|SIMPLE_SEGMENT|3461,3467|false|false|false|C0206046|Zofran|Zofran
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3461,3467|false|false|false|C0206046|Zofran|Zofran
Event|Event|SIMPLE_SEGMENT|3468,3471|false|false|false|||TID
Finding|Gene or Genome|SIMPLE_SEGMENT|3472,3475|false|false|false|C1422467|CIAO3 gene|prn
Event|Event|SIMPLE_SEGMENT|3477,3480|false|false|false|||QTc
Event|Event|SIMPLE_SEGMENT|3492,3495|false|false|false|||EKG
Finding|Intellectual Product|SIMPLE_SEGMENT|3492,3495|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3492,3495|false|false|false|C1623258|Electrocardiography|EKG
Event|Event|SIMPLE_SEGMENT|3508,3518|false|false|false|||continuing
Drug|Organic Chemical|SIMPLE_SEGMENT|3519,3525|false|false|false|C0206046|Zofran|Zofran
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3519,3525|false|false|false|C0206046|Zofran|Zofran
Event|Event|SIMPLE_SEGMENT|3526,3529|false|false|false|||use
Finding|Functional Concept|SIMPLE_SEGMENT|3526,3529|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|SIMPLE_SEGMENT|3526,3529|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|SIMPLE_SEGMENT|3537,3541|false|false|false|C1561540|Transaction counts and value totals - week|week
Event|Event|SIMPLE_SEGMENT|3550,3557|false|false|false|||recheck
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3578,3588|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|3578,3588|false|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|3578,3588|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|SIMPLE_SEGMENT|3592,3601|false|false|false|||prolonged
Finding|Body Substance|SIMPLE_SEGMENT|3606,3613|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|3606,3613|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|3606,3613|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Functional Concept|SIMPLE_SEGMENT|3606,3617|false|false|false|C0332310|Has patient|Patient has
Event|Event|SIMPLE_SEGMENT|3620,3627|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|3620,3627|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|3620,3627|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|3620,3627|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|3620,3630|false|false|false|C0262926|Medical History|history of
Finding|Finding|SIMPLE_SEGMENT|3646,3664|false|false|false|C5687959|Restrained eating behavior|restrictive eating
Event|Event|SIMPLE_SEGMENT|3658,3664|false|false|false|||eating
Finding|Organism Function|SIMPLE_SEGMENT|3658,3664|false|false|false|C0013470|Eating|eating
Finding|Finding|SIMPLE_SEGMENT|3676,3680|false|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|3681,3687|false|false|false|||eating
Event|Event|SIMPLE_SEGMENT|3693,3706|false|false|false|||encouragement
Finding|Social Behavior|SIMPLE_SEGMENT|3693,3706|false|false|false|C0870494|encouragement|encouragement
Event|Event|SIMPLE_SEGMENT|3719,3723|false|false|false|||show
Event|Event|SIMPLE_SEGMENT|3729,3737|false|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|3729,3737|false|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|3729,3740|false|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Event|Event|SIMPLE_SEGMENT|3741,3747|false|false|false|||eating
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3748,3756|false|false|false|C0012634|Disease|disorder
Event|Event|SIMPLE_SEGMENT|3748,3756|false|false|false|||disorder
Event|Event|SIMPLE_SEGMENT|3763,3772|false|false|false|||inpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|3763,3772|false|false|false|C1548438;C1549404|Patient Class - Inpatient;Referral category - Inpatient|inpatient
Procedure|Health Care Activity|SIMPLE_SEGMENT|3763,3772|false|false|false|C1555324|inpatient encounter|inpatient
Event|Event|SIMPLE_SEGMENT|3781,3789|false|false|false|||continue
Event|Event|SIMPLE_SEGMENT|3810,3813|false|false|false|||TID
Event|Event|SIMPLE_SEGMENT|3819,3824|false|false|false|||meals
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|3819,3824|false|false|false|C1998602|Meal (occasion for eating)|meals
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3832,3835|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|3832,3835|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3832,3835|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3832,3835|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|SIMPLE_SEGMENT|3832,3835|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|3832,3835|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|SIMPLE_SEGMENT|3832,3835|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3832,3835|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|SIMPLE_SEGMENT|3832,3835|false|false|false|||PCP
Finding|Gene or Genome|SIMPLE_SEGMENT|3832,3835|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|SIMPLE_SEGMENT|3832,3835|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Body Substance|SIMPLE_SEGMENT|3863,3870|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|3863,3870|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|3863,3870|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|3874,3886|false|false|false|||psychiatrist
Event|Event|SIMPLE_SEGMENT|3899,3908|false|false|false|||titration
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3899,3908|false|false|false|C0162621|Titration Method|titration
Event|Event|SIMPLE_SEGMENT|3913,3924|false|false|false|||psychiatric
Finding|Finding|SIMPLE_SEGMENT|3913,3924|false|false|false|C0205487;C1548428|Psychiatric;Referral type - Psychiatric|psychiatric
Finding|Functional Concept|SIMPLE_SEGMENT|3913,3924|false|false|false|C0205487;C1548428|Psychiatric;Referral type - Psychiatric|psychiatric
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3913,3924|false|false|false|C3526598|Psychiatric service|psychiatric
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3925,3936|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3925,3936|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|3925,3936|false|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|3925,3936|false|false|false|C4284232|Medications|medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3944,3950|false|false|false|C4255046||report
Event|Event|SIMPLE_SEGMENT|3944,3950|false|false|false|||report
Finding|Intellectual Product|SIMPLE_SEGMENT|3944,3950|false|false|false|C0684224|Report (document)|report
Procedure|Health Care Activity|SIMPLE_SEGMENT|3944,3950|false|false|false|C0700287|Reporting|report
Event|Event|SIMPLE_SEGMENT|3963,3974|false|false|false|||sensitivity
Finding|Finding|SIMPLE_SEGMENT|3963,3974|false|false|false|C0020517;C0312418;C0427965|Antimicrobial susceptibility;Hypersensitivity;Sensitivity (Personality)|sensitivity
Finding|Mental Process|SIMPLE_SEGMENT|3963,3974|false|false|false|C0020517;C0312418;C0427965|Antimicrobial susceptibility;Hypersensitivity;Sensitivity (Personality)|sensitivity
Finding|Pathologic Function|SIMPLE_SEGMENT|3963,3974|false|false|false|C0020517;C0312418;C0427965|Antimicrobial susceptibility;Hypersensitivity;Sensitivity (Personality)|sensitivity
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3979,3990|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3979,3990|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|3979,3990|false|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|3979,3990|false|false|false|C4284232|Medications|medications
Event|Event|SIMPLE_SEGMENT|3995,4002|false|false|false|||concern
Finding|Idea or Concept|SIMPLE_SEGMENT|3995,4002|false|false|false|C2699424|Concern|concern
Finding|Finding|SIMPLE_SEGMENT|4007,4015|false|false|false|C0332149|Possible|possible
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|4016,4032|false|true|false|C0005586|Bipolar Disorder|bipolar disorder
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4024,4032|false|true|false|C0012634|Disease|disorder
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4033,4042|false|true|false|C0945731||diagnosis
Event|Event|SIMPLE_SEGMENT|4033,4042|false|false|false|||diagnosis
Finding|Classification|SIMPLE_SEGMENT|4033,4042|false|true|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|4033,4042|false|true|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4033,4042|false|true|false|C0011900|Diagnosis|diagnosis
Event|Event|SIMPLE_SEGMENT|4056,4062|false|false|false|||follow
Finding|Idea or Concept|SIMPLE_SEGMENT|4066,4073|false|true|false|C1691786;C1704475|Pending - Allergy Clinical Status;Pending - referral status|pending
Drug|Organic Chemical|SIMPLE_SEGMENT|4074,4082|false|false|false|C0039840;C3714802|Thiamine Drug Class;thiamine|thiamine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4074,4082|false|false|false|C0039840;C3714802|Thiamine Drug Class;thiamine|thiamine
Drug|Vitamin|SIMPLE_SEGMENT|4074,4082|false|false|false|C0039840;C3714802|Thiamine Drug Class;thiamine|thiamine
Event|Event|SIMPLE_SEGMENT|4074,4082|false|false|false|||thiamine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4074,4082|false|false|false|C0373727|Thiamine measurement|thiamine
Finding|Intellectual Product|SIMPLE_SEGMENT|4092,4097|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|ACUTE
Event|Event|SIMPLE_SEGMENT|4098,4104|false|false|false|||ISSUES
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|4122,4125|false|false|false|C0270549|Generalized Anxiety Disorder|GAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4122,4125|false|false|false|C0017785|Glutamate Decarboxylase|GAD
Drug|Enzyme|SIMPLE_SEGMENT|4122,4125|false|false|false|C0017785|Glutamate Decarboxylase|GAD
Event|Event|SIMPLE_SEGMENT|4122,4125|false|false|false|||GAD
Finding|Gene or Genome|SIMPLE_SEGMENT|4122,4125|false|false|false|C1414925;C5575531|GAD1 gene;GAD1 wt Allele|GAD
Finding|Finding|SIMPLE_SEGMENT|4126,4131|false|false|false|C0030318|Panic|Panic
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|4126,4140|false|false|false|C0030319|Panic Disorder|Panic disorder
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4132,4140|false|false|false|C0012634|Disease|disorder
Event|Event|SIMPLE_SEGMENT|4132,4140|false|false|false|||disorder
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|4143,4153|false|false|false|C0011570;C0011581;C0344315;C0812393|Cancer patients and suicide and depression;Depressed mood;Depressive disorder;Mental Depression|Depression
Event|Event|SIMPLE_SEGMENT|4143,4153|false|false|false|||Depression
Finding|Functional Concept|SIMPLE_SEGMENT|4143,4153|false|false|false|C0460137;C1579931|Depression - motion|Depression
Finding|Sign or Symptom|SIMPLE_SEGMENT|4143,4153|false|false|false|C0460137;C1579931|Depression - motion|Depression
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4156,4160|false|false|false|C0038436;C0878676|6-pyruvoyl-tetrahydropterin synthase deficiency;Post-Traumatic Stress Disorder|PTSD
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|4156,4160|false|false|false|C0038436;C0878676|6-pyruvoyl-tetrahydropterin synthase deficiency;Post-Traumatic Stress Disorder|PTSD
Event|Event|SIMPLE_SEGMENT|4156,4160|false|false|false|||PTSD
Finding|Conceptual Entity|SIMPLE_SEGMENT|4163,4173|false|false|false|C0205245;C0542341;C2700217|Function (attribute);Functional;Functional Relationship|Functional
Finding|Functional Concept|SIMPLE_SEGMENT|4163,4173|false|false|false|C0205245;C0542341;C2700217|Function (attribute);Functional;Functional Relationship|Functional
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|4163,4195|false|false|false|C0009946;C4543816|Conversion disorder;Dissociative neurological symptom disorder (disorder)|Functional neurological disorder
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4174,4195|false|false|false|C0027765|nervous system disorder|neurological disorder
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4187,4195|false|false|false|C0012634|Disease|disorder
Event|Event|SIMPLE_SEGMENT|4187,4195|false|false|false|||disorder
Finding|Body Substance|SIMPLE_SEGMENT|4196,4203|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|4196,4203|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|4196,4203|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|4204,4213|false|false|false|||presented
Event|Event|SIMPLE_SEGMENT|4221,4228|false|false|false|||therapy
Finding|Finding|SIMPLE_SEGMENT|4221,4228|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|SIMPLE_SEGMENT|4221,4228|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4221,4228|false|false|false|C0087111|Therapeutic procedure|therapy
Event|Event|SIMPLE_SEGMENT|4229,4236|false|false|false|||session
Event|Event|SIMPLE_SEGMENT|4229,4236|false|false|false|C1883016|Activity Session|session
Finding|Conceptual Entity|SIMPLE_SEGMENT|4229,4236|false|false|false|C1883017|Session|session
Event|Event|SIMPLE_SEGMENT|4251,4256|false|false|false|||acute
Finding|Intellectual Product|SIMPLE_SEGMENT|4251,4256|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|SIMPLE_SEGMENT|4258,4263|false|false|false|||onset
Event|Event|SIMPLE_SEGMENT|4267,4275|false|false|false|||weakness
Finding|Sign or Symptom|SIMPLE_SEGMENT|4267,4275|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Finding|Finding|SIMPLE_SEGMENT|4277,4285|false|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Finding|Idea or Concept|SIMPLE_SEGMENT|4277,4285|false|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4277,4294|false|false|false|C0013384|Dyskinetic syndrome|abnormal movement
Finding|Finding|SIMPLE_SEGMENT|4277,4294|false|false|false|C0558189|Abnormal movement|abnormal movement
Event|Event|SIMPLE_SEGMENT|4286,4294|false|false|false|||movement
Finding|Organism Function|SIMPLE_SEGMENT|4286,4294|false|false|false|C0026649|Movement|movement
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|4299,4306|false|false|false|C0003537|Aphasia|aphasia
Event|Event|SIMPLE_SEGMENT|4299,4306|false|false|false|||aphasia
Finding|Mental Process|SIMPLE_SEGMENT|4314,4321|false|false|false|C0542559|contextual factors|setting
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4336,4343|false|false|false|C0032930|Precipitating Factors|trigger
Event|Event|SIMPLE_SEGMENT|4336,4343|false|false|false|||trigger
Event|Event|SIMPLE_SEGMENT|4347,4353|false|false|false|||seeing
Event|Event|SIMPLE_SEGMENT|4354,4361|false|false|false|||shadows
Finding|Functional Concept|SIMPLE_SEGMENT|4354,4361|false|false|false|C0332554|Shadow|shadows
Event|Event|SIMPLE_SEGMENT|4389,4398|false|false|false|||therapist
Event|Event|SIMPLE_SEGMENT|4460,4473|false|false|false|||hypervigilant
Event|Event|SIMPLE_SEGMENT|4478,4486|false|false|false|||stressed
Finding|Finding|SIMPLE_SEGMENT|4478,4486|false|false|false|C0038435|Stress|stressed
Event|Event|SIMPLE_SEGMENT|4499,4503|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|4499,4503|false|false|true|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|4499,4503|false|false|true|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|4499,4503|false|false|true|C1553498|home health encounter|home
Event|Event|SIMPLE_SEGMENT|4513,4521|false|false|false|||holidays
Event|Event|SIMPLE_SEGMENT|4513,4521|false|false|false|C0019843|Holidays|holidays
Event|Event|SIMPLE_SEGMENT|4525,4528|false|false|false|||see
Anatomy|Cell Component|SIMPLE_SEGMENT|4533,4536|false|false|false|C3811401|mycolate outer membrane|mom
Finding|Classification|SIMPLE_SEGMENT|4549,4554|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|major
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4555,4562|false|false|false|C0032930|Precipitating Factors|trigger
Event|Event|SIMPLE_SEGMENT|4555,4562|false|false|false|||trigger
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4571,4575|false|false|false|C0038436;C0878676|6-pyruvoyl-tetrahydropterin synthase deficiency;Post-Traumatic Stress Disorder|PTSD
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|4571,4575|false|false|false|C0038436;C0878676|6-pyruvoyl-tetrahydropterin synthase deficiency;Post-Traumatic Stress Disorder|PTSD
Event|Event|SIMPLE_SEGMENT|4571,4575|false|false|false|||PTSD
Event|Event|SIMPLE_SEGMENT|4597,4604|false|false|false|||reports
Event|Event|SIMPLE_SEGMENT|4607,4614|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|4607,4614|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|4607,4614|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|4607,4614|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|4607,4617|false|false|false|C0262926|Medical History|history of
Event|Event|SIMPLE_SEGMENT|4618,4624|false|false|false|||sexual
Finding|Behavior|SIMPLE_SEGMENT|4618,4624|false|false|false|C0036864|Sex Behavior|sexual
Event|Event|SIMPLE_SEGMENT|4625,4633|false|false|false|||physical
Finding|Finding|SIMPLE_SEGMENT|4625,4633|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Finding|Functional Concept|SIMPLE_SEGMENT|4625,4633|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|4625,4633|false|false|false|C0031809|Physical Examination|physical
Event|Event|SIMPLE_SEGMENT|4634,4640|false|false|false|||verbal
Finding|Functional Concept|SIMPLE_SEGMENT|4634,4640|false|false|false|C1548941|Participation Mode - verbal|verbal
Procedure|Health Care Activity|SIMPLE_SEGMENT|4634,4640|false|false|false|C1608381|Consent Mode - Verbal|verbal
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|4642,4647|false|false|false|C0013146|Drug abuse|abuse
Event|Event|SIMPLE_SEGMENT|4642,4647|false|false|false|||abuse
Event|Event|SIMPLE_SEGMENT|4642,4647|false|false|false|C1546935|Abuse|abuse
Finding|Finding|SIMPLE_SEGMENT|4642,4647|false|false|false|C0562381|Victim of abuse (finding)|abuse
Event|Event|SIMPLE_SEGMENT|4652,4659|false|false|false|||patient
Finding|Body Substance|SIMPLE_SEGMENT|4652,4659|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|4652,4659|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|4652,4659|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|4668,4675|false|false|false|||guarded
Event|Event|SIMPLE_SEGMENT|4698,4705|false|false|false|||discuss
Event|Event|SIMPLE_SEGMENT|4714,4726|false|false|false|||presentation
Finding|Idea or Concept|SIMPLE_SEGMENT|4714,4726|false|false|false|C0449450|Presentation|presentation
Finding|Idea or Concept|SIMPLE_SEGMENT|4742,4753|false|false|false|C0750502|Significant|significant
Finding|Intellectual Product|SIMPLE_SEGMENT|4758,4763|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Conceptual Entity|SIMPLE_SEGMENT|4765,4775|false|false|false|C0205245;C0542341;C2700217|Function (attribute);Functional;Functional Relationship|functional
Finding|Functional Concept|SIMPLE_SEGMENT|4765,4775|false|false|false|C0205245;C0542341;C2700217|Function (attribute);Functional;Functional Relationship|functional
Finding|Sign or Symptom|SIMPLE_SEGMENT|4776,4797|false|false|false|C0235031|Neurologic Symptoms|neurological symptoms
Event|Event|SIMPLE_SEGMENT|4789,4797|false|false|false|||symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|4789,4797|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|4789,4797|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|SIMPLE_SEGMENT|4809,4817|false|false|false|||weakness
Finding|Sign or Symptom|SIMPLE_SEGMENT|4809,4817|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Event|Event|SIMPLE_SEGMENT|4819,4827|false|false|false|||abnormal
Finding|Finding|SIMPLE_SEGMENT|4819,4827|false|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Finding|Idea or Concept|SIMPLE_SEGMENT|4819,4827|false|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Event|Event|SIMPLE_SEGMENT|4829,4837|false|false|false|||movement
Finding|Organism Function|SIMPLE_SEGMENT|4829,4837|false|false|false|C0026649|Movement|movement
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|4843,4850|false|false|false|C0003537|Aphasia|aphasia
Event|Event|SIMPLE_SEGMENT|4843,4850|false|false|false|||aphasia
Event|Event|SIMPLE_SEGMENT|4852,4861|false|false|false|||resulting
Finding|Functional Concept|SIMPLE_SEGMENT|4865,4873|false|false|false|C0221099|Impaired|impaired
Event|Event|SIMPLE_SEGMENT|4874,4885|false|false|false|||functioning
Finding|Functional Concept|SIMPLE_SEGMENT|4874,4885|false|false|false|C0205245;C0542341|Function (attribute);Functional|functioning
Event|Event|SIMPLE_SEGMENT|4898,4905|false|false|false|||concern
Finding|Idea or Concept|SIMPLE_SEGMENT|4898,4905|false|false|false|C2699424|Concern|concern
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|4910,4919|false|false|false|C0007398|Catatonia|catatonia
Event|Event|SIMPLE_SEGMENT|4910,4919|false|false|false|||catatonia
Event|Event|SIMPLE_SEGMENT|4928,4936|false|false|false|||improved
Drug|Organic Chemical|SIMPLE_SEGMENT|4951,4957|false|false|false|C0699194|Ativan|ativan
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4951,4957|false|false|false|C0699194|Ativan|ativan
Event|Event|SIMPLE_SEGMENT|4951,4957|false|false|false|||ativan
Event|Event|SIMPLE_SEGMENT|4974,4982|false|false|false|||endorsed
Finding|Idea or Concept|SIMPLE_SEGMENT|4983,4994|false|false|false|C0750502|Significant|significant
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|4995,5002|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Event|Event|SIMPLE_SEGMENT|4995,5002|false|false|false|||anxiety
Finding|Sign or Symptom|SIMPLE_SEGMENT|4995,5002|false|false|false|C0860603|Anxiety symptoms|anxiety
Event|Event|SIMPLE_SEGMENT|5008,5014|false|false|false|||denied
Event|Event|SIMPLE_SEGMENT|5052,5056|false|false|false|||meet
Event|Event|SIMPLE_SEGMENT|5061,5069|false|false|false|||criteria
Finding|Idea or Concept|SIMPLE_SEGMENT|5061,5069|false|false|false|C0243161|criteria|criteria
Event|Event|SIMPLE_SEGMENT|5090,5097|false|false|false|||episode
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|5111,5118|false|false|false|C0082568|ferryl iron|IV iron
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5114,5118|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|5114,5118|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5114,5118|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Event|Event|SIMPLE_SEGMENT|5114,5118|false|false|false|||iron
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5114,5118|false|false|false|C0337439|Iron measurement|iron
Event|Event|SIMPLE_SEGMENT|5119,5127|false|false|false|||infusion
Finding|Functional Concept|SIMPLE_SEGMENT|5119,5127|false|false|false|C1827465|Infusion route|infusion
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5119,5127|false|false|false|C0574032|Infusion procedures|infusion
Event|Event|SIMPLE_SEGMENT|5137,5145|false|false|false|||admitted
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5153,5170|false|false|false|C0587591|neurology services (treatment)|neurology service
Event|Occupational Activity|SIMPLE_SEGMENT|5163,5170|false|false|false|C0557854|Services|service
Finding|Idea or Concept|SIMPLE_SEGMENT|5163,5170|false|false|false|C3245478|ActInformationPrivacyReason - service|service
Event|Event|SIMPLE_SEGMENT|5186,5195|false|false|false|||diagnosed
Finding|Conceptual Entity|SIMPLE_SEGMENT|5202,5212|false|false|false|C0205245;C0542341;C2700217|Function (attribute);Functional;Functional Relationship|functional
Finding|Functional Concept|SIMPLE_SEGMENT|5202,5212|false|false|false|C0205245;C0542341;C2700217|Function (attribute);Functional;Functional Relationship|functional
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|5202,5234|false|false|false|C0009946;C4543816|Conversion disorder;Dissociative neurological symptom disorder (disorder)|functional neurological disorder
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5213,5234|false|false|false|C0027765|nervous system disorder|neurological disorder
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5226,5234|false|false|false|C0012634|Disease|disorder
Event|Event|SIMPLE_SEGMENT|5226,5234|false|false|false|||disorder
Event|Event|SIMPLE_SEGMENT|5243,5251|false|false|false|||improved
Event|Event|SIMPLE_SEGMENT|5266,5271|false|false|false|||rehab
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5266,5271|false|false|false|C0034991|Rehabilitation therapy|rehab
Event|Event|SIMPLE_SEGMENT|5286,5293|false|false|false|||started
Event|Event|SIMPLE_SEGMENT|5297,5310|false|false|false|||nortriptyline
Finding|Finding|SIMPLE_SEGMENT|5330,5334|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|5330,5334|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|5330,5334|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|SIMPLE_SEGMENT|5344,5353|false|false|false|||therapist
Finding|Functional Concept|SIMPLE_SEGMENT|5359,5374|false|false|false|C0332324|Sensitive|is sensitive to
Event|Event|SIMPLE_SEGMENT|5362,5371|false|false|false|||sensitive
Finding|Functional Concept|SIMPLE_SEGMENT|5362,5371|false|false|false|C0332324|Sensitive|sensitive
Finding|Functional Concept|SIMPLE_SEGMENT|5362,5374|false|false|false|C0332324|Sensitive|sensitive to
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5375,5386|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5375,5386|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|5375,5386|false|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|5375,5386|false|false|false|C4284232|Medications|medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5408,5413|false|false|false|C0360105|Selective Serotonin Reuptake Inhibitors|SSRIs
Event|Event|SIMPLE_SEGMENT|5408,5413|false|false|false|||SSRIs
Event|Event|SIMPLE_SEGMENT|5418,5424|false|false|false|||became
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|5425,5430|false|false|false|C0338831|Manic|manic
Event|Event|SIMPLE_SEGMENT|5425,5430|false|false|false|||manic
Finding|Finding|SIMPLE_SEGMENT|5425,5430|false|false|false|C0564408|Manic mood|manic
Event|Event|SIMPLE_SEGMENT|5468,5477|false|false|false|||diagnosed
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|5483,5499|false|false|false|C0005586|Bipolar Disorder|bipolar disorder
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5491,5499|false|false|false|C0012634|Disease|disorder
Event|Event|SIMPLE_SEGMENT|5491,5499|false|false|false|||disorder
Event|Event|SIMPLE_SEGMENT|5506,5514|false|false|false|||admitted
Event|Event|SIMPLE_SEGMENT|5525,5537|false|false|false|||re-evaluated
Event|Event|SIMPLE_SEGMENT|5566,5576|false|false|false|||determined
Event|Event|SIMPLE_SEGMENT|5591,5601|false|false|false|||consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|5591,5601|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|5591,5606|false|false|false|C0332290|Consistent with|consistent with
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|5607,5616|false|false|false|C0007398|Catatonia|catatonia
Event|Event|SIMPLE_SEGMENT|5607,5616|false|false|false|||catatonia
Finding|Finding|SIMPLE_SEGMENT|5633,5639|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|5633,5639|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Conceptual Entity|SIMPLE_SEGMENT|5641,5651|false|false|false|C0205245;C0542341;C2700217|Function (attribute);Functional;Functional Relationship|functional
Finding|Functional Concept|SIMPLE_SEGMENT|5641,5651|false|false|false|C0205245;C0542341;C2700217|Function (attribute);Functional;Functional Relationship|functional
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|5641,5673|false|false|false|C0009946;C4543816|Conversion disorder;Dissociative neurological symptom disorder (disorder)|functional neurological disorder
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5652,5673|false|false|false|C0027765|nervous system disorder|neurological disorder
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5665,5673|false|false|false|C0012634|Disease|disorder
Event|Event|SIMPLE_SEGMENT|5665,5673|false|false|false|||disorder
Event|Event|SIMPLE_SEGMENT|5683,5694|false|false|false|||recommended
Event|Event|SIMPLE_SEGMENT|5699,5704|false|false|false|||acute
Finding|Intellectual Product|SIMPLE_SEGMENT|5699,5704|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|SIMPLE_SEGMENT|5706,5711|false|false|false|||rehab
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5706,5711|false|false|false|C0034991|Rehabilitation therapy|rehab
Event|Event|SIMPLE_SEGMENT|5715,5723|false|false|false|||continue
Event|Event|SIMPLE_SEGMENT|5724,5734|false|false|false|||aggressive
Finding|Individual Behavior|SIMPLE_SEGMENT|5724,5734|false|false|false|C0001807;C1547300;C1548760|Aggressive behavior;Precaution Code - Aggressive;Risk Codes - Aggressive|aggressive
Finding|Intellectual Product|SIMPLE_SEGMENT|5724,5734|false|false|false|C0001807;C1547300;C1548760|Aggressive behavior;Precaution Code - Aggressive;Risk Codes - Aggressive|aggressive
Event|Event|SIMPLE_SEGMENT|5748,5757|false|false|false|||continued
Event|Event|SIMPLE_SEGMENT|5761,5765|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|5761,5765|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|5761,5765|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|5761,5765|false|false|false|C1553498|home health encounter|home
Event|Event|SIMPLE_SEGMENT|5804,5810|false|false|false|||eating
Finding|Organism Function|SIMPLE_SEGMENT|5804,5810|false|false|false|C0013470|Eating|eating
Finding|Finding|SIMPLE_SEGMENT|5812,5830|false|false|false|C5687959|Restrained eating behavior|Restrictive eating
Event|Event|SIMPLE_SEGMENT|5824,5830|false|false|false|||eating
Finding|Organism Function|SIMPLE_SEGMENT|5824,5830|false|false|false|C0013470|Eating|eating
Event|Event|SIMPLE_SEGMENT|5859,5866|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|5859,5866|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|5859,5866|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|5859,5866|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|5859,5869|false|false|false|C0262926|Medical History|history of
Finding|Finding|SIMPLE_SEGMENT|5870,5888|false|false|false|C5687959|Restrained eating behavior|restrictive eating
Event|Event|SIMPLE_SEGMENT|5882,5888|false|false|false|||eating
Finding|Organism Function|SIMPLE_SEGMENT|5882,5888|false|false|false|C0013470|Eating|eating
Event|Event|SIMPLE_SEGMENT|5938,5949|false|false|false|||bradycardia
Finding|Finding|SIMPLE_SEGMENT|5938,5949|false|false|false|C0428977;C3812171|Bradycardia;Bradycardia by ECG Finding|bradycardia
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5954,5965|false|false|false|C0013832;C3536863|Electrolyte [EPC];Electrolytes|electrolyte
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5954,5965|false|false|false|C0013832;C3536863|Electrolyte [EPC];Electrolytes|electrolyte
Event|Event|SIMPLE_SEGMENT|5954,5965|false|false|false|||electrolyte
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|5967,5980|false|false|false|C0000768|Congenital Abnormality|abnormalities
Event|Event|SIMPLE_SEGMENT|5967,5980|false|false|false|||abnormalities
Finding|Functional Concept|SIMPLE_SEGMENT|5967,5980|false|false|false|C0000769|teratologic|abnormalities
Event|Event|SIMPLE_SEGMENT|5990,5999|false|false|false|||therapist
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|6005,6022|false|false|false|C0855228|Eating disorder symptom|disordered eating
Event|Event|SIMPLE_SEGMENT|6016,6022|false|false|false|||eating
Finding|Organism Function|SIMPLE_SEGMENT|6016,6022|false|false|false|C0013470|Eating|eating
Event|Event|SIMPLE_SEGMENT|6028,6034|false|false|false|||become
Finding|Finding|SIMPLE_SEGMENT|6035,6039|false|false|false|C4281574|Much|much
Finding|Finding|SIMPLE_SEGMENT|6035,6045|false|false|false|C3841448|Much worse|much worse
Event|Event|SIMPLE_SEGMENT|6040,6045|false|false|false|||worse
Finding|Finding|SIMPLE_SEGMENT|6040,6045|false|false|false|C1457868;C1550463|Observation Interpretation - worse;Worse|worse
Finding|Idea or Concept|SIMPLE_SEGMENT|6040,6045|false|false|false|C1457868;C1550463|Observation Interpretation - worse;Worse|worse
Finding|Mental Process|SIMPLE_SEGMENT|6078,6085|false|false|false|C0542559|contextual factors|setting
Event|Event|SIMPLE_SEGMENT|6090,6099|false|false|false|||traveling
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|6090,6099|false|false|false|C0040802|travel|traveling
Finding|Finding|SIMPLE_SEGMENT|6100,6105|false|false|false|C2984081|Very Much|a lot
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6102,6105|false|false|false|C0162435;C0175218|Olfactory tract;nucleus of the lateral olfactory tract|lot
Finding|Idea or Concept|SIMPLE_SEGMENT|6102,6105|false|false|false|C1710198|Stock (in-store merchandise)|lot
Event|Event|SIMPLE_SEGMENT|6110,6114|false|false|false|||work
Event|Occupational Activity|SIMPLE_SEGMENT|6110,6114|false|false|false|C0043227|Work|work
Event|Event|SIMPLE_SEGMENT|6120,6127|false|false|false|||started
Event|Event|SIMPLE_SEGMENT|6141,6151|false|false|false|||outpatient
Finding|Classification|SIMPLE_SEGMENT|6141,6151|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|6141,6151|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Drug|Organic Chemical|SIMPLE_SEGMENT|6153,6160|false|false|false|C2728259|Program|program
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6153,6160|false|false|false|C2728259|Program|program
Event|Event|SIMPLE_SEGMENT|6153,6160|false|false|false|||program
Finding|Conceptual Entity|SIMPLE_SEGMENT|6153,6160|false|false|false|C0376691;C1709697;C3484370|Program - framework of goals;Programs;Programs - Publication Format|program
Finding|Functional Concept|SIMPLE_SEGMENT|6153,6160|false|false|false|C0376691;C1709697;C3484370|Program - framework of goals;Programs;Programs - Publication Format|program
Finding|Intellectual Product|SIMPLE_SEGMENT|6153,6160|false|false|false|C0376691;C1709697;C3484370|Program - framework of goals;Programs;Programs - Publication Format|program
Event|Event|SIMPLE_SEGMENT|6196,6205|false|false|false|||therapist
Event|Event|SIMPLE_SEGMENT|6211,6220|false|false|false|||restricts
Event|Event|SIMPLE_SEGMENT|6225,6233|false|false|false|||calories
Finding|Idea or Concept|SIMPLE_SEGMENT|6260,6263|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|6260,6263|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|6268,6282|false|false|false|||over-exercises
Event|Event|SIMPLE_SEGMENT|6290,6294|false|false|false|||good
Finding|Idea or Concept|SIMPLE_SEGMENT|6290,6294|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Event|Event|SIMPLE_SEGMENT|6298,6304|false|false|false|||hiding
Event|Event|SIMPLE_SEGMENT|6327,6333|false|false|false|||review
Finding|Idea or Concept|SIMPLE_SEGMENT|6327,6333|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Finding|Intellectual Product|SIMPLE_SEGMENT|6327,6333|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Finding|Functional Concept|SIMPLE_SEGMENT|6327,6336|false|false|false|C0699752|Review of|review of
Event|Event|SIMPLE_SEGMENT|6337,6340|false|false|false|||OMR
Finding|Gene or Genome|SIMPLE_SEGMENT|6337,6340|false|false|false|C1412647|ATP5F1A gene|OMR
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6346,6349|false|false|false|C1305855;C1542867|Body mass index|BMI
Event|Event|SIMPLE_SEGMENT|6346,6349|false|false|false|||BMI
Finding|Finding|SIMPLE_SEGMENT|6346,6349|false|false|false|C0578022|Finding of body mass index|BMI
Event|Event|SIMPLE_SEGMENT|6362,6368|false|false|false|||normal
Drug|Inorganic Chemical|SIMPLE_SEGMENT|6419,6430|true|false|false|C0013832;C3536863|Electrolyte [EPC];Electrolytes|electrolyte
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6419,6430|true|false|false|C0013832;C3536863|Electrolyte [EPC];Electrolytes|electrolyte
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|6431,6444|true|false|false|C0000768|Congenital Abnormality|abnormalities
Event|Event|SIMPLE_SEGMENT|6431,6444|false|false|false|||abnormalities
Finding|Functional Concept|SIMPLE_SEGMENT|6431,6444|true|false|false|C0000769|teratologic|abnormalities
Event|Event|SIMPLE_SEGMENT|6478,6489|false|false|false|||bradycardic
Event|Event|SIMPLE_SEGMENT|6515,6523|false|false|false|||appetite
Finding|Organism Function|SIMPLE_SEGMENT|6515,6523|false|false|false|C0003618|Desire for food|appetite
Event|Event|SIMPLE_SEGMENT|6524,6532|false|false|false|||improved
Finding|Sign or Symptom|SIMPLE_SEGMENT|6540,6561|false|false|false|C0235031|Neurologic Symptoms|neurological symptoms
Event|Event|SIMPLE_SEGMENT|6553,6561|false|false|false|||symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|6553,6561|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|6553,6561|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|SIMPLE_SEGMENT|6569,6578|false|false|false|||resolving
Event|Event|SIMPLE_SEGMENT|6584,6593|false|false|false|||nutrition
Finding|Finding|SIMPLE_SEGMENT|6584,6593|false|false|false|C0392209;C0518896;C1442959|Nutrition (function);Nutrition outcomes;Nutritional status|nutrition
Finding|Intellectual Product|SIMPLE_SEGMENT|6584,6593|false|false|false|C0392209;C0518896;C1442959|Nutrition (function);Nutrition outcomes;Nutritional status|nutrition
Finding|Organism Function|SIMPLE_SEGMENT|6584,6593|false|false|false|C0392209;C0518896;C1442959|Nutrition (function);Nutrition outcomes;Nutritional status|nutrition
Procedure|Research Activity|SIMPLE_SEGMENT|6584,6593|false|false|false|C0600072;C1521729|Feeding and dietary regimes;Nutritional Study|nutrition
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6584,6593|false|false|false|C0600072;C1521729|Feeding and dietary regimes;Nutritional Study|nutrition
Event|Event|SIMPLE_SEGMENT|6594,6604|false|false|false|||evaluation
Finding|Idea or Concept|SIMPLE_SEGMENT|6594,6604|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|SIMPLE_SEGMENT|6594,6604|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Event|Event|SIMPLE_SEGMENT|6609,6613|false|false|false|||need
Finding|Functional Concept|SIMPLE_SEGMENT|6609,6613|true|false|false|C0686904|Patient need for (contextual qualifier)|need
Finding|Functional Concept|SIMPLE_SEGMENT|6609,6617|true|false|false|C0686904|Patient need for (contextual qualifier)|need for
Finding|Organism Function|SIMPLE_SEGMENT|6618,6624|false|false|false|C0013470|Eating|eating
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|6618,6633|false|false|false|C0013473|Eating Disorders|eating disorder
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6625,6633|false|false|false|C0012634|Disease|disorder
Event|Event|SIMPLE_SEGMENT|6625,6633|false|false|false|||disorder
Event|Event|SIMPLE_SEGMENT|6635,6643|false|false|false|||protocol
Finding|Finding|SIMPLE_SEGMENT|6635,6643|false|false|false|C0442711;C1507394;C1522729;C2348563;C3715209|Clinical trial protocol document;Library Protocol;Protocol - answer to question;Protocols documentation;Study Protocol|protocol
Finding|Intellectual Product|SIMPLE_SEGMENT|6635,6643|false|false|false|C0442711;C1507394;C1522729;C2348563;C3715209|Clinical trial protocol document;Library Protocol;Protocol - answer to question;Protocols documentation;Study Protocol|protocol
Event|Event|SIMPLE_SEGMENT|6650,6659|false|false|false|||inpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|6650,6659|false|false|false|C1548438;C1549404|Patient Class - Inpatient;Referral category - Inpatient|inpatient
Procedure|Health Care Activity|SIMPLE_SEGMENT|6650,6659|false|false|false|C1555324|inpatient encounter|inpatient
Drug|Food|SIMPLE_SEGMENT|6674,6680|false|false|false|C0218063|Ensure (product)|Ensure
Event|Event|SIMPLE_SEGMENT|6681,6692|false|false|false|||supplements
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6694,6699|false|false|false|C0018787;C4037974|Chest>Heart;Heart|Heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6694,6699|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|Heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|6694,6699|false|false|false|C0795691|HEART PROBLEM|Heart
Event|Event|SIMPLE_SEGMENT|6701,6706|false|false|false|||rates
Event|Event|SIMPLE_SEGMENT|6712,6718|false|false|false|||stable
Finding|Intellectual Product|SIMPLE_SEGMENT|6712,6718|false|false|false|C1547311|Patient Condition Code - Stable|stable
Event|Event|SIMPLE_SEGMENT|6720,6731|false|false|false|||bradycardic
Drug|Inorganic Chemical|SIMPLE_SEGMENT|6740,6752|false|false|false|C0013832;C3536863|Electrolyte [EPC];Electrolytes|Electrolytes
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6740,6752|false|false|false|C0013832;C3536863|Electrolyte [EPC];Electrolytes|Electrolytes
Event|Event|SIMPLE_SEGMENT|6759,6768|false|false|false|||monitored
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6770,6773|false|false|false|C2708739||TSH
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6770,6773|false|false|false|C0040160|thyrotropin|TSH
Drug|Hormone|SIMPLE_SEGMENT|6770,6773|false|false|false|C0040160|thyrotropin|TSH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6770,6773|false|false|false|C0040160|thyrotropin|TSH
Event|Event|SIMPLE_SEGMENT|6770,6773|false|false|false|||TSH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6770,6773|false|false|false|C0202230|Thyroid stimulating hormone measurement|TSH
Finding|Gene or Genome|SIMPLE_SEGMENT|6782,6785|false|false|false|C1417635;C1420797;C3538796|NDUFB3 gene;TNFAIP1 gene;TNFAIP1 wt Allele|B12
Event|Event|SIMPLE_SEGMENT|6786,6792|false|false|false|||levels
Event|Event|SIMPLE_SEGMENT|6802,6808|false|false|false|||normal
Event|Event|SIMPLE_SEGMENT|6814,6822|false|false|false|||received
Drug|Organic Chemical|SIMPLE_SEGMENT|6824,6832|false|false|false|C0039840;C3714802|Thiamine Drug Class;thiamine|thiamine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6824,6832|false|false|false|C0039840;C3714802|Thiamine Drug Class;thiamine|thiamine
Drug|Vitamin|SIMPLE_SEGMENT|6824,6832|false|false|false|C0039840;C3714802|Thiamine Drug Class;thiamine|thiamine
Event|Event|SIMPLE_SEGMENT|6824,6832|false|false|false|||thiamine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6824,6832|false|false|false|C0373727|Thiamine measurement|thiamine
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6824,6848|false|false|false|C4524016|Thiamin supplementation|thiamine supplementation
Event|Event|SIMPLE_SEGMENT|6833,6848|false|false|false|||supplementation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6833,6848|false|false|false|C0242297|Dietary Supplementation|supplementation
Drug|Organic Chemical|SIMPLE_SEGMENT|6863,6869|false|false|false|C0206046|Zofran|Zofran
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6863,6869|false|false|false|C0206046|Zofran|Zofran
Event|Event|SIMPLE_SEGMENT|6870,6873|false|false|false|||PRN
Finding|Gene or Genome|SIMPLE_SEGMENT|6870,6873|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6878,6884|false|false|false|C4255480||nausea
Event|Event|SIMPLE_SEGMENT|6878,6884|false|false|false|||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|6878,6884|false|false|false|C0027497|Nausea|nausea
Anatomy|Cell Component|SIMPLE_SEGMENT|6898,6902|false|false|false|C1167518|viral nucleocapsid location|CORE
Finding|Body Substance|SIMPLE_SEGMENT|6898,6902|false|false|false|C3274653|Core Specimen|CORE
Event|Event|SIMPLE_SEGMENT|6903,6911|false|false|false|||MEASURES
Finding|Functional Concept|SIMPLE_SEGMENT|6903,6911|false|false|false|C1879489|Measures (attribute)|MEASURES
Event|Event|SIMPLE_SEGMENT|6927,6931|false|false|false|||CODE
Event|Occupational Activity|SIMPLE_SEGMENT|6927,6931|false|false|false|C0009219|Coding|CODE
Finding|Intellectual Product|SIMPLE_SEGMENT|6927,6931|false|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|CODE
Event|Occupational Activity|SIMPLE_SEGMENT|6938,6942|false|false|false|C0009219|Coding|code
Finding|Intellectual Product|SIMPLE_SEGMENT|6938,6942|false|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|code
Event|Activity|SIMPLE_SEGMENT|6945,6952|false|false|false|C3812666|Personal Contact|CONTACT
Event|Event|SIMPLE_SEGMENT|6945,6952|false|false|false|||CONTACT
Finding|Functional Concept|SIMPLE_SEGMENT|6945,6952|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Finding|Idea or Concept|SIMPLE_SEGMENT|6945,6952|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Finding|Intellectual Product|SIMPLE_SEGMENT|6945,6952|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|6945,6952|false|false|false|C0392367|Physical contact|CONTACT
Finding|Body Substance|SIMPLE_SEGMENT|6958,6965|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|6958,6965|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|6958,6965|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Activity|SIMPLE_SEGMENT|6968,6975|false|false|false|C1272683||request
Event|Event|SIMPLE_SEGMENT|6968,6975|false|false|false|||request
Finding|Idea or Concept|SIMPLE_SEGMENT|6968,6975|false|false|false|C1522634;C1553397;C1553888|Question (inquiry);Request - ActReason;request - ActMood|request
Finding|Intellectual Product|SIMPLE_SEGMENT|6968,6975|false|false|false|C1522634;C1553397;C1553888|Question (inquiry);Request - ActReason;request - ActMood|request
Event|Event|SIMPLE_SEGMENT|6984,6991|false|false|false|||contact
Event|Event|SIMPLE_SEGMENT|6996,7002|false|false|false|||mother
Finding|Idea or Concept|SIMPLE_SEGMENT|6996,7002|false|false|false|C1546508|Relationship - Mother|mother
Event|Event|SIMPLE_SEGMENT|7011,7020|false|false|false|||Emergency
Finding|Finding|SIMPLE_SEGMENT|7011,7020|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Finding|Idea or Concept|SIMPLE_SEGMENT|7011,7020|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Finding|Intellectual Product|SIMPLE_SEGMENT|7011,7020|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Finding|Pathologic Function|SIMPLE_SEGMENT|7011,7020|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|7011,7020|false|false|false|C0013956|Emergency Situation|Emergency
Procedure|Health Care Activity|SIMPLE_SEGMENT|7011,7020|false|false|false|C1553500|emergency encounter|Emergency
Procedure|Health Care Activity|SIMPLE_SEGMENT|7021,7029|false|false|false|C4036459|Contacts|Contacts
Event|Event|SIMPLE_SEGMENT|7096,7107|false|false|false|||coordinates
Finding|Finding|SIMPLE_SEGMENT|7096,7107|false|false|false|C0427184;C0700114|Coordinated|coordinates
Finding|Functional Concept|SIMPLE_SEGMENT|7096,7107|false|false|false|C0427184;C0700114|Coordinated|coordinates
Event|Activity|SIMPLE_SEGMENT|7119,7123|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|7119,7123|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|7119,7123|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|7119,7123|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Event|Event|SIMPLE_SEGMENT|7128,7137|false|false|false|||available
Finding|Functional Concept|SIMPLE_SEGMENT|7128,7137|false|false|false|C0470187|Availability of|available
Event|Event|SIMPLE_SEGMENT|7142,7151|false|false|false|||questions
Event|Event|SIMPLE_SEGMENT|7152,7157|false|false|false|||calls
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7172,7183|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7172,7183|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|7172,7183|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|7172,7183|false|false|false|C4284232|Medications|Medications
Finding|Finding|SIMPLE_SEGMENT|7172,7196|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|SIMPLE_SEGMENT|7187,7196|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|7187,7196|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7215,7225|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|7215,7225|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|7215,7230|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|SIMPLE_SEGMENT|7226,7230|false|false|false|||list
Finding|Intellectual Product|SIMPLE_SEGMENT|7226,7230|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|SIMPLE_SEGMENT|7234,7242|false|false|false|||accurate
Drug|Organic Chemical|SIMPLE_SEGMENT|7247,7255|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7247,7255|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|SIMPLE_SEGMENT|7247,7255|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|SIMPLE_SEGMENT|7247,7255|false|false|false|||complete
Finding|Functional Concept|SIMPLE_SEGMENT|7247,7255|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|SIMPLE_SEGMENT|7247,7255|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Event|Event|SIMPLE_SEGMENT|7291,7300|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|7291,7300|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|7291,7300|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|7291,7300|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|7291,7300|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|7291,7312|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7301,7312|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7301,7312|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|7301,7312|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|7301,7312|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|SIMPLE_SEGMENT|7318,7331|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7318,7331|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|SIMPLE_SEGMENT|7318,7331|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Event|Event|SIMPLE_SEGMENT|7318,7331|false|false|false|||Multivitamins
Drug|Inorganic Chemical|SIMPLE_SEGMENT|7334,7342|false|false|false|C0026162|Minerals|minerals
Event|Event|SIMPLE_SEGMENT|7334,7342|false|false|false|||minerals
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7345,7348|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|SIMPLE_SEGMENT|7345,7348|false|false|false|||TAB
Drug|Organic Chemical|SIMPLE_SEGMENT|7364,7375|false|false|false|C0061851|ondansetron|Ondansetron
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7364,7375|false|false|false|C0061851|ondansetron|Ondansetron
Event|Event|SIMPLE_SEGMENT|7364,7375|false|false|false|||Ondansetron
Event|Event|SIMPLE_SEGMENT|7376,7379|false|false|false|||ODT
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7376,7379|false|false|false|C3898096|Optical Doppler Tomography|ODT
Finding|Gene or Genome|SIMPLE_SEGMENT|7392,7395|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7396,7402|false|false|false|C4255480||Nausea
Event|Event|SIMPLE_SEGMENT|7396,7402|false|false|false|||Nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|7396,7402|false|false|false|C0027497|Nausea|Nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|7396,7411|false|false|false|C0027498|Nausea and vomiting|Nausea/Vomiting
Finding|Sign or Symptom|SIMPLE_SEGMENT|7403,7411|false|false|false|C0042963|Vomiting|Vomiting
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7420,7424|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|Line
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|7420,7424|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|Line
Drug|Substance|SIMPLE_SEGMENT|7420,7424|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|Line
Event|Event|SIMPLE_SEGMENT|7420,7424|false|false|false|||Line
Finding|Intellectual Product|SIMPLE_SEGMENT|7420,7424|false|false|false|C1546701|line source specimen code|Line
Drug|Organic Chemical|SIMPLE_SEGMENT|7432,7440|false|false|false|C0039840;C3714802|Thiamine Drug Class;thiamine|Thiamine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7432,7440|false|false|false|C0039840;C3714802|Thiamine Drug Class;thiamine|Thiamine
Drug|Vitamin|SIMPLE_SEGMENT|7432,7440|false|false|false|C0039840;C3714802|Thiamine Drug Class;thiamine|Thiamine
Event|Event|SIMPLE_SEGMENT|7432,7440|false|false|false|||Thiamine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7432,7440|false|false|false|C0373727|Thiamine measurement|Thiamine
Event|Event|SIMPLE_SEGMENT|7495,7504|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|7495,7504|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|7495,7504|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|7495,7504|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|7495,7504|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7495,7516|false|false|false|C4019243||Discharge Disposition
Finding|Finding|SIMPLE_SEGMENT|7495,7516|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7505,7516|false|false|false|C2926604||Disposition
Event|Event|SIMPLE_SEGMENT|7505,7516|false|false|false|||Disposition
Procedure|Health Care Activity|SIMPLE_SEGMENT|7505,7516|false|false|false|C0184758|Patient disposition|Disposition
Finding|Finding|SIMPLE_SEGMENT|7518,7526|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|SIMPLE_SEGMENT|7518,7526|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Procedure|Health Care Activity|SIMPLE_SEGMENT|7518,7531|false|false|false|C0023977|long-term care|Extended Care
Event|Activity|SIMPLE_SEGMENT|7527,7531|false|false|false|C1947933|care activity|Care
Event|Event|SIMPLE_SEGMENT|7527,7531|false|false|false|||Care
Finding|Finding|SIMPLE_SEGMENT|7527,7531|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|SIMPLE_SEGMENT|7527,7531|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Event|Event|SIMPLE_SEGMENT|7534,7542|false|false|false|||Facility
Finding|Intellectual Product|SIMPLE_SEGMENT|7534,7542|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|SIMPLE_SEGMENT|7550,7559|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|7550,7559|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|7550,7559|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|7550,7559|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|7550,7559|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|7550,7569|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7560,7569|false|false|false|C0945731||Diagnosis
Event|Event|SIMPLE_SEGMENT|7560,7569|false|false|false|||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|7560,7569|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|7560,7569|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7560,7569|false|false|false|C0011900|Diagnosis|Diagnosis
Finding|Conceptual Entity|SIMPLE_SEGMENT|7572,7582|false|false|false|C0205245;C0542341;C2700217|Function (attribute);Functional;Functional Relationship|Functional
Finding|Functional Concept|SIMPLE_SEGMENT|7572,7582|false|false|false|C0205245;C0542341;C2700217|Function (attribute);Functional;Functional Relationship|Functional
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|7572,7604|false|false|false|C0009946;C4543816|Conversion disorder;Dissociative neurological symptom disorder (disorder)|Functional neurological disorder
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7583,7604|false|false|false|C0027765|nervous system disorder|neurological disorder
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7596,7604|false|false|false|C0012634|Disease|disorder
Event|Event|SIMPLE_SEGMENT|7596,7604|false|false|false|||disorder
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|7606,7609|false|false|false|C0270549|Generalized Anxiety Disorder|GAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7606,7609|false|false|false|C0017785|Glutamate Decarboxylase|GAD
Drug|Enzyme|SIMPLE_SEGMENT|7606,7609|false|false|false|C0017785|Glutamate Decarboxylase|GAD
Event|Event|SIMPLE_SEGMENT|7606,7609|false|false|false|||GAD
Finding|Gene or Genome|SIMPLE_SEGMENT|7606,7609|false|false|false|C1414925;C5575531|GAD1 gene;GAD1 wt Allele|GAD
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|7610,7620|false|false|false|C0011570;C0011581;C0344315;C0812393|Cancer patients and suicide and depression;Depressed mood;Depressive disorder;Mental Depression|depression
Event|Event|SIMPLE_SEGMENT|7610,7620|false|false|false|||depression
Finding|Functional Concept|SIMPLE_SEGMENT|7610,7620|false|false|false|C0460137;C1579931|Depression - motion|depression
Finding|Sign or Symptom|SIMPLE_SEGMENT|7610,7620|false|false|false|C0460137;C1579931|Depression - motion|depression
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7622,7626|false|false|false|C0038436;C0878676|6-pyruvoyl-tetrahydropterin synthase deficiency;Post-Traumatic Stress Disorder|PTSD
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|7622,7626|false|false|false|C0038436;C0878676|6-pyruvoyl-tetrahydropterin synthase deficiency;Post-Traumatic Stress Disorder|PTSD
Event|Event|SIMPLE_SEGMENT|7622,7626|false|false|false|||PTSD
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|7632,7649|false|false|false|C0855228|Eating disorder symptom|disordered eating
Event|Event|SIMPLE_SEGMENT|7643,7649|false|false|false|||eating
Finding|Organism Function|SIMPLE_SEGMENT|7643,7649|false|false|false|C0013470|Eating|eating
Event|Event|SIMPLE_SEGMENT|7654,7663|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|7654,7663|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|7654,7663|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|7654,7663|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|7654,7663|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7664,7673|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7664,7673|false|false|false|C0012634|Disease|Condition
Event|Event|SIMPLE_SEGMENT|7664,7673|false|false|false|||Condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|7664,7673|false|false|false|C1705253|Logical Condition|Condition
Finding|Mental Process|SIMPLE_SEGMENT|7675,7681|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7675,7688|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|SIMPLE_SEGMENT|7675,7688|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7682,7688|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|7682,7688|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|7690,7695|false|false|false|||Clear
Finding|Idea or Concept|SIMPLE_SEGMENT|7690,7695|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|SIMPLE_SEGMENT|7700,7708|false|false|false|||coherent
Finding|Finding|SIMPLE_SEGMENT|7700,7708|false|false|false|C4068804|Coherent|coherent
Event|Event|SIMPLE_SEGMENT|7710,7715|false|false|false|||Level
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7710,7732|false|false|false|C4050479||Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|7710,7732|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|SIMPLE_SEGMENT|7719,7732|false|false|false|||Consciousness
Finding|Finding|SIMPLE_SEGMENT|7719,7732|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|SIMPLE_SEGMENT|7719,7732|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7734,7739|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|7734,7739|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7734,7739|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|SIMPLE_SEGMENT|7734,7739|false|false|false|||Alert
Finding|Finding|SIMPLE_SEGMENT|7734,7739|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|7734,7739|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|7734,7739|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|SIMPLE_SEGMENT|7744,7755|false|false|false|||interactive
Finding|Functional Concept|SIMPLE_SEGMENT|7744,7755|false|false|false|C1704675|Interaction|interactive
Event|Activity|SIMPLE_SEGMENT|7757,7765|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|7757,7765|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|SIMPLE_SEGMENT|7757,7765|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7766,7772|false|false|false|C5889824||Status
Event|Event|SIMPLE_SEGMENT|7766,7772|false|false|false|||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|7766,7772|false|false|false|C1546481|What subject filter - Status|Status
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7781,7784|false|false|false|C3159311|BORNHOLM EYE DISEASE|Bed
Event|Event|SIMPLE_SEGMENT|7781,7784|false|false|false|||Bed
Finding|Intellectual Product|SIMPLE_SEGMENT|7781,7784|false|false|false|C2346952|Bachelor of Education|Bed
Event|Event|SIMPLE_SEGMENT|7790,7800|false|false|false|||assistance
Finding|Social Behavior|SIMPLE_SEGMENT|7790,7800|false|false|false|C0018896|Helping Behavior|assistance
Event|Event|SIMPLE_SEGMENT|7814,7824|false|false|false|||wheelchair
Finding|Finding|SIMPLE_SEGMENT|7814,7824|false|false|false|C2135586;C4321408|Wheelchair Usually Used;has wheelchair at home (history)|wheelchair
Event|Event|SIMPLE_SEGMENT|7829,7838|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|7829,7838|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|7829,7838|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|7829,7838|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|7829,7838|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7829,7851|false|false|false|C3669312||Discharge Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|7829,7851|false|false|false|C4282220|Discharge instructions|Discharge Instructions
Procedure|Health Care Activity|SIMPLE_SEGMENT|7829,7851|false|false|false|C2266673|hospital discharge instructions (treatment)|Discharge Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7839,7851|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|7839,7851|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|7839,7851|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Finding|Gene or Genome|SIMPLE_SEGMENT|7853,7857|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Event|Event|SIMPLE_SEGMENT|7877,7886|false|false|false|||privilege
Finding|Conceptual Entity|SIMPLE_SEGMENT|7877,7886|false|false|false|C1547898;C1706335;C1706336|Privilege;Role Privilege;User Privilege|privilege
Finding|Idea or Concept|SIMPLE_SEGMENT|7877,7886|false|false|false|C1547898;C1706335;C1706336|Privilege;Role Privilege;User Privilege|privilege
Event|Activity|SIMPLE_SEGMENT|7894,7898|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|7894,7898|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|7894,7898|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|7894,7898|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|7894,7901|false|false|false|C1555558|care of - AddressPartType|care of
Event|Event|SIMPLE_SEGMENT|7926,7929|false|false|false|||WAS
Event|Event|SIMPLE_SEGMENT|7932,7940|false|false|false|||ADMITTED
Event|Event|SIMPLE_SEGMENT|7948,7956|false|false|false|||HOSPITAL
Finding|Idea or Concept|SIMPLE_SEGMENT|7948,7956|false|false|false|C1547192|Organization unit type - Hospital|HOSPITAL
Event|Event|SIMPLE_SEGMENT|7999,8003|false|false|false|||came
Finding|Idea or Concept|SIMPLE_SEGMENT|8011,8019|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|SIMPLE_SEGMENT|8044,8051|false|false|false|||trouble
Event|Event|SIMPLE_SEGMENT|8064,8072|false|false|false|||speaking
Finding|Individual Behavior|SIMPLE_SEGMENT|8064,8072|false|false|false|C0234856|Speaking (function)|speaking
Event|Activity|SIMPLE_SEGMENT|8081,8089|false|false|false|C1709305|Occur (action)|HAPPENED
Event|Event|SIMPLE_SEGMENT|8098,8101|false|false|false|||WAS
Finding|Idea or Concept|SIMPLE_SEGMENT|8109,8117|false|false|false|C1547192|Organization unit type - Hospital|HOSPITAL
Event|Event|SIMPLE_SEGMENT|8172,8176|false|false|false|||seen
Event|Event|SIMPLE_SEGMENT|8201,8210|false|false|false|||diagnosed
Finding|Conceptual Entity|SIMPLE_SEGMENT|8221,8231|false|false|false|C0205245;C0542341;C2700217|Function (attribute);Functional;Functional Relationship|functional
Finding|Functional Concept|SIMPLE_SEGMENT|8221,8231|false|false|false|C0205245;C0542341;C2700217|Function (attribute);Functional;Functional Relationship|functional
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|8221,8253|false|false|false|C0009946;C4543816|Conversion disorder;Dissociative neurological symptom disorder (disorder)|functional neurological disorder
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8232,8253|false|false|false|C0027765|nervous system disorder|neurological disorder
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8245,8253|false|false|false|C0012634|Disease|disorder
Event|Event|SIMPLE_SEGMENT|8245,8253|false|false|false|||disorder
Event|Event|SIMPLE_SEGMENT|8261,8267|false|false|false|||worked
Event|Event|SIMPLE_SEGMENT|8273,8281|false|false|false|||physical
Finding|Finding|SIMPLE_SEGMENT|8273,8281|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Finding|Functional Concept|SIMPLE_SEGMENT|8273,8281|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|8273,8281|false|false|false|C0031809|Physical Examination|physical
Finding|Functional Concept|SIMPLE_SEGMENT|8286,8298|false|false|false|C0521127|Occupational|occupational
Event|Event|SIMPLE_SEGMENT|8299,8309|false|false|false|||therapists
Event|Event|SIMPLE_SEGMENT|8317,8325|false|false|false|||symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|8317,8325|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|8317,8325|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|SIMPLE_SEGMENT|8326,8331|false|false|false|||began
Event|Event|SIMPLE_SEGMENT|8335,8342|false|false|false|||improve
Event|Event|SIMPLE_SEGMENT|8350,8356|false|false|false|||SHOULD
Event|Event|SIMPLE_SEGMENT|8380,8388|false|false|false|||HOSPITAL
Finding|Idea or Concept|SIMPLE_SEGMENT|8380,8388|false|false|false|C1547192|Organization unit type - Hospital|HOSPITAL
Event|Event|SIMPLE_SEGMENT|8446,8454|false|false|false|||continue
Event|Event|SIMPLE_SEGMENT|8458,8462|false|false|false|||take
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8472,8483|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8472,8483|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|8472,8483|false|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|8472,8483|false|false|false|C4284232|Medications|medications
Event|Event|SIMPLE_SEGMENT|8488,8494|false|false|false|||follow
Event|Event|SIMPLE_SEGMENT|8509,8516|false|false|false|||doctors
Event|Activity|SIMPLE_SEGMENT|8529,8541|false|false|false|C0003629|Appointments|appointments
Event|Event|SIMPLE_SEGMENT|8529,8541|false|false|false|||appointments
Event|Event|SIMPLE_SEGMENT|8554,8562|false|false|false|||continue
Event|Event|SIMPLE_SEGMENT|8566,8570|false|false|false|||work
Event|Event|SIMPLE_SEGMENT|8581,8589|false|false|false|||physical
Finding|Finding|SIMPLE_SEGMENT|8581,8589|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Finding|Functional Concept|SIMPLE_SEGMENT|8581,8589|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|8581,8589|false|false|false|C0031809|Physical Examination|physical
Event|Event|SIMPLE_SEGMENT|8594,8606|false|false|false|||occupational
Finding|Functional Concept|SIMPLE_SEGMENT|8594,8606|false|false|false|C0521127|Occupational|occupational
Event|Event|SIMPLE_SEGMENT|8608,8618|false|false|false|||therapists
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8641,8645|false|false|false|C0339510|Vitelliform Macular Dystrophy|best
Event|Event|SIMPLE_SEGMENT|8641,8645|false|false|false|||best
Finding|Gene or Genome|SIMPLE_SEGMENT|8641,8645|false|false|false|C1826421;C5781213|BEST1 gene;BEST1 wt Allele|best
Event|Activity|SIMPLE_SEGMENT|8671,8675|false|false|false|C1947933|care activity|Care
Finding|Finding|SIMPLE_SEGMENT|8671,8675|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|SIMPLE_SEGMENT|8671,8675|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8671,8680|false|false|false|C4321316||Care Team
Finding|Finding|SIMPLE_SEGMENT|8671,8680|false|false|false|C4321315|Care team|Care Team
Procedure|Health Care Activity|SIMPLE_SEGMENT|8685,8693|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8694,8706|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|8694,8706|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|8694,8706|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

