 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|42,51|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|42,51|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|42,56|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|76,85|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|76,85|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|76,85|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|76,85|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|76,85|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|76,90|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|108,113|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|108,113|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|108,113|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|132,135|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|143,150|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|143,150|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|152,160|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Drug|Indicator, Reagent, or Diagnostic Aid|Allergies|178,181|false|false|false|C0013343|Dyes|Dye
Event|Event|Allergies|178,181|false|false|false|||Dye
Drug|Biologically Active Substance|Allergies|183,189|false|false|false|C0021968;C0885449|Iodine, Homeopathic preparation;iodine|Iodine
Drug|Element, Ion, or Isotope|Allergies|183,189|false|false|false|C0021968;C0885449|Iodine, Homeopathic preparation;iodine|Iodine
Drug|Pharmacologic Substance|Allergies|183,189|false|false|false|C0021968;C0885449|Iodine, Homeopathic preparation;iodine|Iodine
Event|Activity|Allergies|190,200|false|false|false|C2700400|Contain (action)|Containing
Finding|Functional Concept|Allergies|190,200|false|false|false|C0332256|Containing (qualifier value)|Containing
Drug|Indicator, Reagent, or Diagnostic Aid|Allergies|201,209|false|false|false|C0009924|Contrast Media|Contrast
Drug|Indicator, Reagent, or Diagnostic Aid|Allergies|201,215|false|false|false|C0009924|Contrast Media|Contrast Media
Anatomy|Tissue|Allergies|210,215|false|false|false|C0162867;C1254021|Media layer;Tunica Media|Media
Finding|Intellectual Product|Allergies|210,215|false|false|false|C0009458;C0677540|Communications Media;PAMS Media|Media
Drug|Organic Chemical|Allergies|218,227|false|false|false|C0030049|oxycodone|Oxycodone
Drug|Pharmacologic Substance|Allergies|218,227|false|false|false|C0030049|oxycodone|Oxycodone
Event|Event|Allergies|218,227|false|false|false|||Oxycodone
Procedure|Laboratory Procedure|Allergies|218,227|false|false|false|C0524222|Oxycodone measurement|Oxycodone
Drug|Organic Chemical|Allergies|231,241|false|false|false|C0055729|cilostazol|cilostazol
Drug|Pharmacologic Substance|Allergies|231,241|false|false|false|C0055729|cilostazol|cilostazol
Event|Event|Allergies|231,241|false|false|false|||cilostazol
Drug|Organic Chemical|Allergies|244,255|false|false|false|C1569608|varenicline|Varenicline
Drug|Pharmacologic Substance|Allergies|244,255|false|false|false|C1569608|varenicline|Varenicline
Event|Event|Allergies|244,255|false|false|false|||Varenicline
Event|Event|Allergies|258,267|false|false|false|||Attending
Finding|Functional Concept|Allergies|258,267|false|false|false|C1999232|Attending (action)|Attending
Anatomy|Body Location or Region|Chief Complaint|307,312|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|Chief Complaint|307,312|false|false|false|C0741025|Chest problem|Chest
Attribute|Clinical Attribute|Chief Complaint|307,317|false|false|false|C2926613||Chest pain
Finding|Sign or Symptom|Chief Complaint|307,317|false|false|false|C0008031|Chest Pain|Chest pain
Attribute|Clinical Attribute|Chief Complaint|313,317|false|true|false|C2598155||pain
Event|Event|Chief Complaint|313,317|false|false|false|||pain
Finding|Functional Concept|Chief Complaint|313,317|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Chief Complaint|313,317|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Classification|Chief Complaint|320,325|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|326,334|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|326,334|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|338,356|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|347,356|false|false|false|C0945766||Procedure
Event|Event|Chief Complaint|347,356|false|false|false|||Procedure
Event|Occupational Activity|Chief Complaint|347,356|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|347,356|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|347,356|false|false|false|C0184661|Interventional procedure|Procedure
Finding|Idea or Concept|History of Present Illness|408,412|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|History of Present Illness|408,412|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Event|Event|History of Present Illness|413,416|false|false|false|||old
Disorder|Disease or Syndrome|History of Present Illness|434,437|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|434,437|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|History of Present Illness|434,437|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|History of Present Illness|434,437|false|false|false|||CAD
Finding|Gene or Genome|History of Present Illness|434,437|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|History of Present Illness|434,437|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|History of Present Illness|434,437|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|434,437|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Disorder|Disease or Syndrome|History of Present Illness|439,442|false|false|false|C0085096|Peripheral Vascular Diseases|PVD
Event|Event|History of Present Illness|439,442|false|false|false|||PVD
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|439,442|false|false|false|C4521226|Pomalidomide/Bortezomib/Dexamethasone Regimen|PVD
Disorder|Disease or Syndrome|History of Present Illness|447,451|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|History of Present Illness|447,451|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|History of Present Illness|447,451|false|false|false|||COPD
Finding|Gene or Genome|History of Present Illness|447,451|false|false|false|C1412502|ARCN1 gene|COPD
Event|Event|History of Present Illness|453,463|false|false|false|||presenting
Anatomy|Body Location or Region|History of Present Illness|469,474|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|469,474|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|History of Present Illness|469,479|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|History of Present Illness|469,479|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|History of Present Illness|475,479|false|false|false|C2598155||pain
Event|Event|History of Present Illness|475,479|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|475,479|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|475,479|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|History of Present Illness|485,492|false|false|false|||reports
Event|Event|History of Present Illness|502,506|false|false|false|||woke
Event|Event|History of Present Illness|535,543|false|false|false|||pressure
Finding|Finding|History of Present Illness|535,543|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|History of Present Illness|535,543|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|History of Present Illness|535,543|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|History of Present Illness|535,543|false|false|false|C0033095||pressure
Attribute|Clinical Attribute|History of Present Illness|549,553|false|false|false|C2598155||pain
Event|Event|History of Present Illness|549,553|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|549,553|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|549,553|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|History of Present Illness|581,590|false|false|false|||shortness
Attribute|Clinical Attribute|History of Present Illness|581,600|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|History of Present Illness|581,600|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|History of Present Illness|594,600|false|false|false|C0225386|Breath|breath
Event|Event|History of Present Illness|606,611|false|false|false|||rated
Attribute|Clinical Attribute|History of Present Illness|616,620|false|false|false|C2598155||pain
Event|Event|History of Present Illness|616,620|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|616,620|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|616,620|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|History of Present Illness|631,638|false|false|false|||reports
Finding|Intellectual Product|History of Present Illness|631,638|false|false|false|C0684224|Report (document)|reports
Procedure|Health Care Activity|History of Present Illness|631,638|false|false|false|C0700287|Reporting|reports
Event|Event|History of Present Illness|648,654|false|false|false|||lasted
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|665,674|false|false|false|C0886384|5 minutes Office visit|5 minutes
Event|Event|History of Present Illness|667,674|false|false|false|||minutes
Event|Event|History of Present Illness|679,687|false|false|false|||resolved
Event|Event|History of Present Illness|725,733|false|false|false|||episodes
Attribute|Clinical Attribute|History of Present Illness|746,750|false|false|false|C2598155||pain
Event|Event|History of Present Illness|746,750|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|746,750|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|746,750|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|History of Present Illness|751,758|false|false|false|||lasting
Event|Event|History of Present Illness|768,775|false|false|false|||minutes
Finding|Finding|History of Present Illness|781,785|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|History of Present Illness|781,785|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|History of Present Illness|781,785|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Finding|History of Present Illness|824,828|false|false|false|C4281574|Much|much
Event|Event|History of Present Illness|835,841|false|false|false|||severe
Finding|Finding|History of Present Illness|835,841|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|History of Present Illness|835,841|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Event|Event|History of Present Illness|861,868|true|false|false|||episode
Attribute|Clinical Attribute|History of Present Illness|872,876|true|false|false|C2598155||pain
Event|Event|History of Present Illness|872,876|true|false|false|||pain
Finding|Functional Concept|History of Present Illness|872,876|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|872,876|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|History of Present Illness|901,913|true|false|false|||palpitations
Finding|Finding|History of Present Illness|901,913|true|false|false|C0030252|Palpitations|palpitations
Event|Event|History of Present Illness|915,930|true|false|false|||lightheadedness
Finding|Sign or Symptom|History of Present Illness|915,930|true|false|false|C0220870|Lightheadedness|lightheadedness
Event|Event|History of Present Illness|932,941|true|false|false|||dizziness
Finding|Sign or Symptom|History of Present Illness|932,941|true|false|false|C0012833;C0042571|Dizziness;Vertigo|dizziness
Attribute|Clinical Attribute|History of Present Illness|943,949|true|false|false|C4255480||nausea
Event|Event|History of Present Illness|943,949|true|false|false|||nausea
Finding|Sign or Symptom|History of Present Illness|943,949|true|false|false|C0027497|Nausea|nausea
Event|Event|History of Present Illness|952,960|false|false|false|||vomiting
Finding|Sign or Symptom|History of Present Illness|952,960|false|false|false|C0042963|Vomiting|vomiting
Event|Event|History of Present Illness|962,973|false|false|false|||diaphoresis
Finding|Finding|History of Present Illness|962,973|false|false|false|C0700590|Increased sweating|diaphoresis
Finding|Idea or Concept|History of Present Illness|988,995|false|false|false|C1555582|Initial (abbreviation)|initial
Event|Event|History of Present Illness|996,1002|false|false|false|||vitals
Event|Event|History of Present Illness|1035,1039|false|false|false|||Labs
Lab|Laboratory or Test Result|History of Present Illness|1035,1039|false|false|false|C0587081|Laboratory test finding|Labs
Event|Event|History of Present Illness|1045,1056|false|false|false|||significant
Finding|Idea or Concept|History of Present Illness|1045,1056|false|false|false|C0750502|Significant|significant
Drug|Biologically Active Substance|History of Present Illness|1085,1088|false|false|false|C0007012|carbon dioxide|CO2
Drug|Inorganic Chemical|History of Present Illness|1085,1088|false|false|false|C0007012|carbon dioxide|CO2
Event|Event|History of Present Illness|1085,1088|false|false|false|||CO2
Finding|Finding|History of Present Illness|1085,1088|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Finding|Gene or Genome|History of Present Illness|1085,1088|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Drug|Biologically Active Substance|History of Present Illness|1092,1095|false|false|false|C0600137|Blood Urea Nitrogen|BUN
Drug|Inorganic Chemical|History of Present Illness|1092,1095|false|false|false|C0600137|Blood Urea Nitrogen|BUN
Event|Event|History of Present Illness|1092,1095|false|false|false|||BUN
Procedure|Laboratory Procedure|History of Present Illness|1092,1095|false|false|false|C0005845|Blood urea nitrogen measurement|BUN
Anatomy|Cell|History of Present Illness|1138,1141|false|false|false|C0023516|Leukocytes|WBC
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1146,1149|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|History of Present Illness|1146,1149|false|false|false|C0019046|Hemoglobin|Hgb
Event|Event|History of Present Illness|1146,1149|false|false|false|||Hgb
Finding|Gene or Genome|History of Present Illness|1146,1149|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|History of Present Illness|1146,1149|false|false|false|C0019029|Hemoglobin concentration|Hgb
Event|Event|History of Present Illness|1155,1158|false|false|false|||Hct
Procedure|Laboratory Procedure|History of Present Illness|1155,1158|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1155,1158|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Event|Event|History of Present Illness|1164,1167|false|false|false|||Plt
Procedure|Laboratory Procedure|History of Present Illness|1164,1167|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Neoplastic Process|History of Present Illness|1186,1189|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|History of Present Illness|1186,1189|false|false|false|||PTT
Procedure|Laboratory Procedure|History of Present Illness|1186,1189|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Attribute|Clinical Attribute|History of Present Illness|1196,1199|false|false|false|C0368980|Coagulation tissue factor induced.INR|INR
Event|Event|History of Present Illness|1196,1199|false|false|false|||INR
Procedure|Laboratory Procedure|History of Present Illness|1196,1199|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1196,1199|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Drug|Organic Chemical|History of Present Illness|1209,1216|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Drug|Pharmacologic Substance|History of Present Illness|1209,1216|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Event|Event|History of Present Illness|1209,1216|false|false|false|||Lactate
Procedure|Laboratory Procedure|History of Present Illness|1209,1216|false|false|false|C0202115|Lactic acid measurement|Lactate
Event|Event|History of Present Illness|1243,1250|false|false|false|||Imaging
Finding|Finding|History of Present Illness|1243,1250|false|false|false|C0740845|Imaging problem|Imaging
Procedure|Diagnostic Procedure|History of Present Illness|1243,1250|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|Imaging
Event|Event|History of Present Illness|1251,1259|false|false|false|||revealed
Event|Event|History of Present Illness|1265,1268|false|false|false|||CXR
Procedure|Diagnostic Procedure|History of Present Illness|1265,1268|false|false|false|C0039985|Plain chest X-ray|CXR
Finding|Intellectual Product|History of Present Illness|1273,1278|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Anatomy|Body Location or Region|History of Present Illness|1279,1294|true|false|false|C0553534|Cardiopulmonary|cardiopulmonary
Disorder|Disease or Syndrome|History of Present Illness|1279,1294|true|false|false|C4072686|Cardiovascular disease+Pulmonary disease|cardiopulmonary
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1295,1302|true|false|false|C1184743|bony process|process
Drug|Pharmacologic Substance|History of Present Illness|1295,1302|true|false|false|C1951340|Process Pharmacologic Substance|process
Event|Event|History of Present Illness|1295,1302|true|false|false|||process
Finding|Functional Concept|History of Present Illness|1295,1302|true|false|false|C4521054|Process (qualifier value)|process
Phenomenon|Phenomenon or Process|History of Present Illness|1295,1302|true|false|false|C1522240|Process|process
Finding|Body Substance|History of Present Illness|1311,1318|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|1311,1318|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|1311,1318|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Organic Chemical|History of Present Illness|1333,1340|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|History of Present Illness|1333,1340|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|History of Present Illness|1349,1358|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|History of Present Illness|1349,1358|false|false|false|C0001927|albuterol|Albuterol
Event|Event|History of Present Illness|1349,1358|false|false|false|||Albuterol
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1367,1370|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biologically Active Substance|History of Present Illness|1367,1370|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biomedical or Dental Material|History of Present Illness|1367,1370|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Finding|Cell Function|History of Present Illness|1367,1370|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Finding|Gene or Genome|History of Present Illness|1367,1370|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Drug|Organic Chemical|History of Present Illness|1375,1386|false|false|false|C0027235|ipratropium|Ipratropium
Drug|Pharmacologic Substance|History of Present Illness|1375,1386|false|false|false|C0027235|ipratropium|Ipratropium
Event|Event|History of Present Illness|1375,1386|false|false|false|||Ipratropium
Drug|Organic Chemical|History of Present Illness|1375,1394|false|false|false|C0700580|ipratropium bromide|Ipratropium Bromide
Drug|Pharmacologic Substance|History of Present Illness|1375,1394|false|false|false|C0700580|ipratropium bromide|Ipratropium Bromide
Drug|Inorganic Chemical|History of Present Illness|1387,1394|false|false|false|C0006222|Bromides|Bromide
Procedure|Laboratory Procedure|History of Present Illness|1387,1394|false|false|false|C0202341|Bromides measurement|Bromide
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1395,1398|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biologically Active Substance|History of Present Illness|1395,1398|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biomedical or Dental Material|History of Present Illness|1395,1398|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Event|Event|History of Present Illness|1395,1398|false|false|false|||Neb
Finding|Cell Function|History of Present Illness|1395,1398|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Finding|Gene or Genome|History of Present Illness|1395,1398|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Drug|Biologically Active Substance|History of Present Illness|1403,1412|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Element, Ion, or Isotope|History of Present Illness|1403,1412|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Food|History of Present Illness|1403,1412|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Inorganic Chemical|History of Present Illness|1403,1412|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Pharmacologic Substance|History of Present Illness|1403,1412|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Event|Event|History of Present Illness|1403,1412|false|false|false|||Potassium
Finding|Physiologic Function|History of Present Illness|1403,1412|false|false|false|C4553027|Potassium metabolic function|Potassium
Procedure|Laboratory Procedure|History of Present Illness|1403,1412|false|false|false|C0202194|Potassium measurement|Potassium
Drug|Inorganic Chemical|History of Present Illness|1403,1421|false|false|false|C0032825|potassium chloride|Potassium Chloride
Drug|Pharmacologic Substance|History of Present Illness|1403,1421|false|false|false|C0032825|potassium chloride|Potassium Chloride
Drug|Element, Ion, or Isotope|History of Present Illness|1413,1421|false|false|false|C0008203;C0596019|Chlorides;chloride ion|Chloride
Event|Event|History of Present Illness|1413,1421|false|false|false|||Chloride
Finding|Physiologic Function|History of Present Illness|1413,1421|false|false|false|C4553021|Chloride metabolic function|Chloride
Procedure|Laboratory Procedure|History of Present Illness|1413,1421|false|false|false|C0201952|Chloride measurement|Chloride
Drug|Biologically Active Substance|History of Present Illness|1438,1447|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Element, Ion, or Isotope|History of Present Illness|1438,1447|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Food|History of Present Illness|1438,1447|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Inorganic Chemical|History of Present Illness|1438,1447|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Pharmacologic Substance|History of Present Illness|1438,1447|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Event|Event|History of Present Illness|1438,1447|false|false|false|||Potassium
Finding|Physiologic Function|History of Present Illness|1438,1447|false|false|false|C4553027|Potassium metabolic function|Potassium
Procedure|Laboratory Procedure|History of Present Illness|1438,1447|false|false|false|C0202194|Potassium measurement|Potassium
Drug|Inorganic Chemical|History of Present Illness|1438,1456|false|false|false|C0032825|potassium chloride|Potassium Chloride
Drug|Pharmacologic Substance|History of Present Illness|1438,1456|false|false|false|C0032825|potassium chloride|Potassium Chloride
Drug|Element, Ion, or Isotope|History of Present Illness|1448,1456|false|false|false|C0008203;C0596019|Chlorides;chloride ion|Chloride
Event|Event|History of Present Illness|1448,1456|false|false|false|||Chloride
Finding|Physiologic Function|History of Present Illness|1448,1456|false|false|false|C4553021|Chloride metabolic function|Chloride
Procedure|Laboratory Procedure|History of Present Illness|1448,1456|false|false|false|C0201952|Chloride measurement|Chloride
Event|Event|History of Present Illness|1467,1469|false|false|false|||NS
Event|Event|History of Present Illness|1490,1498|false|false|false|||transfer
Finding|Functional Concept|History of Present Illness|1490,1498|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|History of Present Illness|1490,1498|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|History of Present Illness|1490,1498|false|false|false|C4706767|Transfer (immobility management)|transfer
Event|Activity|History of Present Illness|1539,1546|true|false|false|C1706079||arrival
Event|Event|History of Present Illness|1539,1546|true|false|false|||arrival
Finding|Functional Concept|History of Present Illness|1539,1546|true|false|false|C1555577|arrival - ActRelationshipType|arrival
Anatomy|Anatomical Structure|History of Present Illness|1554,1559|true|false|false|C3714591|Floor (anatomic)|floor
Finding|Body Substance|History of Present Illness|1561,1568|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|1561,1568|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|1561,1568|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|1569,1575|false|false|false|||denies
Anatomy|Body Location or Region|History of Present Illness|1576,1581|true|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|1576,1581|true|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|History of Present Illness|1576,1586|true|false|false|C2926613||chest pain
Finding|Sign or Symptom|History of Present Illness|1576,1586|true|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|History of Present Illness|1582,1586|true|false|false|C2598155||pain
Event|Event|History of Present Illness|1582,1586|true|false|false|||pain
Finding|Functional Concept|History of Present Illness|1582,1586|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1582,1586|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|History of Present Illness|1588,1597|true|false|false|||shortness
Finding|Body Substance|History of Present Illness|1602,1608|true|false|false|C0225386|Breath|breath
Event|Event|History of Present Illness|1610,1622|false|false|false|||palpitations
Finding|Finding|History of Present Illness|1610,1622|false|false|false|C0030252|Palpitations|palpitations
Event|Event|History of Present Illness|1624,1639|false|false|false|||lightheadedness
Finding|Sign or Symptom|History of Present Illness|1624,1639|false|false|false|C0220870|Lightheadedness|lightheadedness
Event|Event|History of Present Illness|1641,1650|false|false|false|||dizziness
Finding|Sign or Symptom|History of Present Illness|1641,1650|false|false|false|C0012833;C0042571|Dizziness;Vertigo|dizziness
Event|Event|History of Present Illness|1654,1660|false|false|false|||REVIEW
Finding|Idea or Concept|History of Present Illness|1654,1660|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|REVIEW
Finding|Intellectual Product|History of Present Illness|1654,1660|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|REVIEW
Finding|Functional Concept|History of Present Illness|1654,1663|false|false|false|C0699752|Review of|REVIEW OF
Attribute|Clinical Attribute|History of Present Illness|1654,1671|false|false|false|C0488564;C0488565||REVIEW OF SYSTEMS
Procedure|Health Care Activity|History of Present Illness|1654,1671|false|false|false|C0489633|Review of systems (procedure)|REVIEW OF SYSTEMS
Event|Event|History of Present Illness|1664,1671|false|false|false|||SYSTEMS
Finding|Functional Concept|History of Present Illness|1664,1671|false|false|false|C0449913|System|SYSTEMS
Disorder|Disease or Syndrome|History of Present Illness|1683,1686|false|false|false|C0268529|Proline dehydrogenase deficiency|HPI
Event|Event|History of Present Illness|1683,1686|false|false|false|||HPI
Finding|Finding|History of Present Illness|1683,1686|false|false|false|C0262512;C1323983|History of present illness (finding);allene oxide synthase activity|HPI
Finding|Molecular Function|History of Present Illness|1683,1686|false|false|false|C0262512;C1323983|History of present illness (finding);allene oxide synthase activity|HPI
Disorder|Disease or Syndrome|Past Medical History|1714,1720|false|false|false|C0004096|Asthma|ASTHMA
Event|Event|Past Medical History|1714,1720|false|false|false|||ASTHMA
Disorder|Disease or Syndrome|Past Medical History|1721,1725|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Past Medical History|1721,1725|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Past Medical History|1721,1725|false|false|false|||COPD
Finding|Gene or Genome|Past Medical History|1721,1725|false|false|false|C1412502|ARCN1 gene|COPD
Drug|Hazardous or Poisonous Substance|Past Medical History|1726,1733|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|Tobacco
Drug|Immunologic Factor|Past Medical History|1726,1733|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|Tobacco
Drug|Organic Chemical|Past Medical History|1726,1733|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|Tobacco
Drug|Pharmacologic Substance|Past Medical History|1726,1733|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|Tobacco
Attribute|Clinical Attribute|Past Medical History|1726,1737|false|false|false|C4522050||Tobacco use
Finding|Finding|Past Medical History|1726,1737|false|false|false|C0040335;C0543414;C0841002;C3853727|Encounter due to tobacco use;History of tobacco use;Tobacco use;Tobacco user|Tobacco use
Finding|Individual Behavior|Past Medical History|1726,1737|false|false|false|C0040335;C0543414;C0841002;C3853727|Encounter due to tobacco use;History of tobacco use;Tobacco use;Tobacco user|Tobacco use
Event|Event|Past Medical History|1734,1737|false|false|false|||use
Finding|Functional Concept|Past Medical History|1734,1737|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|Past Medical History|1734,1737|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Disorder|Disease or Syndrome|Past Medical History|1739,1766|false|false|false|C0085096;C1704436|Peripheral Arterial Diseases;Peripheral Vascular Diseases|Peripheral Arterial disease
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1750,1758|false|false|false|C0003842|Arteries|Arterial
Disorder|Disease or Syndrome|Past Medical History|1750,1766|false|false|false|C0852949|Arteriopathic disease|Arterial disease
Disorder|Disease or Syndrome|Past Medical History|1759,1766|false|false|false|C0012634|Disease|disease
Event|Event|Past Medical History|1759,1766|false|false|false|||disease
Finding|Functional Concept|Past Medical History|1779,1785|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Finding|Intellectual Product|Past Medical History|1779,1785|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1786,1791|false|false|false|C0020889|Bone structure of ilium|iliac
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1786,1800|false|false|false|C0850459|iliac stents|iliac stenting
Event|Event|Past Medical History|1792,1800|false|false|false|||stenting
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1792,1800|false|false|false|C2348535|Stenting|stenting
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1802,1808|false|false|false|C0018792|Heart Atrium|ATRIAL
Disorder|Disease or Syndrome|Past Medical History|1802,1820|false|false|false|C0546959|Atrial tachycardia|ATRIAL TACHYCARDIA
Finding|Finding|Past Medical History|1802,1820|false|false|false|C2059391|continuous electrocardiogram atrial tachycardia|ATRIAL TACHYCARDIA
Event|Event|Past Medical History|1809,1820|false|false|false|||TACHYCARDIA
Finding|Finding|Past Medical History|1809,1820|false|false|false|C0039231;C3827868|Tachycardia;Tachycardia by ECG Finding|TACHYCARDIA
Finding|Finding|Past Medical History|1822,1830|false|false|false|C0741302|atypia morphology|ATYPICAL
Finding|Sign or Symptom|Past Medical History|1822,1841|false|false|false|C0262384|Atypical chest pain|ATYPICAL CHEST PAIN
Anatomy|Body Location or Region|Past Medical History|1831,1836|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|CHEST
Finding|Finding|Past Medical History|1831,1836|false|false|false|C0741025|Chest problem|CHEST
Attribute|Clinical Attribute|Past Medical History|1831,1841|false|true|false|C2926613||CHEST PAIN
Finding|Sign or Symptom|Past Medical History|1831,1841|false|true|false|C0008031|Chest Pain|CHEST PAIN
Attribute|Clinical Attribute|Past Medical History|1837,1841|false|true|false|C2598155||PAIN
Event|Event|Past Medical History|1837,1841|false|false|false|||PAIN
Finding|Functional Concept|Past Medical History|1837,1841|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|PAIN
Finding|Sign or Symptom|Past Medical History|1837,1841|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|PAIN
Anatomy|Body Location or Region|Past Medical History|1844,1852|false|false|false|C0027530|Neck|CERVICAL
Disorder|Disease or Syndrome|Past Medical History|1844,1864|false|false|false|C0263884|Cervical radiculitis|CERVICAL RADICULITIS
Disorder|Disease or Syndrome|Past Medical History|1853,1864|false|false|false|C0034544|Radiculitis|RADICULITIS
Event|Event|Past Medical History|1853,1864|false|false|false|||RADICULITIS
Anatomy|Body Location or Region|Past Medical History|1866,1874|false|false|false|C0027530|Neck|CERVICAL
Disorder|Disease or Syndrome|Past Medical History|1866,1886|false|false|false|C0158241;C1384641|Cervical spondylosis;Cervical spondylosis without myelopathy|CERVICAL SPONDYLOSIS
Disorder|Disease or Syndrome|Past Medical History|1875,1886|false|false|false|C0038019|Spondylosis|SPONDYLOSIS
Event|Event|Past Medical History|1875,1886|false|false|false|||SPONDYLOSIS
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1888,1896|false|false|false|C0018787|Heart|CORONARY
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1888,1903|false|false|false|C0205042|Coronary artery|CORONARY ARTERY
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1897,1903|false|false|false|C0003842;C0226004|Arterial system;Arteries|ARTERY
Anatomy|Body System|Past Medical History|1897,1903|false|false|false|C0003842;C0226004|Arterial system;Arteries|ARTERY
Disorder|Disease or Syndrome|Past Medical History|1905,1912|false|false|false|C0012634|Disease|DISEASE
Event|Event|Past Medical History|1905,1912|false|false|false|||DISEASE
Event|Event|Past Medical History|1915,1923|false|false|false|||HEADACHE
Finding|Sign or Symptom|Past Medical History|1915,1923|false|false|false|C0018681|Headache|HEADACHE
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1925,1928|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|HIP
Drug|Amino Acid, Peptide, or Protein|Past Medical History|1925,1928|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|HIP
Drug|Biologically Active Substance|Past Medical History|1925,1928|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|HIP
Drug|Pharmacologic Substance|Past Medical History|1925,1928|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|HIP
Event|Event|Past Medical History|1925,1928|false|false|false|||HIP
Finding|Gene or Genome|Past Medical History|1925,1928|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|HIP
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1925,1928|false|false|false|C1292890|Procedure on hip|HIP
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1925,1940|false|false|false|C0392806|Prosthetic arthroplasty of hip (procedure)|HIP REPLACEMENT
Event|Event|Past Medical History|1929,1940|false|false|false|||REPLACEMENT
Finding|Functional Concept|Past Medical History|1929,1940|false|false|false|C0559956|Replacement|REPLACEMENT
Procedure|Health Care Activity|Past Medical History|1929,1940|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|REPLACEMENT
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1929,1940|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|REPLACEMENT
Disorder|Disease or Syndrome|Past Medical History|1942,1956|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|HYPERLIPIDEMIA
Event|Event|Past Medical History|1942,1956|false|false|false|||HYPERLIPIDEMIA
Finding|Finding|Past Medical History|1942,1956|false|false|false|C0428465|Serum lipids high (finding)|HYPERLIPIDEMIA
Disorder|Disease or Syndrome|Past Medical History|1958,1970|false|false|false|C0020538|Hypertensive disease|HYPERTENSION
Event|Event|Past Medical History|1958,1970|false|false|false|||HYPERTENSION
Disorder|Disease or Syndrome|Past Medical History|1973,1987|false|false|false|C0029408|Degenerative polyarthritis|OSTEOARTHRITIS
Disorder|Disease or Syndrome|Past Medical History|1989,1995|false|false|false|C0019340;C0854331|Herpes simplex dermatitis|HERPES
Disorder|Disease or Syndrome|Past Medical History|1989,2002|false|false|false|C0019360;C0042338|Herpes zoster (disorder);herpesvirus 3, human|HERPES ZOSTER
Disorder|Virus|Past Medical History|1989,2002|false|false|false|C0019360;C0042338|Herpes zoster (disorder);herpesvirus 3, human|HERPES ZOSTER
Disorder|Disease or Syndrome|Past Medical History|1996,2002|false|false|false|C0019360|Herpes zoster (disorder)|ZOSTER
Event|Event|Past Medical History|1996,2002|false|false|false|||ZOSTER
Drug|Hazardous or Poisonous Substance|Past Medical History|2004,2011|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|TOBACCO
Drug|Immunologic Factor|Past Medical History|2004,2011|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|TOBACCO
Drug|Organic Chemical|Past Medical History|2004,2011|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|TOBACCO
Drug|Pharmacologic Substance|Past Medical History|2004,2011|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|TOBACCO
Disorder|Mental or Behavioral Dysfunction|Past Medical History|2004,2017|false|false|false|C0040336|Tobacco Use Disorder|TOBACCO ABUSE
Disorder|Mental or Behavioral Dysfunction|Past Medical History|2012,2017|false|false|false|C0013146|Drug abuse|ABUSE
Event|Event|Past Medical History|2012,2017|false|false|false|||ABUSE
Event|Event|Past Medical History|2012,2017|false|false|false|C1546935|Abuse|ABUSE
Finding|Finding|Past Medical History|2012,2017|false|false|false|C0562381|Victim of abuse (finding)|ABUSE
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2019,2025|false|false|false|C0018792|Heart Atrium|ATRIAL
Disorder|Disease or Syndrome|Past Medical History|2027,2039|false|false|false|C0232197|Fibrillation|FIBRILLATION
Event|Event|Past Medical History|2027,2039|false|false|false|||FIBRILLATION
Disorder|Mental or Behavioral Dysfunction|Past Medical History|2042,2049|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|ANXIETY
Event|Event|Past Medical History|2042,2049|false|false|false|||ANXIETY
Finding|Sign or Symptom|Past Medical History|2042,2049|false|false|false|C0860603|Anxiety symptoms|ANXIETY
Finding|Intellectual Product|Past Medical History|2050,2066|false|false|false|C1314977|Gastrointestinal attachment|GASTROINTESTINAL
Finding|Pathologic Function|Past Medical History|2050,2075|false|false|false|C0017181|Gastrointestinal Hemorrhage|GASTROINTESTINAL BLEEDING
Event|Event|Past Medical History|2067,2075|false|false|false|||BLEEDING
Finding|Pathologic Function|Past Medical History|2067,2075|false|false|false|C0019080|Hemorrhage|BLEEDING
Disorder|Disease or Syndrome|Past Medical History|2077,2091|false|false|false|C0029408|Degenerative polyarthritis|OSTEOARTHRITIS
Event|Event|Past Medical History|2077,2091|false|false|false|||OSTEOARTHRITIS
Finding|Functional Concept|Past Medical History|2094,2109|false|false|false|C0333482|atherosclerotic|ATHEROSCLEROTIC
Disorder|Disease or Syndrome|Past Medical History|2094,2132|false|true|false|C0004153|Atherosclerosis|ATHEROSCLEROTIC CARDIOVASCULAR DISEASE
Anatomy|Body System|Past Medical History|2110,2124|false|false|false|C0007226;C3887460|Cardiovascular;Cardiovascular system|CARDIOVASCULAR
Disorder|Disease or Syndrome|Past Medical History|2110,2132|false|true|false|C0007222|Cardiovascular Diseases|CARDIOVASCULAR DISEASE
Disorder|Disease or Syndrome|Past Medical History|2125,2132|false|true|false|C0012634|Disease|DISEASE
Event|Event|Past Medical History|2125,2132|false|false|false|||DISEASE
Disorder|Disease or Syndrome|Past Medical History|2125,2153|false|false|false|C0085096|Peripheral Vascular Diseases|DISEASE, PERIPHERAL VASCULAR
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2145,2153|false|false|false|C0005847|Blood Vessel|VASCULAR
Disorder|Disease or Syndrome|Past Medical History|2155,2162|false|false|false|C0012634|Disease|DISEASE
Event|Event|Past Medical History|2155,2162|false|false|false|||DISEASE
Disorder|Disease or Syndrome|Past Medical History|2164,2172|false|false|false|C0086543|Cataract|CATARACT
Event|Event|Past Medical History|2164,2172|false|false|false|||CATARACT
Finding|Finding|Past Medical History|2164,2172|false|false|false|C1690964|cataract on exam (physical finding)|CATARACT
Finding|Finding|Past Medical History|2164,2180|false|false|false|C1548833;C2186377|Consent Type - Cataract Surgery;reported history of cataract surgery|CATARACT SURGERY
Finding|Intellectual Product|Past Medical History|2164,2180|false|false|false|C1548833;C2186377|Consent Type - Cataract Surgery;reported history of cataract surgery|CATARACT SURGERY
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2164,2180|false|false|false|C0007389;C2939459|Cataract Extraction;Cataract surgery|CATARACT SURGERY
Event|Event|Past Medical History|2173,2180|false|false|false|||SURGERY
Finding|Finding|Past Medical History|2173,2180|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|SURGERY
Finding|Functional Concept|Past Medical History|2173,2180|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|SURGERY
Finding|Idea or Concept|Past Medical History|2173,2180|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|SURGERY
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2173,2180|false|false|false|C0543467|Operative Surgical Procedures|SURGERY
Finding|Finding|Past Medical History|2187,2194|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|Surgery
Finding|Functional Concept|Past Medical History|2187,2194|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|Surgery
Finding|Idea or Concept|Past Medical History|2187,2194|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|Surgery
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2187,2194|false|false|false|C0543467|Operative Surgical Procedures|Surgery
Finding|Functional Concept|Past Medical History|2208,2214|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|COMMON
Finding|Intellectual Product|Past Medical History|2208,2214|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|COMMON
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2208,2227|false|false|false|C1261084|Common iliac artery structure|COMMON ILIAC ARTERY
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2215,2220|false|false|false|C0020889|Bone structure of ilium|ILIAC
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2215,2227|false|false|false|C0020887|Structure of iliac artery|ILIAC ARTERY
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2221,2227|false|false|false|C0003842;C0226004|Arterial system;Arteries|ARTERY
Anatomy|Body System|Past Medical History|2221,2227|false|false|false|C0003842;C0226004|Arterial system;Arteries|ARTERY
Event|Event|Past Medical History|2228,2236|false|false|false|||STENTING
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2228,2236|false|false|false|C2348535|Stenting|STENTING
Event|Event|Past Medical History|2243,2255|false|false|false|||BUNIONECTOMY
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2243,2255|false|false|false|C1542057|Silver bunionectomy|BUNIONECTOMY
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2258,2261|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|HIP
Drug|Amino Acid, Peptide, or Protein|Past Medical History|2258,2261|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|HIP
Drug|Biologically Active Substance|Past Medical History|2258,2261|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|HIP
Drug|Pharmacologic Substance|Past Medical History|2258,2261|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|HIP
Event|Event|Past Medical History|2258,2261|false|false|false|||HIP
Finding|Gene or Genome|Past Medical History|2258,2261|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|HIP
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2258,2261|false|false|false|C1292890|Procedure on hip|HIP
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2258,2273|false|false|false|C0392806|Prosthetic arthroplasty of hip (procedure)|HIP REPLACEMENT
Event|Event|Past Medical History|2262,2273|false|false|false|||REPLACEMENT
Finding|Functional Concept|Past Medical History|2262,2273|false|false|false|C0559956|Replacement|REPLACEMENT
Procedure|Health Care Activity|Past Medical History|2262,2273|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|REPLACEMENT
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2262,2273|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|REPLACEMENT
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2282,2290|false|false|false|C3841297|Cesarean|CESAREAN
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2282,2298|false|false|false|C0007876|Cesarean section|CESAREAN SECTION
Drug|Substance|Past Medical History|2291,2298|false|false|false|C1522472|section sample|SECTION
Event|Event|Past Medical History|2291,2298|false|false|false|||SECTION
Finding|Intellectual Product|Past Medical History|2291,2298|false|false|false|C1551341;C1552858|Act Class - Section;Html Link Type - section|SECTION
Procedure|Laboratory Procedure|Past Medical History|2291,2298|false|false|false|C0700320|Sectioning technique|SECTION
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2301,2309|false|false|false|C0017067|Ganglia|GANGLION
Disorder|Anatomical Abnormality|Past Medical History|2301,2309|false|false|false|C0085648;C1258666|Myxoid cyst;Synovial Cyst|GANGLION
Disorder|Anatomical Abnormality|Past Medical History|2301,2314|false|false|false|C0085648;C1258666|Myxoid cyst;Synovial Cyst|GANGLION CYST
Disorder|Anatomical Abnormality|Past Medical History|2310,2314|false|false|false|C0010709|Cyst|CYST
Event|Event|Past Medical History|2310,2314|false|false|false|||CYST
Finding|Body Substance|Past Medical History|2310,2314|false|false|false|C1546594;C1550626|SpecimenType - Cyst|CYST
Finding|Intellectual Product|Past Medical History|2310,2314|false|false|false|C1546594;C1550626|SpecimenType - Cyst|CYST
Finding|Idea or Concept|Family Medical History|2353,2359|false|false|false|C1546508|Relationship - Mother|Mother
Disorder|Disease or Syndrome|Family Medical History|2366,2369|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|Family Medical History|2366,2369|false|false|false|||HTN
Finding|Conceptual Entity|Family Medical History|2372,2378|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Idea or Concept|Family Medical History|2372,2378|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Event|Event|Family Medical History|2389,2396|false|false|false|||Brother
Finding|Conceptual Entity|Family Medical History|2389,2396|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Finding|Idea or Concept|Family Medical History|2389,2396|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Event|Event|Family Medical History|2404,2411|false|false|false|||Brother
Finding|Conceptual Entity|Family Medical History|2404,2411|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Finding|Idea or Concept|Family Medical History|2404,2411|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Event|Event|Family Medical History|2420,2428|false|false|false|||Physical
Finding|Finding|Family Medical History|2420,2428|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|Family Medical History|2420,2428|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|Family Medical History|2420,2428|false|false|false|C0031809|Physical Examination|Physical
Event|Event|Family Medical History|2434,2443|false|false|false|||Admission
Procedure|Health Care Activity|Family Medical History|2434,2443|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Event|Event|Family Medical History|2492,2499|false|false|false|||General
Finding|Classification|Family Medical History|2492,2499|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|Family Medical History|2492,2499|false|false|false|C3812897|General medical service|General
Attribute|Clinical Attribute|Family Medical History|2501,2506|true|false|false|C5890168||Alert
Drug|Organic Chemical|Family Medical History|2501,2506|true|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Family Medical History|2501,2506|true|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|Family Medical History|2501,2506|true|false|false|||Alert
Finding|Finding|Family Medical History|2501,2506|true|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Family Medical History|2501,2506|true|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Family Medical History|2501,2506|true|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|Family Medical History|2508,2516|true|false|false|||oriented
Finding|Intellectual Product|Family Medical History|2521,2526|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|Family Medical History|2527,2535|true|false|false|||distress
Finding|Finding|Family Medical History|2527,2535|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|Family Medical History|2527,2535|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Anatomy|Body Location or Region|Family Medical History|2538,2543|true|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2545,2551|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|Family Medical History|2545,2551|false|false|false|C0036412|Scleral Diseases|Sclera
Event|Event|Family Medical History|2545,2551|false|false|false|||Sclera
Procedure|Health Care Activity|Family Medical History|2545,2551|false|false|false|C2228481|examination of sclera|Sclera
Event|Event|Family Medical History|2552,2561|false|false|false|||anicteric
Finding|Finding|Family Medical History|2552,2561|false|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2563,2566|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|Family Medical History|2563,2566|false|false|false|C0026987|Myelofibrosis|MMM
Anatomy|Body Location or Region|Family Medical History|2568,2578|false|false|false|C0521367|Oropharyngeal|oropharynx
Event|Event|Family Medical History|2579,2584|false|false|false|||clear
Finding|Idea or Concept|Family Medical History|2579,2584|false|false|false|C1550016|Remote control command - Clear|clear
Event|Event|Family Medical History|2586,2590|false|false|false|||EOMI
Event|Event|Family Medical History|2592,2597|false|false|false|||PERRL
Finding|Finding|Family Medical History|2592,2597|false|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Anatomy|Body Location or Region|Family Medical History|2600,2604|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Anatomy|Cell Component|Family Medical History|2600,2604|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Finding|Finding|Family Medical History|2600,2604|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|Neck
Event|Event|Family Medical History|2606,2612|true|false|false|||Supple
Finding|Functional Concept|Family Medical History|2606,2612|true|false|false|C0332254|Supple|Supple
Event|Event|Family Medical History|2614,2617|true|false|false|||JVP
Finding|Finding|Family Medical History|2614,2617|true|false|false|C0428897|Jugular venous pressure|JVP
Event|Event|Family Medical History|2622,2630|true|false|false|||elevated
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2635,2638|true|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|Family Medical History|2635,2638|true|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|Family Medical History|2635,2638|true|false|false|||LAD
Finding|Gene or Genome|Family Medical History|2635,2638|true|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Event|Activity|Family Medical History|2653,2657|false|false|false|C0871208|Rating (action)|rate
Event|Event|Family Medical History|2653,2657|false|false|false|||rate
Finding|Idea or Concept|Family Medical History|2653,2657|false|false|false|C1549480|Amount type - Rate|rate
Event|Event|Family Medical History|2662,2668|false|false|false|||rhythm
Finding|Finding|Family Medical History|2662,2668|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|Family Medical History|2662,2668|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Organ or Tissue Function|Family Medical History|2690,2698|false|false|false|C0039155|Systole|systolic
Finding|Finding|Family Medical History|2690,2705|true|false|false|C0232257|Systolic Murmurs|systolic murmur
Event|Event|Family Medical History|2699,2705|true|false|false|||murmur
Finding|Finding|Family Medical History|2699,2705|true|false|false|C0018808|Heart murmur|murmur
Event|Event|Family Medical History|2707,2712|true|false|false|||heard
Event|Event|Family Medical History|2730,2734|true|false|false|||rubs
Finding|Finding|Family Medical History|2730,2734|true|false|false|C0232267|Pericardial friction rub|rubs
Event|Event|Family Medical History|2738,2745|true|false|false|||gallops
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2748,2753|true|false|false|C0024109|Lung|Lungs
Event|Event|Family Medical History|2755,2766|true|false|false|||inspiratory
Finding|Organism Function|Family Medical History|2755,2766|true|false|false|C0004048|Inspiration (function)|inspiratory
Finding|Organism Function|Family Medical History|2771,2781|true|false|false|C0231800|Expiration, Respiratory|expiratory
Finding|Sign or Symptom|Family Medical History|2771,2789|true|false|false|C0231875|Expiratory wheezing|expiratory wheezes
Event|Event|Family Medical History|2782,2789|true|false|false|||wheezes
Finding|Sign or Symptom|Family Medical History|2782,2789|true|false|false|C0043144|Wheezing|wheezes
Event|Event|Family Medical History|2794,2799|true|false|false|||rales
Finding|Finding|Family Medical History|2794,2799|true|false|false|C0034642;C0240859|Basilar Rales;Rales|rales
Event|Event|Family Medical History|2803,2810|true|false|false|||rhonchi
Finding|Finding|Family Medical History|2803,2810|true|false|false|C0035508|Rhonchi|rhonchi
Anatomy|Body Location or Region|Family Medical History|2813,2820|true|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|Family Medical History|2813,2820|true|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Event|Event|Family Medical History|2813,2820|true|false|false|||Abdomen
Finding|Finding|Family Medical History|2813,2820|true|false|false|C0941288|Abdomen problem|Abdomen
Disorder|Disease or Syndrome|Family Medical History|2822,2826|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Event|Event|Family Medical History|2822,2826|false|false|false|||Soft
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2855,2860|true|false|false|C0021853|Intestines|bowel
Finding|Finding|Family Medical History|2855,2867|true|false|false|C0232693|Bowel sounds|bowel sounds
Event|Event|Family Medical History|2861,2867|true|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|Family Medical History|2861,2867|true|false|false|C0037709||sounds
Finding|Finding|Family Medical History|2868,2875|true|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|Family Medical History|2868,2875|true|false|false|C0150312;C0449450|Present;Presentation|present
Event|Event|Family Medical History|2881,2893|true|false|false|||organomegaly
Finding|Finding|Family Medical History|2881,2893|true|false|false|C4054315|Organomegaly|organomegaly
Event|Event|Family Medical History|2898,2905|true|false|false|||rebound
Event|Event|Family Medical History|2909,2917|true|false|false|||guarding
Finding|Finding|Family Medical History|2909,2917|true|false|false|C0427198|Protective muscle spasm|guarding
Disorder|Congenital Abnormality|Family Medical History|2935,2938|true|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Event|Event|Family Medical History|2935,2938|true|false|false|||Ext
Finding|Gene or Genome|Family Medical History|2935,2938|true|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Event|Event|Family Medical History|2940,2944|false|false|false|||Warm
Finding|Finding|Family Medical History|2940,2944|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|Family Medical History|2940,2944|false|false|false|C0687712|warming process|Warm
Finding|Finding|Family Medical History|2946,2950|true|false|false|C5575035|Well (answer to question)|well
Event|Event|Family Medical History|2951,2959|true|false|false|||perfused
Drug|Food|Family Medical History|2964,2970|true|false|false|C5890763||pulses
Event|Event|Family Medical History|2964,2970|true|false|false|||pulses
Finding|Physiologic Function|Family Medical History|2964,2970|true|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|Family Medical History|2964,2970|true|false|false|C0034107|Pulse taking|pulses
Disorder|Anatomical Abnormality|Family Medical History|2975,2983|true|false|false|C0149651|Clubbing|clubbing
Event|Event|Family Medical History|2975,2983|true|false|false|||clubbing
Event|Event|Family Medical History|2985,2993|true|false|false|||cyanosis
Finding|Sign or Symptom|Family Medical History|2985,2993|true|false|false|C0010520|Cyanosis|cyanosis
Attribute|Clinical Attribute|Family Medical History|2998,3003|true|false|false|C1717255||edema
Event|Event|Family Medical History|2998,3003|true|false|false|||edema
Finding|Pathologic Function|Family Medical History|2998,3003|true|false|false|C0013604|Edema|edema
Event|Event|Family Medical History|3005,3014|false|false|false|||Discharge
Finding|Body Substance|Family Medical History|3005,3014|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Family Medical History|3005,3014|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Family Medical History|3005,3014|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Family Medical History|3005,3014|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Family Medical History|3050,3056|false|false|false|C0944911||Weight
Event|Event|Family Medical History|3050,3056|false|false|false|||Weight
Finding|Finding|Family Medical History|3050,3056|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|Weight
Finding|Sign or Symptom|Family Medical History|3050,3056|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|Weight
Procedure|Health Care Activity|Family Medical History|3050,3056|false|false|false|C1305866|Weighing patient|Weight
Attribute|Clinical Attribute|Family Medical History|3063,3069|false|false|false|C0944911||Weight
Event|Event|Family Medical History|3063,3069|false|false|false|||Weight
Finding|Finding|Family Medical History|3063,3069|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|Weight
Finding|Sign or Symptom|Family Medical History|3063,3069|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|Weight
Procedure|Health Care Activity|Family Medical History|3063,3069|false|false|false|C1305866|Weighing patient|Weight
Event|Event|Family Medical History|3073,3082|false|false|false|||admission
Procedure|Health Care Activity|Family Medical History|3073,3082|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|Family Medical History|3089,3096|false|false|false|||General
Finding|Classification|Family Medical History|3089,3096|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|Family Medical History|3089,3096|false|false|false|C3812897|General medical service|General
Disorder|Disease or Syndrome|Family Medical History|3098,3101|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|Family Medical History|3098,3101|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|Family Medical History|3098,3101|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Family Medical History|3098,3101|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|Family Medical History|3098,3101|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|Family Medical History|3098,3101|false|false|false|||NAD
Finding|Finding|Family Medical History|3098,3101|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Location or Region|Family Medical History|3103,3108|false|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|3110,3116|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|Family Medical History|3110,3116|false|false|false|C0036412|Scleral Diseases|Sclera
Event|Event|Family Medical History|3110,3116|false|false|false|||Sclera
Procedure|Health Care Activity|Family Medical History|3110,3116|false|false|false|C2228481|examination of sclera|Sclera
Event|Event|Family Medical History|3117,3126|false|false|false|||anicteric
Finding|Finding|Family Medical History|3117,3126|false|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Location or Region|Family Medical History|3128,3132|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Anatomy|Cell Component|Family Medical History|3128,3132|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Finding|Finding|Family Medical History|3128,3132|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|Neck
Event|Event|Family Medical History|3134,3137|true|false|false|||JVP
Finding|Finding|Family Medical History|3134,3137|true|false|false|C0428897|Jugular venous pressure|JVP
Event|Event|Family Medical History|3142,3150|true|false|false|||elevated
Event|Event|Family Medical History|3165,3171|false|false|false|||rhythm
Finding|Finding|Family Medical History|3165,3171|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|Family Medical History|3165,3171|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Event|Event|Family Medical History|3194,3199|false|false|false|||beats
Finding|Organ or Tissue Function|Family Medical History|3222,3230|true|false|false|C0039155|Systole|systolic
Finding|Finding|Family Medical History|3222,3237|true|false|false|C0232257|Systolic Murmurs|systolic murmur
Event|Event|Family Medical History|3231,3237|true|false|false|||murmur
Finding|Finding|Family Medical History|3231,3237|true|false|false|C0018808|Heart murmur|murmur
Event|Event|Family Medical History|3261,3265|true|false|false|||rubs
Finding|Finding|Family Medical History|3261,3265|true|false|false|C0232267|Pericardial friction rub|rubs
Event|Event|Family Medical History|3269,3276|true|false|false|||gallops
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|3279,3284|true|false|false|C0024109|Lung|Lungs
Finding|Intellectual Product|Family Medical History|3286,3290|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Organism Function|Family Medical History|3291,3301|false|false|false|C0231800|Expiration, Respiratory|expiratory
Finding|Sign or Symptom|Family Medical History|3291,3309|false|false|false|C0231875|Expiratory wheezing|expiratory wheezes
Event|Event|Family Medical History|3302,3309|false|false|false|||wheezes
Finding|Sign or Symptom|Family Medical History|3302,3309|false|false|false|C0043144|Wheezing|wheezes
Finding|Intellectual Product|Family Medical History|3319,3323|false|false|false|C1547225|Mild Severity of Illness Code|mild
Event|Event|Family Medical History|3324,3331|false|false|false|||rhonchi
Finding|Finding|Family Medical History|3324,3331|false|false|false|C0035508|Rhonchi|rhonchi
Anatomy|Body Location or Region|Family Medical History|3350,3357|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|Family Medical History|3350,3357|false|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Event|Event|Family Medical History|3350,3357|false|false|false|||Abdomen
Finding|Finding|Family Medical History|3350,3357|false|false|false|C0941288|Abdomen problem|Abdomen
Disorder|Disease or Syndrome|Family Medical History|3359,3363|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Event|Event|Family Medical History|3359,3363|false|false|false|||Soft
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|3392,3397|true|false|false|C0021853|Intestines|bowel
Finding|Finding|Family Medical History|3392,3404|true|false|false|C0232693|Bowel sounds|bowel sounds
Event|Event|Family Medical History|3398,3404|true|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|Family Medical History|3398,3404|true|false|false|C0037709||sounds
Finding|Finding|Family Medical History|3405,3412|true|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|Family Medical History|3405,3412|true|false|false|C0150312;C0449450|Present;Presentation|present
Event|Event|Family Medical History|3418,3430|true|false|false|||organomegaly
Finding|Finding|Family Medical History|3418,3430|true|false|false|C4054315|Organomegaly|organomegaly
Event|Event|Family Medical History|3435,3442|true|false|false|||rebound
Event|Event|Family Medical History|3446,3454|true|false|false|||guarding
Finding|Finding|Family Medical History|3446,3454|true|false|false|C0427198|Protective muscle spasm|guarding
Disorder|Congenital Abnormality|Family Medical History|3458,3461|true|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Event|Event|Family Medical History|3458,3461|true|false|false|||Ext
Finding|Gene or Genome|Family Medical History|3458,3461|true|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Event|Event|Family Medical History|3463,3467|true|false|false|||Warm
Finding|Finding|Family Medical History|3463,3467|true|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|Family Medical History|3463,3467|true|false|false|C0687712|warming process|Warm
Finding|Finding|Family Medical History|3469,3473|true|false|false|C5575035|Well (answer to question)|well
Event|Event|Family Medical History|3474,3482|true|false|false|||perfused
Attribute|Clinical Attribute|Family Medical History|3487,3492|true|false|false|C1717255||edema
Event|Event|Family Medical History|3487,3492|true|false|false|||edema
Finding|Pathologic Function|Family Medical History|3487,3492|true|false|false|C0013604|Edema|edema
Procedure|Health Care Activity|Family Medical History|3516,3525|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Event|Event|Family Medical History|3526,3530|false|false|false|||Labs
Lab|Laboratory or Test Result|Family Medical History|3526,3530|false|false|false|C0587081|Laboratory test finding|Labs
Disorder|Neoplastic Process|Family Medical History|3552,3555|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|Family Medical History|3552,3555|false|false|false|||PTT
Procedure|Laboratory Procedure|Family Medical History|3552,3555|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Drug|Organic Chemical|Family Medical History|3579,3586|false|false|false|C0022924;C0376261|Lactates;lactate|LACTATE
Drug|Pharmacologic Substance|Family Medical History|3579,3586|false|false|false|C0022924;C0376261|Lactates;lactate|LACTATE
Event|Event|Family Medical History|3579,3586|false|false|false|||LACTATE
Procedure|Laboratory Procedure|Family Medical History|3579,3586|false|false|false|C0202115|Lactic acid measurement|LACTATE
Drug|Biologically Active Substance|Family Medical History|3605,3612|false|false|false|C0017725|glucose|GLUCOSE
Drug|Organic Chemical|Family Medical History|3605,3612|false|false|false|C0017725|glucose|GLUCOSE
Drug|Pharmacologic Substance|Family Medical History|3605,3612|false|false|false|C0017725|glucose|GLUCOSE
Event|Event|Family Medical History|3605,3612|false|false|false|||GLUCOSE
Lab|Laboratory or Test Result|Family Medical History|3605,3612|false|false|false|C5781949|Glucose^1.5H post dose glucagon|GLUCOSE
Procedure|Laboratory Procedure|Family Medical History|3605,3612|false|false|false|C0337438|Glucose measurement|GLUCOSE
Drug|Biologically Active Substance|Family Medical History|3618,3622|false|false|false|C0041942|urea|UREA
Drug|Organic Chemical|Family Medical History|3618,3622|false|false|false|C0041942|urea|UREA
Drug|Pharmacologic Substance|Family Medical History|3618,3622|false|false|false|C0041942|urea|UREA
Event|Event|Family Medical History|3618,3622|false|false|false|||UREA
Procedure|Laboratory Procedure|Family Medical History|3618,3622|false|false|false|C0523961|Urea measurement|UREA
Drug|Biologically Active Substance|Family Medical History|3638,3644|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Element, Ion, or Isotope|Family Medical History|3638,3644|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Pharmacologic Substance|Family Medical History|3638,3644|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Event|Event|Family Medical History|3638,3644|false|false|false|||SODIUM
Finding|Physiologic Function|Family Medical History|3638,3644|false|false|false|C4553025|Sodium metabolic function|SODIUM
Procedure|Laboratory Procedure|Family Medical History|3638,3644|false|false|false|C0337443|Sodium measurement|SODIUM
Drug|Biologically Active Substance|Family Medical History|3650,3659|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Element, Ion, or Isotope|Family Medical History|3650,3659|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Food|Family Medical History|3650,3659|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Inorganic Chemical|Family Medical History|3650,3659|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Pharmacologic Substance|Family Medical History|3650,3659|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Event|Event|Family Medical History|3650,3659|false|false|false|||POTASSIUM
Finding|Physiologic Function|Family Medical History|3650,3659|false|false|false|C4553027|Potassium metabolic function|POTASSIUM
Procedure|Laboratory Procedure|Family Medical History|3650,3659|false|false|false|C0202194|Potassium measurement|POTASSIUM
Drug|Element, Ion, or Isotope|Family Medical History|3665,3673|false|false|false|C0008203;C0596019|Chlorides;chloride ion|CHLORIDE
Event|Event|Family Medical History|3665,3673|false|false|false|||CHLORIDE
Finding|Physiologic Function|Family Medical History|3665,3673|false|false|false|C4553021|Chloride metabolic function|CHLORIDE
Procedure|Laboratory Procedure|Family Medical History|3665,3673|false|false|false|C0201952|Chloride measurement|CHLORIDE
Drug|Biologically Active Substance|Family Medical History|3684,3687|false|false|false|C0007012|carbon dioxide|CO2
Drug|Inorganic Chemical|Family Medical History|3684,3687|false|false|false|C0007012|carbon dioxide|CO2
Event|Event|Family Medical History|3684,3687|false|false|false|||CO2
Finding|Finding|Family Medical History|3684,3687|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Finding|Gene or Genome|Family Medical History|3684,3687|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Drug|Element, Ion, or Isotope|Family Medical History|3691,3696|false|false|false|C0003075|Anions|ANION
Attribute|Clinical Attribute|Family Medical History|3691,3700|false|false|false|C0003074|Anion Gap|ANION GAP
Lab|Laboratory or Test Result|Family Medical History|3691,3700|false|false|false|C1509129|Anion gap result|ANION GAP
Procedure|Laboratory Procedure|Family Medical History|3691,3700|false|false|false|C0201889;C2189246|Anion gap measurement;blood anion gap (lab test)|ANION GAP
Drug|Amino Acid, Peptide, or Protein|Family Medical History|3697,3700|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Drug|Biologically Active Substance|Family Medical History|3697,3700|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Event|Event|Family Medical History|3697,3700|false|false|false|||GAP
Finding|Gene or Genome|Family Medical History|3697,3700|false|false|false|C1419277;C2984552|RASA1 gene;RASA1 wt Allele|GAP
Drug|Biologically Active Substance|Family Medical History|3778,3785|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Element, Ion, or Isotope|Family Medical History|3778,3785|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Inorganic Chemical|Family Medical History|3778,3785|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Pharmacologic Substance|Family Medical History|3778,3785|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Vitamin|Family Medical History|3778,3785|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Event|Event|Family Medical History|3778,3785|false|false|false|||CALCIUM
Finding|Physiologic Function|Family Medical History|3778,3785|false|false|false|C4553026|Calcium metabolic function|CALCIUM
Procedure|Laboratory Procedure|Family Medical History|3778,3785|false|false|false|C0201925|Calcium measurement|CALCIUM
Drug|Element, Ion, or Isotope|Family Medical History|3792,3801|false|false|false|C0031603;C1601799|Phosphates;phosphate ion|PHOSPHATE
Drug|Inorganic Chemical|Family Medical History|3792,3801|false|false|false|C0031603;C1601799|Phosphates;phosphate ion|PHOSPHATE
Drug|Pharmacologic Substance|Family Medical History|3792,3801|false|false|false|C0031603;C1601799|Phosphates;phosphate ion|PHOSPHATE
Procedure|Laboratory Procedure|Family Medical History|3792,3801|false|false|false|C0523826|Phosphate measurement|PHOSPHATE
Drug|Biologically Active Substance|Family Medical History|3806,3815|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Drug|Element, Ion, or Isotope|Family Medical History|3806,3815|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Drug|Inorganic Chemical|Family Medical History|3806,3815|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Drug|Pharmacologic Substance|Family Medical History|3806,3815|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Event|Event|Family Medical History|3806,3815|false|false|false|||MAGNESIUM
Procedure|Laboratory Procedure|Family Medical History|3806,3815|false|false|false|C0373675|Magnesium measurement|MAGNESIUM
Anatomy|Cell|Family Medical History|3834,3837|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|Family Medical History|3842,3845|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|Family Medical History|3842,3845|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|Family Medical History|3842,3845|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|Family Medical History|3851,3854|false|false|false|C0019046|Hemoglobin|HGB
Drug|Biologically Active Substance|Family Medical History|3851,3854|false|false|false|C0019046|Hemoglobin|HGB
Event|Event|Family Medical History|3851,3854|false|false|false|||HGB
Finding|Gene or Genome|Family Medical History|3851,3854|false|false|false|C1424337|CYGB gene|HGB
Lab|Laboratory or Test Result|Family Medical History|3851,3854|false|false|false|C0019029|Hemoglobin concentration|HGB
Event|Event|Family Medical History|3860,3863|false|false|false|||HCT
Procedure|Laboratory Procedure|Family Medical History|3860,3863|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Procedure|Therapeutic or Preventive Procedure|Family Medical History|3860,3863|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Disorder|Virus|Family Medical History|3869,3872|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|Family Medical History|3869,3872|false|false|false|||MCV
Lab|Laboratory or Test Result|Family Medical History|3869,3872|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|Family Medical History|3869,3872|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|Family Medical History|3869,3872|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|Family Medical History|3877,3880|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|Family Medical History|3877,3880|false|false|false|C0600370|methacholine|MCH
Event|Event|Family Medical History|3877,3880|false|false|false|||MCH
Finding|Gene or Genome|Family Medical History|3877,3880|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|Family Medical History|3877,3880|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|Family Medical History|3877,3880|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|Family Medical History|3886,3890|false|false|false|||MCHC
Procedure|Laboratory Procedure|Family Medical History|3886,3890|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Drug|Antibiotic|Family Medical History|3946,3951|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Biomedical or Dental Material|Family Medical History|3946,3951|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Organic Chemical|Family Medical History|3946,3951|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Disorder|Disease or Syndrome|Family Medical History|3956,3959|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|EOS
Event|Event|Family Medical History|3956,3959|false|false|false|||EOS
Finding|Gene or Genome|Family Medical History|3956,3959|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|EOS
Event|Event|Family Medical History|4063,4066|false|false|false|||PLT
Procedure|Laboratory Procedure|Family Medical History|4063,4066|false|false|false|C0201617|Primed lymphocyte test|PLT
Event|Event|Family Medical History|4078,4087|false|false|false|||Discharge
Finding|Body Substance|Family Medical History|4078,4087|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Family Medical History|4078,4087|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Family Medical History|4078,4087|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Family Medical History|4078,4087|false|false|false|C0030685|Patient Discharge|Discharge
Lab|Laboratory or Test Result|Family Medical History|4088,4092|false|false|false|C0587081|Laboratory test finding|Labs
Disorder|Disease or Syndrome|Family Medical History|4107,4112|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|4107,4112|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|4107,4112|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|Family Medical History|4113,4116|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|Family Medical History|4121,4124|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|Family Medical History|4121,4124|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|Family Medical History|4121,4124|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|Family Medical History|4130,4133|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|Family Medical History|4130,4133|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|Family Medical History|4130,4133|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|Family Medical History|4130,4133|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|Family Medical History|4139,4142|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|Family Medical History|4139,4142|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|Family Medical History|4148,4151|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|Family Medical History|4148,4151|false|false|false|||MCV
Lab|Laboratory or Test Result|Family Medical History|4148,4151|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|Family Medical History|4148,4151|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|Family Medical History|4148,4151|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|Family Medical History|4156,4159|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|Family Medical History|4156,4159|false|false|false|C0600370|methacholine|MCH
Event|Event|Family Medical History|4156,4159|false|false|false|||MCH
Finding|Gene or Genome|Family Medical History|4156,4159|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|Family Medical History|4156,4159|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|Family Medical History|4156,4159|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|Family Medical History|4165,4169|false|false|false|||MCHC
Procedure|Laboratory Procedure|Family Medical History|4165,4169|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Event|Event|Family Medical History|4175,4178|false|false|false|||RDW
Procedure|Laboratory Procedure|Family Medical History|4196,4199|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|Family Medical History|4216,4221|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|Family Medical History|4216,4221|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|Family Medical History|4222,4225|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|Family Medical History|4242,4247|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|4242,4247|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|4242,4247|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|Family Medical History|4242,4255|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|Family Medical History|4242,4255|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|Family Medical History|4242,4255|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|Family Medical History|4248,4255|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|Family Medical History|4248,4255|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|Family Medical History|4248,4255|false|false|false|C0017725|glucose|Glucose
Event|Event|Family Medical History|4248,4255|false|false|false|||Glucose
Lab|Laboratory or Test Result|Family Medical History|4248,4255|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|Family Medical History|4248,4255|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|Family Medical History|4298,4302|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|Family Medical History|4298,4302|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|Family Medical History|4298,4302|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|Family Medical History|4327,4332|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|4327,4332|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|4327,4332|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|Family Medical History|4333,4336|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|Family Medical History|4333,4336|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|Family Medical History|4333,4336|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|Family Medical History|4333,4336|false|false|false|||ALT
Finding|Gene or Genome|Family Medical History|4333,4336|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|Family Medical History|4333,4336|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|Family Medical History|4333,4336|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|Family Medical History|4333,4336|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|Family Medical History|4340,4343|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|Family Medical History|4340,4343|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|Family Medical History|4340,4343|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|Family Medical History|4340,4343|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|Family Medical History|4340,4343|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|Family Medical History|4340,4343|false|false|false|||AST
Finding|Gene or Genome|Family Medical History|4340,4343|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|Family Medical History|4350,4353|false|false|false|C0022917|Lactate Dehydrogenase|LDH
Drug|Enzyme|Family Medical History|4350,4353|false|false|false|C0022917|Lactate Dehydrogenase|LDH
Event|Event|Family Medical History|4350,4353|false|false|false|||LDH
Finding|Finding|Family Medical History|4350,4353|false|false|false|C0851148|Lifetime Drinking History|LDH
Procedure|Laboratory Procedure|Family Medical History|4350,4353|false|false|false|C0202113|Lactate dehydrogenase measurement|LDH
Drug|Amino Acid, Peptide, or Protein|Family Medical History|4360,4367|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|Family Medical History|4360,4367|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Disorder|Disease or Syndrome|Family Medical History|4396,4401|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|4396,4401|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|4396,4401|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|Family Medical History|4396,4409|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|Family Medical History|4402,4409|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|Family Medical History|4402,4409|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|Family Medical History|4402,4409|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|Family Medical History|4402,4409|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|Family Medical History|4402,4409|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|Family Medical History|4402,4409|false|false|false|||Calcium
Finding|Physiologic Function|Family Medical History|4402,4409|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|Family Medical History|4402,4409|false|false|false|C0201925|Calcium measurement|Calcium
Event|Event|Family Medical History|4431,4438|false|false|false|||Studies
Procedure|Research Activity|Family Medical History|4431,4438|false|false|false|C0947630|Scientific Study|Studies
Event|Event|Family Medical History|4443,4446|false|false|false|||CXR
Procedure|Diagnostic Procedure|Family Medical History|4443,4446|false|false|false|C0039985|Plain chest X-ray|CXR
Finding|Intellectual Product|Family Medical History|4455,4460|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Anatomy|Body Location or Region|Family Medical History|4461,4476|true|false|false|C0553534|Cardiopulmonary|cardiopulmonary
Disorder|Disease or Syndrome|Family Medical History|4461,4476|true|false|false|C4072686|Cardiovascular disease+Pulmonary disease|cardiopulmonary
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|4477,4484|true|false|false|C1184743|bony process|process
Drug|Pharmacologic Substance|Family Medical History|4477,4484|true|false|false|C1951340|Process Pharmacologic Substance|process
Event|Event|Family Medical History|4477,4484|true|false|false|||process
Finding|Functional Concept|Family Medical History|4477,4484|true|false|false|C4521054|Process (qualifier value)|process
Phenomenon|Phenomenon or Process|Family Medical History|4477,4484|true|false|false|C1522240|Process|process
Event|Event|Family Medical History|4495,4503|false|false|false|||Exercise
Finding|Daily or Recreational Activity|Family Medical History|4495,4503|false|false|false|C0015259|Exercise|Exercise
Procedure|Therapeutic or Preventive Procedure|Family Medical History|4495,4503|false|false|false|C1522704|Exercise Pain Management|Exercise
Procedure|Diagnostic Procedure|Family Medical History|4495,4515|false|false|false|C0015260;C0430120|Exercise stress test;Exercise stress test - endocrine|Exercise stress test
Attribute|Clinical Attribute|Family Medical History|4504,4510|false|false|false|C1718621|W stress|stress
Drug|Organic Chemical|Family Medical History|4504,4510|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|Family Medical History|4504,4510|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Finding|Finding|Family Medical History|4504,4510|false|false|false|C0038435|Stress|stress
Procedure|Diagnostic Procedure|Family Medical History|4504,4515|false|false|false|C0015260;C3494508|Exercise stress test;Stress Test|stress test
Anatomy|Body Location or Region|Family Medical History|4511,4515|false|false|false|C4318744|Test - temporal region|test
Event|Event|Family Medical History|4511,4515|false|false|false|||test
Finding|Functional Concept|Family Medical History|4511,4515|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Finding|Intellectual Product|Family Medical History|4511,4515|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Lab|Laboratory or Test Result|Family Medical History|4511,4515|false|false|false|C0456984|Test Result|test
Procedure|Laboratory Procedure|Family Medical History|4511,4515|false|false|false|C0022885|Laboratory Procedures|test
Attribute|Clinical Attribute|Family Medical History|4518,4532|false|false|false|C3173575||INTERPRETATION
Event|Event|Family Medical History|4518,4532|false|false|false|||INTERPRETATION
Finding|Intellectual Product|Family Medical History|4518,4532|false|false|false|C0459471|Interpretation Process|INTERPRETATION
Finding|Idea or Concept|Family Medical History|4543,4547|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|Family Medical History|4543,4547|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Event|Event|Family Medical History|4565,4572|false|false|false|||history
Finding|Conceptual Entity|Family Medical History|4565,4572|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|4565,4572|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Family Medical History|4565,4572|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|4565,4575|false|false|false|C0262926|Medical History|history of
Anatomy|Anatomical Structure|Family Medical History|4576,4579|false|false|false|C3669270|Strucure of thick cushion of skin|PAD
Disorder|Disease or Syndrome|Family Medical History|4576,4579|false|false|false|C0332568;C1704436|Pad Mass;Peripheral Arterial Diseases|PAD
Disorder|Neoplastic Process|Family Medical History|4576,4579|false|false|false|C0332568;C1704436|Pad Mass;Peripheral Arterial Diseases|PAD
Drug|Biomedical or Dental Material|Family Medical History|4576,4579|false|false|false|C2347441|Pad Dosage Form|PAD
Event|Event|Family Medical History|4576,4579|false|false|false|||PAD
Finding|Gene or Genome|Family Medical History|4576,4579|false|false|false|C1425244;C1425478;C3540603|DHX40 gene;PADI4 gene;PADI4 wt Allele|PAD
Procedure|Therapeutic or Preventive Procedure|Family Medical History|4576,4579|false|false|false|C3814046|PAD Regimen|PAD
Disorder|Disease or Syndrome|Family Medical History|4587,4591|false|false|false|C0023211|Left Bundle-Branch Block|LBBB
Event|Event|Family Medical History|4587,4591|false|false|false|||LBBB
Lab|Laboratory or Test Result|Family Medical History|4587,4591|false|false|false|C0344420||LBBB
Event|Event|Family Medical History|4596,4604|false|false|false|||referred
Finding|Gene or Genome|Family Medical History|4612,4615|true|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|lab
Finding|Intellectual Product|Family Medical History|4612,4615|true|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|lab
Event|Event|Family Medical History|4638,4646|false|false|false|||negative
Finding|Classification|Family Medical History|4638,4646|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Family Medical History|4638,4646|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Family Medical History|4638,4646|false|false|false|C5237010|Expression Negative|negative
Finding|Intellectual Product|Family Medical History|4648,4654|false|false|false|C0031082|Periodicals|serial
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|4657,4664|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|Family Medical History|4657,4664|false|false|false|C1314974|Cardiac attachment|cardiac
Procedure|Laboratory Procedure|Family Medical History|4657,4672|false|false|false|C1271630|Cardiac markers|cardiac markers
Event|Event|Family Medical History|4665,4672|false|false|false|||markers
Event|Event|Family Medical History|4677,4687|false|false|false|||evaluation
Finding|Idea or Concept|Family Medical History|4677,4687|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|Family Medical History|4677,4687|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Anatomy|Body Location or Region|Family Medical History|4691,4696|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Family Medical History|4691,4696|false|false|false|C0741025|Chest problem|chest
Finding|Sign or Symptom|Family Medical History|4691,4707|false|false|false|C0235710|Chest discomfort|chest discomfort
Event|Event|Family Medical History|4697,4707|false|false|false|||discomfort
Finding|Sign or Symptom|Family Medical History|4697,4707|false|false|false|C2364135|Discomfort|discomfort
Finding|Body Substance|Family Medical History|4713,4720|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Family Medical History|4713,4720|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Family Medical History|4713,4720|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Family Medical History|4728,4736|false|false|false|||referred
Drug|Organic Chemical|Family Medical History|4743,4755|false|false|false|C0012582|dipyridamole|dipyridamole
Drug|Pharmacologic Substance|Family Medical History|4743,4755|false|false|false|C0012582|dipyridamole|dipyridamole
Attribute|Clinical Attribute|Family Medical History|4756,4762|false|false|false|C1718621|W stress|stress
Drug|Organic Chemical|Family Medical History|4756,4762|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|Family Medical History|4756,4762|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Event|Event|Family Medical History|4756,4762|false|false|false|||stress
Finding|Finding|Family Medical History|4756,4762|false|false|false|C0038435|Stress|stress
Procedure|Diagnostic Procedure|Family Medical History|4756,4767|false|false|false|C0015260;C3494508|Exercise stress test;Stress Test|stress test
Anatomy|Body Location or Region|Family Medical History|4763,4767|false|false|false|C4318744|Test - temporal region|test
Event|Event|Family Medical History|4763,4767|false|false|false|||test
Finding|Functional Concept|Family Medical History|4763,4767|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Finding|Intellectual Product|Family Medical History|4763,4767|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Lab|Laboratory or Test Result|Family Medical History|4763,4767|false|false|false|C0456984|Test Result|test
Procedure|Laboratory Procedure|Family Medical History|4763,4767|false|false|false|C0022885|Laboratory Procedures|test
Drug|Organic Chemical|Family Medical History|4784,4796|false|false|false|C0039771|theophylline|theophylline
Drug|Pharmacologic Substance|Family Medical History|4784,4796|false|false|false|C0039771|theophylline|theophylline
Event|Event|Family Medical History|4784,4796|false|false|false|||theophylline
Procedure|Laboratory Procedure|Family Medical History|4784,4796|false|false|false|C0039773|Assay of theophylline|theophylline
Event|Event|Family Medical History|4799,4806|false|false|false|||therapy
Finding|Finding|Family Medical History|4799,4806|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|Family Medical History|4799,4806|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|Family Medical History|4799,4806|false|false|false|C0087111|Therapeutic procedure|therapy
Event|Event|Family Medical History|4819,4823|true|false|false|||able
Finding|Finding|Family Medical History|4819,4823|true|false|false|C1299581|Able (qualifier value)|able
Event|Event|Family Medical History|4827,4834|true|false|false|||proceed
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|4856,4862|false|false|false|C0018792|Heart Atrium|atrial
Event|Event|Family Medical History|4874,4879|true|false|false|||chose
Drug|Organic Chemical|Family Medical History|4896,4906|true|false|false|C0012963|dobutamine|dobutamine
Drug|Pharmacologic Substance|Family Medical History|4896,4906|true|false|false|C0012963|dobutamine|dobutamine
Event|Event|Family Medical History|4896,4906|true|false|false|||dobutamine
Finding|Daily or Recreational Activity|Family Medical History|4919,4923|false|false|false|C0080331|Walking (function)|walk
Event|Event|Family Medical History|4932,4941|false|false|false|||treadmill
Finding|Daily or Recreational Activity|Family Medical History|4932,4941|false|false|false|C2712999|Treadmill (physical activity)|treadmill
Procedure|Therapeutic or Preventive Procedure|Family Medical History|4932,4941|false|false|false|C2107089|treadmill conditioning training|treadmill
Event|Event|Family Medical History|4955,4964|false|false|false|||exercised
Event|Event|Family Medical History|4984,4992|false|false|false|||modified
Finding|Functional Concept|Family Medical History|4984,4992|false|false|false|C0392747|Changing|modified
Event|Event|Family Medical History|4998,5006|false|false|false|||protocol
Finding|Finding|Family Medical History|4998,5006|false|false|false|C0442711;C1507394;C1522729;C2348563;C3715209|Clinical trial protocol document;Library Protocol;Protocol - answer to question;Protocols documentation;Study Protocol|protocol
Finding|Intellectual Product|Family Medical History|4998,5006|false|false|false|C0442711;C1507394;C1522729;C2348563;C3715209|Clinical trial protocol document;Library Protocol;Protocol - answer to question;Protocols documentation;Study Protocol|protocol
Event|Event|Family Medical History|5011,5018|false|false|false|||stopped
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|5026,5029|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Disorder|Disease or Syndrome|Family Medical History|5030,5042|false|true|false|C0021775|Intermittent Claudication|claudication
Event|Event|Family Medical History|5030,5042|false|false|false|||claudication
Finding|Finding|Family Medical History|5030,5042|false|true|false|C0311395;C1456822|Claudication (finding);Lameness|claudication
Event|Event|Family Medical History|5068,5076|false|false|false|||capacity
Event|Event|Family Medical History|5091,5101|false|false|false|||represents
Event|Event|Family Medical History|5104,5108|false|false|false|||poor
Finding|Intellectual Product|Family Medical History|5104,5108|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|poor
Finding|Conceptual Entity|Family Medical History|5110,5120|false|false|false|C0205245;C0542341;C2700217|Function (attribute);Functional;Functional Relationship|functional
Finding|Functional Concept|Family Medical History|5110,5120|false|false|false|C0205245;C0542341;C2700217|Function (attribute);Functional;Functional Relationship|functional
Finding|Finding|Family Medical History|5110,5129|false|false|false|C1998319|Functional capacity|functional capacity
Event|Event|Family Medical History|5121,5129|false|false|false|||capacity
Attribute|Clinical Attribute|Family Medical History|5138,5141|false|false|false|C1114365||age
Drug|Biologically Active Substance|Family Medical History|5138,5141|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|Family Medical History|5138,5141|false|false|false|C0162574|Glycation End Products, Advanced|age
Event|Event|Family Medical History|5138,5141|false|false|false|||age
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|5146,5149|true|false|false|C0446516;C1140618;C1269078|Upper Extremity;Upper arm|arm
Disorder|Anatomical Abnormality|Family Medical History|5146,5149|true|false|false|C3495676|Anorectal Malformations|arm
Event|Event|Family Medical History|5146,5149|true|false|false|||arm
Finding|Gene or Genome|Family Medical History|5146,5149|true|false|false|C1824218;C3715044|AKR1A1 wt Allele;ARMC9 gene|arm
Procedure|Diagnostic Procedure|Family Medical History|5146,5149|true|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Research Activity|Family Medical History|5146,5149|true|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Therapeutic or Preventive Procedure|Family Medical History|5146,5149|true|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Anatomy|Body Location or Region|Family Medical History|5151,5155|true|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|Family Medical History|5151,5155|true|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|Family Medical History|5151,5155|true|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Event|Event|Family Medical History|5157,5161|true|false|false|||back
Anatomy|Body Location or Region|Family Medical History|5165,5170|true|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Family Medical History|5165,5170|true|false|false|C0741025|Chest problem|chest
Event|Event|Family Medical History|5172,5182|false|false|false|||discomfort
Finding|Sign or Symptom|Family Medical History|5172,5182|false|false|false|C2364135|Discomfort|discomfort
Event|Event|Family Medical History|5187,5195|false|false|false|||reported
Finding|Body Substance|Family Medical History|5203,5210|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Family Medical History|5203,5210|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Family Medical History|5203,5210|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Family Medical History|5226,5231|false|false|false|||study
Finding|Intellectual Product|Family Medical History|5226,5231|false|false|false|C1705923|Study Object|study
Procedure|Research Activity|Family Medical History|5226,5231|false|false|false|C0008972;C0947630;C2603343|Clinical Research;Scientific Study;Study|study
Event|Event|Family Medical History|5241,5249|false|false|false|||segments
Event|Event|Family Medical History|5254,5269|false|false|false|||uninterpretable
Event|Event|Family Medical History|5274,5282|false|false|false|||ischemia
Finding|Pathologic Function|Family Medical History|5274,5282|false|true|false|C0022116|Ischemia|ischemia
Procedure|Therapeutic or Preventive Procedure|Family Medical History|5274,5282|false|true|false|C4321499|Ischemia Procedure|ischemia
Finding|Mental Process|Family Medical History|5290,5297|false|false|false|C0542559|contextual factors|setting
Drug|Biomedical or Dental Material|Family Medical History|5306,5314|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|Family Medical History|5306,5314|false|false|false|||baseline
Finding|Idea or Concept|Family Medical History|5306,5314|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Disorder|Disease or Syndrome|Family Medical History|5315,5319|false|false|false|C0023211|Left Bundle-Branch Block|LBBB
Event|Event|Family Medical History|5315,5319|false|false|false|||LBBB
Lab|Laboratory or Test Result|Family Medical History|5315,5319|false|false|false|C0344420||LBBB
Event|Event|Family Medical History|5325,5331|false|false|false|||rhythm
Finding|Finding|Family Medical History|5325,5331|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|Family Medical History|5325,5331|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Anatomy|Body Space or Junction|Family Medical History|5336,5341|false|false|false|C0030471;C1305231|Nasal sinus;Sinus - general anatomical term|sinus
Disorder|Anatomical Abnormality|Family Medical History|5336,5341|false|false|false|C0016169|pathologic fistula|sinus
Drug|Organic Chemical|Family Medical History|5336,5341|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Drug|Pharmacologic Substance|Family Medical History|5336,5341|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Event|Event|Family Medical History|5336,5341|false|false|false|||sinus
Event|Event|Family Medical History|5356,5364|false|false|false|||isolated
Finding|Functional Concept|Family Medical History|5356,5364|false|false|false|C0205409;C1548221|Bed Status - Isolated;Isolated|isolated
Finding|Idea or Concept|Family Medical History|5356,5364|false|false|false|C0205409;C1548221|Bed Status - Isolated;Isolated|isolated
Event|Event|Family Medical History|5366,5370|false|false|false|||apbs
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|5383,5389|false|false|false|C0018792|Heart Atrium|atrial
Event|Event|Family Medical History|5390,5398|false|false|false|||couplets
Finding|Finding|Family Medical History|5390,5398|false|false|false|C0429001|Paired ventricular premature complexes|couplets
Finding|Daily or Recreational Activity|Family Medical History|5412,5415|false|false|false|C0035953;C0600140;C1704688;C4722187|Does run (finding);Go Jogging or Running Question;Run action;Running (physical activity)|run
Finding|Finding|Family Medical History|5412,5415|false|false|false|C0035953;C0600140;C1704688;C4722187|Does run (finding);Go Jogging or Running Question;Run action;Running (physical activity)|run
Finding|Functional Concept|Family Medical History|5412,5415|false|false|false|C0035953;C0600140;C1704688;C4722187|Does run (finding);Go Jogging or Running Question;Run action;Running (physical activity)|run
Finding|Intellectual Product|Family Medical History|5412,5415|false|false|false|C0035953;C0600140;C1704688;C4722187|Does run (finding);Go Jogging or Running Question;Run action;Running (physical activity)|run
Disorder|Disease or Syndrome|Family Medical History|5419,5423|false|false|false|C0030590|Paroxysmal supraventricular tachycardia|PSVT
Event|Event|Family Medical History|5419,5423|false|false|false|||PSVT
Finding|Finding|Family Medical History|5419,5423|false|false|false|C2108093|Paroxysmal Supraventricular Tachycardia by ECG Finding|PSVT
Finding|Gene or Genome|Family Medical History|5425,5429|false|false|false|C1514917|Retinoic Acid Response Element|Rare
Finding|Functional Concept|Family Medical History|5431,5439|false|false|false|C0205409;C1548221|Bed Status - Isolated;Isolated|isolated
Finding|Idea or Concept|Family Medical History|5431,5439|false|false|false|C0205409;C1548221|Bed Status - Isolated;Isolated|isolated
Disorder|Disease or Syndrome|Family Medical History|5440,5444|false|false|false|C0151636|Premature ventricular contractions|vpbs
Event|Event|Family Medical History|5440,5444|false|false|false|||vpbs
Event|Event|Family Medical History|5455,5460|false|false|false|||noted
Finding|Daily or Recreational Activity|Family Medical History|5462,5469|false|false|false|C0035253|Rest|Resting
Finding|Intellectual Product|Family Medical History|5470,5474|false|false|false|C1547225|Mild Severity of Illness Code|mild
Event|Event|Family Medical History|5475,5483|false|false|false|||systolic
Finding|Organ or Tissue Function|Family Medical History|5475,5483|false|false|false|C0039155|Systole|systolic
Disorder|Disease or Syndrome|Family Medical History|5485,5497|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|Family Medical History|5485,5497|false|false|false|||hypertension
Event|Event|Family Medical History|5517,5525|false|false|false|||increase
Finding|Functional Concept|Family Medical History|5517,5525|false|false|false|C0442805|Increase|increase
Event|Event|Family Medical History|5537,5545|false|false|false|||exercise
Finding|Daily or Recreational Activity|Family Medical History|5537,5545|false|false|false|C0015259|Exercise|exercise
Procedure|Therapeutic or Preventive Procedure|Family Medical History|5537,5545|false|false|false|C1522704|Exercise Pain Management|exercise
Event|Activity|Family Medical History|5551,5559|false|false|false|C0237820||recovery
Event|Event|Family Medical History|5551,5559|false|false|false|||recovery
Finding|Organism Function|Family Medical History|5551,5559|false|false|false|C2004454|Recovery - healing process|recovery
Event|Event|Family Medical History|5563,5573|false|false|false|||IMPRESSION
Finding|Intellectual Product|Family Medical History|5563,5573|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|Family Medical History|5563,5573|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Gene or Genome|Family Medical History|5586,5590|true|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Finding|Intellectual Product|Family Medical History|5586,5590|true|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Event|Event|Family Medical History|5591,5599|true|false|false|||symptoms
Finding|Functional Concept|Family Medical History|5591,5599|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Family Medical History|5591,5599|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|Family Medical History|5621,5629|false|false|false|||segments
Finding|Finding|Family Medical History|5635,5639|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|Family Medical History|5635,5639|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|Family Medical History|5635,5639|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|5640,5647|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|Family Medical History|5640,5647|false|false|false|C1314974|Cardiac attachment|cardiac
Event|Event|Family Medical History|5648,5654|false|false|false|||demand
Finding|Idea or Concept|Family Medical History|5648,5654|false|false|false|C0699784|Economic demand|demand
Procedure|Therapeutic or Preventive Procedure|Family Medical History|5648,5654|false|false|false|C0441516|Demand (clinical)|demand
Finding|Intellectual Product|Family Medical History|5659,5663|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|poor
Finding|Conceptual Entity|Family Medical History|5664,5674|false|false|false|C0205245;C0542341;C2700217|Function (attribute);Functional;Functional Relationship|functional
Finding|Functional Concept|Family Medical History|5664,5674|false|false|false|C0205245;C0542341;C2700217|Function (attribute);Functional;Functional Relationship|functional
Finding|Finding|Family Medical History|5664,5683|false|false|false|C1998319|Functional capacity|functional capacity
Event|Event|Family Medical History|5675,5683|false|false|false|||capacity
Attribute|Clinical Attribute|Family Medical History|5694,5700|false|false|false|C4255046||report
Event|Event|Family Medical History|5694,5700|false|false|false|||report
Finding|Intellectual Product|Family Medical History|5694,5700|false|false|false|C0684224|Report (document)|report
Procedure|Health Care Activity|Family Medical History|5694,5700|false|false|false|C0700287|Reporting|report
Event|Event|Family Medical History|5701,5705|false|false|false|||sent
Event|Event|Family Medical History|5727,5731|false|false|false|||CATH
Procedure|Therapeutic or Preventive Procedure|Family Medical History|5727,5731|false|false|false|C0007430|Catheterization|CATH
Drug|Organic Chemical|Family Medical History|5735,5739|false|false|false|C2828271|levomefolate calcium|LMCA
Drug|Pharmacologic Substance|Family Medical History|5735,5739|false|false|false|C2828271|levomefolate calcium|LMCA
Drug|Vitamin|Family Medical History|5735,5739|false|false|false|C2828271|levomefolate calcium|LMCA
Event|Event|Family Medical History|5735,5739|false|false|false|||LMCA
Disorder|Disease or Syndrome|Family Medical History|5751,5754|true|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Family Medical History|5751,5754|true|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Family Medical History|5751,5754|true|false|false|C1504769|DFFB protein, human|CAD
Event|Event|Family Medical History|5751,5754|true|false|false|||CAD
Finding|Gene or Genome|Family Medical History|5751,5754|true|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Family Medical History|5751,5754|true|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Family Medical History|5751,5754|true|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Family Medical History|5751,5754|true|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|5756,5759|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|Family Medical History|5756,5759|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|Family Medical History|5756,5759|false|false|false|||LAD
Finding|Gene or Genome|Family Medical History|5756,5759|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Finding|Intellectual Product|Family Medical History|5761,5765|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Finding|Family Medical History|5768,5780|false|false|false|C0449409|Focal origin|focal origin
Finding|Classification|Family Medical History|5774,5780|false|false|false|C0079946;C1550512|National origin;Participation Type - origin|origin
Finding|Intellectual Product|Family Medical History|5774,5780|false|false|false|C0079946;C1550512|National origin;Participation Type - origin|origin
Disorder|Disease or Syndrome|Family Medical History|5781,5788|false|false|false|C0012634|Disease|disease
Event|Event|Family Medical History|5781,5788|false|false|false|||disease
Finding|Intellectual Product|Family Medical History|5799,5803|false|false|false|C1547225|Mild Severity of Illness Code|mild
Attribute|Clinical Attribute|Family Medical History|5804,5812|false|false|false|C4489236|Proximal Resection Margin|proximal
Disorder|Disease or Syndrome|Family Medical History|5813,5820|false|false|false|C0012634|Disease|disease
Event|Event|Family Medical History|5813,5820|false|false|false|||disease
Drug|Amino Acid, Peptide, or Protein|Family Medical History|5828,5831|false|false|false|C2987138|Methylcytosine Dioxygenase TET1|LCX
Drug|Enzyme|Family Medical History|5828,5831|false|false|false|C2987138|Methylcytosine Dioxygenase TET1|LCX
Event|Event|Family Medical History|5828,5831|false|false|false|||LCX
Finding|Gene or Genome|Family Medical History|5828,5831|false|false|false|C1428863;C2987137|TET1 gene;TET1 wt Allele|LCX
Drug|Organic Chemical|Family Medical History|5844,5851|false|false|false|C0699493|Luminal|luminal
Drug|Pharmacologic Substance|Family Medical History|5844,5851|false|false|false|C0699493|Luminal|luminal
Event|Event|Family Medical History|5852,5866|false|false|false|||irregularities
Event|Event|Family Medical History|5868,5871|false|false|false|||RCA
Drug|Amino Acid, Peptide, or Protein|Family Medical History|5883,5886|false|false|false|C0018064|Equine Gonadotropins|ECG
Drug|Hormone|Family Medical History|5883,5886|false|false|false|C0018064|Equine Gonadotropins|ECG
Drug|Pharmacologic Substance|Family Medical History|5883,5886|false|false|false|C0018064|Equine Gonadotropins|ECG
Event|Event|Family Medical History|5883,5886|false|false|false|||ECG
Finding|Intellectual Product|Family Medical History|5883,5886|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|ECG
Procedure|Diagnostic Procedure|Family Medical History|5883,5886|false|false|false|C1623258|Electrocardiography|ECG
Anatomy|Body Space or Junction|Family Medical History|5892,5897|false|false|false|C0030471;C1305231|Nasal sinus;Sinus - general anatomical term|sinus
Disorder|Anatomical Abnormality|Family Medical History|5892,5897|false|false|false|C0016169|pathologic fistula|sinus
Drug|Organic Chemical|Family Medical History|5892,5897|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Drug|Pharmacologic Substance|Family Medical History|5892,5897|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Finding|Finding|Family Medical History|5892,5904|false|false|false|C0232201;C2041122|Sinus rhythm|sinus rhythm
Event|Event|Family Medical History|5898,5904|false|false|false|||rhythm
Finding|Finding|Family Medical History|5898,5904|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|Family Medical History|5898,5904|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Disorder|Disease or Syndrome|Family Medical History|5919,5923|false|false|false|C0033036|Atrial Premature Complexes|PACs
Event|Event|Family Medical History|5919,5923|false|false|false|||PACs
Finding|Intellectual Product|Family Medical History|5919,5923|false|false|false|C0182281|Picture Archiving and Communication Systems|PACs
Finding|Functional Concept|Family Medical History|5925,5929|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|5930,5934|false|false|false|C0004457|Axis vertebra|axis
Disorder|Injury or Poisoning|Family Medical History|5930,5934|false|false|false|C0349013|Fracture of second cervical vertebra|axis
Event|Event|Family Medical History|5936,5945|false|false|false|||deviation
Finding|Finding|Family Medical History|5936,5945|false|false|false|C1705236|Protocol Deviation|deviation
Event|Event|Family Medical History|5947,5950|false|false|false|||old
Disorder|Disease or Syndrome|Family Medical History|5951,5955|false|false|false|C0023211|Left Bundle-Branch Block|LBBB
Event|Event|Family Medical History|5951,5955|false|false|false|||LBBB
Lab|Laboratory or Test Result|Family Medical History|5951,5955|false|false|false|C0344420||LBBB
Drug|Amino Acid, Peptide, or Protein|Family Medical History|5960,5963|true|false|false|C0018064|Equine Gonadotropins|ECG
Drug|Hormone|Family Medical History|5960,5963|true|false|false|C0018064|Equine Gonadotropins|ECG
Drug|Pharmacologic Substance|Family Medical History|5960,5963|true|false|false|C0018064|Equine Gonadotropins|ECG
Event|Event|Family Medical History|5960,5963|false|false|false|||ECG
Finding|Intellectual Product|Family Medical History|5960,5963|true|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|ECG
Procedure|Diagnostic Procedure|Family Medical History|5960,5963|true|false|false|C1623258|Electrocardiography|ECG
Finding|Finding|Family Medical History|5969,5975|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Finding|Idea or Concept|Family Medical History|5969,5975|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|5976,5982|false|false|false|C0018792|Heart Atrium|atrial
Disorder|Disease or Syndrome|Family Medical History|5976,5994|false|true|false|C0546959|Atrial tachycardia|atrial tachycardia
Finding|Finding|Family Medical History|5976,5994|false|true|false|C2059391|continuous electrocardiogram atrial tachycardia|atrial tachycardia
Event|Event|Family Medical History|5983,5994|false|false|false|||tachycardia
Finding|Finding|Family Medical History|5983,5994|false|true|false|C0039231;C3827868|Tachycardia;Tachycardia by ECG Finding|tachycardia
Finding|Functional Concept|Family Medical History|5996,6000|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Drug|Chemical Viewed Structurally|Family Medical History|6008,6014|false|false|false|C1881507|Macromolecular Branch|branch
Event|Event|Family Medical History|6008,6014|false|false|false|||branch
Drug|Biomedical or Dental Material|Family Medical History|6016,6021|false|false|false|C1706085|Block Dosage Form|block
Event|Event|Family Medical History|6016,6021|false|false|false|||block
Finding|Body Substance|Family Medical History|6016,6021|false|false|false|C0028778;C0332206;C1533157|Blocking;Fixed Block;Obstruction|block
Finding|Finding|Family Medical History|6016,6021|false|false|false|C0028778;C0332206;C1533157|Blocking;Fixed Block;Obstruction|block
Finding|Functional Concept|Family Medical History|6016,6021|false|false|false|C0028778;C0332206;C1533157|Blocking;Fixed Block;Obstruction|block
Event|Event|Family Medical History|6023,6031|false|false|false|||Compared
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|6056,6062|false|false|false|C0018792|Heart Atrium|atrial
Disorder|Disease or Syndrome|Family Medical History|6056,6074|false|false|false|C0546959|Atrial tachycardia|atrial tachycardia
Finding|Finding|Family Medical History|6056,6074|false|false|false|C2059391|continuous electrocardiogram atrial tachycardia|atrial tachycardia
Event|Event|Family Medical History|6063,6074|false|false|false|||tachycardia
Finding|Finding|Family Medical History|6063,6074|false|false|false|C0039231;C3827868|Tachycardia;Tachycardia by ECG Finding|tachycardia
Event|Event|Family Medical History|6080,6088|false|false|false|||replaced
Anatomy|Body Space or Junction|Family Medical History|6089,6094|false|false|false|C0030471;C1305231|Nasal sinus;Sinus - general anatomical term|sinus
Disorder|Anatomical Abnormality|Family Medical History|6089,6094|false|false|false|C0016169|pathologic fistula|sinus
Drug|Organic Chemical|Family Medical History|6089,6094|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Drug|Pharmacologic Substance|Family Medical History|6089,6094|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Finding|Finding|Family Medical History|6089,6101|false|false|false|C0232201;C2041122|Sinus rhythm|sinus rhythm
Event|Event|Family Medical History|6095,6101|false|false|false|||rhythm
Finding|Finding|Family Medical History|6095,6101|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|Family Medical History|6095,6101|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Finding|Family Medical History|6107,6116|false|false|false|C0151526;C4018905|Premature Birth;Too early|premature
Finding|Pathologic Function|Family Medical History|6107,6116|false|false|false|C0151526;C4018905|Premature Birth;Too early|premature
Attribute|Clinical Attribute|Family Medical History|6107,6136|false|false|false|C0488348||premature atrial contractions
Disorder|Disease or Syndrome|Family Medical History|6107,6136|false|false|false|C0033036|Atrial Premature Complexes|premature atrial contractions
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|6117,6123|false|false|false|C0018792|Heart Atrium|atrial
Event|Event|Family Medical History|6124,6136|false|false|false|||contractions
Finding|Pathologic Function|Family Medical History|6124,6136|false|false|false|C1140999|Contraction (finding)|contractions
Finding|Functional Concept|Family Medical History|6138,6142|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Disorder|Disease or Syndrome|Family Medical History|6144,6163|false|false|false|C0006384|Bundle-Branch Block|bundle-branch block
Drug|Chemical Viewed Structurally|Family Medical History|6151,6157|false|false|false|C1881507|Macromolecular Branch|branch
Drug|Biomedical or Dental Material|Family Medical History|6158,6163|false|false|false|C1706085|Block Dosage Form|block
Event|Event|Family Medical History|6158,6163|false|false|false|||block
Finding|Body Substance|Family Medical History|6158,6163|false|false|false|C0028778;C0332206;C1533157|Blocking;Fixed Block;Obstruction|block
Finding|Finding|Family Medical History|6158,6163|false|false|false|C0028778;C0332206;C1533157|Blocking;Fixed Block;Obstruction|block
Finding|Functional Concept|Family Medical History|6158,6163|false|false|false|C0028778;C0332206;C1533157|Blocking;Fixed Block;Obstruction|block
Event|Event|Family Medical History|6179,6184|false|false|false|||noted
Event|Event|Family Medical History|6190,6194|false|false|false|||ECHO
Procedure|Health Care Activity|Family Medical History|6190,6194|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Procedure|Therapeutic or Preventive Procedure|Family Medical History|6190,6194|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Event|Event|Family Medical History|6200,6211|false|false|false|||Conclusions
Finding|Idea or Concept|Family Medical History|6200,6211|false|false|false|C1707478|Conclusion|Conclusions
Finding|Functional Concept|Family Medical History|6218,6222|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|6218,6229|false|false|false|C0225860|Left atrial structure|left atrium
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|6223,6229|false|false|false|C0018792|Heart Atrium|atrium
Event|Event|Family Medical History|6233,6239|false|false|false|||normal
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|6252,6258|true|false|false|C0018792|Heart Atrium|atrial
Disorder|Congenital Abnormality|Family Medical History|6252,6272|true|false|false|C0018817|Atrial Septal Defects|atrial septal defect
Disorder|Anatomical Abnormality|Family Medical History|6259,6272|true|false|false|C0018816;C5779791|Congenital septal defect of heart;Heart Septal Defects|septal defect
Disorder|Congenital Abnormality|Family Medical History|6259,6272|true|false|false|C0018816;C5779791|Congenital septal defect of heart;Heart Septal Defects|septal defect
Disorder|Disease or Syndrome|Family Medical History|6266,6272|true|false|false|C1861101|THYROID HORMONE PLASMA MEMBRANE TRANSPORT DEFECT|defect
Event|Event|Family Medical History|6266,6272|true|false|false|||defect
Finding|Functional Concept|Family Medical History|6266,6272|true|false|false|C1457869|Defect|defect
Event|Event|Family Medical History|6277,6281|true|false|false|||seen
Drug|Biomedical or Dental Material|Family Medical History|6291,6296|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|color
Drug|Indicator, Reagent, or Diagnostic Aid|Family Medical History|6291,6296|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|color
Procedure|Diagnostic Procedure|Family Medical History|6291,6304|false|false|false|C0474781|Color doppler ultrasound|color Doppler
Event|Event|Family Medical History|6297,6304|false|false|false|||Doppler
Procedure|Diagnostic Procedure|Family Medical History|6297,6304|false|false|false|C0554756|Doppler studies|Doppler
Finding|Functional Concept|Family Medical History|6320,6325|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Attribute|Clinical Attribute|Family Medical History|6320,6341|false|false|false|C0456165;C4050168|Right atrial pressure|right atrial pressure
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|6326,6332|false|false|false|C0018792|Heart Atrium|atrial
Finding|Finding|Family Medical History|6326,6341|false|false|false|C0428877|Atrial Pressure|atrial pressure
Event|Event|Family Medical History|6333,6341|false|false|false|||pressure
Finding|Finding|Family Medical History|6333,6341|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|Family Medical History|6333,6341|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|Family Medical History|6333,6341|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|Family Medical History|6333,6341|false|false|false|C0033095||pressure
Finding|Functional Concept|Family Medical History|6356,6360|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|6356,6377|false|false|false|C0504053|Wall of left ventricle|Left ventricular wall
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|6361,6372|false|false|false|C0018827|Heart Ventricle|ventricular
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|6361,6377|false|false|false|C0507618|Wall of ventricle|ventricular wall
Finding|Finding|Family Medical History|6361,6387|false|false|false|C2024242|cardiac evaluation of ventricular wall thickness|ventricular wall thickness
Event|Event|Family Medical History|6378,6387|false|false|false|||thickness
Anatomy|Body Space or Junction|Family Medical History|6389,6395|false|false|false|C0333343|Body cavities|cavity
Disorder|Anatomical Abnormality|Family Medical History|6389,6395|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Disorder|Disease or Syndrome|Family Medical History|6389,6395|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Finding|Organ or Tissue Function|Family Medical History|6422,6430|false|false|false|C0039155|Systole|systolic
Event|Event|Family Medical History|6431,6439|false|false|false|||function
Finding|Finding|Family Medical History|6431,6439|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|Family Medical History|6431,6439|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|Family Medical History|6431,6439|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|Family Medical History|6431,6439|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Event|Event|Family Medical History|6444,6450|false|false|false|||normal
Attribute|Clinical Attribute|Family Medical History|6452,6456|false|false|false|C0428772|Left ventricular ejection fraction|LVEF
Event|Event|Family Medical History|6452,6456|false|false|false|||LVEF
Procedure|Diagnostic Procedure|Family Medical History|6452,6456|false|false|false|C3837267|LVEF (procedure)|LVEF
Event|Event|Family Medical History|6487,6491|false|false|false|||beat
Event|Event|Family Medical History|6500,6511|false|false|false|||variability
Finding|Conceptual Entity|Family Medical History|6500,6511|false|false|false|C2827666|Variability|variability
Finding|Functional Concept|Family Medical History|6519,6523|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|6524,6535|false|false|false|C0018827|Heart Ventricle|ventricular
Attribute|Clinical Attribute|Family Medical History|6537,6545|false|false|false|C0812388|Ejection time|ejection
Finding|Daily or Recreational Activity|Family Medical History|6537,6545|false|false|false|C0336969|Ejection as a Sports activity|ejection
Phenomenon|Phenomenon or Process|Family Medical History|6537,6545|false|false|false|C0302131|Ejection as a Circumstance of Injury|ejection
Finding|Finding|Family Medical History|6537,6554|false|false|false|C2020641;C2700378|Ejection fraction;stress echo measurements ejection fraction|ejection fraction
Procedure|Diagnostic Procedure|Family Medical History|6537,6554|false|false|false|C0489482|Ejection fraction (procedure)|ejection fraction
Event|Event|Family Medical History|6546,6554|false|false|false|||fraction
Finding|Intellectual Product|Family Medical History|6546,6554|false|false|false|C1554103|MDFAttributeType - Fraction|fraction
Event|Event|Family Medical History|6575,6581|false|false|false|||rhythm
Finding|Finding|Family Medical History|6575,6581|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|Family Medical History|6575,6581|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Finding|Family Medical History|6582,6591|false|false|false|C0151526;C4018905|Premature Birth;Too early|premature
Finding|Pathologic Function|Family Medical History|6582,6591|false|false|false|C0151526;C4018905|Premature Birth;Too early|premature
Disorder|Disease or Syndrome|Family Medical History|6582,6597|false|false|false|C0340464|Premature Cardiac Complex|premature beats
Event|Event|Family Medical History|6592,6597|false|false|false|||beats
Anatomy|Tissue|Family Medical History|6600,6606|false|false|false|C0040300|Body tissue|Tissue
Finding|Intellectual Product|Family Medical History|6600,6606|false|false|false|C1547928|Tissue Specimen Code|Tissue
Procedure|Diagnostic Procedure|Family Medical History|6607,6614|false|false|false|C0554756|Doppler studies|Doppler
Event|Event|Family Medical History|6615,6622|false|false|false|||imaging
Finding|Finding|Family Medical History|6615,6622|false|false|false|C0740845|Imaging problem|imaging
Procedure|Diagnostic Procedure|Family Medical History|6615,6622|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|imaging
Event|Event|Family Medical History|6623,6631|false|false|false|||suggests
Finding|Functional Concept|Family Medical History|6641,6645|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|6646,6657|false|false|false|C0018827|Heart Ventricle|ventricular
Event|Event|Family Medical History|6667,6675|false|false|false|||pressure
Finding|Finding|Family Medical History|6667,6675|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|Family Medical History|6667,6675|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|Family Medical History|6667,6675|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|Family Medical History|6667,6675|false|false|false|C0033095||pressure
Attribute|Clinical Attribute|Family Medical History|6677,6681|false|false|false|C0034094|Pulmonary Wedge Pressure|PCWP
Finding|Functional Concept|Family Medical History|6691,6696|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|6697,6708|false|false|false|C0018827|Heart Ventricle|ventricular
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|6709,6716|false|false|false|C0935616|chamber [body part]|chamber
Event|Event|Family Medical History|6717,6721|false|false|false|||size
Event|Event|Family Medical History|6727,6731|false|false|false|||free
Finding|Functional Concept|Family Medical History|6727,6731|false|false|false|C0332296|Free of (attribute)|free
Attribute|Clinical Attribute|Family Medical History|6732,6743|false|false|false|C1980023|Wall motion|wall motion
Event|Event|Family Medical History|6737,6743|false|false|false|||motion
Phenomenon|Natural Phenomenon or Process|Family Medical History|6737,6743|false|false|false|C0026597|Motion|motion
Event|Event|Family Medical History|6748,6754|false|false|false|||normal
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|6760,6766|false|false|false|C0003483|Aorta|aortic
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|6760,6772|false|false|false|C0003501;C4533215|Aortic valve structure;Chest>Aortic valve|aortic valve
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|6767,6772|false|false|false|C1186983|Anatomical valve|valve
Event|Event|Family Medical History|6773,6781|false|false|false|||leaflets
Event|Event|Family Medical History|6794,6803|false|false|false|||thickened
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|6822,6828|true|false|false|C0003483|Aorta|aortic
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|6822,6834|true|false|false|C0003501;C4533215|Aortic valve structure;Chest>Aortic valve|aortic valve
Disorder|Congenital Abnormality|Family Medical History|6822,6843|true|false|false|C5193127;C5700069|AORTIC VALVE DISEASE 3;Stenosis of aorta|aortic valve stenosis
Disorder|Disease or Syndrome|Family Medical History|6822,6843|true|false|false|C5193127;C5700069|AORTIC VALVE DISEASE 3;Stenosis of aorta|aortic valve stenosis
Finding|Pathologic Function|Family Medical History|6822,6843|true|false|false|C0003507|Aortic Valve Stenosis|aortic valve stenosis
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|6829,6834|true|false|false|C1186983|Anatomical valve|valve
Event|Event|Family Medical History|6835,6843|true|false|false|||stenosis
Finding|Pathologic Function|Family Medical History|6835,6843|true|false|false|C1261287|Stenosis|stenosis
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|6849,6855|true|false|false|C0003483|Aorta|aortic
Disorder|Disease or Syndrome|Family Medical History|6849,6869|true|false|false|C0003504|Aortic Valve Insufficiency|aortic regurgitation
Event|Event|Family Medical History|6856,6869|true|false|false|||regurgitation
Finding|Finding|Family Medical History|6856,6869|true|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|Family Medical History|6856,6869|true|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|Family Medical History|6856,6869|true|false|false|C0460152|Regurgitation - mechanism|regurgitation
Event|Event|Family Medical History|6873,6877|true|false|false|||seen
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|6883,6895|false|false|false|C0026264|Mitral Valve|mitral valve
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|6890,6895|false|false|false|C1186983|Anatomical valve|valve
Event|Event|Family Medical History|6896,6904|false|false|false|||leaflets
Event|Event|Family Medical History|6917,6926|false|false|false|||thickened
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|6940,6952|true|false|false|C0026264|Mitral Valve|mitral valve
Disorder|Disease or Syndrome|Family Medical History|6940,6961|true|false|false|C0026267|Mitral Valve Prolapse Syndrome|mitral valve prolapse
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|6947,6952|true|false|false|C1186983|Anatomical valve|valve
Disorder|Disease or Syndrome|Family Medical History|6953,6961|true|false|false|C0033377|Ptosis|prolapse
Event|Event|Family Medical History|6953,6961|true|false|false|||prolapse
Finding|Functional Concept|Family Medical History|6963,6974|false|false|false|C0205463|Physiological|Physiologic
Disorder|Disease or Syndrome|Family Medical History|6976,6996|false|false|false|C0026266|Mitral Valve Insufficiency|mitral regurgitation
Event|Event|Family Medical History|6983,6996|false|false|false|||regurgitation
Finding|Finding|Family Medical History|6983,6996|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|Family Medical History|6983,6996|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|Family Medical History|6983,6996|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Event|Event|Family Medical History|7000,7004|false|false|false|||seen
Finding|Finding|Family Medical History|7006,7026|false|false|false|C0442816||within normal limits
Event|Event|Family Medical History|7020,7026|false|false|false|||limits
Finding|Functional Concept|Family Medical History|7020,7026|false|false|false|C0439801|Limited (extensiveness)|limits
Finding|Functional Concept|Family Medical History|7033,7037|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|7039,7050|false|false|false|C0018827|Heart Ventricle|ventricular
Event|Event|Family Medical History|7058,7065|false|false|false|||pattern
Event|Event|Family Medical History|7066,7074|false|false|false|||suggests
Event|Event|Family Medical History|7075,7083|false|false|false|||impaired
Event|Activity|Family Medical History|7084,7094|false|false|false|C0035028|Relaxation|relaxation
Event|Event|Family Medical History|7084,7094|false|false|false|||relaxation
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|7111,7120|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Family Medical History|7111,7120|false|false|false|C2707265||pulmonary
Finding|Finding|Family Medical History|7111,7120|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|7111,7127|false|false|false|C0034052|Pulmonary artery structure|pulmonary artery
Finding|Finding|Family Medical History|7111,7145|false|false|false|C0428643|Pulmonary artery systolic pressure|pulmonary artery systolic pressure
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|7121,7127|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|Family Medical History|7121,7127|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Finding|Organ or Tissue Function|Family Medical History|7128,7136|false|false|false|C0039155|Systole|systolic
Attribute|Clinical Attribute|Family Medical History|7128,7145|false|false|false|C0871470|Systolic Pressure|systolic pressure
Event|Event|Family Medical History|7137,7145|false|false|false|||pressure
Finding|Finding|Family Medical History|7137,7145|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|Family Medical History|7137,7145|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|Family Medical History|7137,7145|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|Family Medical History|7137,7145|false|false|false|C0033095||pressure
Event|Event|Family Medical History|7149,7155|false|false|false|||normal
Anatomy|Body Location or Region|Family Medical History|7170,7181|true|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|7170,7181|true|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Disorder|Disease or Syndrome|Family Medical History|7170,7190|true|false|false|C0031039|Pericardial effusion|pericardial effusion
Finding|Body Substance|Family Medical History|7170,7190|true|false|false|C1253937|Pericardial effusion body substance|pericardial effusion
Event|Event|Family Medical History|7182,7190|true|false|false|||effusion
Finding|Body Substance|Family Medical History|7182,7190|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|Family Medical History|7182,7190|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|Family Medical History|7182,7190|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Event|Event|Family Medical History|7217,7222|false|false|false|||study
Finding|Intellectual Product|Family Medical History|7217,7222|false|false|false|C1705923|Study Object|study
Procedure|Research Activity|Family Medical History|7217,7222|false|false|false|C0008972;C0947630;C2603343|Clinical Research;Scientific Study;Study|study
Event|Event|Family Medical History|7231,7239|false|false|false|||reviewed
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|7259,7265|false|false|false|C0018792|Heart Atrium|atrial
Finding|Pathologic Function|Family Medical History|7259,7272|false|false|false|C0085611|Atrial arrhythmia|atrial ectopy
Event|Event|Family Medical History|7266,7272|false|false|false|||ectopy
Event|Event|Family Medical History|7276,7280|false|false|false|||seen
Finding|Finding|Family Medical History|7296,7304|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|Family Medical History|7296,7304|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|Family Medical History|7296,7304|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|Family Medical History|7296,7304|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Event|Event|Family Medical History|7305,7312|false|false|false|||appears
Event|Event|Family Medical History|7314,7321|false|false|false|||similar
Event|Event|Family Medical History|7327,7332|false|false|false|||Micro
Finding|Conceptual Entity|Family Medical History|7327,7332|false|false|false|C3811161;C4049106|Micro (prefix);Microbiology - Laboratory Class|Micro
Finding|Intellectual Product|Family Medical History|7327,7332|false|false|false|C3811161;C4049106|Micro (prefix);Microbiology - Laboratory Class|Micro
Procedure|Laboratory Procedure|Family Medical History|7327,7332|false|false|false|C0085672|Microbiology procedure|Micro
Event|Event|Family Medical History|7343,7350|false|false|false|||pending
Finding|Idea or Concept|Family Medical History|7343,7350|false|false|false|C1691786;C1704475|Pending - Allergy Clinical Status;Pending - referral status|pending
Event|Event|Hospital Course|7462,7465|false|false|false|||PMH
Finding|Finding|Hospital Course|7462,7465|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|PMH
Disorder|Disease or Syndrome|Hospital Course|7469,7472|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7469,7472|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Hospital Course|7469,7472|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|Hospital Course|7469,7472|false|false|false|||CAD
Finding|Gene or Genome|Hospital Course|7469,7472|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Hospital Course|7469,7472|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Hospital Course|7469,7472|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7469,7472|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Disorder|Disease or Syndrome|Hospital Course|7474,7477|false|false|false|C0085096|Peripheral Vascular Diseases|PVD
Event|Event|Hospital Course|7474,7477|false|false|false|||PVD
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7474,7477|false|false|false|C4521226|Pomalidomide/Bortezomib/Dexamethasone Regimen|PVD
Disorder|Disease or Syndrome|Hospital Course|7483,7487|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Hospital Course|7483,7487|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Hospital Course|7483,7487|false|false|false|||COPD
Finding|Gene or Genome|Hospital Course|7483,7487|false|false|false|C1412502|ARCN1 gene|COPD
Event|Event|Hospital Course|7488,7498|false|false|false|||presenting
Event|Event|Hospital Course|7504,7513|false|false|false|||recurrent
Finding|Sign or Symptom|Hospital Course|7530,7551|false|false|false|C0151826|Retrosternal pain|substernal chest pain
Anatomy|Body Location or Region|Hospital Course|7541,7546|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Hospital Course|7541,7546|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Hospital Course|7541,7551|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|Hospital Course|7541,7551|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Hospital Course|7547,7551|false|true|false|C2598155||pain
Event|Event|Hospital Course|7547,7551|false|false|false|||pain
Finding|Functional Concept|Hospital Course|7547,7551|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|7547,7551|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Body Substance|Hospital Course|7557,7564|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|7557,7564|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|7557,7564|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|Hospital Course|7557,7568|false|false|false|C0332310|Has patient|patient has
Event|Event|Hospital Course|7571,7578|false|false|false|||history
Finding|Conceptual Entity|Hospital Course|7571,7578|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|7571,7578|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Hospital Course|7571,7578|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Intellectual Product|Hospital Course|7583,7587|false|false|false|C1547225|Mild Severity of Illness Code|mild
Disorder|Disease or Syndrome|Hospital Course|7588,7591|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7588,7591|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Hospital Course|7588,7591|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|Hospital Course|7588,7591|false|false|false|||CAD
Finding|Gene or Genome|Hospital Course|7588,7591|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Hospital Course|7588,7591|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Hospital Course|7588,7591|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7588,7591|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Event|Event|Hospital Course|7596,7600|false|false|false|||labs
Lab|Laboratory or Test Result|Hospital Course|7596,7600|false|false|false|C0587081|Laboratory test finding|labs
Event|Event|Hospital Course|7606,7617|false|false|false|||significant
Finding|Idea or Concept|Hospital Course|7606,7617|false|false|false|C0750502|Significant|significant
Finding|Finding|Hospital Course|7618,7630|true|false|false|C0205160|Negative|for negative
Finding|Classification|Hospital Course|7622,7630|true|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|7622,7630|true|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|7622,7630|true|false|false|C5237010|Expression Negative|negative
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7631,7640|true|false|false|C0041199|Troponin|troponins
Drug|Biologically Active Substance|Hospital Course|7631,7640|true|false|false|C0041199|Troponin|troponins
Event|Event|Hospital Course|7631,7640|true|false|false|||troponins
Event|Event|Hospital Course|7646,7649|true|false|false|||EKG
Finding|Intellectual Product|Hospital Course|7646,7649|true|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|Hospital Course|7646,7649|true|false|false|C1623258|Electrocardiography|EKG
Finding|Functional Concept|Hospital Course|7662,7670|true|false|false|C0475224|Ischemic|ischemic
Event|Event|Hospital Course|7671,7678|true|false|false|||changes
Finding|Functional Concept|Hospital Course|7671,7678|true|false|false|C0392747|Changing|changes
Event|Event|Hospital Course|7691,7700|false|false|false|||admission
Procedure|Health Care Activity|Hospital Course|7691,7700|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|Hospital Course|7712,7721|false|false|false|||developed
Event|Event|Hospital Course|7731,7739|false|false|false|||episodes
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7743,7749|false|false|false|C0018792|Heart Atrium|atrial
Disorder|Disease or Syndrome|Hospital Course|7743,7761|false|false|false|C0546959|Atrial tachycardia|atrial tachycardia
Finding|Finding|Hospital Course|7743,7761|false|false|false|C2059391|continuous electrocardiogram atrial tachycardia|atrial tachycardia
Event|Event|Hospital Course|7750,7761|false|false|false|||tachycardia
Finding|Finding|Hospital Course|7750,7761|false|false|false|C0039231;C3827868|Tachycardia;Tachycardia by ECG Finding|tachycardia
Disorder|Disease or Syndrome|Hospital Course|7763,7767|false|false|false|C0004238|Atrial Fibrillation|AFib
Event|Event|Hospital Course|7763,7767|false|false|false|||AFib
Lab|Laboratory or Test Result|Hospital Course|7763,7767|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|AFib
Event|Event|Hospital Course|7791,7798|false|false|false|||started
Drug|Organic Chemical|Hospital Course|7802,7812|false|false|false|C0002598|amiodarone|Amiodarone
Drug|Pharmacologic Substance|Hospital Course|7802,7812|false|false|false|C0002598|amiodarone|Amiodarone
Event|Event|Hospital Course|7802,7812|false|false|false|||Amiodarone
Procedure|Laboratory Procedure|Hospital Course|7802,7812|false|false|false|C5399868|Drug assay amiodarone|Amiodarone
Event|Activity|Hospital Course|7817,7821|false|false|false|C0871208|Rating (action)|rate
Event|Event|Hospital Course|7817,7821|false|false|false|||rate
Finding|Idea or Concept|Hospital Course|7817,7821|false|false|false|C1549480|Amount type - Rate|rate
Finding|Finding|Hospital Course|7822,7828|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|Hospital Course|7822,7828|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Drug|Organic Chemical|Hospital Course|7829,7836|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Pharmacologic Substance|Hospital Course|7829,7836|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Substance|Hospital Course|7829,7836|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Event|Event|Hospital Course|7829,7836|false|false|false|||control
Finding|Conceptual Entity|Hospital Course|7829,7836|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Functional Concept|Hospital Course|7829,7836|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Idea or Concept|Hospital Course|7829,7836|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Drug|Organic Chemical|Hospital Course|7842,7853|false|false|false|C1739768|rivaroxaban|Rivaroxaban
Drug|Pharmacologic Substance|Hospital Course|7842,7853|false|false|false|C1739768|rivaroxaban|Rivaroxaban
Event|Event|Hospital Course|7842,7853|false|false|false|||Rivaroxaban
Event|Event|Hospital Course|7858,7873|false|false|false|||anticoagulation
Finding|Finding|Hospital Course|7858,7873|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Finding|Physiologic Function|Hospital Course|7858,7873|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7858,7873|false|false|false|C0003281|Anticoagulation Therapy|anticoagulation
Event|Event|Hospital Course|7879,7883|false|false|false|||kept
Finding|Idea or Concept|Hospital Course|7887,7891|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|7887,7891|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|7887,7891|false|false|false|C1553498|home health encounter|home
Event|Event|Hospital Course|7892,7896|false|false|false|||dose
Drug|Organic Chemical|Hospital Course|7901,7910|false|false|false|C0012373|diltiazem|Diltiazem
Drug|Pharmacologic Substance|Hospital Course|7901,7910|false|false|false|C0012373|diltiazem|Diltiazem
Event|Activity|Hospital Course|7920,7924|false|false|false|C0871208|Rating (action)|rate
Finding|Idea or Concept|Hospital Course|7920,7924|false|false|false|C1549480|Amount type - Rate|rate
Finding|Functional Concept|Hospital Course|7920,7932|false|false|false|C0489879|rate control|rate control
Drug|Organic Chemical|Hospital Course|7925,7932|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Pharmacologic Substance|Hospital Course|7925,7932|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Substance|Hospital Course|7925,7932|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Event|Event|Hospital Course|7925,7932|false|false|false|||control
Finding|Conceptual Entity|Hospital Course|7925,7932|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Functional Concept|Hospital Course|7925,7932|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Idea or Concept|Hospital Course|7925,7932|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Event|Event|Hospital Course|7955,7963|true|false|false|||episodes
Anatomy|Body Location or Region|Hospital Course|7968,7973|true|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Hospital Course|7968,7973|true|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Hospital Course|7968,7978|true|false|false|C2926613||chest pain
Finding|Sign or Symptom|Hospital Course|7968,7978|true|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Hospital Course|7974,7978|true|false|false|C2598155||pain
Event|Event|Hospital Course|7974,7978|true|false|false|||pain
Finding|Functional Concept|Hospital Course|7974,7978|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|7974,7978|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|7986,8001|true|false|false|||hospitalization
Procedure|Health Care Activity|Hospital Course|7986,8001|true|false|false|C0019993|Hospitalization|hospitalization
Event|Event|Hospital Course|8010,8020|false|false|false|||discharged
Finding|Intellectual Product|Hospital Course|8021,8025|false|false|false|C1720092|Once - dosing instruction fragment|once
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8027,8033|false|false|false|C0018792|Heart Atrium|atrial
Attribute|Clinical Attribute|Hospital Course|8027,8046|false|false|false|C2926591||atrial fibrillation
Disorder|Disease or Syndrome|Hospital Course|8027,8046|false|false|false|C0004238|Atrial Fibrillation|atrial fibrillation
Lab|Laboratory or Test Result|Hospital Course|8027,8046|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|atrial fibrillation
Finding|Pathologic Function|Hospital Course|8027,8054|false|false|false|C0155709|Atrial fibrillation and flutter|atrial fibrillation/flutter
Disorder|Disease or Syndrome|Hospital Course|8034,8046|false|false|false|C0232197|Fibrillation|fibrillation
Event|Event|Hospital Course|8034,8046|false|false|false|||fibrillation
Event|Event|Hospital Course|8047,8054|false|false|false|||flutter
Finding|Pathologic Function|Hospital Course|8047,8054|false|false|false|C0016385|Cardiac Flutter|flutter
Event|Event|Hospital Course|8059,8069|false|false|false|||controlled
Event|Event|Hospital Course|8080,8084|false|false|false|||need
Event|Event|Hospital Course|8089,8095|false|false|false|||follow
Finding|Intellectual Product|Hospital Course|8108,8120|false|false|false|C1547426|Location Service Code - Primary Care|primary care
Procedure|Health Care Activity|Hospital Course|8108,8120|false|false|false|C0033137|Primary Health Care|primary care
Event|Activity|Hospital Course|8116,8120|false|false|false|C1947933|care activity|care
Event|Event|Hospital Course|8116,8120|false|false|false|||care
Finding|Finding|Hospital Course|8116,8120|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Hospital Course|8116,8120|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Hospital Course|8121,8127|false|false|false|C2348314|Doctor - Title|doctor
Anatomy|Body Location or Region|Hospital Course|8144,8149|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Hospital Course|8144,8149|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Hospital Course|8151,8155|false|false|false|C2598155||pain
Event|Event|Hospital Course|8151,8155|false|false|false|||pain
Finding|Functional Concept|Hospital Course|8151,8155|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|8151,8155|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|8169,8178|false|false|false|||admission
Procedure|Health Care Activity|Hospital Course|8169,8178|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Intellectual Product|Hospital Course|8181,8186|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|Acute
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8253,8259|false|false|false|C0018792|Heart Atrium|Atrial
Disorder|Disease or Syndrome|Hospital Course|8253,8271|false|false|false|C0546959|Atrial tachycardia|Atrial Tachycardia
Finding|Finding|Hospital Course|8253,8271|false|false|false|C2059391|continuous electrocardiogram atrial tachycardia|Atrial Tachycardia
Event|Event|Hospital Course|8260,8271|false|false|false|||Tachycardia
Finding|Finding|Hospital Course|8260,8271|false|false|false|C0039231;C3827868|Tachycardia;Tachycardia by ECG Finding|Tachycardia
Event|Event|Hospital Course|8280,8289|false|false|false|||admission
Procedure|Health Care Activity|Hospital Course|8280,8289|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|Hospital Course|8297,8301|false|false|false|||runs
Finding|Finding|Hospital Course|8297,8301|false|false|false|C0600140|Does run (finding)|runs
Drug|Chemical Viewed Structurally|Hospital Course|8311,8318|false|false|false|C1704241|complex (molecular entity)|complex
Event|Event|Hospital Course|8319,8333|false|false|false|||tachyarrythmia
Finding|Idea or Concept|Hospital Course|8335,8342|false|false|false|C0039869;C4319827|Thought|thought
Finding|Mental Process|Hospital Course|8335,8342|false|false|false|C0039869;C4319827|Thought|thought
Finding|Finding|Hospital Course|8343,8349|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Hospital Course|8343,8349|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|Hospital Course|8371,8377|false|false|false|||origin
Finding|Classification|Hospital Course|8371,8377|false|false|false|C0079946;C1550512|National origin;Participation Type - origin|origin
Finding|Intellectual Product|Hospital Course|8371,8377|false|false|false|C0079946;C1550512|National origin;Participation Type - origin|origin
Disorder|Disease or Syndrome|Hospital Course|8379,8404|false|false|false|C1281999|Rapid atrial fibrillation|rapid Atrial Fibrillation
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8385,8391|false|false|false|C0018792|Heart Atrium|Atrial
Attribute|Clinical Attribute|Hospital Course|8385,8404|false|false|false|C2926591||Atrial Fibrillation
Disorder|Disease or Syndrome|Hospital Course|8385,8404|false|false|false|C0004238|Atrial Fibrillation|Atrial Fibrillation
Lab|Laboratory or Test Result|Hospital Course|8385,8404|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Atrial Fibrillation
Finding|Pathologic Function|Hospital Course|8385,8413|false|false|false|C0155709|Atrial fibrillation and flutter|Atrial Fibrillation/ Flutter
Disorder|Disease or Syndrome|Hospital Course|8392,8404|false|false|false|C0232197|Fibrillation|Fibrillation
Event|Event|Hospital Course|8392,8404|false|false|false|||Fibrillation
Finding|Pathologic Function|Hospital Course|8406,8413|false|false|false|C0016385|Cardiac Flutter|Flutter
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8418,8424|false|false|false|C0018792|Heart Atrium|atrial
Event|Event|Hospital Course|8426,8437|false|false|false|||tachycardia
Finding|Finding|Hospital Course|8426,8437|false|false|false|C0039231;C3827868|Tachycardia;Tachycardia by ECG Finding|tachycardia
Drug|Chemical Viewed Structurally|Hospital Course|8455,8464|false|false|false|C1704241|complex (molecular entity)|complexes
Event|Event|Hospital Course|8455,8464|false|false|false|||complexes
Event|Event|Hospital Course|8478,8488|false|false|false|||morphology
Finding|Finding|Hospital Course|8478,8488|false|false|false|C0700329|Physical shape|morphology
Finding|Functional Concept|Hospital Course|8493,8499|false|false|false|C0302891|Native (qualifier value)|native
Disorder|Disease or Syndrome|Hospital Course|8500,8504|false|false|false|C0023211|Left Bundle-Branch Block|LBBB
Event|Event|Hospital Course|8500,8504|false|false|false|||LBBB
Lab|Laboratory or Test Result|Hospital Course|8500,8504|false|false|false|C0344420||LBBB
Event|Event|Hospital Course|8515,8522|false|false|false|||treated
Drug|Organic Chemical|Hospital Course|8528,8537|false|false|false|C0012373|diltiazem|Diltiazem
Drug|Pharmacologic Substance|Hospital Course|8528,8537|false|false|false|C0012373|diltiazem|Diltiazem
Event|Event|Hospital Course|8528,8537|false|false|false|||Diltiazem
Drug|Organic Chemical|Hospital Course|8542,8552|false|false|false|C0002598|amiodarone|Amiodarone
Drug|Pharmacologic Substance|Hospital Course|8542,8552|false|false|false|C0002598|amiodarone|Amiodarone
Event|Event|Hospital Course|8542,8552|false|false|false|||Amiodarone
Procedure|Laboratory Procedure|Hospital Course|8542,8552|false|false|false|C5399868|Drug assay amiodarone|Amiodarone
Event|Event|Hospital Course|8568,8576|false|false|false|||episodes
Event|Event|Hospital Course|8580,8591|false|false|false|||tachycardia
Finding|Finding|Hospital Course|8580,8591|false|false|false|C0039231;C3827868|Tachycardia;Tachycardia by ECG Finding|tachycardia
Event|Event|Hospital Course|8601,8610|false|false|false|||evaluated
Finding|Body Substance|Hospital Course|8611,8618|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|8611,8618|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|8611,8618|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|8624,8635|false|false|false|||recommended
Event|Event|Hospital Course|8636,8651|false|false|false|||anticoagulation
Finding|Finding|Hospital Course|8636,8651|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Finding|Physiologic Function|Hospital Course|8636,8651|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8636,8651|false|false|false|C0003281|Anticoagulation Therapy|anticoagulation
Finding|Classification|Hospital Course|8656,8666|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|8656,8666|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|Hospital Course|8667,8673|false|false|false|||follow
Finding|Functional Concept|Hospital Course|8667,8673|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|Hospital Course|8667,8673|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|Hospital Course|8667,8676|false|false|false|C0589120|Follow-up status|follow up
Procedure|Health Care Activity|Hospital Course|8667,8676|false|false|false|C1522577|follow-up|follow up
Event|Event|Hospital Course|8681,8689|false|false|false|||consider
Procedure|Diagnostic Procedure|Hospital Course|8690,8698|false|false|false|C5551547|Cardiac electrophysiology study|EP study
Event|Event|Hospital Course|8693,8698|false|false|false|||study
Finding|Intellectual Product|Hospital Course|8693,8698|false|false|false|C1705923|Study Object|study
Procedure|Research Activity|Hospital Course|8693,8698|false|false|false|C0008972;C0947630;C2603343|Clinical Research;Scientific Study;Study|study
Finding|Finding|Hospital Course|8703,8711|false|false|false|C0332149|Possible|possible
Event|Event|Hospital Course|8712,8720|false|false|false|||ablation
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8712,8720|false|false|false|C0547070;C1261381|Ablation;Destructive procedure (surgical)|ablation
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8724,8730|false|false|false|C0018792|Heart Atrium|Atrial
Finding|Pathologic Function|Hospital Course|8724,8738|false|false|false|C0004239|Atrial Flutter|Atrial Flutter
Lab|Laboratory or Test Result|Hospital Course|8724,8738|false|false|false|C0344423|Atrial Flutter by ECG Finding|Atrial Flutter
Event|Event|Hospital Course|8731,8738|false|false|false|||Flutter
Finding|Pathologic Function|Hospital Course|8731,8738|false|false|false|C0016385|Cardiac Flutter|Flutter
Finding|Body Substance|Hospital Course|8741,8748|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|8741,8748|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|8741,8748|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Hospital Course|8753,8763|false|false|false|||discharged
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8776,8782|false|false|false|C0018787|Heart|Hearts
Drug|Hazardous or Poisonous Substance|Hospital Course|8783,8790|false|false|false|C0728873|Monitor brand of insecticide|monitor
Drug|Organic Chemical|Hospital Course|8783,8790|false|false|false|C0728873|Monitor brand of insecticide|monitor
Event|Event|Hospital Course|8783,8790|false|false|false|||monitor
Drug|Organic Chemical|Hospital Course|8792,8802|false|false|false|C0002598|amiodarone|Amiodarone
Drug|Pharmacologic Substance|Hospital Course|8792,8802|false|false|false|C0002598|amiodarone|Amiodarone
Event|Event|Hospital Course|8792,8802|false|false|false|||Amiodarone
Procedure|Laboratory Procedure|Hospital Course|8792,8802|false|false|false|C5399868|Drug assay amiodarone|Amiodarone
Event|Event|Hospital Course|8826,8830|false|false|false|||week
Finding|Intellectual Product|Hospital Course|8826,8830|false|false|false|C1561540|Transaction counts and value totals - week|week
Drug|Organic Chemical|Hospital Course|8869,8878|false|false|false|C0012373|diltiazem|Diltiazem
Drug|Pharmacologic Substance|Hospital Course|8869,8878|false|false|false|C0012373|diltiazem|Diltiazem
Event|Event|Hospital Course|8879,8888|false|false|false|||continued
Finding|Finding|Hospital Course|8889,8896|false|false|false|C4534363|At home|at home
Finding|Idea or Concept|Hospital Course|8892,8896|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|8892,8896|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|8892,8896|false|false|false|C1553498|home health encounter|home
Event|Event|Hospital Course|8897,8901|false|false|false|||dose
Drug|Organic Chemical|Hospital Course|8903,8914|false|false|false|C1739768|rivaroxaban|Rivaroxaban
Drug|Pharmacologic Substance|Hospital Course|8903,8914|false|false|false|C1739768|rivaroxaban|Rivaroxaban
Event|Event|Hospital Course|8915,8920|false|false|false|||added
Event|Event|Hospital Course|8926,8941|false|false|false|||anticoagulation
Finding|Finding|Hospital Course|8926,8941|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Finding|Physiologic Function|Hospital Course|8926,8941|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8926,8941|false|false|false|C0003281|Anticoagulation Therapy|anticoagulation
Finding|Classification|Hospital Course|8950,8960|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|8950,8960|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|Hospital Course|8961,8973|false|false|false|||cardiologist
Drug|Organic Chemical|Hospital Course|8985,8991|false|false|false|C0633084|Plavix|plavix
Drug|Pharmacologic Substance|Hospital Course|8985,8991|false|false|false|C0633084|Plavix|plavix
Event|Event|Hospital Course|8985,8991|false|false|false|||plavix
Event|Event|Hospital Course|8996,9008|false|false|false|||discontinued
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9012,9017|false|false|false|C1570446|TNFSF14 protein, human|light
Drug|Biologically Active Substance|Hospital Course|9012,9017|false|false|false|C1570446|TNFSF14 protein, human|light
Event|Event|Hospital Course|9012,9017|false|false|false|||light
Finding|Finding|Hospital Course|9012,9017|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Functional Concept|Hospital Course|9012,9017|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Gene or Genome|Hospital Course|9012,9017|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Phenomenon|Natural Phenomenon or Process|Hospital Course|9012,9017|false|false|false|C0023693|Light|light
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9012,9017|false|false|false|C0031765|Phototherapy|light
Event|Event|Hospital Course|9021,9029|false|false|false|||addition
Finding|Functional Concept|Hospital Course|9021,9029|false|false|false|C0332287;C1883712|Add - instruction imperative;In addition to|addition
Drug|Organic Chemical|Hospital Course|9033,9044|false|false|false|C1739768|rivaroxaban|Rivaroxaban
Drug|Pharmacologic Substance|Hospital Course|9033,9044|false|false|false|C1739768|rivaroxaban|Rivaroxaban
Event|Event|Hospital Course|9050,9058|false|false|false|||interest
Finding|Mental Process|Hospital Course|9050,9058|false|false|false|C0543488|Interested|interest
Event|Event|Hospital Course|9078,9085|false|false|false|||therapy
Finding|Finding|Hospital Course|9078,9085|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|Hospital Course|9078,9085|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9078,9085|false|false|false|C0087111|Therapeutic procedure|therapy
Finding|Body Substance|Hospital Course|9094,9101|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|9094,9101|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|9094,9101|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|9117,9123|false|false|false|||follow
Event|Activity|Hospital Course|9127,9139|false|false|false|C0003629|Appointments|appointments
Event|Event|Hospital Course|9127,9139|false|false|false|||appointments
Event|Event|Hospital Course|9164,9173|false|false|false|||scheduled
Event|Event|Hospital Course|9177,9180|false|false|false|||see
Event|Event|Hospital Course|9192,9202|false|false|false|||evaluation
Finding|Idea or Concept|Hospital Course|9192,9202|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|Hospital Course|9192,9202|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Anatomy|Body Location or Region|Hospital Course|9218,9223|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|Hospital Course|9218,9223|false|false|false|C0741025|Chest problem|Chest
Attribute|Clinical Attribute|Hospital Course|9218,9228|false|false|false|C2926613||Chest pain
Finding|Sign or Symptom|Hospital Course|9218,9228|false|false|false|C0008031|Chest Pain|Chest pain
Attribute|Clinical Attribute|Hospital Course|9224,9228|false|false|false|C2598155||pain
Event|Event|Hospital Course|9224,9228|false|false|false|||pain
Finding|Functional Concept|Hospital Course|9224,9228|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|9224,9228|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|9233,9242|false|false|false|||presented
Finding|Sign or Symptom|Hospital Course|9248,9269|false|false|false|C0151826|Retrosternal pain|substernal chest pain
Anatomy|Body Location or Region|Hospital Course|9259,9264|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Hospital Course|9259,9264|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Hospital Course|9259,9269|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|Hospital Course|9259,9269|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Hospital Course|9265,9269|false|true|false|C2598155||pain
Event|Event|Hospital Course|9265,9269|false|false|false|||pain
Finding|Functional Concept|Hospital Course|9265,9269|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|9265,9269|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|9276,9284|true|false|false|||occurred
Finding|Functional Concept|Hospital Course|9285,9292|true|false|false|C0443144|At rest (qualifier value)|at rest
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9288,9292|true|false|false|C1742913|REST protein, human|rest
Drug|Biologically Active Substance|Hospital Course|9288,9292|true|false|false|C1742913|REST protein, human|rest
Finding|Daily or Recreational Activity|Hospital Course|9288,9292|true|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Gene or Genome|Hospital Course|9288,9292|true|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Molecular Function|Hospital Course|9288,9292|true|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Event|Event|Hospital Course|9301,9306|true|false|false|||ruled
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9326,9334|true|false|false|C0041199|Troponin|troponin
Drug|Biologically Active Substance|Hospital Course|9326,9334|true|false|false|C0041199|Troponin|troponin
Event|Event|Hospital Course|9326,9334|true|false|false|||troponin
Procedure|Laboratory Procedure|Hospital Course|9326,9334|true|false|false|C0523952|Troponin measurement|troponin
Event|Event|Hospital Course|9336,9345|true|false|false|||elevation
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9336,9345|true|false|false|C0439775|Elevation procedure|elevation
Event|Event|Hospital Course|9349,9360|true|false|false|||significant
Finding|Idea or Concept|Hospital Course|9349,9360|true|false|false|C0750502|Significant|significant
Finding|Finding|Hospital Course|9361,9364|true|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Hospital Course|9361,9364|true|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9365,9368|true|false|false|C0018064|Equine Gonadotropins|ECG
Drug|Hormone|Hospital Course|9365,9368|true|false|false|C0018064|Equine Gonadotropins|ECG
Drug|Pharmacologic Substance|Hospital Course|9365,9368|true|false|false|C0018064|Equine Gonadotropins|ECG
Event|Event|Hospital Course|9365,9368|true|false|false|||ECG
Finding|Intellectual Product|Hospital Course|9365,9368|true|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|ECG
Procedure|Diagnostic Procedure|Hospital Course|9365,9368|true|false|false|C1623258|Electrocardiography|ECG
Event|Event|Hospital Course|9369,9376|false|false|false|||changes
Finding|Functional Concept|Hospital Course|9369,9376|false|false|false|C0392747|Changing|changes
Anatomy|Body Location or Region|Hospital Course|9389,9394|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Hospital Course|9389,9394|false|true|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Hospital Course|9389,9399|false|true|false|C2926613||chest pain
Finding|Sign or Symptom|Hospital Course|9389,9399|false|true|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Hospital Course|9395,9399|false|true|false|C2598155||pain
Event|Event|Hospital Course|9395,9399|false|false|false|||pain
Finding|Functional Concept|Hospital Course|9395,9399|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|9395,9399|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|9405,9412|false|false|false|||related
Event|Event|Hospital Course|9416,9423|false|false|false|||periods
Finding|Organism Function|Hospital Course|9416,9423|false|false|false|C0025344|Menstruation|periods
Event|Event|Hospital Course|9427,9438|false|false|false|||tachycardia
Finding|Finding|Hospital Course|9427,9438|false|false|false|C0039231;C3827868|Tachycardia;Tachycardia by ECG Finding|tachycardia
Finding|Idea or Concept|Hospital Course|9463,9471|true|false|false|C1547192|Organization unit type - Hospital|hospital
Finding|Sign or Symptom|Hospital Course|9472,9480|true|false|false|C0011991|Diarrhea|the runs
Finding|Finding|Hospital Course|9476,9480|true|false|false|C0600140|Does run (finding)|runs
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9484,9490|true|false|false|C0018792|Heart Atrium|atrial
Disorder|Disease or Syndrome|Hospital Course|9484,9502|true|false|false|C0546959|Atrial tachycardia|atrial tachycardia
Finding|Finding|Hospital Course|9484,9502|true|false|false|C2059391|continuous electrocardiogram atrial tachycardia|atrial tachycardia
Event|Event|Hospital Course|9491,9502|true|false|false|||tachycardia
Finding|Finding|Hospital Course|9491,9502|true|false|false|C0039231;C3827868|Tachycardia;Tachycardia by ECG Finding|tachycardia
Event|Event|Hospital Course|9511,9520|true|false|false|||reproduce
Anatomy|Body Location or Region|Hospital Course|9521,9526|true|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Hospital Course|9521,9526|true|true|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Hospital Course|9528,9532|true|false|false|C2598155||pain
Event|Event|Hospital Course|9528,9532|true|false|false|||pain
Finding|Functional Concept|Hospital Course|9528,9532|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|9528,9532|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|9555,9563|true|false|false|||episodes
Anatomy|Body Location or Region|Hospital Course|9567,9572|true|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Hospital Course|9567,9572|true|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Hospital Course|9567,9577|true|false|false|C2926613||chest pain
Finding|Sign or Symptom|Hospital Course|9567,9577|true|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Hospital Course|9573,9577|true|false|false|C2598155||pain
Event|Event|Hospital Course|9573,9577|true|false|false|||pain
Finding|Functional Concept|Hospital Course|9573,9577|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|9573,9577|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|9586,9601|true|false|false|||hospitalization
Procedure|Health Care Activity|Hospital Course|9586,9601|true|false|false|C0019993|Hospitalization|hospitalization
Event|Event|Hospital Course|9610,9620|false|false|false|||discharged
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9626,9632|false|false|false|C0018792|Heart Atrium|atrial
Disorder|Disease or Syndrome|Hospital Course|9634,9646|false|false|false|C0232197|Fibrillation|fibrillation
Event|Event|Hospital Course|9634,9646|false|false|false|||fibrillation
Event|Event|Hospital Course|9647,9654|false|false|false|||flutter
Finding|Pathologic Function|Hospital Course|9647,9654|false|false|false|C0016385|Cardiac Flutter|flutter
Event|Event|Hospital Course|9659,9669|false|false|false|||controlled
Event|Event|Hospital Course|9680,9684|false|false|false|||need
Event|Event|Hospital Course|9688,9694|false|false|false|||follow
Finding|Intellectual Product|Hospital Course|9708,9720|false|false|false|C1547426|Location Service Code - Primary Care|primary care
Procedure|Health Care Activity|Hospital Course|9708,9720|false|false|false|C0033137|Primary Health Care|primary care
Event|Activity|Hospital Course|9716,9720|false|false|false|C1947933|care activity|care
Event|Event|Hospital Course|9716,9720|false|false|false|||care
Finding|Finding|Hospital Course|9716,9720|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Hospital Course|9716,9720|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Hospital Course|9721,9727|false|false|false|C2348314|Doctor - Title|doctor
Anatomy|Body Location or Region|Hospital Course|9744,9749|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Hospital Course|9744,9749|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Hospital Course|9744,9754|false|true|false|C2926613||chest pain
Finding|Sign or Symptom|Hospital Course|9744,9754|false|true|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Hospital Course|9750,9754|false|true|false|C2598155||pain
Event|Event|Hospital Course|9750,9754|false|false|false|||pain
Finding|Functional Concept|Hospital Course|9750,9754|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|9750,9754|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|9762,9765|false|false|false|||led
Event|Event|Hospital Course|9769,9778|false|false|false|||admission
Procedure|Health Care Activity|Hospital Course|9769,9778|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Disorder|Disease or Syndrome|Hospital Course|9782,9790|false|false|false|C0013238;C0022575|Dry Eye Syndromes;Keratoconjunctivitis Sicca|Dry eyes
Drug|Pharmacologic Substance|Hospital Course|9782,9790|false|false|false|C0720056|Dry Eyes brand of ocular lubricant|Dry eyes
Finding|Sign or Symptom|Hospital Course|9782,9790|false|false|false|C0314719|Dryness of eye|Dry eyes
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9786,9790|false|false|false|C0015392|Eye|eyes
Attribute|Clinical Attribute|Hospital Course|9786,9790|false|false|false|C5848506||eyes
Event|Event|Hospital Course|9786,9790|false|false|false|||eyes
Disorder|Disease or Syndrome|Hospital Course|9799,9807|false|false|false|C0041834|Erythema|erythema
Event|Event|Hospital Course|9799,9807|false|false|false|||erythema
Attribute|Clinical Attribute|Hospital Course|9812,9816|false|false|false|C2598155||pain
Event|Event|Hospital Course|9812,9816|false|false|false|||pain
Finding|Functional Concept|Hospital Course|9812,9816|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|9812,9816|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|Hospital Course|9820,9825|false|false|false|C5886197||R eye
Anatomy|Body Location or Region|Hospital Course|9822,9825|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|eye
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9822,9825|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|eye
Disorder|Disease or Syndrome|Hospital Course|9822,9825|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|eye
Disorder|Neoplastic Process|Hospital Course|9822,9825|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|eye
Finding|Body Substance|Hospital Course|9822,9825|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Finding|Hospital Course|9822,9825|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Intellectual Product|Hospital Course|9822,9825|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Event|Event|Hospital Course|9827,9832|false|false|false|||found
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9846,9850|false|false|false|C0015392|Eye|eyes
Attribute|Clinical Attribute|Hospital Course|9846,9850|false|false|false|C5848506||eyes
Event|Event|Hospital Course|9855,9867|false|false|false|||optholmology
Event|Event|Hospital Course|9869,9873|false|false|false|||Sent
Drug|Pharmacologic Substance|Hospital Course|9883,9899|false|false|false|C0003921;C2608262;C3853661|Artificial Tears;Lubricant Eye Drops;artificial tears (medication)|Artificial tears
Event|Event|Hospital Course|9894,9899|false|false|false|||tears
Finding|Body Substance|Hospital Course|9894,9899|false|false|false|C0039409;C1547924;C1611838|Tears (substance);Tears specimen|tears
Finding|Intellectual Product|Hospital Course|9894,9899|false|false|false|C0039409;C1547924;C1611838|Tears (substance);Tears specimen|tears
Drug|Antibiotic|Hospital Course|9905,9917|false|false|false|C0014806|erythromycin|erythromycin
Drug|Organic Chemical|Hospital Course|9905,9917|false|false|false|C0014806|erythromycin|erythromycin
Event|Event|Hospital Course|9905,9917|false|false|false|||erythromycin
Anatomy|Body Location or Region|Hospital Course|9918,9921|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|eye
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9918,9921|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|eye
Disorder|Disease or Syndrome|Hospital Course|9918,9921|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|eye
Disorder|Neoplastic Process|Hospital Course|9918,9921|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|eye
Finding|Body Substance|Hospital Course|9918,9921|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Finding|Hospital Course|9918,9921|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Intellectual Product|Hospital Course|9918,9921|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Drug|Biomedical or Dental Material|Hospital Course|9918,9927|false|false|false|C0015399;C1154269|Eye Drops;Eye drops brand of Tetrahydrozoline|eye drops
Drug|Organic Chemical|Hospital Course|9918,9927|false|false|false|C0015399;C1154269|Eye Drops;Eye drops brand of Tetrahydrozoline|eye drops
Drug|Pharmacologic Substance|Hospital Course|9918,9927|false|false|false|C0015399;C1154269|Eye Drops;Eye drops brand of Tetrahydrozoline|eye drops
Drug|Biomedical or Dental Material|Hospital Course|9922,9927|false|false|false|C0991568|Drops - Drug Form|drops
Event|Event|Hospital Course|9922,9927|false|false|false|||drops
Finding|Body Substance|Hospital Course|9929,9936|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|9929,9936|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|9929,9936|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Hospital Course|9941,9947|false|false|false|||follow
Event|Activity|Hospital Course|9951,9962|false|false|false|C0003629|Appointments|appointment
Event|Event|Hospital Course|9951,9962|false|false|false|||appointment
Event|Event|Hospital Course|9972,9981|false|false|false|||scheduled
Event|Event|Hospital Course|10008,10018|false|false|false|||instructed
Event|Event|Hospital Course|10022,10028|false|false|false|||attend
Finding|Functional Concept|Hospital Course|10022,10028|false|false|false|C1999232|Attending (action)|attend
Event|Activity|Hospital Course|10030,10041|false|false|false|C0003629|Appointments|appointment
Event|Event|Hospital Course|10030,10041|false|false|false|||appointment
Finding|Intellectual Product|Hospital Course|10044,10051|false|false|false|C1547296|Chronic - Admission Level of Care Code|Chronic
Procedure|Health Care Activity|Hospital Course|10044,10051|false|false|false|C1555457|Provision of recurring care for chronic illness|Chronic
Disorder|Disease or Syndrome|Hospital Course|10124,10128|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Hospital Course|10124,10128|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Hospital Course|10124,10128|false|false|false|||COPD
Finding|Gene or Genome|Hospital Course|10124,10128|false|false|false|C1412502|ARCN1 gene|COPD
Event|Event|Hospital Course|10130,10132|false|false|false|||Pt
Drug|Biomedical or Dental Material|Hospital Course|10151,10159|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|Hospital Course|10151,10159|false|false|false|||baseline
Finding|Idea or Concept|Hospital Course|10151,10159|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Attribute|Clinical Attribute|Hospital Course|10160,10171|false|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|Hospital Course|10160,10171|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|Hospital Course|10160,10171|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|Hospital Course|10160,10171|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Attribute|Clinical Attribute|Hospital Course|10160,10178|false|false|false|C2598168||respiratory status
Finding|Finding|Hospital Course|10160,10178|false|false|false|C1998827|Respiratory Status|respiratory status
Attribute|Clinical Attribute|Hospital Course|10172,10178|false|false|false|C5889824||status
Event|Event|Hospital Course|10172,10178|false|false|false|||status
Finding|Idea or Concept|Hospital Course|10172,10178|false|false|false|C1546481|What subject filter - Status|status
Event|Event|Hospital Course|10189,10193|false|false|false|||sent
Event|Event|Hospital Course|10194,10198|false|false|false|||home
Finding|Idea or Concept|Hospital Course|10194,10198|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|10194,10198|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|10194,10198|false|false|false|C1553498|home health encounter|home
Finding|Idea or Concept|Hospital Course|10208,10212|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|10208,10212|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|10208,10212|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Hospital Course|10213,10222|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|Hospital Course|10213,10222|false|false|false|C0001927|albuterol|albuterol
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10223,10226|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|neb
Drug|Biologically Active Substance|Hospital Course|10223,10226|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|neb
Drug|Biomedical or Dental Material|Hospital Course|10223,10226|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|neb
Event|Event|Hospital Course|10223,10226|false|false|false|||neb
Finding|Cell Function|Hospital Course|10223,10226|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|neb
Finding|Gene or Genome|Hospital Course|10223,10226|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|neb
Drug|Organic Chemical|Hospital Course|10228,10237|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|Hospital Course|10228,10237|false|false|false|C0001927|albuterol|albuterol
Event|Event|Hospital Course|10238,10245|false|false|false|||inhaler
Finding|Functional Concept|Hospital Course|10238,10245|false|false|false|C4319647|Inhaler (unit of presentation)|inhaler
Drug|Organic Chemical|Hospital Course|10248,10259|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Hospital Course|10248,10259|false|false|false|C0082607|fluticasone|Fluticasone
Event|Event|Hospital Course|10248,10259|false|false|false|||Fluticasone
Drug|Clinical Drug|Hospital Course|10248,10265|false|false|false|C0360577||Fluticasone nasal
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10260,10265|false|false|false|C0028429||nasal
Drug|Biomedical or Dental Material|Hospital Course|10260,10265|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Organic Chemical|Hospital Course|10260,10265|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Pharmacologic Substance|Hospital Course|10260,10265|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Finding|Finding|Hospital Course|10260,10265|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Functional Concept|Hospital Course|10260,10265|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Drug|Pharmacologic Substance|Hospital Course|10260,10271|false|false|false|C2608294|Nasal Spray brand of phenylephrine|nasal spray
Drug|Biomedical or Dental Material|Hospital Course|10266,10271|false|false|false|C1154182|Spray Dosage Form|spray
Event|Activity|Hospital Course|10266,10271|false|false|false|C2003858|Spray (action)|spray
Event|Event|Hospital Course|10266,10271|false|false|false|||spray
Finding|Functional Concept|Hospital Course|10266,10271|false|false|false|C4521772|Spray (administration method)|spray
Drug|Organic Chemical|Hospital Course|10273,10284|false|false|false|C0082607|fluticasone|fluticasone
Drug|Pharmacologic Substance|Hospital Course|10273,10284|false|false|false|C0082607|fluticasone|fluticasone
Event|Event|Hospital Course|10273,10284|false|false|false|||fluticasone
Drug|Pharmacologic Substance|Hospital Course|10273,10295|false|false|false|C0939232|fluticasone / salmeterol|fluticasone-salmeterol
Drug|Organic Chemical|Hospital Course|10273,10302|false|false|false|C4762496|Fluticasone-Salmeterol Diskus|fluticasone-salmeterol diskus
Drug|Pharmacologic Substance|Hospital Course|10273,10302|false|false|false|C4762496|Fluticasone-Salmeterol Diskus|fluticasone-salmeterol diskus
Drug|Organic Chemical|Hospital Course|10285,10295|false|false|false|C0073992|salmeterol|salmeterol
Drug|Pharmacologic Substance|Hospital Course|10285,10295|false|false|false|C0073992|salmeterol|salmeterol
Event|Event|Hospital Course|10296,10302|false|false|false|||diskus
Drug|Organic Chemical|Hospital Course|10305,10315|false|false|false|C0213771|tiotropium|tiotropium
Drug|Pharmacologic Substance|Hospital Course|10305,10315|false|false|false|C0213771|tiotropium|tiotropium
Event|Event|Hospital Course|10305,10315|false|false|false|||tiotropium
Drug|Organic Chemical|Hospital Course|10305,10323|false|false|false|C1306772|tiotropium bromide|tiotropium bromide
Drug|Pharmacologic Substance|Hospital Course|10305,10323|false|false|false|C1306772|tiotropium bromide|tiotropium bromide
Drug|Inorganic Chemical|Hospital Course|10316,10323|false|false|false|C0006222|Bromides|bromide
Event|Event|Hospital Course|10316,10323|false|false|false|||bromide
Procedure|Laboratory Procedure|Hospital Course|10316,10323|false|false|false|C0202341|Bromides measurement|bromide
Drug|Biomedical or Dental Material|Hospital Course|10324,10328|false|false|false|C1300458|Nebulizer solution|nebs
Event|Event|Hospital Course|10324,10328|false|false|false|||nebs
Drug|Organic Chemical|Hospital Course|10334,10346|false|false|false|C0039771|theophylline|theophylline
Drug|Pharmacologic Substance|Hospital Course|10334,10346|false|false|false|C0039771|theophylline|theophylline
Event|Event|Hospital Course|10334,10346|false|false|false|||theophylline
Procedure|Laboratory Procedure|Hospital Course|10334,10346|false|false|false|C0039773|Assay of theophylline|theophylline
Anatomy|Anatomical Structure|Hospital Course|10350,10353|false|false|false|C3669270|Strucure of thick cushion of skin|PAD
Disorder|Disease or Syndrome|Hospital Course|10350,10353|false|false|false|C0332568;C1704436|Pad Mass;Peripheral Arterial Diseases|PAD
Disorder|Neoplastic Process|Hospital Course|10350,10353|false|false|false|C0332568;C1704436|Pad Mass;Peripheral Arterial Diseases|PAD
Drug|Biomedical or Dental Material|Hospital Course|10350,10353|false|false|false|C2347441|Pad Dosage Form|PAD
Event|Event|Hospital Course|10350,10353|false|false|false|||PAD
Finding|Gene or Genome|Hospital Course|10350,10353|false|false|false|C1425244;C1425478;C3540603|DHX40 gene;PADI4 gene;PADI4 wt Allele|PAD
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10350,10353|false|false|false|C3814046|PAD Regimen|PAD
Finding|Idea or Concept|Hospital Course|10359,10364|false|false|false|C1552828|Table Frame - above|above
Event|Event|Hospital Course|10369,10376|false|false|false|||stopped
Drug|Organic Chemical|Hospital Course|10377,10388|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Pharmacologic Substance|Hospital Course|10377,10388|false|false|false|C0070166|clopidogrel|Clopidogrel
Event|Event|Hospital Course|10377,10388|false|false|false|||Clopidogrel
Finding|Body Substance|Hospital Course|10392,10399|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|10392,10399|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|10392,10399|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Organic Chemical|Hospital Course|10411,10422|false|false|false|C1739768|rivaroxaban|Rivaroxaban
Drug|Pharmacologic Substance|Hospital Course|10411,10422|false|false|false|C1739768|rivaroxaban|Rivaroxaban
Event|Event|Hospital Course|10427,10433|false|false|false|||wanted
Event|Event|Hospital Course|10437,10442|false|false|false|||avoid
Event|Event|Hospital Course|10450,10457|false|false|false|||therapy
Finding|Finding|Hospital Course|10450,10457|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|Hospital Course|10450,10457|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10450,10457|false|false|false|C0087111|Therapeutic procedure|therapy
Finding|Idea or Concept|Hospital Course|10493,10505|false|false|false|C1548597|Marketing basis - Transitional|Transitional
Finding|Body Substance|Hospital Course|10580,10587|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|10580,10587|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|10580,10587|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Hospital Course|10592,10602|false|false|false|||discharged
Drug|Organic Chemical|Hospital Course|10606,10616|false|false|false|C0002598|amiodarone|Amiodarone
Drug|Pharmacologic Substance|Hospital Course|10606,10616|false|false|false|C0002598|amiodarone|Amiodarone
Event|Event|Hospital Course|10606,10616|false|false|false|||Amiodarone
Procedure|Laboratory Procedure|Hospital Course|10606,10616|false|false|false|C5399868|Drug assay amiodarone|Amiodarone
Finding|Intellectual Product|Hospital Course|10648,10652|false|false|false|C1561540|Transaction counts and value totals - week|week
Finding|Intellectual Product|Hospital Course|10667,10671|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Activity|Hospital Course|10712,10723|false|false|false|C0003629|Appointments|appointment
Event|Event|Hospital Course|10712,10723|false|false|false|||appointment
Event|Event|Hospital Course|10774,10784|false|false|false|||discharged
Drug|Organic Chemical|Hospital Course|10788,10799|false|false|false|C1739768|rivaroxaban|Rivaroxaban
Drug|Pharmacologic Substance|Hospital Course|10788,10799|false|false|false|C1739768|rivaroxaban|Rivaroxaban
Event|Event|Hospital Course|10788,10799|false|false|false|||Rivaroxaban
Event|Event|Hospital Course|10815,10821|false|false|false|||dinner
Finding|Daily or Recreational Activity|Hospital Course|10815,10821|false|false|false|C4048877|Dinner|dinner
Event|Event|Hospital Course|10828,10838|false|false|false|||discharged
Event|Event|Hospital Course|10844,10854|false|false|false|||outpatient
Finding|Classification|Hospital Course|10844,10854|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|10844,10854|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10862,10868|false|false|false|C0018787|Heart|Hearts
Drug|Hazardous or Poisonous Substance|Hospital Course|10869,10876|false|false|false|C0728873|Monitor brand of insecticide|monitor
Drug|Organic Chemical|Hospital Course|10869,10876|false|false|false|C0728873|Monitor brand of insecticide|monitor
Event|Event|Hospital Course|10883,10890|false|false|false|||results
Event|Event|Hospital Course|10897,10908|false|false|false|||interpreted
Event|Event|Hospital Course|10933,10942|false|false|false|||presented
Anatomy|Body Location or Region|Hospital Course|10948,10953|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Hospital Course|10948,10953|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Hospital Course|10948,10958|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|Hospital Course|10948,10958|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Hospital Course|10954,10958|false|false|false|C2598155||pain
Event|Event|Hospital Course|10954,10958|false|false|false|||pain
Finding|Functional Concept|Hospital Course|10954,10958|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|10954,10958|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|Hospital Course|10986,10996|true|false|false|C0005516|Biological Markers|biomarkers
Event|Event|Hospital Course|10986,10996|true|false|false|||biomarkers
Event|Event|Hospital Course|11000,11003|true|false|false|||EKG
Finding|Intellectual Product|Hospital Course|11000,11003|true|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|Hospital Course|11000,11003|true|false|false|C1623258|Electrocardiography|EKG
Event|Event|Hospital Course|11004,11011|true|false|false|||changes
Finding|Functional Concept|Hospital Course|11004,11011|true|false|false|C0392747|Changing|changes
Anatomy|Tissue|Hospital Course|11027,11037|false|false|false|C0027061|Myocardium|myocardial
Disorder|Injury or Poisoning|Hospital Course|11038,11044|false|false|false|C0010957|Tissue damage|damage
Event|Event|Hospital Course|11038,11044|false|false|false|||damage
Finding|Functional Concept|Hospital Course|11038,11044|false|false|false|C1883709;C2681922|Damage;MAGEE1 gene|damage
Finding|Gene or Genome|Hospital Course|11038,11044|false|false|false|C1883709;C2681922|Damage;MAGEE1 gene|damage
Event|Event|Hospital Course|11060,11068|false|false|false|||remained
Event|Event|Hospital Course|11069,11081|false|false|false|||asymptomatic
Finding|Finding|Hospital Course|11069,11081|false|false|false|C0231221;C0332151|Asymptomatic (finding);Asymptomatic diagnosis of|asymptomatic
Event|Event|Hospital Course|11089,11096|false|false|false|||periods
Finding|Organism Function|Hospital Course|11089,11096|false|false|false|C0025344|Menstruation|periods
Disorder|Disease or Syndrome|Hospital Course|11101,11129|false|false|false|C0039240|Supraventricular tachycardia|supraventricular tachycardia
Finding|Finding|Hospital Course|11101,11129|false|false|false|C3815188|Supraventricular Tachycardia by ECG Finding|supraventricular tachycardia
Event|Event|Hospital Course|11118,11129|false|false|false|||tachycardia
Finding|Finding|Hospital Course|11118,11129|false|false|false|C0039231;C3827868|Tachycardia;Tachycardia by ECG Finding|tachycardia
Event|Event|Hospital Course|11144,11156|false|false|false|||hospitalized
Finding|Body Substance|Hospital Course|11158,11165|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|11158,11165|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|11158,11165|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Hospital Course|11171,11178|false|false|false|||benefit
Finding|Classification|Hospital Course|11184,11194|false|true|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|11184,11194|false|true|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Attribute|Clinical Attribute|Hospital Course|11195,11201|false|false|false|C1718621|W stress|stress
Drug|Organic Chemical|Hospital Course|11195,11201|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|Hospital Course|11195,11201|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Finding|Finding|Hospital Course|11195,11201|false|false|false|C0038435|Stress|stress
Procedure|Diagnostic Procedure|Hospital Course|11195,11206|false|false|false|C0015260;C3494508|Exercise stress test;Stress Test|stress test
Anatomy|Body Location or Region|Hospital Course|11202,11206|false|false|false|C4318744|Test - temporal region|test
Event|Event|Hospital Course|11202,11206|false|false|false|||test
Finding|Functional Concept|Hospital Course|11202,11206|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Finding|Intellectual Product|Hospital Course|11202,11206|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Lab|Laboratory or Test Result|Hospital Course|11202,11206|false|false|false|C0456984|Test Result|test
Procedure|Laboratory Procedure|Hospital Course|11202,11206|false|false|false|C0022885|Laboratory Procedures|test
Event|Event|Hospital Course|11215,11223|false|false|false|||symptoms
Finding|Functional Concept|Hospital Course|11215,11223|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Hospital Course|11215,11223|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|Hospital Course|11224,11230|false|false|false|||return
Finding|Idea or Concept|Hospital Course|11238,11241|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|11238,11241|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Hospital Course|11245,11254|false|false|false|||discharge
Finding|Body Substance|Hospital Course|11245,11254|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|11245,11254|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|11245,11254|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|11245,11254|false|false|false|C0030685|Patient Discharge|discharge
Finding|Idea or Concept|Hospital Course|11263,11274|false|false|false|C0750502|Significant|significant
Attribute|Clinical Attribute|Hospital Course|11275,11280|false|false|false|C5886197||R eye
Anatomy|Body Location or Region|Hospital Course|11277,11280|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|eye
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11277,11280|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|eye
Disorder|Disease or Syndrome|Hospital Course|11277,11280|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|eye
Disorder|Neoplastic Process|Hospital Course|11277,11280|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|eye
Finding|Body Substance|Hospital Course|11277,11280|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Finding|Hospital Course|11277,11280|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Intellectual Product|Hospital Course|11277,11280|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Sign or Symptom|Hospital Course|11277,11285|false|false|false|C0151827|Eye pain|eye pain
Attribute|Clinical Attribute|Hospital Course|11281,11285|false|false|false|C2598155||pain
Event|Event|Hospital Course|11281,11285|false|false|false|||pain
Finding|Functional Concept|Hospital Course|11281,11285|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|11281,11285|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Disorder|Disease or Syndrome|Hospital Course|11291,11298|false|false|false|C0041834|Erythema|redness
Event|Event|Hospital Course|11291,11298|false|false|false|||redness
Finding|Finding|Hospital Course|11291,11298|false|false|false|C0332575|Redness|redness
Event|Event|Hospital Course|11304,11313|false|false|false|||evaluated
Event|Event|Hospital Course|11335,11339|false|false|false|||felt
Disorder|Disease or Syndrome|Hospital Course|11358,11366|false|false|false|C0013238;C0022575|Dry Eye Syndromes;Keratoconjunctivitis Sicca|dry eyes
Drug|Pharmacologic Substance|Hospital Course|11358,11366|false|false|false|C0720056|Dry Eyes brand of ocular lubricant|dry eyes
Finding|Sign or Symptom|Hospital Course|11358,11366|false|false|false|C0314719|Dryness of eye|dry eyes
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11362,11366|false|false|false|C0015392|Eye|eyes
Attribute|Clinical Attribute|Hospital Course|11362,11366|false|false|false|C5848506||eyes
Event|Event|Hospital Course|11362,11366|false|false|false|||eyes
Event|Event|Hospital Course|11368,11375|false|false|false|||treated
Drug|Antibiotic|Hospital Course|11381,11393|false|false|false|C0014806|erythromycin|erythromycin
Drug|Organic Chemical|Hospital Course|11381,11393|false|false|false|C0014806|erythromycin|erythromycin
Drug|Biomedical or Dental Material|Hospital Course|11394,11399|false|false|false|C0991568|Drops - Drug Form|drops
Event|Event|Hospital Course|11394,11399|false|false|false|||drops
Event|Event|Hospital Course|11404,11414|false|false|false|||artifiical
Event|Event|Hospital Course|11416,11421|false|false|false|||tears
Finding|Body Substance|Hospital Course|11416,11421|false|false|false|C0039409;C1547924;C1611838|Tears (substance);Tears specimen|tears
Finding|Intellectual Product|Hospital Course|11416,11421|false|false|false|C0039409;C1547924;C1611838|Tears (substance);Tears specimen|tears
Finding|Body Substance|Hospital Course|11423,11430|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|11423,11430|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|11423,11430|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Biologically Active Substance|Hospital Course|11443,11447|false|false|false|C0245203|4-azido-7-phenylpyrazolo-(1,5a)-1,3,5-triazine|appt
Drug|Organic Chemical|Hospital Course|11443,11447|false|false|false|C0245203|4-azido-7-phenylpyrazolo-(1,5a)-1,3,5-triazine|appt
Event|Event|Hospital Course|11443,11447|false|false|false|||appt
Event|Event|Hospital Course|11489,11493|false|false|false|||need
Event|Event|Hospital Course|11497,11503|false|false|false|||attend
Event|Event|Hospital Course|11511,11515|false|false|false|||Code
Event|Occupational Activity|Hospital Course|11511,11515|false|false|false|C0009219|Coding|Code
Finding|Intellectual Product|Hospital Course|11511,11515|false|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|Code
Event|Activity|Hospital Course|11516,11523|false|false|false|C3812666|Personal Contact|Contact
Event|Event|Hospital Course|11516,11523|false|false|false|||Contact
Finding|Functional Concept|Hospital Course|11516,11523|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|Contact
Finding|Idea or Concept|Hospital Course|11516,11523|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|Contact
Finding|Intellectual Product|Hospital Course|11516,11523|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|Contact
Phenomenon|Phenomenon or Process|Hospital Course|11516,11523|false|false|false|C0392367|Physical contact|Contact
Event|Activity|Hospital Course|11525,11532|false|false|false|C3812666|Personal Contact|CONTACT
Event|Event|Hospital Course|11525,11532|false|false|false|||CONTACT
Finding|Functional Concept|Hospital Course|11525,11532|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Finding|Idea or Concept|Hospital Course|11525,11532|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Finding|Intellectual Product|Hospital Course|11525,11532|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Phenomenon|Phenomenon or Process|Hospital Course|11525,11532|false|false|false|C0392367|Physical contact|CONTACT
Attribute|Clinical Attribute|Hospital Course|11576,11587|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|11576,11587|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|11576,11587|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|11576,11587|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|11576,11600|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|Hospital Course|11591,11600|false|false|false|||Admission
Procedure|Health Care Activity|Hospital Course|11591,11600|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|Hospital Course|11619,11629|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|Hospital Course|11619,11629|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|Hospital Course|11619,11634|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|Hospital Course|11630,11634|false|false|false|||list
Finding|Intellectual Product|Hospital Course|11630,11634|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|Hospital Course|11638,11646|false|false|false|||accurate
Drug|Organic Chemical|Hospital Course|11651,11659|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|Hospital Course|11651,11659|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|Hospital Course|11651,11659|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|Hospital Course|11651,11659|false|false|false|||complete
Finding|Functional Concept|Hospital Course|11651,11659|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|Hospital Course|11651,11659|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Organic Chemical|Hospital Course|11664,11677|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Hospital Course|11664,11677|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|Hospital Course|11664,11677|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|Hospital Course|11664,11677|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|Hospital Course|11692,11695|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|11696,11700|false|false|false|C2598155||pain
Event|Event|Hospital Course|11696,11700|false|false|false|||pain
Finding|Functional Concept|Hospital Course|11696,11700|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|11696,11700|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|Hospital Course|11705,11714|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|Hospital Course|11705,11714|false|false|false|C0001927|albuterol|Albuterol
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11722,11725|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biologically Active Substance|Hospital Course|11722,11725|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biomedical or Dental Material|Hospital Course|11722,11725|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Finding|Cell Function|Hospital Course|11722,11725|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Finding|Gene or Genome|Hospital Course|11722,11725|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11733,11736|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biologically Active Substance|Hospital Course|11733,11736|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biomedical or Dental Material|Hospital Course|11733,11736|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Event|Event|Hospital Course|11733,11736|false|false|false|||NEB
Finding|Cell Function|Hospital Course|11733,11736|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|Hospital Course|11733,11736|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|Hospital Course|11744,11747|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|Hospital Course|11748,11757|false|false|false|||shortness
Finding|Body Substance|Hospital Course|11762,11768|false|false|false|C0225386|Breath|breath
Drug|Organic Chemical|Hospital Course|11773,11780|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|Hospital Course|11773,11780|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|Hospital Course|11800,11812|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|Hospital Course|11800,11812|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|Hospital Course|11830,11841|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Pharmacologic Substance|Hospital Course|11830,11841|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Organic Chemical|Hospital Course|11861,11870|false|false|false|C0012373|diltiazem|Diltiazem
Drug|Pharmacologic Substance|Hospital Course|11861,11870|false|false|false|C0012373|diltiazem|Diltiazem
Finding|Finding|Hospital Course|11871,11879|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|11871,11879|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|Hospital Course|11880,11887|false|false|false|||Release
Finding|Functional Concept|Hospital Course|11880,11887|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|11880,11887|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|11880,11887|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|Hospital Course|11908,11919|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Hospital Course|11908,11919|false|false|false|C0082607|fluticasone|Fluticasone
Event|Event|Hospital Course|11908,11919|false|false|false|||Fluticasone
Drug|Organic Chemical|Hospital Course|11908,11930|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Pharmacologic Substance|Hospital Course|11908,11930|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Organic Chemical|Hospital Course|11920,11930|false|false|false|C0033474;C0392214|Propionates;propionate|Propionate
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11931,11936|false|false|false|C0028429||NASAL
Drug|Biomedical or Dental Material|Hospital Course|11931,11936|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Drug|Organic Chemical|Hospital Course|11931,11936|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Drug|Pharmacologic Substance|Hospital Course|11931,11936|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Finding|Finding|Hospital Course|11931,11936|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|NASAL
Finding|Functional Concept|Hospital Course|11931,11936|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|NASAL
Event|Event|Hospital Course|11939,11943|false|false|false|||SPRY
Finding|Gene or Genome|Hospital Course|11953,11956|false|false|false|C1422467|CIAO3 gene|PRN
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11957,11962|false|false|false|C0028429||nasal
Drug|Biomedical or Dental Material|Hospital Course|11957,11962|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Organic Chemical|Hospital Course|11957,11962|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Pharmacologic Substance|Hospital Course|11957,11962|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Event|Event|Hospital Course|11957,11962|false|false|false|||nasal
Finding|Finding|Hospital Course|11957,11962|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Functional Concept|Hospital Course|11957,11962|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Event|Event|Hospital Course|11964,11974|false|false|false|||congestion
Finding|Pathologic Function|Hospital Course|11964,11974|false|false|false|C0700148|Congestion|congestion
Drug|Organic Chemical|Hospital Course|11979,11990|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Hospital Course|11979,11990|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Hospital Course|11979,12001|false|false|false|C0939232|fluticasone / salmeterol|Fluticasone-Salmeterol
Drug|Organic Chemical|Hospital Course|11979,12008|false|false|false|C4762496|Fluticasone-Salmeterol Diskus|Fluticasone-Salmeterol Diskus
Drug|Pharmacologic Substance|Hospital Course|11979,12008|false|false|false|C4762496|Fluticasone-Salmeterol Diskus|Fluticasone-Salmeterol Diskus
Drug|Organic Chemical|Hospital Course|11991,12001|false|false|false|C0073992|salmeterol|Salmeterol
Drug|Pharmacologic Substance|Hospital Course|11991,12001|false|false|false|C0073992|salmeterol|Salmeterol
Event|Event|Hospital Course|12002,12008|false|false|false|||Diskus
Drug|Biomedical or Dental Material|Hospital Course|12021,12024|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Organic Chemical|Hospital Course|12021,12024|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Pharmacologic Substance|Hospital Course|12021,12024|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Event|Event|Hospital Course|12021,12024|false|false|false|||INH
Finding|Functional Concept|Hospital Course|12021,12024|false|false|false|C0205535|Inhalation Route of Administration|INH
Disorder|Mental or Behavioral Dysfunction|Hospital Course|12028,12031|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12028,12031|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|12028,12031|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|12028,12031|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|12028,12031|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|12036,12055|false|false|false|C0020261|hydrochlorothiazide|Hydrochlorothiazide
Drug|Pharmacologic Substance|Hospital Course|12036,12055|false|false|false|C0020261|hydrochlorothiazide|Hydrochlorothiazide
Drug|Organic Chemical|Hospital Course|12076,12086|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Pharmacologic Substance|Hospital Course|12076,12086|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Organic Chemical|Hospital Course|12076,12098|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Drug|Pharmacologic Substance|Hospital Course|12076,12098|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Event|Event|Hospital Course|12087,12098|false|false|false|||Mononitrate
Finding|Finding|Hospital Course|12100,12108|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|12100,12108|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|Hospital Course|12109,12116|false|false|false|||Release
Finding|Functional Concept|Hospital Course|12109,12116|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|12109,12116|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|12109,12116|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|Hospital Course|12139,12150|false|false|false|C0090306|latanoprost|Latanoprost
Drug|Pharmacologic Substance|Hospital Course|12139,12150|false|false|false|C0090306|latanoprost|Latanoprost
Finding|Functional Concept|Hospital Course|12158,12163|false|false|false|C1522230|Ophthalmic Route of Administration|Ophth
Drug|Biomedical or Dental Material|Hospital Course|12173,12177|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|Hospital Course|12173,12177|false|false|false|C1705648|Dropping|DROP
Event|Event|Hospital Course|12178,12182|false|false|false|||LEFT
Finding|Functional Concept|Hospital Course|12178,12182|false|false|false|C1552822|Table Cell Horizontal Align - left|LEFT
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|12178,12186|false|false|false|C0229090|Left eye structure|LEFT EYE
Procedure|Diagnostic Procedure|Hospital Course|12178,12186|false|false|false|C2141124|examination of left eye|LEFT EYE
Anatomy|Body Location or Region|Hospital Course|12183,12186|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|EYE
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|12183,12186|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|EYE
Disorder|Disease or Syndrome|Hospital Course|12183,12186|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|EYE
Disorder|Neoplastic Process|Hospital Course|12183,12186|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|EYE
Event|Event|Hospital Course|12183,12186|false|false|false|||EYE
Finding|Body Substance|Hospital Course|12183,12186|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|EYE
Finding|Finding|Hospital Course|12183,12186|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|EYE
Finding|Intellectual Product|Hospital Course|12183,12186|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|EYE
Drug|Organic Chemical|Hospital Course|12195,12204|false|false|false|C0024002|lorazepam|Lorazepam
Drug|Pharmacologic Substance|Hospital Course|12195,12204|false|false|false|C0024002|lorazepam|Lorazepam
Event|Event|Hospital Course|12215,12218|false|false|false|||QHS
Finding|Gene or Genome|Hospital Course|12219,12222|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Pharmacologic Substance|Hospital Course|12223,12231|false|false|false|C1950154|Insomnia homeopathic medication|insomnia
Event|Event|Hospital Course|12223,12231|false|false|false|||insomnia
Finding|Sign or Symptom|Hospital Course|12223,12231|false|false|false|C0917801|Sleeplessness|insomnia
Drug|Organic Chemical|Hospital Course|12237,12250|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|Hospital Course|12237,12250|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|Hospital Course|12237,12250|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Event|Event|Hospital Course|12237,12250|false|false|false|||Multivitamins
Drug|Inorganic Chemical|Hospital Course|12253,12261|false|false|false|C0026162|Minerals|minerals
Event|Event|Hospital Course|12253,12261|false|false|false|||minerals
Drug|Biomedical or Dental Material|Hospital Course|12264,12267|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|Hospital Course|12264,12267|false|false|false|||TAB
Drug|Organic Chemical|Hospital Course|12282,12292|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Pharmacologic Substance|Hospital Course|12282,12292|false|false|false|C0034665|ranitidine|Ranitidine
Disorder|Mental or Behavioral Dysfunction|Hospital Course|12303,12306|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12303,12306|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|12303,12306|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|12303,12306|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|12303,12306|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|12312,12320|false|false|false|C0040610|tramadol|TraMADOL
Drug|Pharmacologic Substance|Hospital Course|12312,12320|false|false|false|C0040610|tramadol|TraMADOL
Event|Event|Hospital Course|12312,12320|false|false|false|||TraMADOL
Procedure|Laboratory Procedure|Hospital Course|12312,12320|false|false|false|C1266765|Tramadol measurement (procedure)|TraMADOL
Drug|Organic Chemical|Hospital Course|12322,12328|false|false|false|C0724054|Ultram|Ultram
Drug|Pharmacologic Substance|Hospital Course|12322,12328|false|false|false|C0724054|Ultram|Ultram
Finding|Gene or Genome|Hospital Course|12343,12346|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|12347,12351|false|false|false|C2598155||pain
Event|Event|Hospital Course|12347,12351|false|false|false|||pain
Finding|Functional Concept|Hospital Course|12347,12351|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|12347,12351|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|Hospital Course|12357,12369|false|false|false|C0039771|theophylline|Theophylline
Drug|Pharmacologic Substance|Hospital Course|12357,12369|false|false|false|C0039771|theophylline|Theophylline
Event|Event|Hospital Course|12357,12369|false|false|false|||Theophylline
Procedure|Laboratory Procedure|Hospital Course|12357,12369|false|false|false|C0039773|Assay of theophylline|Theophylline
Drug|Organic Chemical|Hospital Course|12357,12372|false|false|false|C2241157|Theophylline ER|Theophylline ER
Drug|Pharmacologic Substance|Hospital Course|12357,12372|false|false|false|C2241157|Theophylline ER|Theophylline ER
Disorder|Mental or Behavioral Dysfunction|Hospital Course|12383,12386|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12383,12386|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|12383,12386|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|12383,12386|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|12383,12386|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|12392,12402|false|false|false|C0213771|tiotropium|Tiotropium
Drug|Pharmacologic Substance|Hospital Course|12392,12402|false|false|false|C0213771|tiotropium|Tiotropium
Event|Event|Hospital Course|12392,12402|false|false|false|||Tiotropium
Drug|Organic Chemical|Hospital Course|12392,12410|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Pharmacologic Substance|Hospital Course|12392,12410|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Inorganic Chemical|Hospital Course|12403,12410|false|false|false|C0006222|Bromides|Bromide
Event|Event|Hospital Course|12403,12410|false|false|false|||Bromide
Procedure|Laboratory Procedure|Hospital Course|12403,12410|false|false|false|C0202341|Bromides measurement|Bromide
Disorder|Congenital Abnormality|Hospital Course|12413,12416|false|false|false|C1855179|CATARACT, ANTERIOR POLAR|CAP
Drug|Biomedical or Dental Material|Hospital Course|12413,12416|false|false|false|C0006935|capsule (pharmacologic)|CAP
Event|Event|Hospital Course|12413,12416|false|false|false|||CAP
Finding|Gene or Genome|Hospital Course|12413,12416|false|false|false|C1416891;C1418551;C1419093;C1422073;C1422760;C2985259;C4522312|BRD4 gene;BRD4 wt Allele;CAP1 gene;HACD1 gene;LNPEP gene;SERPINB6 gene;SORBS1 gene|CAP
Procedure|Therapeutic or Preventive Procedure|Hospital Course|12413,12416|false|false|false|C0278651;C0280547;C1879916|CAP Regimen;cisplatin/cyclophosphamide/doxorubicin protocol;cyclophosphamide/doxorubicin/prednisone protocol|CAP
Drug|Organic Chemical|Hospital Course|12431,12442|false|false|false|C0018305|guaifenesin|Guaifenesin
Drug|Pharmacologic Substance|Hospital Course|12431,12442|false|false|false|C0018305|guaifenesin|Guaifenesin
Event|Event|Hospital Course|12431,12442|false|false|false|||Guaifenesin
Drug|Organic Chemical|Hospital Course|12443,12450|false|false|false|C0009214|codeine|CODEINE
Drug|Pharmacologic Substance|Hospital Course|12443,12450|false|false|false|C0009214|codeine|CODEINE
Event|Event|Hospital Course|12443,12450|false|false|false|||CODEINE
Drug|Organic Chemical|Hospital Course|12443,12460|false|false|false|C0009217|codeine phosphate|CODEINE Phosphate
Drug|Pharmacologic Substance|Hospital Course|12443,12460|false|false|false|C0009217|codeine phosphate|CODEINE Phosphate
Drug|Element, Ion, or Isotope|Hospital Course|12451,12460|false|false|false|C0031603;C1601799|Phosphates;phosphate ion|Phosphate
Drug|Inorganic Chemical|Hospital Course|12451,12460|false|false|false|C0031603;C1601799|Phosphates;phosphate ion|Phosphate
Drug|Pharmacologic Substance|Hospital Course|12451,12460|false|false|false|C0031603;C1601799|Phosphates;phosphate ion|Phosphate
Event|Event|Hospital Course|12451,12460|false|false|false|||Phosphate
Procedure|Laboratory Procedure|Hospital Course|12451,12460|false|false|false|C0523826|Phosphate measurement|Phosphate
Finding|Gene or Genome|Hospital Course|12473,12476|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Organic Chemical|Hospital Course|12477,12482|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|Hospital Course|12477,12482|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|Hospital Course|12477,12482|false|false|false|||cough
Finding|Sign or Symptom|Hospital Course|12477,12482|false|false|false|C0010200|Coughing|cough
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12488,12491|false|false|false|C0056632;C0459207;C2702357;C3488428|Cyclophosphamide/Dacarbazine/Vincristine;cod, unspecified preparation;codfish allergenic extract|cod
Drug|Food|Hospital Course|12488,12491|false|false|false|C0056632;C0459207;C2702357;C3488428|Cyclophosphamide/Dacarbazine/Vincristine;cod, unspecified preparation;codfish allergenic extract|cod
Drug|Immunologic Factor|Hospital Course|12488,12491|false|false|false|C0056632;C0459207;C2702357;C3488428|Cyclophosphamide/Dacarbazine/Vincristine;cod, unspecified preparation;codfish allergenic extract|cod
Drug|Pharmacologic Substance|Hospital Course|12488,12491|false|false|false|C0056632;C0459207;C2702357;C3488428|Cyclophosphamide/Dacarbazine/Vincristine;cod, unspecified preparation;codfish allergenic extract|cod
Finding|Finding|Hospital Course|12488,12491|false|false|false|C0007465;C0457523;C1420285;C5444130|Cancerization of Pancreatic Ducts;Cause of Death;Cemento-osseous dysplasia;SNRPB gene|cod
Finding|Gene or Genome|Hospital Course|12488,12491|false|false|false|C0007465;C0457523;C1420285;C5444130|Cancerization of Pancreatic Ducts;Cause of Death;Cemento-osseous dysplasia;SNRPB gene|cod
Finding|Pathologic Function|Hospital Course|12488,12491|false|false|false|C0007465;C0457523;C1420285;C5444130|Cancerization of Pancreatic Ducts;Cause of Death;Cemento-osseous dysplasia;SNRPB gene|cod
Drug|Food|Hospital Course|12488,12501|false|false|false|C0009213|cod liver oil|cod liver oil
Drug|Organic Chemical|Hospital Course|12488,12501|false|false|false|C0009213|cod liver oil|cod liver oil
Drug|Pharmacologic Substance|Hospital Course|12488,12501|false|false|false|C0009213|cod liver oil|cod liver oil
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|12492,12497|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|Hospital Course|12492,12497|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|Hospital Course|12492,12497|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|Hospital Course|12492,12497|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|Hospital Course|12492,12497|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|Hospital Course|12492,12497|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|Hospital Course|12492,12497|false|false|false|||liver
Finding|Finding|Hospital Course|12492,12497|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|Hospital Course|12492,12497|false|false|false|C0872387|Procedures on liver|liver
Drug|Biomedical or Dental Material|Hospital Course|12498,12501|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|oil
Drug|Food|Hospital Course|12498,12501|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|oil
Drug|Organic Chemical|Hospital Course|12498,12501|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|oil
Drug|Pharmacologic Substance|Hospital Course|12498,12501|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|oil
Anatomy|Body Space or Junction|Hospital Course|12517,12521|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|12517,12521|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|12517,12521|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|12517,12521|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Disorder|Mental or Behavioral Dysfunction|Hospital Course|12522,12525|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12522,12525|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|12522,12525|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|12522,12525|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|12522,12525|false|false|false|C1332410|BID gene|BID
Drug|Inorganic Chemical|Hospital Course|12531,12538|false|false|false|C0719084|CalCarb|Calcarb
Event|Event|Hospital Course|12531,12538|false|false|false|||Calcarb
Drug|Organic Chemical|Hospital Course|12548,12555|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|Hospital Course|12548,12555|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|Hospital Course|12548,12555|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|Hospital Course|12548,12557|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|Hospital Course|12548,12557|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|Hospital Course|12548,12557|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|Hospital Course|12548,12557|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|Hospital Course|12548,12557|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Drug|Biologically Active Substance|Hospital Course|12559,12566|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Element, Ion, or Isotope|Hospital Course|12559,12566|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Inorganic Chemical|Hospital Course|12559,12566|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Pharmacologic Substance|Hospital Course|12559,12566|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Vitamin|Hospital Course|12559,12566|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Event|Event|Hospital Course|12559,12566|false|false|false|||calcium
Finding|Physiologic Function|Hospital Course|12559,12566|false|false|false|C4553026|Calcium metabolic function|calcium
Procedure|Laboratory Procedure|Hospital Course|12559,12566|false|false|false|C0201925|Calcium measurement|calcium
Drug|Inorganic Chemical|Hospital Course|12559,12576|false|false|false|C0006681|calcium carbonate|calcium carbonate
Drug|Pharmacologic Substance|Hospital Course|12559,12576|false|false|false|C0006681|calcium carbonate|calcium carbonate
Drug|Element, Ion, or Isotope|Hospital Course|12567,12576|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|carbonate
Drug|Organic Chemical|Hospital Course|12567,12576|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|carbonate
Drug|Pharmacologic Substance|Hospital Course|12567,12576|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|carbonate
Event|Event|Hospital Course|12567,12576|false|false|false|||carbonate
Drug|Organic Chemical|Hospital Course|12577,12584|false|false|false|C0042890|Vitamins|vitamin
Drug|Pharmacologic Substance|Hospital Course|12577,12584|false|false|false|C0042890|Vitamins|vitamin
Drug|Vitamin|Hospital Course|12577,12584|false|false|false|C0042890|Vitamins|vitamin
Event|Event|Hospital Course|12577,12584|false|false|false|||vitamin
Drug|Organic Chemical|Hospital Course|12577,12587|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Drug|Pharmacologic Substance|Hospital Course|12577,12587|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Drug|Vitamin|Hospital Course|12577,12587|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Anatomy|Body Space or Junction|Hospital Course|12601,12605|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|12601,12605|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|12601,12605|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|12601,12605|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Event|Event|Hospital Course|12616,12625|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|12616,12625|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|12616,12625|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|12616,12625|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|12616,12625|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|12616,12637|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|12626,12637|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|12626,12637|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|12626,12637|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|12626,12637|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Hospital Course|12642,12652|false|false|false|C0002598|amiodarone|Amiodarone
Drug|Pharmacologic Substance|Hospital Course|12642,12652|false|false|false|C0002598|amiodarone|Amiodarone
Event|Event|Hospital Course|12642,12652|false|false|false|||Amiodarone
Procedure|Laboratory Procedure|Hospital Course|12642,12652|false|false|false|C5399868|Drug assay amiodarone|Amiodarone
Disorder|Mental or Behavioral Dysfunction|Hospital Course|12663,12666|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12663,12666|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|12663,12666|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|12663,12666|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|12663,12666|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|12672,12682|false|false|false|C0002598|amiodarone|amiodarone
Drug|Pharmacologic Substance|Hospital Course|12672,12682|false|false|false|C0002598|amiodarone|amiodarone
Event|Event|Hospital Course|12672,12682|false|false|false|||amiodarone
Procedure|Laboratory Procedure|Hospital Course|12672,12682|false|false|false|C5399868|Drug assay amiodarone|amiodarone
Drug|Biomedical or Dental Material|Hospital Course|12692,12698|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|Hospital Course|12702,12710|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|12705,12710|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|12705,12710|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Idea or Concept|Hospital Course|12719,12722|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|12719,12722|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Biomedical or Dental Material|Hospital Course|12734,12740|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|12741,12748|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|12741,12748|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|12755,12766|false|false|false|C1739768|rivaroxaban|Rivaroxaban
Drug|Pharmacologic Substance|Hospital Course|12755,12766|false|false|false|C1739768|rivaroxaban|Rivaroxaban
Event|Event|Hospital Course|12776,12782|false|false|false|||DINNER
Finding|Daily or Recreational Activity|Hospital Course|12776,12782|false|false|false|C4048877|Dinner|DINNER
Event|Event|Hospital Course|12784,12786|false|false|false|||RX
Drug|Organic Chemical|Hospital Course|12788,12799|false|false|false|C1739768|rivaroxaban|rivaroxaban
Drug|Pharmacologic Substance|Hospital Course|12788,12799|false|false|false|C1739768|rivaroxaban|rivaroxaban
Event|Event|Hospital Course|12788,12799|false|false|false|||rivaroxaban
Drug|Organic Chemical|Hospital Course|12801,12808|false|false|false|C3159309|Xarelto|Xarelto
Drug|Pharmacologic Substance|Hospital Course|12801,12808|false|false|false|C3159309|Xarelto|Xarelto
Drug|Biomedical or Dental Material|Hospital Course|12818,12824|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|Hospital Course|12828,12836|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|12831,12836|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|12831,12836|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Event|Activity|Hospital Course|12841,12845|false|false|false|C1880359|Dispense (activity)|Disp
Finding|Gene or Genome|Hospital Course|12841,12845|false|false|false|C2828567|PRSS30P gene|Disp
Drug|Biomedical or Dental Material|Hospital Course|12852,12858|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|12859,12866|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|12859,12866|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|12873,12886|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Hospital Course|12873,12886|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|Hospital Course|12873,12886|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|Hospital Course|12873,12886|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|Hospital Course|12901,12904|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|12905,12909|false|false|false|C2598155||pain
Event|Event|Hospital Course|12905,12909|false|false|false|||pain
Finding|Functional Concept|Hospital Course|12905,12909|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|12905,12909|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|Hospital Course|12914,12923|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|Hospital Course|12914,12923|false|false|false|C0001927|albuterol|Albuterol
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12931,12934|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biologically Active Substance|Hospital Course|12931,12934|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biomedical or Dental Material|Hospital Course|12931,12934|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Finding|Cell Function|Hospital Course|12931,12934|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Finding|Gene or Genome|Hospital Course|12931,12934|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12942,12945|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biologically Active Substance|Hospital Course|12942,12945|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biomedical or Dental Material|Hospital Course|12942,12945|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Event|Event|Hospital Course|12942,12945|false|false|false|||NEB
Finding|Cell Function|Hospital Course|12942,12945|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|Hospital Course|12942,12945|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|Hospital Course|12953,12956|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|Hospital Course|12957,12966|false|false|false|||shortness
Finding|Body Substance|Hospital Course|12971,12977|false|false|false|C0225386|Breath|breath
Drug|Organic Chemical|Hospital Course|12982,12989|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|Hospital Course|12982,12989|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|Hospital Course|13009,13021|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|Hospital Course|13009,13021|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|Hospital Course|13039,13048|false|false|false|C0012373|diltiazem|Diltiazem
Drug|Pharmacologic Substance|Hospital Course|13039,13048|false|false|false|C0012373|diltiazem|Diltiazem
Finding|Finding|Hospital Course|13049,13057|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|13049,13057|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|Hospital Course|13058,13065|false|false|false|||Release
Finding|Functional Concept|Hospital Course|13058,13065|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|13058,13065|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|13058,13065|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|Hospital Course|13086,13097|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Hospital Course|13086,13097|false|false|false|C0082607|fluticasone|Fluticasone
Event|Event|Hospital Course|13086,13097|false|false|false|||Fluticasone
Drug|Organic Chemical|Hospital Course|13086,13108|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Pharmacologic Substance|Hospital Course|13086,13108|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Organic Chemical|Hospital Course|13098,13108|false|false|false|C0033474;C0392214|Propionates;propionate|Propionate
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|13109,13114|false|false|false|C0028429||NASAL
Drug|Biomedical or Dental Material|Hospital Course|13109,13114|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Drug|Organic Chemical|Hospital Course|13109,13114|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Drug|Pharmacologic Substance|Hospital Course|13109,13114|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Finding|Finding|Hospital Course|13109,13114|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|NASAL
Finding|Functional Concept|Hospital Course|13109,13114|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|NASAL
Event|Event|Hospital Course|13117,13121|false|false|false|||SPRY
Finding|Gene or Genome|Hospital Course|13131,13134|false|false|false|C1422467|CIAO3 gene|PRN
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|13135,13140|false|false|false|C0028429||nasal
Drug|Biomedical or Dental Material|Hospital Course|13135,13140|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Organic Chemical|Hospital Course|13135,13140|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Pharmacologic Substance|Hospital Course|13135,13140|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Event|Event|Hospital Course|13135,13140|false|false|false|||nasal
Finding|Finding|Hospital Course|13135,13140|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Functional Concept|Hospital Course|13135,13140|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Event|Event|Hospital Course|13142,13152|false|false|false|||congestion
Finding|Pathologic Function|Hospital Course|13142,13152|false|false|false|C0700148|Congestion|congestion
Drug|Organic Chemical|Hospital Course|13157,13168|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Hospital Course|13157,13168|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Hospital Course|13157,13179|false|false|false|C0939232|fluticasone / salmeterol|Fluticasone-Salmeterol
Drug|Organic Chemical|Hospital Course|13157,13186|false|false|false|C4762496|Fluticasone-Salmeterol Diskus|Fluticasone-Salmeterol Diskus
Drug|Pharmacologic Substance|Hospital Course|13157,13186|false|false|false|C4762496|Fluticasone-Salmeterol Diskus|Fluticasone-Salmeterol Diskus
Drug|Organic Chemical|Hospital Course|13169,13179|false|false|false|C0073992|salmeterol|Salmeterol
Drug|Pharmacologic Substance|Hospital Course|13169,13179|false|false|false|C0073992|salmeterol|Salmeterol
Event|Event|Hospital Course|13180,13186|false|false|false|||Diskus
Drug|Biomedical or Dental Material|Hospital Course|13199,13202|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Organic Chemical|Hospital Course|13199,13202|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Pharmacologic Substance|Hospital Course|13199,13202|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Event|Event|Hospital Course|13199,13202|false|false|false|||INH
Finding|Functional Concept|Hospital Course|13199,13202|false|false|false|C0205535|Inhalation Route of Administration|INH
Disorder|Mental or Behavioral Dysfunction|Hospital Course|13206,13209|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|13206,13209|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|13206,13209|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|13206,13209|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|13206,13209|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|13215,13226|false|false|false|C0018305|guaifenesin|Guaifenesin
Drug|Pharmacologic Substance|Hospital Course|13215,13226|false|false|false|C0018305|guaifenesin|Guaifenesin
Event|Event|Hospital Course|13215,13226|false|false|false|||Guaifenesin
Drug|Organic Chemical|Hospital Course|13227,13234|false|false|false|C0009214|codeine|CODEINE
Drug|Pharmacologic Substance|Hospital Course|13227,13234|false|false|false|C0009214|codeine|CODEINE
Event|Event|Hospital Course|13227,13234|false|false|false|||CODEINE
Drug|Organic Chemical|Hospital Course|13227,13244|false|false|false|C0009217|codeine phosphate|CODEINE Phosphate
Drug|Pharmacologic Substance|Hospital Course|13227,13244|false|false|false|C0009217|codeine phosphate|CODEINE Phosphate
Drug|Element, Ion, or Isotope|Hospital Course|13235,13244|false|false|false|C0031603;C1601799|Phosphates;phosphate ion|Phosphate
Drug|Inorganic Chemical|Hospital Course|13235,13244|false|false|false|C0031603;C1601799|Phosphates;phosphate ion|Phosphate
Drug|Pharmacologic Substance|Hospital Course|13235,13244|false|false|false|C0031603;C1601799|Phosphates;phosphate ion|Phosphate
Event|Event|Hospital Course|13235,13244|false|false|false|||Phosphate
Procedure|Laboratory Procedure|Hospital Course|13235,13244|false|false|false|C0523826|Phosphate measurement|Phosphate
Finding|Gene or Genome|Hospital Course|13257,13260|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Organic Chemical|Hospital Course|13261,13266|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|Hospital Course|13261,13266|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|Hospital Course|13261,13266|false|false|false|||cough
Finding|Sign or Symptom|Hospital Course|13261,13266|false|false|false|C0010200|Coughing|cough
Drug|Organic Chemical|Hospital Course|13272,13291|false|false|false|C0020261|hydrochlorothiazide|Hydrochlorothiazide
Drug|Pharmacologic Substance|Hospital Course|13272,13291|false|false|false|C0020261|hydrochlorothiazide|Hydrochlorothiazide
Drug|Organic Chemical|Hospital Course|13312,13322|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Pharmacologic Substance|Hospital Course|13312,13322|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Organic Chemical|Hospital Course|13312,13334|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Drug|Pharmacologic Substance|Hospital Course|13312,13334|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Event|Event|Hospital Course|13323,13334|false|false|false|||Mononitrate
Finding|Finding|Hospital Course|13336,13344|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|13336,13344|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|Hospital Course|13345,13352|false|false|false|||Release
Finding|Functional Concept|Hospital Course|13345,13352|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|13345,13352|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|13345,13352|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|Hospital Course|13375,13386|false|false|false|C0090306|latanoprost|Latanoprost
Drug|Pharmacologic Substance|Hospital Course|13375,13386|false|false|false|C0090306|latanoprost|Latanoprost
Finding|Functional Concept|Hospital Course|13394,13399|false|false|false|C1522230|Ophthalmic Route of Administration|Ophth
Drug|Biomedical or Dental Material|Hospital Course|13409,13413|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|Hospital Course|13409,13413|false|false|false|C1705648|Dropping|DROP
Event|Event|Hospital Course|13414,13418|false|false|false|||LEFT
Finding|Functional Concept|Hospital Course|13414,13418|false|false|false|C1552822|Table Cell Horizontal Align - left|LEFT
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|13414,13422|false|false|false|C0229090|Left eye structure|LEFT EYE
Procedure|Diagnostic Procedure|Hospital Course|13414,13422|false|false|false|C2141124|examination of left eye|LEFT EYE
Anatomy|Body Location or Region|Hospital Course|13419,13422|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|EYE
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|13419,13422|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|EYE
Disorder|Disease or Syndrome|Hospital Course|13419,13422|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|EYE
Disorder|Neoplastic Process|Hospital Course|13419,13422|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|EYE
Event|Event|Hospital Course|13419,13422|false|false|false|||EYE
Finding|Body Substance|Hospital Course|13419,13422|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|EYE
Finding|Finding|Hospital Course|13419,13422|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|EYE
Finding|Intellectual Product|Hospital Course|13419,13422|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|EYE
Drug|Organic Chemical|Hospital Course|13431,13440|false|false|false|C0024002|lorazepam|Lorazepam
Drug|Pharmacologic Substance|Hospital Course|13431,13440|false|false|false|C0024002|lorazepam|Lorazepam
Event|Event|Hospital Course|13451,13454|false|false|false|||QHS
Finding|Gene or Genome|Hospital Course|13455,13458|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Pharmacologic Substance|Hospital Course|13459,13467|false|false|false|C1950154|Insomnia homeopathic medication|insomnia
Event|Event|Hospital Course|13459,13467|false|false|false|||insomnia
Finding|Sign or Symptom|Hospital Course|13459,13467|false|false|false|C0917801|Sleeplessness|insomnia
Drug|Organic Chemical|Hospital Course|13473,13486|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|Hospital Course|13473,13486|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|Hospital Course|13473,13486|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Event|Event|Hospital Course|13473,13486|false|false|false|||Multivitamins
Drug|Inorganic Chemical|Hospital Course|13489,13497|false|false|false|C0026162|Minerals|minerals
Event|Event|Hospital Course|13489,13497|false|false|false|||minerals
Drug|Biomedical or Dental Material|Hospital Course|13500,13503|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|Hospital Course|13500,13503|false|false|false|||TAB
Drug|Organic Chemical|Hospital Course|13518,13528|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Pharmacologic Substance|Hospital Course|13518,13528|false|false|false|C0034665|ranitidine|Ranitidine
Disorder|Mental or Behavioral Dysfunction|Hospital Course|13539,13542|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|13539,13542|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|13539,13542|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|13539,13542|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|13539,13542|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|13548,13560|false|false|false|C0039771|theophylline|Theophylline
Drug|Pharmacologic Substance|Hospital Course|13548,13560|false|false|false|C0039771|theophylline|Theophylline
Event|Event|Hospital Course|13548,13560|false|false|false|||Theophylline
Procedure|Laboratory Procedure|Hospital Course|13548,13560|false|false|false|C0039773|Assay of theophylline|Theophylline
Drug|Organic Chemical|Hospital Course|13548,13563|false|false|false|C2241157|Theophylline ER|Theophylline ER
Drug|Pharmacologic Substance|Hospital Course|13548,13563|false|false|false|C2241157|Theophylline ER|Theophylline ER
Event|Event|Hospital Course|13561,13563|false|false|false|||ER
Disorder|Mental or Behavioral Dysfunction|Hospital Course|13574,13577|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|13574,13577|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|13574,13577|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|13574,13577|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|13574,13577|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|13583,13593|false|false|false|C0213771|tiotropium|Tiotropium
Drug|Pharmacologic Substance|Hospital Course|13583,13593|false|false|false|C0213771|tiotropium|Tiotropium
Event|Event|Hospital Course|13583,13593|false|false|false|||Tiotropium
Drug|Organic Chemical|Hospital Course|13583,13601|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Pharmacologic Substance|Hospital Course|13583,13601|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Inorganic Chemical|Hospital Course|13594,13601|false|false|false|C0006222|Bromides|Bromide
Event|Event|Hospital Course|13594,13601|false|false|false|||Bromide
Procedure|Laboratory Procedure|Hospital Course|13594,13601|false|false|false|C0202341|Bromides measurement|Bromide
Disorder|Congenital Abnormality|Hospital Course|13604,13607|false|false|false|C1855179|CATARACT, ANTERIOR POLAR|CAP
Drug|Biomedical or Dental Material|Hospital Course|13604,13607|false|false|false|C0006935|capsule (pharmacologic)|CAP
Event|Event|Hospital Course|13604,13607|false|false|false|||CAP
Finding|Gene or Genome|Hospital Course|13604,13607|false|false|false|C1416891;C1418551;C1419093;C1422073;C1422760;C2985259;C4522312|BRD4 gene;BRD4 wt Allele;CAP1 gene;HACD1 gene;LNPEP gene;SERPINB6 gene;SORBS1 gene|CAP
Procedure|Therapeutic or Preventive Procedure|Hospital Course|13604,13607|false|false|false|C0278651;C0280547;C1879916|CAP Regimen;cisplatin/cyclophosphamide/doxorubicin protocol;cyclophosphamide/doxorubicin/prednisone protocol|CAP
Drug|Organic Chemical|Hospital Course|13622,13630|false|false|false|C0040610|tramadol|TraMADOL
Drug|Pharmacologic Substance|Hospital Course|13622,13630|false|false|false|C0040610|tramadol|TraMADOL
Event|Event|Hospital Course|13622,13630|false|false|false|||TraMADOL
Procedure|Laboratory Procedure|Hospital Course|13622,13630|false|false|false|C1266765|Tramadol measurement (procedure)|TraMADOL
Drug|Organic Chemical|Hospital Course|13632,13638|false|false|false|C0724054|Ultram|Ultram
Drug|Pharmacologic Substance|Hospital Course|13632,13638|false|false|false|C0724054|Ultram|Ultram
Finding|Gene or Genome|Hospital Course|13653,13656|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|13657,13661|false|false|false|C2598155||pain
Event|Event|Hospital Course|13657,13661|false|false|false|||pain
Finding|Functional Concept|Hospital Course|13657,13661|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|13657,13661|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Pharmacologic Substance|Hospital Course|13667,13683|false|false|false|C0003921;C2608262;C3853661|Artificial Tears;Lubricant Eye Drops;artificial tears (medication)|Artificial Tears
Finding|Body Substance|Hospital Course|13678,13683|false|false|false|C0039409;C1547924;C1611838|Tears (substance);Tears specimen|Tears
Finding|Intellectual Product|Hospital Course|13678,13683|false|false|false|C0039409;C1547924;C1611838|Tears (substance);Tears specimen|Tears
Event|Event|Hospital Course|13684,13691|false|false|false|||Preserv
Finding|Functional Concept|Hospital Course|13684,13691|false|false|false|C0728887|Preserving|Preserv
Procedure|Laboratory Procedure|Hospital Course|13684,13691|false|false|false|C0033085|Biologic Preservation|Preserv
Finding|Functional Concept|Hospital Course|13693,13697|false|false|false|C0332296|Free of (attribute)|Free
Drug|Biomedical or Dental Material|Hospital Course|13702,13706|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|Hospital Course|13702,13706|false|false|false|C1705648|Dropping|DROP
Event|Event|Hospital Course|13702,13706|false|false|false|||DROP
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|13707,13716|false|false|false|C0229118|Structure of both eyes|BOTH EYES
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|13712,13716|false|false|false|C0015392|Eye|EYES
Attribute|Clinical Attribute|Hospital Course|13712,13716|false|false|false|C5848506||EYES
Finding|Gene or Genome|Hospital Course|13717,13720|false|false|false|C1422467|CIAO3 gene|PRN
Anatomy|Body Location or Region|Hospital Course|13721,13724|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|eye
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|13721,13724|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|eye
Disorder|Disease or Syndrome|Hospital Course|13721,13724|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|eye
Disorder|Neoplastic Process|Hospital Course|13721,13724|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|eye
Event|Event|Hospital Course|13721,13724|false|false|false|||eye
Finding|Body Substance|Hospital Course|13721,13724|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Finding|Hospital Course|13721,13724|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Intellectual Product|Hospital Course|13721,13724|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Event|Event|Hospital Course|13726,13736|false|false|false|||irritation
Finding|Intellectual Product|Hospital Course|13726,13736|false|false|false|C1706307;C2700617;C5575347|Have Vulvar Irritation question;Irritability - emotion;Irritation (finding)|irritation
Finding|Mental Process|Hospital Course|13726,13736|false|false|false|C1706307;C2700617;C5575347|Have Vulvar Irritation question;Irritability - emotion;Irritation (finding)|irritation
Finding|Pathologic Function|Hospital Course|13726,13736|false|false|false|C1706307;C2700617;C5575347|Have Vulvar Irritation question;Irritability - emotion;Irritation (finding)|irritation
Phenomenon|Phenomenon or Process|Hospital Course|13726,13736|false|false|false|C0441723|Irritation|irritation
Drug|Organic Chemical|Hospital Course|13742,13749|false|false|false|C0011806;C0086140|Dextrans;dextran|dextran
Drug|Pharmacologic Substance|Hospital Course|13742,13749|false|false|false|C0011806;C0086140|Dextrans;dextran|dextran
Event|Event|Hospital Course|13742,13749|false|false|false|||dextran
Drug|Organic Chemical|Hospital Course|13742,13752|false|false|false|C0011795|dextran 70|dextran 70
Drug|Pharmacologic Substance|Hospital Course|13742,13752|false|false|false|C0011795|dextran 70|dextran 70
Drug|Organic Chemical|Hospital Course|13753,13765|false|false|false|C0063242|hypromellose|hypromellose
Drug|Pharmacologic Substance|Hospital Course|13753,13765|false|false|false|C0063242|hypromellose|hypromellose
Drug|Pharmacologic Substance|Hospital Course|13767,13783|false|false|false|C0003921;C2608262;C3853661|Artificial Tears;Lubricant Eye Drops;artificial tears (medication)|Artificial Tears
Event|Event|Hospital Course|13778,13783|false|false|false|||Tears
Finding|Body Substance|Hospital Course|13778,13783|false|false|false|C0039409;C1547924;C1611838|Tears (substance);Tears specimen|Tears
Finding|Intellectual Product|Hospital Course|13778,13783|false|false|false|C0039409;C1547924;C1611838|Tears (substance);Tears specimen|Tears
Drug|Biomedical or Dental Material|Hospital Course|13788,13792|false|false|false|C0991568|Drops - Drug Form|drop
Event|Activity|Hospital Course|13788,13792|false|false|false|C1705648|Dropping|drop
Event|Event|Hospital Course|13793,13797|false|false|false|||OPTH
Finding|Gene or Genome|Hospital Course|13803,13806|false|false|false|C1422467|CIAO3 gene|prn
Event|Event|Hospital Course|13807,13814|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|13807,13814|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|13822,13829|false|false|false|C0011806;C0086140|Dextrans;dextran|dextran
Drug|Pharmacologic Substance|Hospital Course|13822,13829|false|false|false|C0011806;C0086140|Dextrans;dextran|dextran
Event|Event|Hospital Course|13822,13829|false|false|false|||dextran
Drug|Organic Chemical|Hospital Course|13822,13832|false|false|false|C0011795|dextran 70|dextran 70
Drug|Pharmacologic Substance|Hospital Course|13822,13832|false|false|false|C0011795|dextran 70|dextran 70
Drug|Organic Chemical|Hospital Course|13833,13845|false|false|false|C0063242|hypromellose|hypromellose
Drug|Pharmacologic Substance|Hospital Course|13833,13845|false|false|false|C0063242|hypromellose|hypromellose
Drug|Pharmacologic Substance|Hospital Course|13847,13863|false|false|false|C0003921;C2608262;C3853661|Artificial Tears;Lubricant Eye Drops;artificial tears (medication)|Artificial Tears
Finding|Body Substance|Hospital Course|13858,13863|false|false|false|C0039409;C1547924;C1611838|Tears (substance);Tears specimen|Tears
Finding|Intellectual Product|Hospital Course|13858,13863|false|false|false|C0039409;C1547924;C1611838|Tears (substance);Tears specimen|Tears
Drug|Biomedical or Dental Material|Hospital Course|13875,13880|false|false|false|C0991568|Drops - Drug Form|drops
Event|Event|Hospital Course|13875,13880|false|false|false|||drops
Anatomy|Body Location or Region|Hospital Course|13882,13885|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|eye
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|13882,13885|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|eye
Disorder|Disease or Syndrome|Hospital Course|13882,13885|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|eye
Disorder|Neoplastic Process|Hospital Course|13882,13885|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|eye
Finding|Body Substance|Hospital Course|13882,13885|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Finding|Hospital Course|13882,13885|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Intellectual Product|Hospital Course|13882,13885|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Event|Event|Hospital Course|13889,13895|false|false|false|||needed
Finding|Intellectual Product|Hospital Course|13905,13912|false|false|false|C1704709|Computer program package|Package
Event|Event|Hospital Course|13913,13920|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|13913,13920|false|false|false|C0807726|refill|Refills
Drug|Antibiotic|Hospital Course|13928,13940|false|false|false|C0014806|erythromycin|Erythromycin
Drug|Organic Chemical|Hospital Course|13928,13940|false|false|false|C0014806|erythromycin|Erythromycin
Finding|Functional Concept|Hospital Course|13946,13951|false|false|false|C1522230|Ophthalmic Route of Administration|Ophth
Drug|Biomedical or Dental Material|Hospital Course|13952,13956|false|false|false|C0028912|Ointments|Oint
Event|Event|Hospital Course|13952,13956|false|false|false|||Oint
Finding|Functional Concept|Hospital Course|13964,13969|false|false|false|C1552823|Table Cell Horizontal Align - right|RIGHT
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|13964,13973|false|false|false|C0229089|Right eye|RIGHT EYE
Procedure|Diagnostic Procedure|Hospital Course|13964,13973|false|false|false|C2177784|examination of right eye|RIGHT EYE
Anatomy|Body Location or Region|Hospital Course|13970,13973|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|EYE
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|13970,13973|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|EYE
Disorder|Disease or Syndrome|Hospital Course|13970,13973|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|EYE
Disorder|Neoplastic Process|Hospital Course|13970,13973|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|EYE
Finding|Body Substance|Hospital Course|13970,13973|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|EYE
Finding|Finding|Hospital Course|13970,13973|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|EYE
Finding|Intellectual Product|Hospital Course|13970,13973|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|EYE
Event|Event|Hospital Course|13974,13977|false|false|false|||TID
Event|Event|Hospital Course|13979,13981|false|false|false|||RX
Drug|Antibiotic|Hospital Course|13983,13995|false|false|false|C0014806|erythromycin|erythromycin
Drug|Organic Chemical|Hospital Course|13983,13995|false|false|false|C0014806|erythromycin|erythromycin
Event|Event|Hospital Course|13983,13995|false|false|false|||erythromycin
Event|Event|Hospital Course|14034,14038|false|false|false|||OPTH
Event|Event|Hospital Course|14040,14043|false|false|false|||TID
Finding|Gene or Genome|Hospital Course|14044,14047|false|false|false|C1422467|CIAO3 gene|prn
Event|Event|Hospital Course|14048,14055|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|14048,14055|false|false|false|C0807726|refill|Refills
Drug|Inorganic Chemical|Hospital Course|14063,14070|false|false|false|C0719084|CalCarb|Calcarb
Event|Event|Hospital Course|14063,14070|false|false|false|||Calcarb
Drug|Organic Chemical|Hospital Course|14080,14087|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|Hospital Course|14080,14087|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|Hospital Course|14080,14087|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|Hospital Course|14080,14089|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|Hospital Course|14080,14089|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|Hospital Course|14080,14089|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|Hospital Course|14080,14089|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|Hospital Course|14080,14089|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Drug|Biologically Active Substance|Hospital Course|14091,14098|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Element, Ion, or Isotope|Hospital Course|14091,14098|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Inorganic Chemical|Hospital Course|14091,14098|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Pharmacologic Substance|Hospital Course|14091,14098|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Vitamin|Hospital Course|14091,14098|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Event|Event|Hospital Course|14091,14098|false|false|false|||calcium
Finding|Physiologic Function|Hospital Course|14091,14098|false|false|false|C4553026|Calcium metabolic function|calcium
Procedure|Laboratory Procedure|Hospital Course|14091,14098|false|false|false|C0201925|Calcium measurement|calcium
Drug|Inorganic Chemical|Hospital Course|14091,14108|false|false|false|C0006681|calcium carbonate|calcium carbonate
Drug|Pharmacologic Substance|Hospital Course|14091,14108|false|false|false|C0006681|calcium carbonate|calcium carbonate
Drug|Element, Ion, or Isotope|Hospital Course|14099,14108|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|carbonate
Drug|Organic Chemical|Hospital Course|14099,14108|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|carbonate
Drug|Pharmacologic Substance|Hospital Course|14099,14108|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|carbonate
Event|Event|Hospital Course|14099,14108|false|false|false|||carbonate
Drug|Organic Chemical|Hospital Course|14109,14116|false|false|false|C0042890|Vitamins|vitamin
Drug|Pharmacologic Substance|Hospital Course|14109,14116|false|false|false|C0042890|Vitamins|vitamin
Drug|Vitamin|Hospital Course|14109,14116|false|false|false|C0042890|Vitamins|vitamin
Event|Event|Hospital Course|14109,14116|false|false|false|||vitamin
Drug|Organic Chemical|Hospital Course|14109,14119|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Drug|Pharmacologic Substance|Hospital Course|14109,14119|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Drug|Vitamin|Hospital Course|14109,14119|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Anatomy|Body Space or Junction|Hospital Course|14133,14137|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|14133,14137|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|14133,14137|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|14133,14137|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Drug|Amino Acid, Peptide, or Protein|Hospital Course|14149,14152|false|false|false|C0056632;C0459207;C2702357;C3488428|Cyclophosphamide/Dacarbazine/Vincristine;cod, unspecified preparation;codfish allergenic extract|cod
Drug|Food|Hospital Course|14149,14152|false|false|false|C0056632;C0459207;C2702357;C3488428|Cyclophosphamide/Dacarbazine/Vincristine;cod, unspecified preparation;codfish allergenic extract|cod
Drug|Immunologic Factor|Hospital Course|14149,14152|false|false|false|C0056632;C0459207;C2702357;C3488428|Cyclophosphamide/Dacarbazine/Vincristine;cod, unspecified preparation;codfish allergenic extract|cod
Drug|Pharmacologic Substance|Hospital Course|14149,14152|false|false|false|C0056632;C0459207;C2702357;C3488428|Cyclophosphamide/Dacarbazine/Vincristine;cod, unspecified preparation;codfish allergenic extract|cod
Finding|Finding|Hospital Course|14149,14152|false|false|false|C0007465;C0457523;C1420285;C5444130|Cancerization of Pancreatic Ducts;Cause of Death;Cemento-osseous dysplasia;SNRPB gene|cod
Finding|Gene or Genome|Hospital Course|14149,14152|false|false|false|C0007465;C0457523;C1420285;C5444130|Cancerization of Pancreatic Ducts;Cause of Death;Cemento-osseous dysplasia;SNRPB gene|cod
Finding|Pathologic Function|Hospital Course|14149,14152|false|false|false|C0007465;C0457523;C1420285;C5444130|Cancerization of Pancreatic Ducts;Cause of Death;Cemento-osseous dysplasia;SNRPB gene|cod
Drug|Food|Hospital Course|14149,14162|false|false|false|C0009213|cod liver oil|cod liver oil
Drug|Organic Chemical|Hospital Course|14149,14162|false|false|false|C0009213|cod liver oil|cod liver oil
Drug|Pharmacologic Substance|Hospital Course|14149,14162|false|false|false|C0009213|cod liver oil|cod liver oil
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|14153,14158|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|Hospital Course|14153,14158|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|Hospital Course|14153,14158|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|Hospital Course|14153,14158|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|Hospital Course|14153,14158|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|Hospital Course|14153,14158|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|Hospital Course|14153,14158|false|false|false|||liver
Finding|Finding|Hospital Course|14153,14158|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|Hospital Course|14153,14158|false|false|false|C0872387|Procedures on liver|liver
Drug|Biomedical or Dental Material|Hospital Course|14159,14162|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|oil
Drug|Food|Hospital Course|14159,14162|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|oil
Drug|Organic Chemical|Hospital Course|14159,14162|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|oil
Drug|Pharmacologic Substance|Hospital Course|14159,14162|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|oil
Anatomy|Body Space or Junction|Hospital Course|14178,14182|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|14178,14182|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|14178,14182|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|14178,14182|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Disorder|Mental or Behavioral Dysfunction|Hospital Course|14183,14186|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|14183,14186|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|14183,14186|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|14183,14186|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|14183,14186|false|false|false|C1332410|BID gene|BID
Event|Event|Hospital Course|14191,14200|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|14191,14200|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|14191,14200|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|14191,14200|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|14191,14200|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|14191,14212|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|14191,14212|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|14201,14212|false|false|false|C2926604||Disposition
Event|Event|Hospital Course|14201,14212|false|false|false|||Disposition
Procedure|Health Care Activity|Hospital Course|14201,14212|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|Hospital Course|14214,14218|false|false|false|||Home
Finding|Idea or Concept|Hospital Course|14214,14218|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|14214,14218|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|14214,14218|false|false|false|C1553498|home health encounter|Home
Event|Event|Hospital Course|14221,14230|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|14221,14230|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|14221,14230|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|14221,14230|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|14221,14230|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|14221,14240|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|14231,14240|false|false|false|C0945731||Diagnosis
Event|Event|Hospital Course|14231,14240|false|false|false|||Diagnosis
Finding|Classification|Hospital Course|14231,14240|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|14231,14240|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|14231,14240|false|false|false|C0011900|Diagnosis|Diagnosis
Disorder|Disease or Syndrome|Hospital Course|14242,14267|false|false|false|C1281999|Rapid atrial fibrillation|Rapid Atrial Fibrillation
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|14248,14254|false|false|false|C0018792|Heart Atrium|Atrial
Attribute|Clinical Attribute|Hospital Course|14248,14267|false|false|false|C2926591||Atrial Fibrillation
Disorder|Disease or Syndrome|Hospital Course|14248,14267|false|false|false|C0004238|Atrial Fibrillation|Atrial Fibrillation
Lab|Laboratory or Test Result|Hospital Course|14248,14267|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Atrial Fibrillation
Finding|Pathologic Function|Hospital Course|14248,14275|false|false|false|C0155709|Atrial fibrillation and flutter|Atrial Fibrillation/Flutter
Disorder|Disease or Syndrome|Hospital Course|14255,14267|false|false|false|C0232197|Fibrillation|Fibrillation
Event|Event|Hospital Course|14255,14267|false|false|false|||Fibrillation
Finding|Pathologic Function|Hospital Course|14268,14275|false|false|false|C0016385|Cardiac Flutter|Flutter
Disorder|Disease or Syndrome|Hospital Course|14276,14280|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Hospital Course|14276,14280|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Hospital Course|14276,14280|false|false|false|||COPD
Finding|Gene or Genome|Hospital Course|14276,14280|false|false|false|C1412502|ARCN1 gene|COPD
Finding|Mental Process|Discharge Condition|14305,14311|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|14305,14318|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|14305,14318|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|14312,14318|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|14312,14318|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|14320,14325|false|false|false|||Clear
Finding|Idea or Concept|Discharge Condition|14320,14325|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|Discharge Condition|14330,14338|false|false|false|||coherent
Finding|Finding|Discharge Condition|14330,14338|false|false|false|C4068804|Coherent|coherent
Event|Event|Discharge Condition|14340,14345|false|false|false|||Level
Attribute|Clinical Attribute|Discharge Condition|14340,14362|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|14340,14362|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|Discharge Condition|14349,14362|false|false|false|||Consciousness
Finding|Finding|Discharge Condition|14349,14362|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|14349,14362|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|14364,14369|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|14364,14369|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|14364,14369|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|Discharge Condition|14364,14369|false|false|false|||Alert
Finding|Finding|Discharge Condition|14364,14369|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|14364,14369|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|14364,14369|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|Discharge Condition|14374,14385|false|false|false|||interactive
Finding|Functional Concept|Discharge Condition|14374,14385|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|14387,14395|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|14387,14395|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|14387,14395|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|14396,14402|false|false|false|C5889824||Status
Event|Event|Discharge Condition|14396,14402|false|false|false|||Status
Finding|Idea or Concept|Discharge Condition|14396,14402|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|14404,14414|false|false|false|||Ambulatory
Finding|Functional Concept|Discharge Condition|14404,14414|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|Discharge Condition|14404,14414|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|Discharge Condition|14404,14414|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|Discharge Condition|14404,14414|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|Discharge Condition|14417,14428|false|false|false|||Independent
Finding|Finding|Discharge Condition|14417,14428|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|Discharge Condition|14417,14428|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Gene or Genome|Discharge Instructions|14457,14461|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Event|Event|Discharge Instructions|14481,14489|false|false|false|||admitted
Anatomy|Body Location or Region|Discharge Instructions|14515,14520|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Discharge Instructions|14515,14520|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Discharge Instructions|14515,14525|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|Discharge Instructions|14515,14525|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Discharge Instructions|14521,14525|false|true|false|C2598155||pain
Finding|Functional Concept|Discharge Instructions|14521,14525|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|14521,14525|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|14521,14534|false|false|false|C0030193|Pain|pain symptoms
Event|Event|Discharge Instructions|14526,14534|false|false|false|||symptoms
Finding|Functional Concept|Discharge Instructions|14526,14534|false|true|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Discharge Instructions|14526,14534|false|true|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|Discharge Instructions|14573,14579|false|false|false|||bursts
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|14591,14596|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Discharge Instructions|14591,14596|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Event|Event|Discharge Instructions|14591,14596|false|false|false|||heart
Finding|Sign or Symptom|Discharge Instructions|14591,14596|false|false|false|C0795691|HEART PROBLEM|heart
Event|Activity|Discharge Instructions|14598,14602|false|false|false|C0871208|Rating (action)|rate
Event|Event|Discharge Instructions|14598,14602|false|false|false|||rate
Finding|Idea or Concept|Discharge Instructions|14598,14602|false|false|false|C1549480|Amount type - Rate|rate
Event|Activity|Discharge Instructions|14620,14624|false|false|false|C0871208|Rating (action)|rate
Event|Event|Discharge Instructions|14620,14624|false|false|false|||rate
Finding|Idea or Concept|Discharge Instructions|14620,14624|false|false|false|C1549480|Amount type - Rate|rate
Event|Event|Discharge Instructions|14625,14630|false|false|false|||makes
Finding|Finding|Discharge Instructions|14638,14652|false|false|false|C4699158|Increased risk|increased risk
Event|Event|Discharge Instructions|14648,14652|false|false|false|||risk
Finding|Idea or Concept|Discharge Instructions|14648,14652|false|false|false|C0035647|Risk|risk
Disorder|Disease or Syndrome|Discharge Instructions|14658,14664|false|false|false|C0038454|Cerebrovascular accident|stroke
Event|Event|Discharge Instructions|14658,14664|false|false|false|||stroke
Finding|Finding|Discharge Instructions|14658,14664|false|false|false|C5977286|Stroke (heart beat)|stroke
Event|Event|Discharge Instructions|14675,14682|false|false|false|||started
Disorder|Disease or Syndrome|Discharge Instructions|14688,14693|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Discharge Instructions|14688,14693|false|false|false|||blood
Finding|Body Substance|Discharge Instructions|14688,14693|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Sign or Symptom|Discharge Instructions|14694,14702|false|false|false|C0851184|Thinning Weight Loss|thinning
Drug|Pharmacologic Substance|Discharge Instructions|14703,14713|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Discharge Instructions|14703,14713|false|false|false|||medication
Finding|Intellectual Product|Discharge Instructions|14703,14713|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|Discharge Instructions|14714,14720|false|false|false|||called
Drug|Organic Chemical|Discharge Instructions|14722,14733|false|false|false|C1739768|rivaroxaban|Rivaroxaban
Drug|Pharmacologic Substance|Discharge Instructions|14722,14733|false|false|false|C1739768|rivaroxaban|Rivaroxaban
Event|Event|Discharge Instructions|14749,14753|false|false|false|||need
Event|Event|Discharge Instructions|14757,14761|false|false|false|||take
Finding|Idea or Concept|Discharge Instructions|14768,14771|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Discharge Instructions|14768,14771|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Conceptual Entity|Discharge Instructions|14778,14789|false|false|false|C1704211|Specialized|specialized
Event|Event|Discharge Instructions|14790,14803|false|false|false|||cardiologists
Event|Event|Discharge Instructions|14808,14812|false|false|false|||deal
Finding|Functional Concept|Discharge Instructions|14836,14846|false|false|false|C0442828|Electrical (qualifier value)|electrical
Phenomenon|Natural Phenomenon or Process|Discharge Instructions|14836,14846|false|false|false|C0013790|Electricity|electrical
Event|Event|Discharge Instructions|14847,14853|false|false|false|||rhythm
Finding|Finding|Discharge Instructions|14847,14853|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|Discharge Instructions|14847,14853|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|14861,14866|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Discharge Instructions|14861,14866|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Discharge Instructions|14861,14866|false|false|false|C0795691|HEART PROBLEM|heart
Event|Event|Discharge Instructions|14867,14876|false|false|false|||evaluated
Event|Event|Discharge Instructions|14885,14889|false|false|false|||felt
Event|Event|Discharge Instructions|14906,14913|false|false|false|||benefit
Drug|Pharmacologic Substance|Discharge Instructions|14921,14931|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Discharge Instructions|14921,14931|false|false|false|||medication
Finding|Intellectual Product|Discharge Instructions|14921,14931|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|Discharge Instructions|14932,14938|false|false|false|||called
Drug|Organic Chemical|Discharge Instructions|14939,14949|false|false|false|C0002598|amiodarone|amiodarone
Drug|Pharmacologic Substance|Discharge Instructions|14939,14949|false|false|false|C0002598|amiodarone|amiodarone
Event|Event|Discharge Instructions|14939,14949|false|false|false|||amiodarone
Procedure|Laboratory Procedure|Discharge Instructions|14939,14949|false|false|false|C5399868|Drug assay amiodarone|amiodarone
Event|Event|Discharge Instructions|14966,14973|false|false|false|||started
Event|Event|Discharge Instructions|14984,14988|false|false|false|||need
Event|Event|Discharge Instructions|14992,14998|false|false|false|||follow
Finding|Finding|Discharge Instructions|15044,15052|false|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Finding|Idea or Concept|Discharge Instructions|15044,15052|false|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Event|Event|Discharge Instructions|15053,15059|false|false|false|||rhythm
Finding|Finding|Discharge Instructions|15053,15059|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|Discharge Instructions|15053,15059|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Event|Event|Discharge Instructions|15088,15097|false|false|false|||outfitted
Procedure|Diagnostic Procedure|Discharge Instructions|15105,15119|false|false|false|C0013801|Holter Electrocardiography|Holter monitor
Drug|Hazardous or Poisonous Substance|Discharge Instructions|15112,15119|false|false|false|C0728873|Monitor brand of insecticide|monitor
Drug|Organic Chemical|Discharge Instructions|15112,15119|false|false|false|C0728873|Monitor brand of insecticide|monitor
Event|Event|Discharge Instructions|15112,15119|false|false|false|||monitor
Event|Event|Discharge Instructions|15123,15129|false|false|false|||record
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|15135,15140|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Discharge Instructions|15135,15140|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Discharge Instructions|15135,15140|false|false|false|C0795691|HEART PROBLEM|heart
Attribute|Clinical Attribute|Discharge Instructions|15135,15145|false|false|false|C0018810;C0488794|heart rate|heart rate
Finding|Finding|Discharge Instructions|15135,15145|false|false|false|C2041121||heart rate
Procedure|Health Care Activity|Discharge Instructions|15135,15145|false|false|false|C2197023|examination of heart rate|heart rate
Event|Activity|Discharge Instructions|15141,15145|false|false|false|C0871208|Rating (action)|rate
Event|Event|Discharge Instructions|15141,15145|false|false|false|||rate
Finding|Idea or Concept|Discharge Instructions|15141,15145|false|false|false|C1549480|Amount type - Rate|rate
Event|Event|Discharge Instructions|15150,15154|false|false|false|||home
Finding|Idea or Concept|Discharge Instructions|15150,15154|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Discharge Instructions|15150,15154|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Discharge Instructions|15150,15154|false|false|false|C1553498|home health encounter|home
Finding|Finding|Discharge Instructions|15162,15176|false|false|false|C3844729|Very Important|very important
Event|Event|Discharge Instructions|15167,15176|false|false|false|||important
Event|Event|Discharge Instructions|15186,15192|false|false|false|||follow
Event|Event|Discharge Instructions|15215,15227|false|false|false|||cardiologist
Disorder|Disease or Syndrome|Discharge Instructions|15250,15254|false|false|false|C0339510|Vitelliform Macular Dystrophy|best
Event|Event|Discharge Instructions|15250,15254|false|false|false|||best
Finding|Gene or Genome|Discharge Instructions|15250,15254|false|false|false|C1826421;C5781213|BEST1 gene;BEST1 wt Allele|best
Event|Activity|Discharge Instructions|15273,15277|false|false|false|C1947933|care activity|care
Finding|Finding|Discharge Instructions|15273,15277|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|15273,15277|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Attribute|Clinical Attribute|Discharge Instructions|15273,15282|false|false|false|C4321316||care team
Finding|Finding|Discharge Instructions|15273,15282|false|false|false|C4321315|Care team|care team
Procedure|Health Care Activity|Discharge Instructions|15292,15300|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|15301,15313|false|false|false|C3263700||Instructions
Event|Event|Discharge Instructions|15301,15313|false|false|false|||Instructions
Finding|Intellectual Product|Discharge Instructions|15301,15313|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

