 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|26,30
No|31,33
:|33,34
_|37,38
_|38,39
_|39,40
<EOL>|40,41
<EOL>|42,43
Admission|43,52
Date|53,57
:|57,58
_|60,61
_|61,62
_|62,63
Discharge|77,86
Date|87,91
:|91,92
_|95,96
_|96,97
_|97,98
<EOL>|98,99
<EOL>|100,101
Date|101,105
of|106,108
Birth|109,114
:|114,115
_|117,118
_|118,119
_|119,120
Sex|133,136
:|136,137
M|140,141
<EOL>|141,142
<EOL>|143,144
Service|144,151
:|151,152
SURGERY|153,160
<EOL>|160,161
<EOL>|162,163
Allergies|163,172
:|172,173
<EOL>|174,175
Corgard|175,182
/|183,184
Vasotec|185,192
<EOL>|192,193
<EOL>|194,195
Attending|195,204
:|204,205
_|206,207
_|207,208
_|208,209
.|209,210
<EOL>|210,211
<EOL>|212,213
Chief|213,218
Complaint|219,228
:|228,229
<EOL>|229,230
incarcerated|230,242
inguinal|243,251
hernia|252,258
<EOL>|258,259
<EOL>|260,261
Major|261,266
Surgical|267,275
or|276,278
Invasive|279,287
Procedure|288,297
:|297,298
<EOL>|298,299
Left|299,303
inguinal|304,312
hernia|313,319
repair|320,326
<EOL>|326,327
<EOL>|328,329
History|329,336
of|337,339
Present|340,347
Illness|348,355
:|355,356
<EOL>|356,357
_|357,358
_|358,359
_|359,360
with|361,365
afib|366,370
on|371,373
apixiban|374,382
,|382,383
CAD|384,387
s|388,389
/|389,390
p|390,391
CABG|392,396
,|396,397
b|398,399
/|399,400
l|400,401
carotid|402,409
disease|410,417
,|417,418
<EOL>|419,420
COPD|420,424
/|424,425
emphysema|425,434
with|435,439
recent|440,446
pneumonia|447,456
presents|457,465
for|466,469
elective|470,478
left|479,483
<EOL>|484,485
inguinal|485,493
hernia|494,500
repair|501,507
(|508,509
large|509,514
,|514,515
with|516,520
incarcerated|521,533
sigmoid|534,541
colon|542,547
)|547,548
<EOL>|548,549
<EOL>|549,550
<EOL>|551,552
Past|552,556
Medical|557,564
History|565,572
:|572,573
<EOL>|573,574
Past|574,578
Medical|579,586
History|587,594
:|594,595
<EOL>|595,596
BILATERAL|596,605
MODERATE|606,614
CAROTID|615,622
DISEASE|623,630
<EOL>|631,632
CONGESTIVE|632,642
HEART|643,648
FAILURE|649,656
<EOL>|657,658
CORONARY|658,666
ARTERY|667,673
DISEASE|674,681
<EOL>|682,683
GASTROESOPHAGEAL|683,699
REFLUX|700,706
<EOL>|707,708
HYPERTENSION|708,720
<EOL>|721,722
SEVERE|722,728
EMPHYSEMA|729,738
<EOL>|739,740
PULMONARY|740,749
HYPERTENSION|750,762
<EOL>|763,764
RIGHT|764,769
BUNDLE|770,776
BRANCH|777,783
BLOCK|784,789
<EOL>|790,791
BENIGN|791,797
PROSTATIC|798,807
HYPERTROPHY|808,819
<EOL>|820,821
HYPERLIPIDEMIA|821,835
<EOL>|836,837
PAROXYSMAL|837,847
ATRIAL|848,854
FIBRILLATION|855,867
<EOL>|868,869
H|869,870
/|870,871
O|871,872
HISTIOPLASMOSIS|873,888
<EOL>|889,890
<EOL>|890,891
Past|891,895
Surgical|896,904
History|905,912
:|912,913
<EOL>|913,914
CARDIOVERSION|914,927
_|928,929
_|929,930
_|930,931
<EOL>|932,933
RIGHT|933,938
LOWER|939,944
LOBE|945,949
LOBECTOMY|950,959
_|960,961
_|961,962
_|962,963
<EOL>|964,965
CORONARY|965,973
BYPASS|974,980
SURGERY|981,988
_|989,990
_|990,991
_|991,992
<EOL>|993,994
<EOL>|994,995
<EOL>|996,997
Social|997,1003
History|1004,1011
:|1011,1012
<EOL>|1012,1013
_|1013,1014
_|1014,1015
_|1015,1016
<EOL>|1016,1017
Family|1017,1023
History|1024,1031
:|1031,1032
<EOL>|1032,1033
Non-contributory|1033,1049
<EOL>|1049,1050
<EOL>|1051,1052
Physical|1052,1060
Exam|1061,1065
:|1065,1066
<EOL>|1066,1067
Gen|1067,1070
:|1070,1071
Awake|1072,1077
and|1078,1081
alert|1082,1087
<EOL>|1087,1088
CV|1088,1090
:|1090,1091
Irregularly|1092,1103
irregular|1104,1113
rhythm|1114,1120
,|1120,1121
normal|1122,1128
rate|1129,1133
<EOL>|1133,1134
Resp|1134,1138
:|1138,1139
CTAB|1140,1144
<EOL>|1144,1145
GI|1145,1147
:|1147,1148
Soft|1149,1153
,|1153,1154
appropriately|1155,1168
tender|1169,1175
near|1176,1180
incision|1181,1189
,|1189,1190
non-distended|1191,1204
<EOL>|1204,1205
Incision|1205,1213
clean|1214,1219
,|1219,1220
dry|1221,1224
,|1224,1225
and|1226,1229
intact|1230,1236
with|1237,1241
no|1242,1244
erythema|1245,1253
<EOL>|1253,1254
Ext|1254,1257
:|1257,1258
Warm|1259,1263
and|1264,1267
well|1268,1272
perfused|1273,1281
<EOL>|1281,1282
<EOL>|1283,1284
Pertinent|1284,1293
Results|1294,1301
:|1301,1302
<EOL>|1302,1303
<EOL>|1304,1305
<EOL>|1306,1307
Brief|1307,1312
Hospital|1313,1321
Course|1322,1328
:|1328,1329
<EOL>|1329,1330
Mr.|1330,1333
_|1334,1335
_|1335,1336
_|1336,1337
was|1338,1341
admitted|1342,1350
to|1351,1353
_|1354,1355
_|1355,1356
_|1356,1357
<EOL>|1358,1359
_|1359,1360
_|1360,1361
_|1361,1362
on|1363,1365
_|1366,1367
_|1367,1368
_|1368,1369
after|1370,1375
undergoing|1376,1386
repair|1387,1393
of|1394,1396
a|1397,1398
left|1399,1403
<EOL>|1404,1405
incarcerated|1405,1417
inguinal|1418,1426
hernia|1427,1433
.|1433,1434
For|1435,1438
details|1439,1446
of|1447,1449
the|1450,1453
procedure|1454,1463
,|1463,1464
<EOL>|1465,1466
please|1466,1472
refer|1473,1478
to|1479,1481
the|1482,1485
operative|1486,1495
report|1496,1502
.|1502,1503
His|1504,1507
postoperative|1508,1521
course|1522,1528
<EOL>|1529,1530
was|1530,1533
uncomplicated|1534,1547
.|1547,1548
After|1549,1554
a|1555,1556
brief|1557,1562
stay|1563,1567
in|1568,1570
the|1571,1574
PACU|1575,1579
,|1579,1580
he|1581,1583
was|1584,1587
<EOL>|1588,1589
transferred|1589,1600
to|1601,1603
the|1604,1607
regular|1608,1615
nursing|1616,1623
floor|1624,1629
.|1629,1630
His|1631,1634
pain|1635,1639
was|1640,1643
<EOL>|1644,1645
controlled|1645,1655
with|1656,1660
IV|1661,1663
medication|1664,1674
.|1674,1675
On|1676,1678
POD|1679,1682
#|1683,1684
1|1684,1685
,|1685,1686
he|1687,1689
was|1690,1693
started|1694,1701
on|1702,1704
a|1705,1706
<EOL>|1707,1708
regular|1708,1715
diet|1716,1720
,|1720,1721
and|1722,1725
his|1726,1729
pain|1730,1734
was|1735,1738
controlled|1739,1749
with|1750,1754
PO|1755,1757
pain|1758,1762
<EOL>|1763,1764
medication|1764,1774
.|1774,1775
He|1776,1778
voided|1779,1785
without|1786,1793
issue|1794,1799
.|1799,1800
He|1801,1803
was|1804,1807
ambulating|1808,1818
<EOL>|1819,1820
independently|1820,1833
in|1834,1836
the|1837,1840
halls|1841,1846
.|1846,1847
He|1848,1850
was|1851,1854
given|1855,1860
a|1861,1862
bowel|1863,1868
regimen|1869,1876
,|1876,1877
and|1878,1881
<EOL>|1882,1883
passed|1883,1889
flatus|1890,1896
.|1896,1897
On|1898,1900
POD|1901,1904
#|1905,1906
2|1906,1907
,|1907,1908
he|1909,1911
continued|1912,1921
to|1922,1924
tolerate|1925,1933
his|1934,1937
diet|1938,1942
,|1942,1943
his|1944,1947
<EOL>|1948,1949
pain|1949,1953
was|1954,1957
well|1958,1962
-|1962,1963
controlled|1963,1973
on|1974,1976
oral|1977,1981
medication|1982,1992
,|1992,1993
and|1994,1997
he|1998,2000
continued|2001,2010
to|2011,2013
<EOL>|2014,2015
ambulate|2015,2023
independently|2024,2037
.|2037,2038
He|2039,2041
was|2042,2045
discharged|2046,2056
home|2057,2061
in|2062,2064
stable|2065,2071
<EOL>|2072,2073
condition|2073,2082
on|2083,2085
POD|2086,2089
#|2090,2091
2|2091,2092
with|2093,2097
plans|2098,2103
to|2104,2106
follow|2107,2113
-|2113,2114
up|2114,2116
with|2117,2121
Dr.|2122,2125
_|2126,2127
_|2127,2128
_|2128,2129
.|2129,2130
<EOL>|2131,2132
<EOL>|2133,2134
Discharge|2134,2143
Medications|2144,2155
:|2155,2156
<EOL>|2156,2157
1.|2157,2159
Amiodarone|2160,2170
200|2171,2174
mg|2175,2177
PO|2178,2180
DAILY|2181,2186
<EOL>|2187,2188
2.|2188,2190
Apixaban|2191,2199
5|2200,2201
mg|2202,2204
PO|2205,2207
BID|2208,2211
<EOL>|2212,2213
3.|2213,2215
Aspirin|2216,2223
81|2224,2226
mg|2227,2229
PO|2230,2232
DAILY|2233,2238
<EOL>|2239,2240
4.|2240,2242
Docusate|2243,2251
Sodium|2252,2258
100|2259,2262
mg|2263,2265
PO|2266,2268
BID|2269,2272
<EOL>|2273,2274
5.|2274,2276
Losartan|2277,2285
Potassium|2286,2295
25|2296,2298
mg|2299,2301
PO|2302,2304
DAILY|2305,2310
<EOL>|2311,2312
6.|2312,2314
Omeprazole|2315,2325
10|2326,2328
mg|2329,2331
PO|2332,2334
DAILY|2335,2340
<EOL>|2341,2342
7.|2342,2344
Triamterene|2345,2356
-|2356,2357
HCTZ|2357,2361
(|2362,2363
37.5|2363,2367
/|2367,2368
25|2368,2370
)|2370,2371
1|2372,2373
CAP|2374,2377
PO|2378,2380
DAILY|2381,2386
<EOL>|2387,2388
8.|2388,2390
Acetaminophen|2391,2404
1000|2405,2409
mg|2410,2412
PO|2413,2415
Q6H|2416,2419
:|2419,2420
PRN|2420,2423
pain|2424,2428
or|2429,2431
fever|2432,2437
<EOL>|2438,2439
Do|2439,2441
not|2442,2445
exceed|2446,2452
4|2453,2454
grams|2455,2460
per|2461,2464
day|2465,2468
.|2468,2469
<EOL>|2470,2471
RX|2471,2473
*|2474,2475
acetaminophen|2475,2488
500|2489,2492
mg|2493,2495
_|2496,2497
_|2497,2498
_|2498,2499
tablet|2500,2506
(|2506,2507
s|2507,2508
)|2508,2509
by|2510,2512
mouth|2513,2518
every|2519,2524
6|2525,2526
hours|2527,2532
<EOL>|2533,2534
Disp|2534,2538
#|2539,2540
*|2540,2541
60|2541,2543
Tablet|2544,2550
Refills|2551,2558
:|2558,2559
*|2559,2560
0|2560,2561
<EOL>|2561,2562
9.|2562,2564
OxycoDONE|2565,2574
(|2575,2576
Immediate|2576,2585
Release|2586,2593
)|2593,2594
5|2596,2597
mg|2598,2600
PO|2601,2603
Q4H|2604,2607
:|2607,2608
PRN|2608,2611
pain|2612,2616
<EOL>|2617,2618
RX|2618,2620
*|2621,2622
oxycodone|2622,2631
5|2632,2633
mg|2634,2636
_|2637,2638
_|2638,2639
_|2639,2640
tablet|2641,2647
(|2647,2648
s|2648,2649
)|2649,2650
by|2651,2653
mouth|2654,2659
every|2660,2665
4|2666,2667
hours|2668,2673
Disp|2674,2678
<EOL>|2679,2680
#|2680,2681
*|2681,2682
40|2682,2684
Tablet|2685,2691
Refills|2692,2699
:|2699,2700
*|2700,2701
0|2701,2702
<EOL>|2702,2703
10.|2703,2706
Senna|2707,2712
17.2|2713,2717
mg|2718,2720
PO|2721,2723
HS|2724,2726
<EOL>|2727,2728
Take|2728,2732
this|2733,2737
while|2738,2743
you|2744,2747
are|2748,2751
taking|2752,2758
oxycodone|2759,2768
.|2768,2769
<EOL>|2770,2771
RX|2771,2773
*|2774,2775
sennosides|2775,2785
[|2786,2787
Evac|2787,2791
-|2791,2792
U-Gen|2792,2797
(|2798,2799
sennosides|2799,2809
)|2809,2810
]|2810,2811
8.6|2812,2815
mg|2816,2818
1|2819,2820
capsule|2821,2828
by|2829,2831
<EOL>|2832,2833
mouth|2833,2838
daily|2839,2844
Disp|2845,2849
#|2850,2851
*|2851,2852
30|2852,2854
Tablet|2855,2861
Refills|2862,2869
:|2869,2870
*|2870,2871
0|2871,2872
<EOL>|2872,2873
11.|2873,2876
Align|2877,2882
(|2883,2884
bifidobacterium|2884,2899
infantis|2900,2908
)|2908,2909
4|2910,2911
mg|2912,2914
oral|2915,2919
DAILY|2920,2925
<EOL>|2926,2927
12.|2927,2930
coenzyme|2931,2939
Q10|2940,2943
100|2944,2947
mg|2948,2950
oral|2951,2955
DAILY|2956,2961
<EOL>|2962,2963
13.|2963,2966
Rosuvastatin|2967,2979
Calcium|2980,2987
40|2988,2990
mg|2991,2993
PO|2994,2996
QPM|2997,3000
<EOL>|3001,3002
14.|3002,3005
Vitamin|3006,3013
D|3014,3015
1000|3016,3020
UNIT|3021,3025
PO|3026,3028
DAILY|3029,3034
<EOL>|3035,3036
<EOL>|3036,3037
<EOL>|3038,3039
Discharge|3039,3048
Disposition|3049,3060
:|3060,3061
<EOL>|3061,3062
Home|3062,3066
With|3067,3071
Service|3072,3079
<EOL>|3079,3080
<EOL>|3081,3082
Facility|3082,3090
:|3090,3091
<EOL>|3091,3092
_|3092,3093
_|3093,3094
_|3094,3095
<EOL>|3095,3096
<EOL>|3097,3098
Discharge|3098,3107
Diagnosis|3108,3117
:|3117,3118
<EOL>|3118,3119
Inguinal|3119,3127
hernia|3128,3134
<EOL>|3134,3135
<EOL>|3136,3137
Discharge|3137,3146
Condition|3147,3156
:|3156,3157
<EOL>|3157,3158
Mental|3158,3164
Status|3165,3171
:|3171,3172
Clear|3173,3178
and|3179,3182
coherent|3183,3191
.|3191,3192
<EOL>|3192,3193
Level|3193,3198
of|3199,3201
Consciousness|3202,3215
:|3215,3216
Alert|3217,3222
and|3223,3226
interactive|3227,3238
.|3238,3239
<EOL>|3239,3240
Activity|3240,3248
Status|3249,3255
:|3255,3256
Ambulatory|3257,3267
-|3268,3269
Independent|3270,3281
.|3281,3282
<EOL>|3282,3283
<EOL>|3284,3285
Discharge|3285,3294
Instructions|3295,3307
:|3307,3308
<EOL>|3308,3309
Dear|3309,3313
Mr.|3314,3317
_|3318,3319
_|3319,3320
_|3320,3321
,|3321,3322
<EOL>|3322,3323
It|3323,3325
was|3326,3329
a|3330,3331
pleasure|3332,3340
taking|3341,3347
care|3348,3352
of|3353,3355
you|3356,3359
here|3360,3364
at|3365,3367
_|3368,3369
_|3369,3370
_|3370,3371
<EOL>|3372,3373
_|3373,3374
_|3374,3375
_|3375,3376
.|3376,3377
You|3378,3381
were|3382,3386
admitted|3387,3395
to|3396,3398
our|3399,3402
hospital|3403,3411
<EOL>|3412,3413
after|3413,3418
undergoing|3419,3429
repair|3430,3436
of|3437,3439
your|3440,3444
inguinal|3445,3453
hernia|3454,3460
.|3460,3461
You|3462,3465
have|3466,3470
<EOL>|3471,3472
recovered|3472,3481
from|3482,3486
surgery|3487,3494
and|3495,3498
are|3499,3502
now|3503,3506
ready|3507,3512
to|3513,3515
be|3516,3518
discharged|3519,3529
home|3530,3534
.|3534,3535
<EOL>|3536,3537
Please|3537,3543
follow|3544,3550
the|3551,3554
recommendations|3555,3570
below|3571,3576
to|3577,3579
ensure|3580,3586
a|3587,3588
speedy|3589,3595
and|3596,3599
<EOL>|3600,3601
uneventful|3601,3611
recovery|3612,3620
.|3620,3621
<EOL>|3622,3623
<EOL>|3624,3625
ACTIVITY|3625,3633
:|3633,3634
<EOL>|3634,3635
-|3635,3636
Do|3637,3639
not|3640,3643
drive|3644,3649
until|3650,3655
you|3656,3659
have|3660,3664
stopped|3665,3672
taking|3673,3679
pain|3680,3684
medicine|3685,3693
and|3694,3697
<EOL>|3698,3699
feel|3699,3703
you|3704,3707
could|3708,3713
respond|3714,3721
in|3722,3724
an|3725,3727
emergency|3728,3737
.|3737,3738
<EOL>|3738,3739
-|3739,3740
You|3741,3744
may|3745,3748
climb|3749,3754
stairs|3755,3761
.|3761,3762
<EOL>|3763,3764
-|3764,3765
You|3766,3769
may|3770,3773
go|3774,3776
outside|3777,3784
,|3784,3785
but|3786,3789
avoid|3790,3795
traveling|3796,3805
long|3806,3810
distances|3811,3820
until|3821,3826
<EOL>|3827,3828
you|3828,3831
see|3832,3835
your|3836,3840
surgeon|3841,3848
at|3849,3851
your|3852,3856
next|3857,3861
visit|3862,3867
.|3867,3868
<EOL>|3868,3869
-|3869,3870
Do|3871,3873
n't|3873,3876
lift|3877,3881
more|3882,3886
than|3887,3891
10|3892,3894
lbs|3895,3898
for|3899,3902
6|3903,3904
weeks|3905,3910
.|3910,3911
(|3912,3913
This|3913,3917
is|3918,3920
about|3921,3926
the|3927,3930
<EOL>|3931,3932
weight|3932,3938
of|3939,3941
a|3942,3943
briefcase|3944,3953
or|3954,3956
a|3957,3958
bag|3959,3962
of|3963,3965
groceries|3966,3975
.|3975,3976
)|3976,3977
This|3978,3982
applies|3983,3990
to|3991,3993
<EOL>|3994,3995
lifting|3995,4002
children|4003,4011
,|4011,4012
but|4013,4016
they|4017,4021
may|4022,4025
sit|4026,4029
on|4030,4032
your|4033,4037
lap|4038,4041
.|4041,4042
<EOL>|4042,4043
-|4043,4044
You|4045,4048
may|4049,4052
start|4053,4058
some|4059,4063
light|4064,4069
exercise|4070,4078
when|4079,4083
you|4084,4087
feel|4088,4092
comfortable|4093,4104
.|4104,4105
<EOL>|4105,4106
-|4106,4107
You|4108,4111
will|4112,4116
need|4117,4121
to|4122,4124
stay|4125,4129
out|4130,4133
of|4134,4136
bathtubs|4137,4145
or|4146,4148
swimming|4149,4157
pools|4158,4163
for|4164,4167
a|4168,4169
<EOL>|4170,4171
time|4171,4175
while|4176,4181
your|4182,4186
incision|4187,4195
is|4196,4198
healing|4199,4206
.|4206,4207
Ask|4208,4211
your|4212,4216
doctor|4217,4223
when|4224,4228
you|4229,4232
<EOL>|4233,4234
can|4234,4237
resume|4238,4244
tub|4245,4248
baths|4249,4254
or|4255,4257
swimming|4258,4266
.|4266,4267
<EOL>|4267,4268
-|4268,4269
Heavy|4270,4275
exercise|4276,4284
may|4285,4288
be|4289,4291
started|4292,4299
after|4300,4305
6|4306,4307
weeks|4308,4313
,|4313,4314
but|4315,4318
use|4319,4322
common|4323,4329
<EOL>|4330,4331
sense|4331,4336
and|4337,4340
go|4341,4343
slowly|4344,4350
at|4351,4353
first|4354,4359
.|4359,4360
<EOL>|4360,4361
-|4361,4362
You|4363,4366
may|4367,4370
resume|4371,4377
sexual|4378,4384
activity|4385,4393
unless|4394,4400
your|4401,4405
doctor|4406,4412
has|4413,4416
told|4417,4421
you|4422,4425
<EOL>|4426,4427
otherwise|4427,4436
.|4436,4437
<EOL>|4437,4438
<EOL>|4439,4440
HOW|4440,4443
YOU|4444,4447
MAY|4448,4451
FEEL|4452,4456
:|4456,4457
<EOL>|4458,4459
-|4459,4460
You|4461,4464
may|4465,4468
feel|4469,4473
weak|4474,4478
or|4479,4481
"|4482,4483
washed|4483,4489
out|4490,4493
"|4493,4494
for|4495,4498
6|4499,4500
weeks|4501,4506
.|4506,4507
You|4508,4511
might|4512,4517
want|4518,4522
<EOL>|4523,4524
to|4524,4526
nap|4527,4530
often|4531,4536
.|4536,4537
Simple|4538,4544
tasks|4545,4550
may|4551,4554
exhaust|4555,4562
you|4563,4566
.|4566,4567
<EOL>|4567,4568
-|4568,4569
You|4570,4573
may|4574,4577
have|4578,4582
a|4583,4584
sore|4585,4589
throat|4590,4596
because|4597,4604
of|4605,4607
a|4608,4609
tube|4610,4614
that|4615,4619
was|4620,4623
in|4624,4626
your|4627,4631
<EOL>|4632,4633
throat|4633,4639
during|4640,4646
surgery|4647,4654
.|4654,4655
<EOL>|4655,4656
-|4656,4657
You|4658,4661
might|4662,4667
have|4668,4672
trouble|4673,4680
concentrating|4681,4694
or|4695,4697
difficulty|4698,4708
sleeping|4709,4717
.|4717,4718
<EOL>|4719,4720
You|4720,4723
might|4724,4729
feel|4730,4734
somewhat|4735,4743
depressed|4744,4753
.|4753,4754
<EOL>|4754,4755
-|4755,4756
You|4757,4760
could|4761,4766
have|4767,4771
a|4772,4773
poor|4774,4778
appetite|4779,4787
for|4788,4791
a|4792,4793
while|4794,4799
.|4799,4800
Food|4801,4805
may|4806,4809
seem|4810,4814
<EOL>|4815,4816
unappealing|4816,4827
.|4827,4828
<EOL>|4828,4829
-|4829,4830
All|4831,4834
of|4835,4837
these|4838,4843
feelings|4844,4852
and|4853,4856
reactions|4857,4866
are|4867,4870
normal|4871,4877
and|4878,4881
should|4882,4888
go|4889,4891
<EOL>|4892,4893
away|4893,4897
in|4898,4900
a|4901,4902
short|4903,4908
time|4909,4913
.|4913,4914
If|4915,4917
they|4918,4922
do|4923,4925
not|4926,4929
,|4929,4930
tell|4931,4935
your|4936,4940
surgeon|4941,4948
.|4948,4949
<EOL>|4949,4950
<EOL>|4951,4952
YOUR|4952,4956
INCISION|4957,4965
:|4965,4966
<EOL>|4966,4967
-|4967,4968
Your|4969,4973
incision|4974,4982
may|4983,4986
be|4987,4989
slightly|4990,4998
red|4999,5002
around|5003,5009
the|5010,5013
edges|5014,5019
.|5019,5020
This|5021,5025
is|5026,5028
<EOL>|5029,5030
normal|5030,5036
.|5036,5037
<EOL>|5037,5038
-|5038,5039
If|5040,5042
you|5043,5046
have|5047,5051
steri|5052,5057
strips|5058,5064
,|5064,5065
do|5066,5068
not|5069,5072
remove|5073,5079
them|5080,5084
for|5085,5088
2|5089,5090
weeks|5091,5096
.|5096,5097
<EOL>|5098,5099
(|5099,5100
These|5100,5105
are|5106,5109
the|5110,5113
thin|5114,5118
paper|5119,5124
strips|5125,5131
that|5132,5136
are|5137,5140
on|5141,5143
your|5144,5148
incision|5149,5157
.|5157,5158
)|5158,5159
But|5160,5163
<EOL>|5164,5165
if|5165,5167
they|5168,5172
fall|5173,5177
off|5178,5181
before|5182,5188
that|5189,5193
that|5194,5198
's|5198,5200
okay|5201,5205
)|5205,5206
.|5206,5207
<EOL>|5207,5208
-|5208,5209
You|5210,5213
may|5214,5217
gently|5218,5224
wash|5225,5229
away|5230,5234
dried|5235,5240
material|5241,5249
around|5250,5256
your|5257,5261
incision|5262,5270
.|5270,5271
<EOL>|5271,5272
-|5272,5273
It|5274,5276
is|5277,5279
normal|5280,5286
to|5287,5289
feel|5290,5294
a|5295,5296
firm|5297,5301
ridge|5302,5307
along|5308,5313
the|5314,5317
incision|5318,5326
.|5326,5327
This|5328,5332
<EOL>|5333,5334
will|5334,5338
go|5339,5341
away|5342,5346
.|5346,5347
<EOL>|5347,5348
-|5348,5349
Avoid|5350,5355
direct|5356,5362
sun|5363,5366
exposure|5367,5375
to|5376,5378
the|5379,5382
incision|5383,5391
area|5392,5396
.|5396,5397
<EOL>|5397,5398
-|5398,5399
Do|5400,5402
not|5403,5406
use|5407,5410
any|5411,5414
ointments|5415,5424
on|5425,5427
the|5428,5431
incision|5432,5440
unless|5441,5447
you|5448,5451
were|5452,5456
told|5457,5461
<EOL>|5462,5463
otherwise|5463,5472
.|5472,5473
<EOL>|5473,5474
-|5474,5475
You|5476,5479
may|5480,5483
see|5484,5487
a|5488,5489
small|5490,5495
amount|5496,5502
of|5503,5505
clear|5506,5511
or|5512,5514
light|5515,5520
red|5521,5524
fluid|5525,5530
<EOL>|5531,5532
staining|5532,5540
your|5541,5545
dressing|5546,5554
or|5555,5557
clothes|5558,5565
.|5565,5566
If|5567,5569
the|5570,5573
staining|5574,5582
is|5583,5585
severe|5586,5592
,|5592,5593
<EOL>|5594,5595
please|5595,5601
call|5602,5606
your|5607,5611
surgeon|5612,5619
.|5619,5620
<EOL>|5620,5621
-|5621,5622
You|5623,5626
may|5627,5630
shower|5631,5637
.|5637,5638
As|5639,5641
noted|5642,5647
above|5648,5653
,|5653,5654
ask|5655,5658
your|5659,5663
doctor|5664,5670
when|5671,5675
you|5676,5679
may|5680,5683
<EOL>|5684,5685
resume|5685,5691
tub|5692,5695
baths|5696,5701
or|5702,5704
swimming|5705,5713
.|5713,5714
<EOL>|5714,5715
-|5715,5716
Over|5717,5721
the|5722,5725
next|5726,5730
_|5731,5732
_|5732,5733
_|5733,5734
months|5735,5741
,|5741,5742
your|5743,5747
incision|5748,5756
will|5757,5761
fade|5762,5766
and|5767,5770
become|5771,5777
<EOL>|5778,5779
less|5779,5783
prominent|5784,5793
.|5793,5794
<EOL>|5794,5795
<EOL>|5796,5797
YOUR|5797,5801
BOWELS|5802,5808
:|5808,5809
<EOL>|5809,5810
-|5810,5811
Constipation|5812,5824
is|5825,5827
a|5828,5829
common|5830,5836
side|5837,5841
effect|5842,5848
of|5849,5851
medicine|5852,5860
such|5861,5865
as|5866,5868
<EOL>|5869,5870
Percocet|5870,5878
or|5879,5881
codeine|5882,5889
.|5889,5890
If|5891,5893
needed|5894,5900
,|5900,5901
you|5902,5905
may|5906,5909
take|5910,5914
a|5915,5916
stool|5917,5922
softener|5923,5931
<EOL>|5932,5933
(|5933,5934
such|5934,5938
as|5939,5941
Colace|5942,5948
,|5948,5949
one|5950,5953
capsule|5954,5961
)|5961,5962
or|5963,5965
gentle|5966,5972
laxative|5973,5981
(|5982,5983
such|5983,5987
as|5988,5990
milk|5991,5995
<EOL>|5996,5997
of|5997,5999
magnesia|6000,6008
,|6008,6009
1|6010,6011
tbs|6012,6015
)|6015,6016
twice|6017,6022
a|6023,6024
day|6025,6028
.|6028,6029
You|6030,6033
can|6034,6037
get|6038,6041
both|6042,6046
of|6047,6049
these|6050,6055
<EOL>|6056,6057
medicines|6057,6066
without|6067,6074
a|6075,6076
prescription|6077,6089
.|6089,6090
<EOL>|6090,6091
-|6091,6092
If|6093,6095
you|6096,6099
go|6100,6102
48|6103,6105
hours|6106,6111
without|6112,6119
a|6120,6121
bowel|6122,6127
movement|6128,6136
,|6136,6137
or|6138,6140
have|6141,6145
pain|6146,6150
<EOL>|6151,6152
moving|6152,6158
your|6159,6163
bowels|6164,6170
,|6170,6171
call|6172,6176
your|6177,6181
surgeon|6182,6189
.|6189,6190
<EOL>|6190,6191
-|6191,6192
After|6193,6198
some|6199,6203
operations|6204,6214
,|6214,6215
diarrhea|6216,6224
can|6225,6228
occur|6229,6234
.|6234,6235
If|6236,6238
you|6239,6242
get|6243,6246
<EOL>|6247,6248
diarrhea|6248,6256
,|6256,6257
do|6258,6260
n't|6260,6263
take|6264,6268
anti-diarrhea|6269,6282
medicines|6283,6292
.|6292,6293
Drink|6294,6299
plenty|6300,6306
of|6307,6309
<EOL>|6310,6311
fluids|6311,6317
and|6318,6321
see|6322,6325
if|6326,6328
it|6329,6331
goes|6332,6336
away|6337,6341
.|6341,6342
If|6343,6345
it|6346,6348
does|6349,6353
not|6354,6357
go|6358,6360
away|6361,6365
,|6365,6366
or|6367,6369
is|6370,6372
<EOL>|6373,6374
severe|6374,6380
and|6381,6384
you|6385,6388
feel|6389,6393
ill|6394,6397
,|6397,6398
please|6399,6405
call|6406,6410
your|6411,6415
surgeon|6416,6423
.|6423,6424
<EOL>|6424,6425
<EOL>|6426,6427
PAIN|6427,6431
MANAGEMENT|6432,6442
:|6442,6443
<EOL>|6443,6444
-|6444,6445
It|6446,6448
is|6449,6451
normal|6452,6458
to|6459,6461
feel|6462,6466
some|6467,6471
discomfort|6472,6482
/|6482,6483
pain|6483,6487
following|6488,6497
abdominal|6498,6507
<EOL>|6508,6509
surgery|6509,6516
.|6516,6517
This|6518,6522
pain|6523,6527
is|6528,6530
often|6531,6536
described|6537,6546
as|6547,6549
"|6550,6551
soreness|6551,6559
"|6559,6560
.|6560,6561
<EOL>|6562,6563
-|6563,6564
Your|6565,6569
pain|6570,6574
should|6575,6581
get|6582,6585
better|6586,6592
day|6593,6596
by|6597,6599
day|6600,6603
.|6603,6604
If|6605,6607
you|6608,6611
find|6612,6616
the|6617,6620
pain|6621,6625
<EOL>|6626,6627
is|6627,6629
getting|6630,6637
worse|6638,6643
instead|6644,6651
of|6652,6654
better|6655,6661
,|6661,6662
please|6663,6669
contact|6670,6677
your|6678,6682
surgeon|6683,6690
.|6690,6691
<EOL>|6691,6692
-|6692,6693
You|6693,6696
will|6697,6701
receive|6702,6709
a|6710,6711
prescription|6712,6724
from|6725,6729
your|6730,6734
surgeon|6735,6742
for|6743,6746
pain|6747,6751
<EOL>|6752,6753
medicine|6753,6761
to|6762,6764
take|6765,6769
by|6770,6772
mouth|6773,6778
.|6778,6779
It|6780,6782
is|6783,6785
important|6786,6795
to|6796,6798
take|6799,6803
this|6804,6808
medicine|6809,6817
<EOL>|6818,6819
as|6819,6821
directed|6822,6830
.|6830,6831
<EOL>|6832,6833
-|6833,6834
Do|6835,6837
not|6838,6841
take|6842,6846
it|6847,6849
more|6850,6854
frequently|6855,6865
than|6866,6870
prescribed|6871,6881
.|6881,6882
Do|6883,6885
not|6886,6889
take|6890,6894
<EOL>|6895,6896
more|6896,6900
medicine|6901,6909
at|6910,6912
one|6913,6916
time|6917,6921
than|6922,6926
prescribed|6927,6937
.|6937,6938
<EOL>|6938,6939
-|6939,6940
Your|6941,6945
pain|6946,6950
medicine|6951,6959
will|6960,6964
work|6965,6969
better|6970,6976
if|6977,6979
you|6980,6983
take|6984,6988
it|6989,6991
before|6992,6998
your|6999,7003
<EOL>|7004,7005
pain|7005,7009
gets|7010,7014
too|7015,7018
severe|7019,7025
.|7025,7026
<EOL>|7027,7028
-|7028,7029
If|7030,7032
you|7033,7036
are|7037,7040
experiencing|7041,7053
no|7054,7056
pain|7057,7061
,|7061,7062
it|7063,7065
is|7066,7068
okay|7069,7073
to|7074,7076
skip|7077,7081
a|7082,7083
dose|7084,7088
of|7089,7091
<EOL>|7092,7093
pain|7093,7097
medicine|7098,7106
.|7106,7107
<EOL>|7107,7108
If|7108,7110
you|7111,7114
experience|7115,7125
any|7126,7129
of|7130,7132
the|7133,7136
folloiwng|7137,7146
,|7146,7147
please|7148,7154
contact|7155,7162
your|7163,7167
<EOL>|7168,7169
surgeon|7169,7176
:|7176,7177
<EOL>|7177,7178
-|7178,7179
sharp|7180,7185
pain|7186,7190
or|7191,7193
any|7194,7197
severe|7198,7204
pain|7205,7209
that|7210,7214
lasts|7215,7220
several|7221,7228
hours|7229,7234
<EOL>|7234,7235
-|7235,7236
pain|7237,7241
that|7242,7246
is|7247,7249
getting|7250,7257
worse|7258,7263
over|7264,7268
time|7269,7273
<EOL>|7273,7274
-|7274,7275
pain|7276,7280
accompanied|7281,7292
by|7293,7295
fever|7296,7301
of|7302,7304
more|7305,7309
than|7310,7314
101|7315,7318
<EOL>|7318,7319
-|7319,7320
a|7321,7322
drastic|7323,7330
change|7331,7337
in|7338,7340
nature|7341,7347
or|7348,7350
quality|7351,7358
of|7359,7361
your|7362,7366
pain|7367,7371
<EOL>|7371,7372
<EOL>|7373,7374
MEDICATIONS|7374,7385
:|7385,7386
<EOL>|7386,7387
-|7387,7388
Take|7389,7393
all|7394,7397
the|7398,7401
medicines|7402,7411
you|7412,7415
were|7416,7420
on|7421,7423
before|7424,7430
the|7431,7434
operation|7435,7444
just|7445,7449
<EOL>|7450,7451
as|7451,7453
you|7454,7457
did|7458,7461
before|7462,7468
,|7468,7469
unless|7470,7476
you|7477,7480
have|7481,7485
been|7486,7490
told|7491,7495
differently|7496,7507
.|7507,7508
<EOL>|7508,7509
-|7509,7510
If|7511,7513
you|7514,7517
have|7518,7522
any|7523,7526
questions|7527,7536
about|7537,7542
what|7543,7547
medicine|7548,7556
to|7557,7559
take|7560,7564
or|7565,7567
not|7568,7571
<EOL>|7572,7573
to|7573,7575
take|7576,7580
,|7580,7581
please|7582,7588
call|7589,7593
your|7594,7598
surgeon|7599,7606
.|7606,7607
<EOL>|7607,7608
<EOL>|7608,7609
<EOL>|7610,7611
Followup|7611,7619
Instructions|7620,7632
:|7632,7633
<EOL>|7633,7634
_|7634,7635
_|7635,7636
_|7636,7637
<EOL>|7637,7638

