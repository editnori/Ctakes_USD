 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|46,55|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|46,55|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|46,60|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|80,89|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|80,89|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|80,94|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|136,139|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|147,154|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|147,154|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|156,164|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|SIMPLE_SEGMENT|167,176|false|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|167,176|false|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|167,176|false|false|false|C0020517|Hypersensitivity|Allergies
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|179,189|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|179,189|false|false|false|C0065374|lisinopril|lisinopril
Event|Event|SIMPLE_SEGMENT|179,189|false|false|false|||lisinopril
Event|Event|SIMPLE_SEGMENT|192,201|false|false|false|||Attending
Finding|Functional Concept|SIMPLE_SEGMENT|192,201|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|SIMPLE_SEGMENT|210,225|false|false|false|C0277786|Chief complaint (finding)|Chief Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|216,225|false|false|false|C3864418||Complaint
Event|Event|SIMPLE_SEGMENT|216,225|false|false|false|||Complaint
Finding|Finding|SIMPLE_SEGMENT|216,225|false|false|false|C5441521|Complaint (finding)|Complaint
Anatomy|Body Location or Region|SIMPLE_SEGMENT|227,232|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|227,232|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|227,237|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|227,237|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|233,237|false|true|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|233,237|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|233,237|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|233,237|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Classification|SIMPLE_SEGMENT|240,245|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|SIMPLE_SEGMENT|246,254|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|246,254|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|258,276|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|267,276|false|false|false|C0945766||Procedure
Event|Event|SIMPLE_SEGMENT|267,276|false|false|false|||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|267,276|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|267,276|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|267,276|false|false|false|C0184661|Interventional procedure|Procedure
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|278,285|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|278,285|false|false|false|C1314974|Cardiac attachment|cardiac
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|278,301|false|false|false|C0261588|Cardiac catheterisation as the cause of abnormal reaction of the patient, or of later complication, without mention of misadventure at the time of the procedure|cardiac catheterization
Finding|Intellectual Product|SIMPLE_SEGMENT|278,301|false|false|false|C1547981|Diagnostic Service Section ID - Cardiac Catheterization|cardiac catheterization
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|278,301|false|false|false|C0018795;C1548828|Cardiac Catheterization Procedures;Consent Type - Cardiac Catheterization|cardiac catheterization
Procedure|Health Care Activity|SIMPLE_SEGMENT|278,301|false|false|false|C0018795;C1548828|Cardiac Catheterization Procedures;Consent Type - Cardiac Catheterization|cardiac catheterization
Event|Event|SIMPLE_SEGMENT|286,301|false|false|false|||catheterization
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|286,301|false|false|false|C0007430|Catheterization|catheterization
Event|Event|SIMPLE_SEGMENT|305,312|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|305,312|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|305,312|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|305,312|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|305,315|false|false|false|C0262926|Medical History|History of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|305,331|false|false|false|C0488508||History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|305,331|false|false|false|C0262512|History of present illness (finding)|History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|316,323|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Idea or Concept|SIMPLE_SEGMENT|316,323|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Finding|SIMPLE_SEGMENT|316,331|false|false|false|C4264312|Present illness|Present Illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|324,331|false|false|false|C0221423|Illness (finding)|Illness
Event|Event|SIMPLE_SEGMENT|335,336|false|false|false|||_
Event|Event|SIMPLE_SEGMENT|340,343|false|false|false|||PMH
Finding|Finding|SIMPLE_SEGMENT|340,343|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|PMH
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|347,350|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|347,350|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|347,350|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|347,350|false|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|347,350|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|347,350|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|347,350|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|347,350|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|355,358|false|false|false|C2713669|SERPINA5 protein, human|PCI
Drug|Biologically Active Substance|SIMPLE_SEGMENT|355,358|false|false|false|C2713669|SERPINA5 protein, human|PCI
Event|Event|SIMPLE_SEGMENT|355,358|false|false|false|||PCI
Finding|Gene or Genome|SIMPLE_SEGMENT|355,358|false|false|false|C1418370;C1705930;C4049621|Peritoneal Cancer Index;SERPINA5 gene;SERPINA5 wt Allele|PCI
Finding|Intellectual Product|SIMPLE_SEGMENT|355,358|false|false|false|C1418370;C1705930;C4049621|Peritoneal Cancer Index;SERPINA5 gene;SERPINA5 wt Allele|PCI
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|355,358|false|false|false|C1514496;C1532338;C4724254|Percutaneous Coronary Intervention;Prophylactic Cranial Irradiation;photochemical internalization|PCI
Event|Event|SIMPLE_SEGMENT|359,361|false|false|false|||x3
Finding|Molecular Function|SIMPLE_SEGMENT|371,375|false|false|false|C1150186|matrix metalloproteinase 7 activity|pump
Event|Event|SIMPLE_SEGMENT|376,380|false|false|false|||CABG
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|376,380|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|396,399|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|396,399|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|SIMPLE_SEGMENT|396,399|false|false|false|||LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|396,399|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Event|Event|SIMPLE_SEGMENT|408,412|false|false|false|||diag
Finding|Functional Concept|SIMPLE_SEGMENT|408,412|false|false|false|C1704338|diagnosis aspects|diag
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|408,412|false|false|false|C0011900|Diagnosis|diag
Event|Event|SIMPLE_SEGMENT|419,423|false|false|false|||type
Finding|Gene or Genome|SIMPLE_SEGMENT|419,423|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Finding|Intellectual Product|SIMPLE_SEGMENT|419,423|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Finding|Classification|SIMPLE_SEGMENT|419,425|false|false|false|C0441730|Type 2|type 2
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|432,439|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|SIMPLE_SEGMENT|432,439|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|432,439|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|SIMPLE_SEGMENT|432,439|false|false|false|||insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|432,439|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|432,439|false|false|false|C0202098|Insulin measurement|insulin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|441,444|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|SIMPLE_SEGMENT|441,444|false|false|false|||HTN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|447,461|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|hyperlipidemia
Event|Event|SIMPLE_SEGMENT|447,461|false|false|false|||hyperlipidemia
Finding|Finding|SIMPLE_SEGMENT|447,461|false|false|false|C0428465|Serum lipids high (finding)|hyperlipidemia
Event|Event|SIMPLE_SEGMENT|462,470|false|false|false|||presents
Finding|Idea or Concept|SIMPLE_SEGMENT|480,483|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|480,483|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|484,491|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|484,491|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|484,491|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|484,491|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|484,494|false|false|false|C0262926|Medical History|history of
Event|Event|SIMPLE_SEGMENT|499,504|false|false|false|||sharp
Finding|Finding|SIMPLE_SEGMENT|499,504|false|false|false|C1444775;C1539835;C3890003|SPEN gene;SPEN wt Allele;Sharp sensation quality|sharp
Finding|Gene or Genome|SIMPLE_SEGMENT|499,504|false|false|false|C1444775;C1539835;C3890003|SPEN gene;SPEN wt Allele;Sharp sensation quality|sharp
Finding|Functional Concept|SIMPLE_SEGMENT|507,511|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|SIMPLE_SEGMENT|518,523|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|518,523|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|518,528|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|518,528|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|524,528|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|524,528|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|524,528|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|524,528|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|533,536|false|false|false|||SOB
Finding|Sign or Symptom|SIMPLE_SEGMENT|533,536|false|false|false|C0013404|Dyspnea|SOB
Event|Event|SIMPLE_SEGMENT|542,551|false|false|false|||describes
Anatomy|Body Location or Region|SIMPLE_SEGMENT|556,561|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|556,561|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|556,566|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|556,566|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|562,566|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|562,566|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|562,566|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|562,566|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|572,580|false|false|false|C0418416|Pinched|pinching
Event|Event|SIMPLE_SEGMENT|572,580|false|false|false|||pinching
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|605,609|false|false|false|C0262950;C1442209|Skeletal bone;XXX bone|bone
Finding|Body Substance|SIMPLE_SEGMENT|605,609|false|false|false|C1546560;C1550616|Specimen Type - Bone|bone
Finding|Intellectual Product|SIMPLE_SEGMENT|605,609|false|false|false|C1546560;C1550616|Specimen Type - Bone|bone
Event|Event|SIMPLE_SEGMENT|616,624|false|false|false|||endorses
Event|Event|SIMPLE_SEGMENT|630,638|false|false|false|||episodes
Attribute|Clinical Attribute|SIMPLE_SEGMENT|642,646|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|642,646|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|642,646|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|642,646|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Idea or Concept|SIMPLE_SEGMENT|647,650|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|647,650|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|652,658|false|false|false|||always
Finding|Finding|SIMPLE_SEGMENT|652,658|false|false|false|C1549493;C3812891|All of the Time;Always - AcknowledgementCondition|always
Finding|Idea or Concept|SIMPLE_SEGMENT|652,658|false|false|false|C1549493;C3812891|All of the Time;Always - AcknowledgementCondition|always
Finding|Functional Concept|SIMPLE_SEGMENT|659,666|false|false|false|C0443144|At rest (qualifier value)|at rest
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|662,666|false|false|false|C1742913|REST protein, human|rest
Drug|Biologically Active Substance|SIMPLE_SEGMENT|662,666|false|false|false|C1742913|REST protein, human|rest
Event|Event|SIMPLE_SEGMENT|662,666|false|false|false|||rest
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|662,666|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Gene or Genome|SIMPLE_SEGMENT|662,666|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Molecular Function|SIMPLE_SEGMENT|662,666|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Event|Event|SIMPLE_SEGMENT|672,680|false|false|false|||episodes
Attribute|Clinical Attribute|SIMPLE_SEGMENT|684,688|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|684,688|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|684,688|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|684,688|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|709,718|false|false|false|C0886384|5 minutes Office visit|5 minutes
Event|Event|SIMPLE_SEGMENT|711,718|false|false|false|||minutes
Event|Event|SIMPLE_SEGMENT|727,735|false|false|false|||relieved
Drug|Organic Chemical|SIMPLE_SEGMENT|739,752|false|false|false|C0017887|nitroglycerin|nitroglycerin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|739,752|false|false|false|C0017887|nitroglycerin|nitroglycerin
Event|Event|SIMPLE_SEGMENT|739,752|false|false|false|||nitroglycerin
Attribute|Clinical Attribute|SIMPLE_SEGMENT|759,763|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|759,763|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|759,763|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|759,763|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|771,779|false|false|false|||worsened
Event|Event|SIMPLE_SEGMENT|783,791|false|false|false|||exertion
Finding|Organism Function|SIMPLE_SEGMENT|783,791|true|true|false|C0015264|Exertion|exertion
Event|Event|SIMPLE_SEGMENT|795,801|false|false|false|||eating
Finding|Organism Function|SIMPLE_SEGMENT|795,801|false|false|false|C0013470|Eating|eating
Event|Event|SIMPLE_SEGMENT|807,816|false|false|false|||described
Event|Event|SIMPLE_SEGMENT|822,830|false|false|false|||symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|822,830|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|822,830|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|838,841|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|838,841|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|838,841|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|838,841|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|SIMPLE_SEGMENT|838,841|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|838,841|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|SIMPLE_SEGMENT|838,841|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|838,841|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|SIMPLE_SEGMENT|838,841|false|false|false|||PCP
Finding|Gene or Genome|SIMPLE_SEGMENT|838,841|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|SIMPLE_SEGMENT|838,841|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Event|SIMPLE_SEGMENT|851,856|false|false|false|||phone
Finding|Idea or Concept|SIMPLE_SEGMENT|851,856|false|false|false|C1515258;C1547567;C1548343;C1576870|Authorization Mode - Phone;MDFAttributeType - Phone;Telephone Number;Visit User Code - Phone|phone
Finding|Intellectual Product|SIMPLE_SEGMENT|851,856|false|false|false|C1515258;C1547567;C1548343;C1576870|Authorization Mode - Phone;MDFAttributeType - Phone;Telephone Number;Visit User Code - Phone|phone
Event|Event|SIMPLE_SEGMENT|862,866|false|false|false|||told
Event|Event|SIMPLE_SEGMENT|874,878|false|false|false|||come
Event|Event|SIMPLE_SEGMENT|887,889|false|false|false|||ED
Event|Event|SIMPLE_SEGMENT|905,909|false|false|false|||feel
Event|Event|SIMPLE_SEGMENT|910,917|false|false|false|||similar
Event|Event|SIMPLE_SEGMENT|951,959|false|false|false|||endorsed
Event|Event|SIMPLE_SEGMENT|960,968|false|false|false|||vomiting
Finding|Sign or Symptom|SIMPLE_SEGMENT|960,968|false|false|false|C0042963|Vomiting|vomiting
Event|Event|SIMPLE_SEGMENT|985,991|false|false|false|||denies
Event|Event|SIMPLE_SEGMENT|996,1007|false|false|false|||diaphoresis
Finding|Finding|SIMPLE_SEGMENT|996,1007|true|false|false|C0700590|Increased sweating|diaphoresis
Event|Event|SIMPLE_SEGMENT|1019,1027|false|false|false|||endorses
Drug|Organic Chemical|SIMPLE_SEGMENT|1030,1035|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1030,1035|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|SIMPLE_SEGMENT|1030,1035|false|false|false|||cough
Finding|Sign or Symptom|SIMPLE_SEGMENT|1030,1035|false|false|false|C0010200|Coughing|cough
Finding|Body Substance|SIMPLE_SEGMENT|1043,1050|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1043,1050|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1043,1050|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|SIMPLE_SEGMENT|1043,1054|false|false|false|C0332310|Has patient|patient has
Event|Event|SIMPLE_SEGMENT|1055,1064|false|false|false|||developed
Finding|Sign or Symptom|SIMPLE_SEGMENT|1065,1094|false|false|false|C0574066|Increasing breathlessness|increased shortness of breath
Event|Event|SIMPLE_SEGMENT|1075,1084|false|false|false|||shortness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1075,1094|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|SIMPLE_SEGMENT|1075,1094|false|false|false|C0013404|Dyspnea|shortness of breath
Event|Event|SIMPLE_SEGMENT|1088,1094|false|false|false|||breath
Finding|Body Substance|SIMPLE_SEGMENT|1088,1094|false|false|false|C0225386|Breath|breath
Event|Event|SIMPLE_SEGMENT|1140,1149|false|false|false|||orthopnea
Finding|Finding|SIMPLE_SEGMENT|1140,1149|false|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|1140,1149|false|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Event|Event|SIMPLE_SEGMENT|1179,1185|false|false|false|||denies
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1186,1189|false|false|false|C1956415|Paroxysmal nocturnal dyspnea|PND
Event|Event|SIMPLE_SEGMENT|1186,1189|false|false|false|||PND
Finding|Gene or Genome|SIMPLE_SEGMENT|1186,1189|false|false|false|C1417807;C4552608|NPPA gene;NPPA wt Allele|PND
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1194,1199|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|1194,1199|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1194,1209|false|false|false|C0023216|Lower Extremity|lower extremity
Finding|Pathologic Function|SIMPLE_SEGMENT|1194,1215|true|false|false|C0239340|Edema of lower extremity|lower extremity edema
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1200,1209|false|false|false|C0015385|Limb structure|extremity
Finding|Pathologic Function|SIMPLE_SEGMENT|1200,1215|false|false|false|C0085649|Peripheral edema|extremity edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1210,1215|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|1210,1215|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|1210,1215|false|false|false|C0013604|Edema|edema
Event|Event|SIMPLE_SEGMENT|1220,1224|false|false|false|||exam
Finding|Functional Concept|SIMPLE_SEGMENT|1220,1224|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|1220,1224|false|false|false|C0582103|Medical Examination|exam
Event|Event|SIMPLE_SEGMENT|1244,1255|false|false|false|||tachycardic
Event|Event|SIMPLE_SEGMENT|1270,1276|false|false|false|||rhythm
Finding|Finding|SIMPLE_SEGMENT|1270,1276|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|SIMPLE_SEGMENT|1270,1276|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1278,1283|false|false|false|C0024109|Lung|Lungs
Drug|Organic Chemical|SIMPLE_SEGMENT|1289,1293|false|false|false|C0951233|cetrimonium bromide|CTAB
Event|Event|SIMPLE_SEGMENT|1289,1293|false|false|false|||CTAB
Finding|Functional Concept|SIMPLE_SEGMENT|1304,1309|false|false|false|C1883002|Sequence Chromatogram|trace
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1310,1315|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|1310,1315|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|1310,1315|false|false|false|C0013604|Edema|edema
Finding|Functional Concept|SIMPLE_SEGMENT|1323,1327|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1323,1343|false|false|false|C0230416|Left lower extremity|left lower extremity
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1328,1333|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|1328,1333|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1328,1343|false|false|false|C0023216|Lower Extremity|lower extremity
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1334,1343|false|false|false|C0015385|Limb structure|extremity
Finding|Functional Concept|SIMPLE_SEGMENT|1358,1363|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1358,1367|false|false|false|C0230415;C0230442|Right lower extremity;Structure of right lower leg|right leg
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1364,1367|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Finding|Idea or Concept|SIMPLE_SEGMENT|1384,1391|false|false|false|C1555582|Initial (abbreviation)|initial
Event|Event|SIMPLE_SEGMENT|1392,1398|false|false|false|||vitals
Event|Event|SIMPLE_SEGMENT|1428,1432|false|false|false|||Labs
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1428,1432|false|false|false|C0587081|Laboratory test finding|Labs
Event|Event|SIMPLE_SEGMENT|1438,1445|false|false|false|||imaging
Finding|Finding|SIMPLE_SEGMENT|1438,1445|false|false|false|C0740845|Imaging problem|imaging
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1438,1445|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|imaging
Event|Event|SIMPLE_SEGMENT|1446,1457|false|false|false|||significant
Finding|Idea or Concept|SIMPLE_SEGMENT|1446,1457|false|false|false|C0750502|Significant|significant
Event|Event|SIMPLE_SEGMENT|1464,1467|false|false|false|||CXR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1464,1467|false|false|false|C0039985|Plain chest X-ray|CXR
Finding|Finding|SIMPLE_SEGMENT|1473,1476|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|1473,1476|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Finding|SIMPLE_SEGMENT|1477,1485|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|SIMPLE_SEGMENT|1477,1485|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Functional Concept|SIMPLE_SEGMENT|1486,1490|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Tissue|SIMPLE_SEGMENT|1491,1498|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1491,1498|false|false|false|C0032226|Pleural Diseases|pleural
Event|Event|SIMPLE_SEGMENT|1500,1508|false|false|false|||effusion
Finding|Body Substance|SIMPLE_SEGMENT|1500,1508|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|SIMPLE_SEGMENT|1500,1508|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|1500,1508|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Event|Event|SIMPLE_SEGMENT|1523,1534|false|false|false|||atelectasis
Finding|Pathologic Function|SIMPLE_SEGMENT|1523,1534|false|false|false|C0004144|Atelectasis|atelectasis
Finding|Functional Concept|SIMPLE_SEGMENT|1542,1546|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1542,1551|false|false|false|C0225730|Left lung|left lung
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1542,1556|false|false|false|C0225732|Structure of base of left lung|left lung base
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1547,1551|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1547,1551|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1547,1551|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|SIMPLE_SEGMENT|1547,1551|false|false|false|C0740941|Lung Problem|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1547,1556|false|false|false|C0225704|Basal segment of lung|lung base
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1552,1556|false|false|false|C2987514|Anatomical base|base
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|1552,1556|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Chemical Viewed Functionally|SIMPLE_SEGMENT|1552,1556|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|1552,1556|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Finding|Gene or Genome|SIMPLE_SEGMENT|1552,1556|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Finding|Idea or Concept|SIMPLE_SEGMENT|1552,1556|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Anatomy|Cell Component|SIMPLE_SEGMENT|1558,1561|false|false|false|C2263086|Nuclear cap binding complex location|CBC
Event|Event|SIMPLE_SEGMENT|1558,1561|false|false|false|||CBC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1558,1561|false|false|false|C0009555|Complete Blood Count|CBC
Finding|Finding|SIMPLE_SEGMENT|1563,1583|false|false|false|C0442816||within normal limits
Event|Event|SIMPLE_SEGMENT|1577,1583|false|false|false|||limits
Finding|Functional Concept|SIMPLE_SEGMENT|1577,1583|false|false|false|C0439801|Limited (extensiveness)|limits
Drug|Inorganic Chemical|SIMPLE_SEGMENT|1585,1597|false|false|false|C0013832;C3536863|Electrolyte [EPC];Electrolytes|electrolytes
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1585,1597|false|false|false|C0013832;C3536863|Electrolyte [EPC];Electrolytes|electrolytes
Event|Event|SIMPLE_SEGMENT|1585,1597|false|false|false|||electrolytes
Finding|Finding|SIMPLE_SEGMENT|1598,1618|false|false|false|C0442816||within normal limits
Event|Event|SIMPLE_SEGMENT|1612,1618|false|false|false|||limits
Finding|Functional Concept|SIMPLE_SEGMENT|1612,1618|false|false|false|C0439801|Limited (extensiveness)|limits
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1630,1638|false|false|false|C0041199|Troponin|troponin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1630,1638|false|false|false|C0041199|Troponin|troponin
Event|Event|SIMPLE_SEGMENT|1630,1638|false|false|false|||troponin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1630,1638|false|false|false|C0523952|Troponin measurement|troponin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1648,1655|false|false|false|C0060323|Fibrin fragment D|D-dimer
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1648,1655|false|false|false|C0060323|Fibrin fragment D|D-dimer
Drug|Chemical Viewed Structurally|SIMPLE_SEGMENT|1650,1655|false|false|false|C0596448|dimer|dimer
Event|Event|SIMPLE_SEGMENT|1650,1655|false|false|false|||dimer
Event|Event|SIMPLE_SEGMENT|1664,1666|false|false|false|||CT
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1674,1679|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|1674,1679|false|false|false|C0741025|Chest problem|chest
Event|Event|SIMPLE_SEGMENT|1702,1708|false|false|false|||showed
Event|Event|SIMPLE_SEGMENT|1715,1723|false|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|1715,1723|false|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|1715,1727|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence for
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1728,1737|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1728,1737|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|1728,1737|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|SIMPLE_SEGMENT|1728,1745|true|false|false|C0034065|Pulmonary Embolism|pulmonary embolus
Event|Event|SIMPLE_SEGMENT|1738,1745|false|false|false|||embolus
Finding|Finding|SIMPLE_SEGMENT|1738,1745|true|false|false|C1704212;C2046122|Embolus|embolus
Finding|Functional Concept|SIMPLE_SEGMENT|1758,1762|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Tissue|SIMPLE_SEGMENT|1763,1770|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1763,1770|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Body Substance|SIMPLE_SEGMENT|1763,1779|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Finding|Finding|SIMPLE_SEGMENT|1763,1779|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|1763,1779|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Event|Event|SIMPLE_SEGMENT|1771,1779|false|false|false|||effusion
Finding|Body Substance|SIMPLE_SEGMENT|1771,1779|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|SIMPLE_SEGMENT|1771,1779|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|1771,1779|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Event|Event|SIMPLE_SEGMENT|1794,1805|false|false|false|||atelectasis
Finding|Pathologic Function|SIMPLE_SEGMENT|1794,1805|false|false|false|C0004144|Atelectasis|atelectasis
Finding|Body Substance|SIMPLE_SEGMENT|1809,1816|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1809,1816|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1809,1816|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Organic Chemical|SIMPLE_SEGMENT|1823,1830|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1823,1830|false|false|false|C0004057|aspirin|aspirin
Drug|Organic Chemical|SIMPLE_SEGMENT|1844,1857|false|false|false|C0017887|nitroglycerin|nitroglycerin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1844,1857|false|false|false|C0017887|nitroglycerin|nitroglycerin
Event|Event|SIMPLE_SEGMENT|1844,1857|false|false|false|||nitroglycerin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1866,1873|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Organic Chemical|SIMPLE_SEGMENT|1866,1873|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1866,1873|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Event|Event|SIMPLE_SEGMENT|1866,1873|false|false|false|||heparin
Event|Event|SIMPLE_SEGMENT|1875,1880|false|false|false|||bolus
Finding|Body Substance|SIMPLE_SEGMENT|1875,1880|false|false|false|C1186706;C1550436|Bolus of ingested food;Response Modality - Bolus|bolus
Finding|Intellectual Product|SIMPLE_SEGMENT|1875,1880|false|false|false|C1186706;C1550436|Bolus of ingested food;Response Modality - Bolus|bolus
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1875,1880|false|false|false|C1511237|bolus infusion|bolus
Event|Event|SIMPLE_SEGMENT|1884,1890|false|false|false|||Vitals
Event|Event|SIMPLE_SEGMENT|1894,1902|false|false|false|||transfer
Finding|Functional Concept|SIMPLE_SEGMENT|1894,1902|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|SIMPLE_SEGMENT|1894,1902|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|SIMPLE_SEGMENT|1894,1902|false|false|false|C4706767|Transfer (immobility management)|transfer
Event|Activity|SIMPLE_SEGMENT|1939,1946|false|false|false|C1706079||arrival
Event|Event|SIMPLE_SEGMENT|1939,1946|false|false|false|||arrival
Finding|Functional Concept|SIMPLE_SEGMENT|1939,1946|false|false|false|C1555577|arrival - ActRelationshipType|arrival
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|1954,1959|false|false|false|C3714591|Floor (anatomic)|floor
Finding|Body Substance|SIMPLE_SEGMENT|1961,1968|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1961,1968|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1961,1968|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|1972,1977|false|false|false|||AAOx3
Event|Event|SIMPLE_SEGMENT|1983,1994|false|false|false|||comfortable
Finding|Finding|SIMPLE_SEGMENT|1983,1994|false|false|false|C5546696|Feeling comfortable|comfortable
Event|Event|SIMPLE_SEGMENT|2000,2006|false|false|false|||REVIEW
Finding|Idea or Concept|SIMPLE_SEGMENT|2000,2006|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|REVIEW
Finding|Intellectual Product|SIMPLE_SEGMENT|2000,2006|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|REVIEW
Finding|Functional Concept|SIMPLE_SEGMENT|2000,2009|false|false|false|C0699752|Review of|REVIEW OF
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2000,2017|false|false|false|C0488564;C0488565||REVIEW OF SYSTEMS
Procedure|Health Care Activity|SIMPLE_SEGMENT|2000,2017|false|false|false|C0489633|Review of systems (procedure)|REVIEW OF SYSTEMS
Event|Event|SIMPLE_SEGMENT|2010,2017|false|false|false|||SYSTEMS
Finding|Functional Concept|SIMPLE_SEGMENT|2010,2017|false|false|false|C0449913|System|SYSTEMS
Event|Event|SIMPLE_SEGMENT|2023,2029|false|false|false|||review
Finding|Idea or Concept|SIMPLE_SEGMENT|2023,2029|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Finding|Intellectual Product|SIMPLE_SEGMENT|2023,2029|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Finding|Functional Concept|SIMPLE_SEGMENT|2023,2032|false|false|false|C0699752|Review of|review of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2023,2040|false|false|false|C0488564;C0488565||review of systems
Procedure|Health Care Activity|SIMPLE_SEGMENT|2023,2040|false|false|false|C0489633|Review of systems (procedure)|review of systems
Event|Event|SIMPLE_SEGMENT|2033,2040|false|false|false|||systems
Finding|Functional Concept|SIMPLE_SEGMENT|2033,2040|false|false|false|C0449913|System|systems
Event|Event|SIMPLE_SEGMENT|2046,2052|false|false|false|||denies
Event|Event|SIMPLE_SEGMENT|2063,2070|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|2063,2070|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|2063,2070|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|2063,2070|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|2063,2073|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2074,2080|true|false|false|C0038454|Cerebrovascular accident|stroke
Event|Event|SIMPLE_SEGMENT|2074,2080|false|false|false|||stroke
Finding|Finding|SIMPLE_SEGMENT|2074,2080|true|false|false|C5977286|Stroke (heart beat)|stroke
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2083,2086|false|false|false|C0007787;C0917805|Transient Cerebral Ischemia;Transient Ischemic Attack|TIA
Event|Event|SIMPLE_SEGMENT|2083,2086|false|false|false|||TIA
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2088,2092|false|false|false|C4318566|Deep Resection Margin|deep
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2088,2110|false|false|false|C0149871|Deep Vein Thrombosis|deep venous thrombosis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2093,2099|false|false|false|C0042449|Veins|venous
Finding|Finding|SIMPLE_SEGMENT|2093,2110|false|false|false|C0042487;C0517555|Venous Thrombosis;Venous thrombosis after immobility|venous thrombosis
Finding|Pathologic Function|SIMPLE_SEGMENT|2093,2110|false|false|false|C0042487;C0517555|Venous Thrombosis;Venous thrombosis after immobility|venous thrombosis
Event|Event|SIMPLE_SEGMENT|2100,2110|false|false|false|||thrombosis
Finding|Pathologic Function|SIMPLE_SEGMENT|2100,2110|false|false|false|C0040053|Thrombosis|thrombosis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2112,2121|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2112,2121|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|2112,2121|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|SIMPLE_SEGMENT|2112,2130|false|false|false|C0034065|Pulmonary Embolism|pulmonary embolism
Event|Event|SIMPLE_SEGMENT|2122,2130|false|false|false|||embolism
Finding|Finding|SIMPLE_SEGMENT|2122,2130|false|false|false|C0013922;C1704212|Embolism;Embolus|embolism
Finding|Pathologic Function|SIMPLE_SEGMENT|2122,2130|false|false|false|C0013922;C1704212|Embolism;Embolus|embolism
Event|Event|SIMPLE_SEGMENT|2132,2140|false|false|false|||bleeding
Finding|Pathologic Function|SIMPLE_SEGMENT|2132,2140|false|false|false|C0019080|Hemorrhage|bleeding
Finding|Finding|SIMPLE_SEGMENT|2149,2153|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|2149,2153|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|2149,2153|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|SIMPLE_SEGMENT|2157,2164|false|false|false|||surgery
Finding|Finding|SIMPLE_SEGMENT|2157,2164|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|SIMPLE_SEGMENT|2157,2164|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|SIMPLE_SEGMENT|2157,2164|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2157,2164|false|false|false|C0543467|Operative Surgical Procedures|surgery
Event|Event|SIMPLE_SEGMENT|2166,2174|false|false|false|||myalgias
Finding|Sign or Symptom|SIMPLE_SEGMENT|2166,2174|false|false|false|C0231528|Myalgia|myalgias
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|2176,2181|false|false|false|C0022417;C0392905;C1269611|Articular system;Joints|joint
Anatomy|Body System|SIMPLE_SEGMENT|2176,2181|false|false|false|C0022417;C0392905;C1269611|Articular system;Joints|joint
Finding|Finding|SIMPLE_SEGMENT|2176,2181|false|false|false|C0575044|Joint problem|joint
Finding|Sign or Symptom|SIMPLE_SEGMENT|2176,2187|false|false|false|C0003862|Arthralgia|joint pains
Event|Event|SIMPLE_SEGMENT|2182,2187|false|false|false|||pains
Finding|Sign or Symptom|SIMPLE_SEGMENT|2182,2187|false|false|false|C0030193|Pain|pains
Drug|Organic Chemical|SIMPLE_SEGMENT|2189,2194|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2189,2194|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|SIMPLE_SEGMENT|2189,2194|false|false|false|||cough
Finding|Sign or Symptom|SIMPLE_SEGMENT|2189,2194|false|false|false|C0010200|Coughing|cough
Event|Event|SIMPLE_SEGMENT|2196,2206|false|false|false|||hemoptysis
Finding|Sign or Symptom|SIMPLE_SEGMENT|2196,2206|false|false|false|C0019079|Hemoptysis|hemoptysis
Event|Event|SIMPLE_SEGMENT|2208,2213|false|false|false|||black
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2215,2221|false|false|false|C0489144||stools
Event|Event|SIMPLE_SEGMENT|2215,2221|false|false|false|||stools
Finding|Body Substance|SIMPLE_SEGMENT|2215,2221|false|false|false|C0015733|Feces|stools
Finding|Finding|SIMPLE_SEGMENT|2225,2228|false|false|false|C0332575;C1414207;C1416378|DYRK3 gene;IK gene;Redness|red
Finding|Gene or Genome|SIMPLE_SEGMENT|2225,2228|false|false|false|C0332575;C1414207;C1416378|DYRK3 gene;IK gene;Redness|red
Finding|Sign or Symptom|SIMPLE_SEGMENT|2225,2235|false|false|false|C0278012|Red stools|red stools
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2229,2235|false|false|false|C0489144||stools
Event|Event|SIMPLE_SEGMENT|2229,2235|false|false|false|||stools
Finding|Body Substance|SIMPLE_SEGMENT|2229,2235|false|false|false|C0015733|Feces|stools
Event|Event|SIMPLE_SEGMENT|2241,2247|false|false|false|||denies
Event|Event|SIMPLE_SEGMENT|2255,2261|false|false|false|||fevers
Finding|Sign or Symptom|SIMPLE_SEGMENT|2255,2261|true|false|false|C0015967|Fever|fevers
Event|Event|SIMPLE_SEGMENT|2263,2269|false|false|false|||chills
Finding|Sign or Symptom|SIMPLE_SEGMENT|2263,2269|true|false|false|C0085593|Chills|chills
Event|Event|SIMPLE_SEGMENT|2274,2280|false|false|false|||rigors
Finding|Sign or Symptom|SIMPLE_SEGMENT|2274,2280|false|false|false|C0424790|Rigor - Temperature-associated observation|rigors
Event|Event|SIMPLE_SEGMENT|2286,2292|false|false|false|||denies
Finding|Sign or Symptom|SIMPLE_SEGMENT|2293,2303|false|false|false|C0239313|exercise induced|exertional
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2304,2311|false|false|false|C0006497|Buttocks|buttock
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2315,2319|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2315,2319|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Finding|Sign or Symptom|SIMPLE_SEGMENT|2315,2324|true|false|false|C0236040|Pain in calf|calf pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2320,2324|false|true|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|2320,2324|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|2320,2324|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|2320,2324|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|2344,2350|false|false|false|||review
Finding|Idea or Concept|SIMPLE_SEGMENT|2344,2350|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Finding|Intellectual Product|SIMPLE_SEGMENT|2344,2350|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Finding|Functional Concept|SIMPLE_SEGMENT|2344,2353|false|false|false|C0699752|Review of|review of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2344,2361|false|false|false|C0488564;C0488565||review of systems
Procedure|Health Care Activity|SIMPLE_SEGMENT|2344,2361|false|false|false|C0489633|Review of systems (procedure)|review of systems
Event|Event|SIMPLE_SEGMENT|2354,2361|false|false|false|||systems
Finding|Functional Concept|SIMPLE_SEGMENT|2354,2361|false|false|false|C0449913|System|systems
Event|Event|SIMPLE_SEGMENT|2367,2375|false|false|false|||negative
Finding|Classification|SIMPLE_SEGMENT|2367,2375|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|2367,2375|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2367,2375|false|false|false|C5237010|Expression Negative|negative
Finding|Finding|SIMPLE_SEGMENT|2382,2402|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Event|Event|SIMPLE_SEGMENT|2387,2394|false|false|false|||Medical
Finding|Functional Concept|SIMPLE_SEGMENT|2387,2394|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|2387,2394|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|2387,2394|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|2387,2394|false|false|false|C0199168|Medical service|Medical
Finding|Finding|SIMPLE_SEGMENT|2387,2402|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2395,2402|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2395,2402|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2395,2402|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2407,2414|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|SIMPLE_SEGMENT|2407,2414|false|false|false|C1314974|Cardiac attachment|CARDIAC
Finding|Finding|SIMPLE_SEGMENT|2407,2419|false|false|false|C3176821|CARD.RISK|CARDIAC RISK
Finding|Finding|SIMPLE_SEGMENT|2407,2427|false|false|false|C2024776|cardiac risk factors|CARDIAC RISK FACTORS
Event|Event|SIMPLE_SEGMENT|2415,2419|false|false|false|||RISK
Finding|Idea or Concept|SIMPLE_SEGMENT|2415,2419|false|false|false|C0035647|Risk|RISK
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2415,2427|false|false|false|C1830376||RISK FACTORS
Finding|Finding|SIMPLE_SEGMENT|2415,2427|false|false|false|C0035648;C0455624;C1553898|History of - risk factor;risk factors;risk factors - observation list|RISK FACTORS
Finding|Intellectual Product|SIMPLE_SEGMENT|2415,2427|false|false|false|C0035648;C0455624;C1553898|History of - risk factor;risk factors;risk factors - observation list|RISK FACTORS
Event|Event|SIMPLE_SEGMENT|2420,2427|false|false|false|||FACTORS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2432,2440|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|Diabetes
Event|Event|SIMPLE_SEGMENT|2432,2440|false|false|false|||Diabetes
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2445,2457|false|false|false|C0242339|Dyslipidemias|Dyslipidemia
Event|Event|SIMPLE_SEGMENT|2445,2457|false|false|false|||Dyslipidemia
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2462,2465|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|SIMPLE_SEGMENT|2462,2465|false|false|false|||HTN
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2471,2478|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|SIMPLE_SEGMENT|2471,2478|true|false|false|C1314974|Cardiac attachment|CARDIAC
Event|Event|SIMPLE_SEGMENT|2479,2486|false|false|false|||HISTORY
Finding|Conceptual Entity|SIMPLE_SEGMENT|2479,2486|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|HISTORY
Finding|Finding|SIMPLE_SEGMENT|2479,2486|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|HISTORY
Finding|Functional Concept|SIMPLE_SEGMENT|2479,2486|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|HISTORY
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2491,2499|false|false|false|C0018787|Heart|Coronary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2491,2506|false|false|false|C0205042|Coronary artery|Coronary artery
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2491,2514|false|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|Coronary artery disease
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2500,2506|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|SIMPLE_SEGMENT|2500,2506|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2500,2514|false|false|false|C0852949|Arteriopathic disease|artery disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2507,2514|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|2507,2514|false|false|false|||disease
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2518,2527|false|false|false|C0012000|Diastole|Diastolic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2518,2552|false|false|false|C2183328|diastolic congestive heart failure|Diastolic congestive heart failure
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2528,2552|false|false|false|C0018802|Congestive heart failure|congestive heart failure
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2539,2544|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2539,2544|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|2539,2544|false|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2539,2552|false|false|false|C0018801;C0018802|Congestive heart failure;Heart failure|heart failure
Event|Event|SIMPLE_SEGMENT|2545,2552|false|false|false|||failure
Finding|Functional Concept|SIMPLE_SEGMENT|2545,2552|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|SIMPLE_SEGMENT|2545,2552|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|SIMPLE_SEGMENT|2545,2552|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Event|Event|SIMPLE_SEGMENT|2556,2560|false|false|false|||CABG
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2556,2560|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Event|Event|SIMPLE_SEGMENT|2562,2566|false|false|false|||CABG
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2562,2566|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2572,2603|false|false|false|C1449706|Coronary Artery Bypass, Off-Pump|Off pump coronary artery bypass
Finding|Molecular Function|SIMPLE_SEGMENT|2576,2580|false|false|false|C1150186|matrix metalloproteinase 7 activity|pump
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2581,2589|false|false|false|C0018787|Heart|coronary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2581,2596|false|false|false|C0205042|Coronary artery|coronary artery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2581,2603|false|false|false|C0010055|Coronary Artery Bypass Surgery|coronary artery bypass
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2581,2609|false|false|false|C0010055|Coronary Artery Bypass Surgery|coronary artery bypass graft
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2590,2596|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|SIMPLE_SEGMENT|2590,2596|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2590,2609|false|false|false|C5886769|Arterial bypass graft|artery bypass graft
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2597,2603|false|false|false|C0813207|Creation of shunt|bypass
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2597,2609|false|false|false|C0185098|Bypass graft|bypass graft
Anatomy|Tissue|SIMPLE_SEGMENT|2604,2609|false|false|false|C0332835|Transplanted tissue|graft
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|2604,2609|false|false|false|C0181074;C1705210|Graft Dosage Form;Graft material|graft
Event|Event|SIMPLE_SEGMENT|2604,2609|false|false|false|||graft
Finding|Intellectual Product|SIMPLE_SEGMENT|2604,2609|false|false|false|C1546653|Graft - Specimen Source Codes|graft
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2604,2609|false|false|false|C1961139;C3683798|Graft Procedures on the Head;Grafting procedure|graft
Finding|Functional Concept|SIMPLE_SEGMENT|2614,2618|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2622,2645|false|false|false|C0226276|Structure of internal thoracic artery|internal mammary artery
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2631,2638|false|false|false|C0006141;C0929301|Breast;Mammary gland|mammary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2631,2645|false|false|false|C0024661|Mammary Arteries|mammary artery
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2639,2645|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|SIMPLE_SEGMENT|2639,2645|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Finding|Functional Concept|SIMPLE_SEGMENT|2649,2653|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2649,2680|false|false|false|C0226032;C1321506|Anterior descending branch of left coronary artery|left anterior descending artery
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2654,2662|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Finding|Functional Concept|SIMPLE_SEGMENT|2663,2673|false|false|false|C1547177|Sequencing - Descending|descending
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2674,2680|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|SIMPLE_SEGMENT|2674,2680|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2687,2701|false|false|false|C0036186;C0392907|Great saphenous vein structure;Saphenous Vein|saphenous vein
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2697,2701|false|false|false|C0042449|Veins|vein
Anatomy|Tissue|SIMPLE_SEGMENT|2702,2708|false|false|false|C0332835|Transplanted tissue|grafts
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|2702,2708|false|false|false|C0181074|Graft material|grafts
Event|Event|SIMPLE_SEGMENT|2702,2708|false|false|false|||grafts
Finding|Finding|SIMPLE_SEGMENT|2733,2741|false|false|false|C1550517|Target Awareness - marginal|marginal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2742,2750|false|false|false|C0003842;C0226004|Arterial system;Arteries|arteries
Anatomy|Body System|SIMPLE_SEGMENT|2742,2750|false|false|false|C0003842;C0226004|Arterial system;Arteries|arteries
Procedure|Health Care Activity|SIMPLE_SEGMENT|2742,2750|false|false|false|C0397581|Procedure on artery|arteries
Finding|Functional Concept|SIMPLE_SEGMENT|2756,2768|false|false|false|C1522243|Percutaneous Route of Drug Administration|PERCUTANEOUS
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2756,2791|false|false|false|C1532338|Percutaneous Coronary Intervention|PERCUTANEOUS CORONARY INTERVENTIONS
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2769,2777|false|false|false|C0018787|Heart|CORONARY
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2778,2791|false|false|false|C2979881||INTERVENTIONS
Event|Event|SIMPLE_SEGMENT|2778,2791|false|false|false|||INTERVENTIONS
Procedure|Health Care Activity|SIMPLE_SEGMENT|2778,2791|false|false|false|C0886296;C1273869|Intervention regimes;Nursing interventions|INTERVENTIONS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2793,2796|false|false|false|C0006430|Burning Mouth Syndrome|BMS
Event|Event|SIMPLE_SEGMENT|2793,2796|false|false|false|||BMS
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2800,2808|false|false|false|C4489236|Proximal Resection Margin|proximal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2809,2812|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2809,2812|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|SIMPLE_SEGMENT|2809,2812|false|false|false|||LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|2809,2812|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2820,2823|false|false|false|C4551552|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|DES
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2820,2823|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2820,2823|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Hormone|SIMPLE_SEGMENT|2820,2823|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Organic Chemical|SIMPLE_SEGMENT|2820,2823|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2820,2823|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Event|Event|SIMPLE_SEGMENT|2820,2823|false|false|false|||DES
Finding|Gene or Genome|SIMPLE_SEGMENT|2820,2823|false|false|false|C1413980|DES gene|DES
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2831,2834|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2831,2834|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|SIMPLE_SEGMENT|2831,2834|false|false|false|||LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|2831,2834|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2840,2843|false|false|false|C4551552|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|DES
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2840,2843|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2840,2843|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Hormone|SIMPLE_SEGMENT|2840,2843|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Organic Chemical|SIMPLE_SEGMENT|2840,2843|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2840,2843|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Event|Event|SIMPLE_SEGMENT|2840,2843|false|false|false|||DES
Finding|Gene or Genome|SIMPLE_SEGMENT|2840,2843|false|false|false|C1413980|DES gene|DES
Event|Event|SIMPLE_SEGMENT|2847,2851|false|false|false|||edge
Finding|Conceptual Entity|SIMPLE_SEGMENT|2847,2851|false|false|false|C2697523|Graph Edge|edge
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2863,2866|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2863,2866|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|2863,2866|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2867,2870|false|false|false|C4551552|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|DES
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2867,2870|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2867,2870|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Hormone|SIMPLE_SEGMENT|2867,2870|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Organic Chemical|SIMPLE_SEGMENT|2867,2870|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2867,2870|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Event|Event|SIMPLE_SEGMENT|2867,2870|false|false|false|||DES
Finding|Gene or Genome|SIMPLE_SEGMENT|2867,2870|false|false|false|C1413980|DES gene|DES
Event|Event|SIMPLE_SEGMENT|2877,2885|false|false|false|||stenosis
Finding|Pathologic Function|SIMPLE_SEGMENT|2877,2885|false|false|false|C1261287|Stenosis|stenosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2886,2892|false|false|false|C4522154|Distal Resection Margin|distal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2907,2910|false|false|false|C4551552|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|DES
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2907,2910|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2907,2910|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Hormone|SIMPLE_SEGMENT|2907,2910|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Organic Chemical|SIMPLE_SEGMENT|2907,2910|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2907,2910|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Event|Event|SIMPLE_SEGMENT|2907,2910|false|false|false|||DES
Finding|Gene or Genome|SIMPLE_SEGMENT|2907,2910|false|false|false|C1413980|DES gene|DES
Finding|Individual Behavior|SIMPLE_SEGMENT|2926,2932|false|false|false|C0562458|Pacing up and down|PACING
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2933,2936|false|false|false|C0020725;C0021122|Disruptive, Impulse Control, and Conduct Disorders;Type II Mucolipidosis|ICD
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|2933,2936|false|false|false|C0020725;C0021122|Disruptive, Impulse Control, and Conduct Disorders;Type II Mucolipidosis|ICD
Event|Event|SIMPLE_SEGMENT|2933,2936|false|false|false|||ICD
Finding|Gene or Genome|SIMPLE_SEGMENT|2933,2936|false|false|false|C0870733;C5891008|GNPTAB wt Allele;International Classification of Diseases|ICD
Finding|Intellectual Product|SIMPLE_SEGMENT|2933,2936|false|false|false|C0870733;C5891008|GNPTAB wt Allele;International Classification of Diseases|ICD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2933,2936|false|false|false|C5575277|Icd Regimen|ICD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2944,2958|false|false|false|C0028756|Morbid obesity|Morbid obesity
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2951,2958|false|false|false|C0028754|Obesity|obesity
Event|Event|SIMPLE_SEGMENT|2951,2958|false|false|false|||obesity
Finding|Finding|SIMPLE_SEGMENT|2951,2958|false|false|false|C4759928|BODY MASS INDEX QUANTITATIVE TRAIT LOCUS 20|obesity
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2962,2966|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2962,2966|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|SIMPLE_SEGMENT|2962,2966|false|false|false|||COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|2962,2966|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2969,2973|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Event|Event|SIMPLE_SEGMENT|2969,2973|false|false|false|||GERD
Finding|Functional Concept|SIMPLE_SEGMENT|2976,2981|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2976,2994|false|false|false|C0828608|Right tendinous cuff|Right rotator cuff
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2982,2994|false|false|false|C0085515|Rotator Cuff|rotator cuff
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|2982,3001|false|false|false|C0851122|Rotator Cuff Injuries|rotator cuff injury
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2990,2994|false|false|false|C1550244|Cuff - body part|cuff
Finding|Pathologic Function|SIMPLE_SEGMENT|2990,2994|false|false|false|C3668885|Cuffing (morphologic abnormality)|cuff
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|2995,3001|false|false|false|C3263722;C3263723|Traumatic AND/OR non-traumatic injury;Traumatic injury|injury
Event|Event|SIMPLE_SEGMENT|2995,3001|false|false|false|||injury
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3002,3010|false|false|false|C0006444|Bursitis|bursitis
Event|Event|SIMPLE_SEGMENT|3002,3010|false|false|false|||bursitis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3013,3022|false|false|false|C0149931|Migraine Disorders|Migraines
Event|Event|SIMPLE_SEGMENT|3013,3022|false|false|false|||Migraines
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|3025,3035|false|false|false|C0011570;C0011581;C0344315;C0812393|Cancer patients and suicide and depression;Depressed mood;Depressive disorder;Mental Depression|Depression
Event|Event|SIMPLE_SEGMENT|3025,3035|false|false|false|||Depression
Finding|Functional Concept|SIMPLE_SEGMENT|3025,3035|false|false|false|C0460137;C1579931|Depression - motion|Depression
Finding|Sign or Symptom|SIMPLE_SEGMENT|3025,3035|false|false|false|C0460137;C1579931|Depression - motion|Depression
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3038,3041|false|false|false|C0029408|Degenerative polyarthritis|DJD
Event|Event|SIMPLE_SEGMENT|3038,3041|false|false|false|||DJD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3044,3055|false|false|false|C0019112|Hemorrhoids|Hemorrhoids
Event|Event|SIMPLE_SEGMENT|3044,3055|false|false|false|||Hemorrhoids
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3058,3065|false|false|false|C0035854|Rosacea|Rosacea
Event|Event|SIMPLE_SEGMENT|3058,3065|false|false|false|||Rosacea
Finding|Functional Concept|SIMPLE_SEGMENT|3071,3077|false|false|false|C0728831|Social|Social
Finding|Finding|SIMPLE_SEGMENT|3071,3085|false|false|false|C0424945;C3714536|Social History;Social and personal history|Social History
Event|Event|SIMPLE_SEGMENT|3078,3085|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|3078,3085|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|3078,3085|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|3078,3085|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Classification|SIMPLE_SEGMENT|3091,3097|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|SIMPLE_SEGMENT|3091,3097|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|SIMPLE_SEGMENT|3091,3097|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|SIMPLE_SEGMENT|3091,3097|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Finding|SIMPLE_SEGMENT|3091,3105|false|false|false|C0241889|Family Medical History|Family History
Event|Event|SIMPLE_SEGMENT|3098,3105|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|3098,3105|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|3098,3105|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|3098,3105|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Event|Event|SIMPLE_SEGMENT|3146,3150|false|false|false|||know
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3151,3161|false|true|false|C3812393|ErbB Receptors|her family
Drug|Enzyme|SIMPLE_SEGMENT|3151,3161|false|true|false|C3812393|ErbB Receptors|her family
Finding|Receptor|SIMPLE_SEGMENT|3151,3161|false|true|false|C3812393|ErbB Receptors|her family
Event|Event|SIMPLE_SEGMENT|3155,3161|false|false|false|||family
Finding|Classification|SIMPLE_SEGMENT|3155,3161|true|true|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|3155,3161|true|true|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|3155,3161|true|true|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|3155,3161|true|true|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Event|Event|SIMPLE_SEGMENT|3168,3176|false|false|false|||Physical
Finding|Finding|SIMPLE_SEGMENT|3168,3176|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|3168,3176|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|3168,3176|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|3168,3181|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|3168,3181|false|false|false|C0031809|Physical Examination|Physical Exam
Event|Event|SIMPLE_SEGMENT|3177,3181|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|3177,3181|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|3177,3181|false|false|false|C0582103|Medical Examination|Exam
Event|Event|SIMPLE_SEGMENT|3183,3192|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|3183,3192|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Event|Event|SIMPLE_SEGMENT|3237,3244|false|false|false|||GENERAL
Finding|Classification|SIMPLE_SEGMENT|3237,3244|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|3237,3244|false|false|false|C3812897|General medical service|GENERAL
Event|Event|SIMPLE_SEGMENT|3246,3250|false|false|false|||WDWN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3256,3259|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3256,3259|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3256,3259|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|3256,3259|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3256,3259|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|SIMPLE_SEGMENT|3256,3259|false|false|false|||NAD
Finding|Finding|SIMPLE_SEGMENT|3256,3259|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Finding|Finding|SIMPLE_SEGMENT|3261,3269|false|false|false|C1961028|Oriented to place|Oriented
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3274,3278|false|false|false|C2713234||Mood
Event|Event|SIMPLE_SEGMENT|3274,3278|false|false|false|||Mood
Finding|Conceptual Entity|SIMPLE_SEGMENT|3274,3278|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|Mood
Finding|Finding|SIMPLE_SEGMENT|3274,3278|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|Mood
Finding|Mental Process|SIMPLE_SEGMENT|3274,3278|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|Mood
Event|Event|SIMPLE_SEGMENT|3280,3286|false|false|false|||affect
Event|Event|SIMPLE_SEGMENT|3287,3298|false|false|false|||appropriate
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3302,3307|false|false|false|C1512338|HEENT|HEENT
Event|Event|SIMPLE_SEGMENT|3309,3313|false|false|false|||NCAT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3315,3321|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3315,3321|false|false|false|C0036412|Scleral Diseases|Sclera
Event|Event|SIMPLE_SEGMENT|3315,3321|false|false|false|||Sclera
Procedure|Health Care Activity|SIMPLE_SEGMENT|3315,3321|false|false|false|C2228481|examination of sclera|Sclera
Event|Event|SIMPLE_SEGMENT|3322,3331|false|false|false|||anicteric
Finding|Finding|SIMPLE_SEGMENT|3322,3331|false|false|false|C0205180|Anicteric|anicteric
Event|Event|SIMPLE_SEGMENT|3333,3338|false|false|false|||PERRL
Finding|Finding|SIMPLE_SEGMENT|3333,3338|false|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Event|Event|SIMPLE_SEGMENT|3340,3344|false|false|false|||EOMI
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3346,3357|false|false|false|C0009758;C0229274|Structure of palpebral conjunctiva;conjunctiva|Conjunctiva
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3346,3357|false|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|Conjunctiva
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3346,3357|false|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|Conjunctiva
Event|Event|SIMPLE_SEGMENT|3346,3357|false|false|false|||Conjunctiva
Finding|Body Substance|SIMPLE_SEGMENT|3346,3357|false|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|Conjunctiva
Finding|Intellectual Product|SIMPLE_SEGMENT|3346,3357|false|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|Conjunctiva
Procedure|Health Care Activity|SIMPLE_SEGMENT|3346,3357|false|false|false|C0872390;C2228431|Procedure on conjunctiva;examination of conjunctiva|Conjunctiva
Event|Event|SIMPLE_SEGMENT|3373,3379|false|false|false|||pallor
Finding|Finding|SIMPLE_SEGMENT|3373,3379|true|false|false|C0241137|Pallor of skin|pallor
Event|Event|SIMPLE_SEGMENT|3383,3391|false|false|false|||cyanosis
Finding|Sign or Symptom|SIMPLE_SEGMENT|3383,3391|true|false|false|C0010520|Cyanosis|cyanosis
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|3399,3403|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3399,3403|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|3399,3403|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|3399,3403|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3399,3410|false|false|false|C0026639|Oral mucous membrane structure|oral mucosa
Anatomy|Tissue|SIMPLE_SEGMENT|3404,3410|false|false|false|C0026724|Mucous Membrane|mucosa
Finding|Intellectual Product|SIMPLE_SEGMENT|3404,3410|false|false|false|C1561514||mucosa
Event|Event|SIMPLE_SEGMENT|3415,3426|false|false|false|||xanthalesma
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3431,3435|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|SIMPLE_SEGMENT|3431,3435|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|SIMPLE_SEGMENT|3431,3435|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Event|Event|SIMPLE_SEGMENT|3437,3443|false|false|false|||Supple
Finding|Functional Concept|SIMPLE_SEGMENT|3437,3443|false|false|false|C0332254|Supple|Supple
Event|Event|SIMPLE_SEGMENT|3452,3455|false|false|false|||JVP
Finding|Finding|SIMPLE_SEGMENT|3452,3455|true|false|false|C0428897|Jugular venous pressure|JVP
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3458,3465|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|SIMPLE_SEGMENT|3458,3465|false|false|false|C1314974|Cardiac attachment|CARDIAC
Event|Event|SIMPLE_SEGMENT|3467,3470|false|false|false|||PMI
Finding|Finding|SIMPLE_SEGMENT|3467,3470|false|false|false|C1417244;C1418674;C1823304;C5238618;C5780972|MPI gene;PMM2 gene;PMM2 wt Allele;Point of Maximum Impulse;TMEM11 gene|PMI
Finding|Gene or Genome|SIMPLE_SEGMENT|3467,3470|false|false|false|C1417244;C1418674;C1823304;C5238618;C5780972|MPI gene;PMM2 gene;PMM2 wt Allele;Point of Maximum Impulse;TMEM11 gene|PMI
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|3486,3503|false|false|false|C0230136;C4085247|Space of intercostal compartment;Structure of intercostal space|intercostal space
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3498,3503|false|false|false|C0282173|Space (Astronomy)|space
Event|Event|SIMPLE_SEGMENT|3505,3518|false|false|false|||midclavicular
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3520,3524|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|3520,3524|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Substance|SIMPLE_SEGMENT|3520,3524|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Event|Event|SIMPLE_SEGMENT|3520,3524|false|false|false|||line
Finding|Intellectual Product|SIMPLE_SEGMENT|3520,3524|false|false|false|C1546701|line source specimen code|line
Event|Event|SIMPLE_SEGMENT|3526,3529|false|false|false|||RRR
Anatomy|Cell Component|SIMPLE_SEGMENT|3540,3547|false|false|false|C1660780|midline cell component|Midline
Event|Event|SIMPLE_SEGMENT|3548,3552|false|false|false|||scar
Finding|Finding|SIMPLE_SEGMENT|3548,3552|false|false|false|C0241158;C1419736;C2004491|Cicatrix;RPS4X gene;Scar Tissue|scar
Finding|Gene or Genome|SIMPLE_SEGMENT|3548,3552|false|false|false|C0241158;C1419736;C2004491|Cicatrix;RPS4X gene;Scar Tissue|scar
Finding|Pathologic Function|SIMPLE_SEGMENT|3548,3552|false|false|false|C0241158;C1419736;C2004491|Cicatrix;RPS4X gene;Scar Tissue|scar
Finding|Finding|SIMPLE_SEGMENT|3558,3572|false|false|false|C2169607|recent surgery|recent surgery
Event|Event|SIMPLE_SEGMENT|3565,3572|false|false|false|||surgery
Finding|Finding|SIMPLE_SEGMENT|3565,3572|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|SIMPLE_SEGMENT|3565,3572|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|SIMPLE_SEGMENT|3565,3572|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3565,3572|false|false|false|C0543467|Operative Surgical Procedures|surgery
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3581,3586|false|false|false|C0024109|Lung|LUNGS
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3592,3597|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|3592,3597|false|false|false|C0741025|Chest problem|chest
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3592,3602|false|false|false|C0205076;C4266615|Chest wall structure;Chest>Chest wall|chest wall
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3592,3602|false|false|false|C0205076;C4266615|Chest wall structure;Chest>Chest wall|chest wall
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|3592,3614|true|false|false|C3164427|Deformity of chest wall|chest wall deformities
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|3603,3614|true|false|false|C0000768|Congenital Abnormality|deformities
Event|Event|SIMPLE_SEGMENT|3603,3614|false|false|false|||deformities
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|3616,3625|true|false|false|C0036439;C0559260;C0700208|Acquired scoliosis;Congenital scoliosis|scoliosis
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|3616,3625|true|false|false|C0036439;C0559260;C0700208|Acquired scoliosis;Congenital scoliosis|scoliosis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3616,3625|true|false|false|C0036439;C0559260;C0700208|Acquired scoliosis;Congenital scoliosis|scoliosis
Event|Event|SIMPLE_SEGMENT|3616,3625|false|false|false|||scoliosis
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|3629,3637|true|false|false|C0022821;C0022822;C0265673|Acquired kyphosis;Congenital kyphosis;Kyphosis deformity of spine|kyphosis
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|3629,3637|true|false|false|C0022821;C0022822;C0265673|Acquired kyphosis;Congenital kyphosis;Kyphosis deformity of spine|kyphosis
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|3629,3637|true|false|false|C0022821;C0022822;C0265673|Acquired kyphosis;Congenital kyphosis;Kyphosis deformity of spine|kyphosis
Event|Event|SIMPLE_SEGMENT|3629,3637|false|false|false|||kyphosis
Finding|Finding|SIMPLE_SEGMENT|3629,3637|true|false|false|C2115817|kyphosis|kyphosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3639,3643|false|false|false|C0231832|Respiratory rate|Resp
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3639,3643|false|false|false|C0851355|Respiratory, thoracic and mediastinal disorders|Resp
Event|Event|SIMPLE_SEGMENT|3639,3643|false|false|false|||Resp
Event|Event|SIMPLE_SEGMENT|3650,3659|false|false|false|||unlabored
Finding|Functional Concept|SIMPLE_SEGMENT|3650,3659|false|false|false|C2983702|Unlabored|unlabored
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|3664,3680|true|false|false|C0158784|Accessory skeletal muscle|accessory muscle
Finding|Finding|SIMPLE_SEGMENT|3664,3684|true|false|false|C1821466|Use of accessory muscles|accessory muscle use
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3674,3680|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Anatomy|Tissue|SIMPLE_SEGMENT|3674,3680|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Event|Event|SIMPLE_SEGMENT|3681,3684|false|false|false|||use
Finding|Functional Concept|SIMPLE_SEGMENT|3681,3684|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|SIMPLE_SEGMENT|3681,3684|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Drug|Organic Chemical|SIMPLE_SEGMENT|3686,3690|false|false|false|C0951233|cetrimonium bromide|CTAB
Event|Event|SIMPLE_SEGMENT|3686,3690|false|false|false|||CTAB
Event|Event|SIMPLE_SEGMENT|3695,3703|false|false|false|||crackles
Finding|Finding|SIMPLE_SEGMENT|3695,3703|true|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Event|Event|SIMPLE_SEGMENT|3706,3713|false|false|false|||wheezes
Finding|Sign or Symptom|SIMPLE_SEGMENT|3706,3713|false|false|false|C0043144|Wheezing|wheezes
Event|Event|SIMPLE_SEGMENT|3717,3724|false|false|false|||rhonchi
Finding|Finding|SIMPLE_SEGMENT|3717,3724|false|false|false|C0035508|Rhonchi|rhonchi
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3728,3735|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3728,3735|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Event|Event|SIMPLE_SEGMENT|3728,3735|false|false|false|||ABDOMEN
Finding|Finding|SIMPLE_SEGMENT|3728,3735|false|false|false|C0941288|Abdomen problem|ABDOMEN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3737,3741|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Event|Event|SIMPLE_SEGMENT|3737,3741|false|false|false|||Soft
Event|Event|SIMPLE_SEGMENT|3743,3747|false|false|false|||NTND
Event|Event|SIMPLE_SEGMENT|3752,3755|false|false|false|||HSM
Finding|Gene or Genome|SIMPLE_SEGMENT|3752,3755|true|false|false|C1537594|LRRC4B gene|HSM
Event|Event|SIMPLE_SEGMENT|3759,3769|false|false|false|||tenderness
Finding|Mental Process|SIMPLE_SEGMENT|3759,3769|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|SIMPLE_SEGMENT|3759,3769|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3773,3784|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Event|Event|SIMPLE_SEGMENT|3789,3790|false|false|false|||c
Event|Event|SIMPLE_SEGMENT|3798,3807|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|3798,3807|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|3798,3807|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|3798,3807|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|3798,3807|false|false|false|C0030685|Patient Discharge|Discharge
Event|Event|SIMPLE_SEGMENT|3860,3866|false|false|false|||Intake
Finding|Functional Concept|SIMPLE_SEGMENT|3860,3866|false|false|false|C1512806|Intake|Intake
Procedure|Health Care Activity|SIMPLE_SEGMENT|3860,3866|false|false|false|C3251814;C4521161|Intake (treatment);Measurement of fluid intake|Intake
Event|Event|SIMPLE_SEGMENT|3876,3882|false|false|false|||Output
Finding|Conceptual Entity|SIMPLE_SEGMENT|3876,3882|false|false|false|C1709366|system output|Output
Procedure|Health Care Activity|SIMPLE_SEGMENT|3876,3882|false|false|false|C3251815|Measurement of fluid output|Output
Event|Event|SIMPLE_SEGMENT|3899,3907|false|false|false|||recorded
Event|Event|SIMPLE_SEGMENT|3910,3917|false|false|false|||GENERAL
Finding|Classification|SIMPLE_SEGMENT|3910,3917|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|3910,3917|false|false|false|C3812897|General medical service|GENERAL
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3920,3925|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|3920,3925|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3920,3925|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|SIMPLE_SEGMENT|3920,3925|false|false|false|||Alert
Finding|Finding|SIMPLE_SEGMENT|3920,3925|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|3920,3925|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|3920,3925|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|SIMPLE_SEGMENT|3927,3938|false|false|false|||interactive
Finding|Functional Concept|SIMPLE_SEGMENT|3927,3938|false|false|false|C1704675|Interaction|interactive
Finding|Finding|SIMPLE_SEGMENT|3940,3944|false|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|3945,3954|false|false|false|||appearing
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3958,3961|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3958,3961|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3958,3961|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|3958,3961|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3958,3961|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|SIMPLE_SEGMENT|3958,3961|false|false|false|||NAD
Finding|Finding|SIMPLE_SEGMENT|3958,3961|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3964,3969|false|false|false|C1512338|HEENT|HEENT
Event|Event|SIMPLE_SEGMENT|3972,3978|false|false|false|||PERRLA
Finding|Finding|SIMPLE_SEGMENT|3972,3978|false|false|false|C2143306|PERRLA|PERRLA
Event|Event|SIMPLE_SEGMENT|3980,3984|false|false|false|||EOMI
Event|Event|SIMPLE_SEGMENT|3994,4003|false|false|false|||anicteric
Finding|Finding|SIMPLE_SEGMENT|3994,4003|false|false|false|C0205180|Anicteric|anicteric
Finding|Finding|SIMPLE_SEGMENT|4005,4025|false|false|false|C1999162|dry mucous membranes|dry mucous membranes
Finding|Body Substance|SIMPLE_SEGMENT|4009,4015|false|false|false|C0026727;C2753459|Mucus (substance);mucus layer|mucous
Anatomy|Tissue|SIMPLE_SEGMENT|4009,4025|false|false|false|C0026724|Mucous Membrane|mucous membranes
Finding|Finding|SIMPLE_SEGMENT|4009,4025|false|false|false|C2230150|moisture of mucous membranes (physical finding)|mucous membranes
Anatomy|Tissue|SIMPLE_SEGMENT|4016,4025|false|false|false|C0025255|Membrane Tissue|membranes
Event|Event|SIMPLE_SEGMENT|4031,4036|false|false|false|||clear
Finding|Idea or Concept|SIMPLE_SEGMENT|4031,4036|false|false|false|C1550016|Remote control command - Clear|clear
Event|Event|SIMPLE_SEGMENT|4041,4044|false|false|false|||JVP
Finding|Finding|SIMPLE_SEGMENT|4041,4044|true|false|false|C0428897|Jugular venous pressure|JVP
Event|Event|SIMPLE_SEGMENT|4045,4055|false|false|false|||visualized
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4059,4064|false|false|false|C0018787;C4037974|Chest>Heart;Heart|HEART
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4059,4064|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|HEART
Event|Event|SIMPLE_SEGMENT|4059,4064|false|false|false|||HEART
Finding|Sign or Symptom|SIMPLE_SEGMENT|4059,4064|false|false|false|C0795691|HEART PROBLEM|HEART
Event|Event|SIMPLE_SEGMENT|4067,4070|false|false|false|||RRR
Event|Event|SIMPLE_SEGMENT|4085,4088|false|false|false|||MRG
Finding|Gene or Genome|SIMPLE_SEGMENT|4085,4088|true|false|false|C1422304|MAS1L gene|MRG
Event|Event|SIMPLE_SEGMENT|4090,4094|false|false|false|||Scar
Finding|Finding|SIMPLE_SEGMENT|4090,4094|false|false|false|C0241158;C1419736;C2004491|Cicatrix;RPS4X gene;Scar Tissue|Scar
Finding|Gene or Genome|SIMPLE_SEGMENT|4090,4094|false|false|false|C0241158;C1419736;C2004491|Cicatrix;RPS4X gene;Scar Tissue|Scar
Finding|Pathologic Function|SIMPLE_SEGMENT|4090,4094|false|false|false|C0241158;C1419736;C2004491|Cicatrix;RPS4X gene;Scar Tissue|Scar
Finding|Finding|SIMPLE_SEGMENT|4100,4114|false|false|false|C2169607|recent surgery|recent surgery
Event|Event|SIMPLE_SEGMENT|4107,4114|false|false|false|||surgery
Finding|Finding|SIMPLE_SEGMENT|4107,4114|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|SIMPLE_SEGMENT|4107,4114|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|SIMPLE_SEGMENT|4107,4114|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4107,4114|false|false|false|C0543467|Operative Surgical Procedures|surgery
Event|Event|SIMPLE_SEGMENT|4115,4122|false|false|false|||present
Finding|Finding|SIMPLE_SEGMENT|4115,4122|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|SIMPLE_SEGMENT|4115,4122|false|false|false|C0150312;C0449450|Present;Presentation|present
Anatomy|Cell Component|SIMPLE_SEGMENT|4127,4134|false|false|false|C1660780|midline cell component|midline
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|4136,4141|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|Wound
Event|Event|SIMPLE_SEGMENT|4136,4141|false|false|false|||Wound
Finding|Body Substance|SIMPLE_SEGMENT|4136,4141|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|Wound
Finding|Functional Concept|SIMPLE_SEGMENT|4136,4141|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|Wound
Finding|Intellectual Product|SIMPLE_SEGMENT|4136,4141|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|Wound
Event|Event|SIMPLE_SEGMENT|4145,4152|false|false|false|||healing
Finding|Finding|SIMPLE_SEGMENT|4153,4157|false|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|4162,4172|false|false|false|||tenderness
Finding|Mental Process|SIMPLE_SEGMENT|4162,4172|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|SIMPLE_SEGMENT|4162,4172|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Event|Event|SIMPLE_SEGMENT|4179,4183|false|false|false|||scar
Finding|Finding|SIMPLE_SEGMENT|4179,4183|false|false|false|C0241158;C1419736;C2004491|Cicatrix;RPS4X gene;Scar Tissue|scar
Finding|Gene or Genome|SIMPLE_SEGMENT|4179,4183|false|false|false|C0241158;C1419736;C2004491|Cicatrix;RPS4X gene;Scar Tissue|scar
Finding|Pathologic Function|SIMPLE_SEGMENT|4179,4183|false|false|false|C0241158;C1419736;C2004491|Cicatrix;RPS4X gene;Scar Tissue|scar
Finding|Finding|SIMPLE_SEGMENT|4186,4192|false|false|false|C5202796|Intensity and Distress 1|Slight
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4193,4201|false|false|false|C0041834|Erythema|erythema
Event|Event|SIMPLE_SEGMENT|4193,4201|false|false|false|||erythema
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4205,4209|false|false|false|C2987514|Anatomical base|base
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4205,4209|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Chemical Viewed Functionally|SIMPLE_SEGMENT|4205,4209|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|4205,4209|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Finding|Gene or Genome|SIMPLE_SEGMENT|4205,4209|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Finding|Idea or Concept|SIMPLE_SEGMENT|4205,4209|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Event|Governmental or Regulatory Activity|SIMPLE_SEGMENT|4218,4222|false|false|false|C1510751|Academic Research Enhancement Awards|area
Event|Event|SIMPLE_SEGMENT|4232,4236|false|false|false|||scar
Finding|Finding|SIMPLE_SEGMENT|4232,4236|false|false|false|C0241158;C1419736;C2004491|Cicatrix;RPS4X gene;Scar Tissue|scar
Finding|Gene or Genome|SIMPLE_SEGMENT|4232,4236|false|false|false|C0241158;C1419736;C2004491|Cicatrix;RPS4X gene;Scar Tissue|scar
Finding|Pathologic Function|SIMPLE_SEGMENT|4232,4236|false|false|false|C0241158;C1419736;C2004491|Cicatrix;RPS4X gene;Scar Tissue|scar
Event|Event|SIMPLE_SEGMENT|4240,4247|false|false|false|||present
Finding|Finding|SIMPLE_SEGMENT|4240,4247|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|SIMPLE_SEGMENT|4240,4247|false|false|false|C0150312;C0449450|Present;Presentation|present
Event|Event|SIMPLE_SEGMENT|4263,4274|false|false|false|||debridement
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4263,4274|false|false|false|C0011079;C3245462|Debridement;Sterile maggot wound debridement|debridement
Event|Event|SIMPLE_SEGMENT|4278,4286|false|false|false|||reported
Event|Event|SIMPLE_SEGMENT|4291,4299|false|false|false|||patinent
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4305,4310|false|false|false|C0024109|Lung|LUNGS
Event|Event|SIMPLE_SEGMENT|4323,4331|false|false|false|||crackles
Finding|Finding|SIMPLE_SEGMENT|4323,4331|false|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Event|Event|SIMPLE_SEGMENT|4332,4339|false|false|false|||present
Finding|Finding|SIMPLE_SEGMENT|4332,4339|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|SIMPLE_SEGMENT|4332,4339|false|false|false|C0150312;C0449450|Present;Presentation|present
Drug|Chemical Viewed Functionally|SIMPLE_SEGMENT|4343,4348|false|false|false|C0178499|Base|bases
Event|Event|SIMPLE_SEGMENT|4343,4348|false|false|false|||bases
Event|Event|SIMPLE_SEGMENT|4353,4360|false|false|false|||wheezes
Finding|Sign or Symptom|SIMPLE_SEGMENT|4353,4360|true|false|false|C0043144|Wheezing|wheezes
Event|Event|SIMPLE_SEGMENT|4365,4371|false|false|false|||rhonci
Event|Event|SIMPLE_SEGMENT|4373,4385|false|false|false|||Respirations
Finding|Physiologic Function|SIMPLE_SEGMENT|4373,4385|false|false|false|C0035203|Respiration|Respirations
Event|Event|SIMPLE_SEGMENT|4386,4395|false|false|false|||unlabored
Finding|Functional Concept|SIMPLE_SEGMENT|4386,4395|false|false|false|C2983702|Unlabored|unlabored
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4399,4406|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4399,4406|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Finding|Finding|SIMPLE_SEGMENT|4399,4406|false|false|false|C0941288|Abdomen problem|ABDOMEN
Event|Event|SIMPLE_SEGMENT|4409,4413|false|false|false|||NABS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4415,4419|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|SIMPLE_SEGMENT|4415,4419|false|false|false|||soft
Event|Event|SIMPLE_SEGMENT|4430,4436|false|false|false|||masses
Event|Event|SIMPLE_SEGMENT|4440,4443|false|false|false|||HSM
Finding|Gene or Genome|SIMPLE_SEGMENT|4440,4443|true|false|false|C1537594|LRRC4B gene|HSM
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4446,4457|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Event|Event|SIMPLE_SEGMENT|4460,4463|false|false|false|||WWP
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|4478,4495|false|false|false|C0232139|Peripheral pulse|peripheral pulses
Drug|Food|SIMPLE_SEGMENT|4489,4495|false|false|false|C5890763||pulses
Event|Event|SIMPLE_SEGMENT|4489,4495|false|false|false|||pulses
Finding|Physiologic Function|SIMPLE_SEGMENT|4489,4495|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|SIMPLE_SEGMENT|4489,4495|false|false|false|C0034107|Pulse taking|pulses
Event|Event|SIMPLE_SEGMENT|4506,4511|false|false|false|||awake
Finding|Finding|SIMPLE_SEGMENT|4506,4511|false|false|false|C0234422|Awake (finding)|awake
Anatomy|Body System|SIMPLE_SEGMENT|4520,4523|false|false|false|C3714787|Central Nervous System|CNs
Event|Event|SIMPLE_SEGMENT|4539,4545|false|false|false|||intact
Finding|Finding|SIMPLE_SEGMENT|4539,4545|false|false|false|C1554187|Gender Status - Intact|intact
Procedure|Health Care Activity|SIMPLE_SEGMENT|4569,4578|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4579,4583|false|false|false|C0587081|Laboratory test finding|labs
Anatomy|Cell|SIMPLE_SEGMENT|4599,4602|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|4607,4610|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4607,4610|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4607,4610|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4617,4620|false|false|false|C0019046|Hemoglobin|HGB
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4617,4620|false|false|false|C0019046|Hemoglobin|HGB
Event|Event|SIMPLE_SEGMENT|4617,4620|false|false|false|||HGB
Finding|Gene or Genome|SIMPLE_SEGMENT|4617,4620|false|false|false|C1424337|CYGB gene|HGB
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4617,4620|false|false|false|C0019029|Hemoglobin concentration|HGB
Event|Event|SIMPLE_SEGMENT|4626,4629|false|false|false|||HCT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4626,4629|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4626,4629|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Disorder|Virus|SIMPLE_SEGMENT|4636,4639|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|4636,4639|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4636,4639|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4636,4639|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4636,4639|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|4644,4647|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4644,4647|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|4644,4647|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|4644,4647|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|4644,4647|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4644,4647|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4654,4658|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Drug|Antibiotic|SIMPLE_SEGMENT|4703,4708|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4703,4708|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Organic Chemical|SIMPLE_SEGMENT|4703,4708|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4713,4716|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|EOS
Event|Event|SIMPLE_SEGMENT|4713,4716|false|false|false|||EOS
Finding|Gene or Genome|SIMPLE_SEGMENT|4713,4716|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|EOS
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4746,4753|false|false|false|C0017725|glucose|GLUCOSE
Drug|Organic Chemical|SIMPLE_SEGMENT|4746,4753|false|false|false|C0017725|glucose|GLUCOSE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4746,4753|false|false|false|C0017725|glucose|GLUCOSE
Event|Event|SIMPLE_SEGMENT|4746,4753|false|false|false|||GLUCOSE
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4746,4753|false|false|false|C5781949|Glucose^1.5H post dose glucagon|GLUCOSE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4746,4753|false|false|false|C0337438|Glucose measurement|GLUCOSE
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4759,4763|false|false|false|C0041942|urea|UREA
Drug|Organic Chemical|SIMPLE_SEGMENT|4759,4763|false|false|false|C0041942|urea|UREA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4759,4763|false|false|false|C0041942|urea|UREA
Event|Event|SIMPLE_SEGMENT|4759,4763|false|false|false|||UREA
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4759,4763|false|false|false|C0523961|Urea measurement|UREA
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4780,4786|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4780,4786|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4780,4786|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Event|Event|SIMPLE_SEGMENT|4780,4786|false|false|false|||SODIUM
Finding|Physiologic Function|SIMPLE_SEGMENT|4780,4786|false|false|false|C4553025|Sodium metabolic function|SODIUM
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4780,4786|false|false|false|C0337443|Sodium measurement|SODIUM
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4792,4801|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4792,4801|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Food|SIMPLE_SEGMENT|4792,4801|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4792,4801|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4792,4801|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Event|Event|SIMPLE_SEGMENT|4792,4801|false|false|false|||POTASSIUM
Finding|Physiologic Function|SIMPLE_SEGMENT|4792,4801|false|false|false|C4553027|Potassium metabolic function|POTASSIUM
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4792,4801|false|false|false|C0202194|Potassium measurement|POTASSIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4806,4814|false|false|false|C0008203;C0596019|Chlorides;chloride ion|CHLORIDE
Event|Event|SIMPLE_SEGMENT|4806,4814|false|false|false|||CHLORIDE
Finding|Physiologic Function|SIMPLE_SEGMENT|4806,4814|false|false|false|C4553021|Chloride metabolic function|CHLORIDE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4806,4814|false|false|false|C0201952|Chloride measurement|CHLORIDE
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4825,4828|false|false|false|C0007012|carbon dioxide|CO2
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4825,4828|false|false|false|C0007012|carbon dioxide|CO2
Finding|Finding|SIMPLE_SEGMENT|4825,4828|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Finding|Gene or Genome|SIMPLE_SEGMENT|4825,4828|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4832,4837|false|false|false|C0003075|Anions|ANION
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4832,4841|false|false|false|C0003074|Anion Gap|ANION GAP
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4832,4841|false|false|false|C1509129|Anion gap result|ANION GAP
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4832,4841|false|false|false|C0201889;C2189246|Anion gap measurement;blood anion gap (lab test)|ANION GAP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4838,4841|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4838,4841|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Event|Event|SIMPLE_SEGMENT|4838,4841|false|false|false|||GAP
Finding|Gene or Genome|SIMPLE_SEGMENT|4838,4841|false|false|false|C1419277;C2984552|RASA1 gene;RASA1 wt Allele|GAP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4863,4866|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|SIMPLE_SEGMENT|4863,4866|false|false|false|||PTT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4863,4866|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4921,4924|false|false|false|C0010287|Creatine Kinase|CPK
Drug|Enzyme|SIMPLE_SEGMENT|4921,4924|false|false|false|C0010287|Creatine Kinase|CPK
Event|Event|SIMPLE_SEGMENT|4921,4924|false|false|false|||CPK
Finding|Gene or Genome|SIMPLE_SEGMENT|4921,4924|false|false|false|C1418571|PIK3C2A gene|CPK
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4921,4924|false|false|false|C0201973|Creatine kinase measurement|CPK
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4943,4950|false|false|false|C0060323|Fibrin fragment D|D-DIMER
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4943,4950|false|false|false|C0060323|Fibrin fragment D|D-DIMER
Drug|Chemical Viewed Structurally|SIMPLE_SEGMENT|4945,4950|false|false|false|C0596448|dimer|DIMER
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4968,4972|false|false|false|C0587081|Laboratory test finding|labs
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4986,4991|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4986,4991|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4986,4991|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5018,5023|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5018,5023|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5018,5023|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5024,5029|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|SIMPLE_SEGMENT|5024,5029|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|SIMPLE_SEGMENT|5024,5029|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5024,5029|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Drug|Organic Chemical|SIMPLE_SEGMENT|5027,5031|false|false|false|C0602254|MB 3|MB-3
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5058,5063|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5058,5063|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5058,5063|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5064,5069|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|SIMPLE_SEGMENT|5064,5069|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|SIMPLE_SEGMENT|5064,5069|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5064,5069|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Drug|Organic Chemical|SIMPLE_SEGMENT|5067,5071|false|false|false|C0602254|MB 3|MB-3
Event|Event|SIMPLE_SEGMENT|5087,5094|false|false|false|||Imaging
Finding|Finding|SIMPLE_SEGMENT|5087,5094|false|false|false|C0740845|Imaging problem|Imaging
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5087,5094|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|Imaging
Event|Event|SIMPLE_SEGMENT|5095,5102|false|false|false|||studies
Procedure|Research Activity|SIMPLE_SEGMENT|5095,5102|false|false|false|C0947630|Scientific Study|studies
Event|Event|SIMPLE_SEGMENT|5104,5107|false|false|false|||EKG
Finding|Intellectual Product|SIMPLE_SEGMENT|5104,5107|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5104,5107|false|false|false|C1623258|Electrocardiography|EKG
Event|Event|SIMPLE_SEGMENT|5111,5120|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|5111,5120|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5122,5127|false|false|false|C0030471;C1305231|Nasal sinus;Sinus - general anatomical term|Sinus
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|5122,5127|false|false|false|C0016169|pathologic fistula|Sinus
Drug|Organic Chemical|SIMPLE_SEGMENT|5122,5127|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|Sinus
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5122,5127|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|Sinus
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5122,5139|false|false|false|C0039239|Sinus Tachycardia|Sinus tachycardia
Finding|Finding|SIMPLE_SEGMENT|5122,5139|false|false|false|C2108109;C5235163|Sinus Tachycardia by ECG Finding;continuous electrocardiogram sinus tachycardia|Sinus tachycardia
Event|Event|SIMPLE_SEGMENT|5128,5139|false|false|false|||tachycardia
Finding|Finding|SIMPLE_SEGMENT|5128,5139|false|false|false|C0039231;C3827868|Tachycardia;Tachycardia by ECG Finding|tachycardia
Finding|Finding|SIMPLE_SEGMENT|5151,5161|false|false|false|C0429029|ST segment|ST segment
Event|Event|SIMPLE_SEGMENT|5163,5170|false|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|5163,5170|false|false|false|C0392747|Changing|changes
Event|Event|SIMPLE_SEGMENT|5185,5193|false|false|false|||ischemia
Finding|Pathologic Function|SIMPLE_SEGMENT|5185,5193|false|true|false|C0022116|Ischemia|ischemia
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5185,5193|false|true|false|C4321499|Ischemia Procedure|ischemia
Event|Event|SIMPLE_SEGMENT|5220,5227|false|false|false|||tracing
Event|Event|SIMPLE_SEGMENT|5232,5238|false|false|false|||change
Finding|Functional Concept|SIMPLE_SEGMENT|5232,5238|true|false|false|C0392747|Changing|change
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5232,5238|true|false|false|C4319952|Change - procedure|change
Event|Event|SIMPLE_SEGMENT|5243,5246|false|false|false|||CXR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5243,5246|false|false|false|C0039985|Plain chest X-ray|CXR
Finding|Finding|SIMPLE_SEGMENT|5252,5255|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|New
Finding|Idea or Concept|SIMPLE_SEGMENT|5252,5255|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|New
Finding|Finding|SIMPLE_SEGMENT|5256,5264|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|SIMPLE_SEGMENT|5256,5264|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Functional Concept|SIMPLE_SEGMENT|5265,5269|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Tissue|SIMPLE_SEGMENT|5270,5277|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5270,5277|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Body Substance|SIMPLE_SEGMENT|5270,5286|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Finding|Finding|SIMPLE_SEGMENT|5270,5286|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|5270,5286|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Event|Event|SIMPLE_SEGMENT|5278,5286|false|false|false|||effusion
Finding|Body Substance|SIMPLE_SEGMENT|5278,5286|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|SIMPLE_SEGMENT|5278,5286|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|5278,5286|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Event|Event|SIMPLE_SEGMENT|5302,5313|false|false|false|||atelectasis
Finding|Pathologic Function|SIMPLE_SEGMENT|5302,5313|false|false|false|C0004144|Atelectasis|atelectasis
Finding|Functional Concept|SIMPLE_SEGMENT|5321,5325|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5321,5330|false|false|false|C0225730|Left lung|left lung
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5321,5335|false|false|false|C0225732|Structure of base of left lung|left lung base
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5326,5330|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5326,5330|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5326,5330|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|SIMPLE_SEGMENT|5326,5330|false|false|false|C0740941|Lung Problem|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5326,5335|false|false|false|C0225704|Basal segment of lung|lung base
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5331,5335|false|false|false|C2987514|Anatomical base|base
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5331,5335|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Chemical Viewed Functionally|SIMPLE_SEGMENT|5331,5335|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|5331,5335|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Finding|Gene or Genome|SIMPLE_SEGMENT|5331,5335|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Finding|Idea or Concept|SIMPLE_SEGMENT|5331,5335|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5341,5344|false|false|false|C3813556|Cancer/Testis Antigen|CTA
Event|Event|SIMPLE_SEGMENT|5341,5344|false|false|false|||CTA
Finding|Gene or Genome|SIMPLE_SEGMENT|5341,5344|false|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5341,5344|false|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5345,5350|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|SIMPLE_SEGMENT|5345,5350|false|false|false|C0741025|Chest problem|Chest
Event|Event|SIMPLE_SEGMENT|5363,5371|false|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|5363,5371|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|5363,5375|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence for
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5376,5385|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5376,5385|true|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|5376,5385|true|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|SIMPLE_SEGMENT|5376,5393|true|false|false|C0034065|Pulmonary Embolism|pulmonary embolus
Event|Event|SIMPLE_SEGMENT|5386,5393|false|false|false|||embolus
Finding|Finding|SIMPLE_SEGMENT|5386,5393|true|false|false|C1704212;C2046122|Embolus|embolus
Finding|Functional Concept|SIMPLE_SEGMENT|5406,5410|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Tissue|SIMPLE_SEGMENT|5411,5418|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5411,5418|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Body Substance|SIMPLE_SEGMENT|5411,5427|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Finding|Finding|SIMPLE_SEGMENT|5411,5427|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|5411,5427|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Event|Event|SIMPLE_SEGMENT|5419,5427|false|false|false|||effusion
Finding|Body Substance|SIMPLE_SEGMENT|5419,5427|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|SIMPLE_SEGMENT|5419,5427|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|5419,5427|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Event|Event|SIMPLE_SEGMENT|5442,5453|false|false|false|||atelectasis
Finding|Pathologic Function|SIMPLE_SEGMENT|5442,5453|false|false|false|C0004144|Atelectasis|atelectasis
Finding|Finding|SIMPLE_SEGMENT|5461,5469|false|false|false|C0332149|Possible|Possible
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5480,5487|false|false|false|C0037993|Spleen|splenic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5480,5494|false|false|false|C0037996;C4482214|Abdomen>Splenic artery;Structure of splenic artery|splenic artery
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5480,5503|false|true|false|C0155747|Aneurysm of splenic artery|splenic artery aneurysm
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5488,5494|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|SIMPLE_SEGMENT|5488,5494|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Event|Event|SIMPLE_SEGMENT|5495,5503|false|false|false|||aneurysm
Finding|Pathologic Function|SIMPLE_SEGMENT|5495,5503|false|false|false|C0002940|Aneurysm|aneurysm
Drug|Amino Acid Sequence|SIMPLE_SEGMENT|5511,5517|false|false|false|C1514562|Protein Domain|region
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5526,5531|false|false|false|C0929176|Hilum|hilum
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5535,5542|false|false|false|C0018787|Heart|Cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|5535,5542|false|false|false|C1314974|Cardiac attachment|Cardiac
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|5535,5558|false|false|false|C0261588|Cardiac catheterisation as the cause of abnormal reaction of the patient, or of later complication, without mention of misadventure at the time of the procedure|Cardiac catheterization
Finding|Intellectual Product|SIMPLE_SEGMENT|5535,5558|false|false|false|C1547981|Diagnostic Service Section ID - Cardiac Catheterization|Cardiac catheterization
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5535,5558|false|false|false|C0018795;C1548828|Cardiac Catheterization Procedures;Consent Type - Cardiac Catheterization|Cardiac catheterization
Procedure|Health Care Activity|SIMPLE_SEGMENT|5535,5558|false|false|false|C0018795;C1548828|Cardiac Catheterization Procedures;Consent Type - Cardiac Catheterization|Cardiac catheterization
Event|Event|SIMPLE_SEGMENT|5543,5558|false|false|false|||catheterization
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5543,5558|false|false|false|C0007430|Catheterization|catheterization
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5574,5582|false|false|false|C0018787|Heart|coronary
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5574,5594|false|false|false|C0085532;C1548829|Consent Type - Coronary Angiography;Coronary angiography|coronary angiography
Procedure|Health Care Activity|SIMPLE_SEGMENT|5574,5594|false|false|false|C0085532;C1548829|Consent Type - Coronary Angiography;Coronary angiography|coronary angiography
Event|Event|SIMPLE_SEGMENT|5583,5594|false|false|false|||angiography
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5583,5594|false|false|false|C0002978|angiogram|angiography
Finding|Functional Concept|SIMPLE_SEGMENT|5603,5608|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Finding|Functional Concept|SIMPLE_SEGMENT|5609,5617|false|false|false|C1527180|Dominant|dominant
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5618,5624|false|false|false|C5671121|System (basic dose form)|system
Event|Event|SIMPLE_SEGMENT|5618,5624|false|false|false|||system
Finding|Functional Concept|SIMPLE_SEGMENT|5618,5624|false|false|false|C0449913;C5441654|System;System, LOINC Axis 4|system
Event|Event|SIMPLE_SEGMENT|5626,5638|false|false|false|||demonstrated
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5641,5647|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5641,5647|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5641,5656|false|false|false|C0010075|Coronary Vessels|vessel coronary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5648,5656|false|false|false|C0018787|Heart|coronary
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5648,5664|false|false|false|C0010068;C1956346|Coronary Artery Disease;Coronary heart disease|coronary disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5657,5664|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|5657,5664|false|false|false|||disease
Finding|Functional Concept|SIMPLE_SEGMENT|5672,5678|false|false|false|C0302891|Native (qualifier value)|native
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5679,5686|false|false|false|C0005847|Blood Vessel|vessels
Finding|Idea or Concept|SIMPLE_SEGMENT|5723,5731|false|false|false|C0750489|apparent|apparent
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5732,5739|true|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|5732,5739|false|false|false|||disease
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5746,5749|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5746,5749|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|SIMPLE_SEGMENT|5746,5749|false|false|false|||LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|5746,5749|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Event|Event|SIMPLE_SEGMENT|5761,5767|false|false|false|||lesion
Finding|Finding|SIMPLE_SEGMENT|5761,5767|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|SIMPLE_SEGMENT|5761,5767|false|false|false|C0221198;C1546698|Lesion|lesion
Event|Event|SIMPLE_SEGMENT|5780,5785|false|false|false|||stent
Event|Event|SIMPLE_SEGMENT|5819,5824|false|false|false|||small
Finding|Intellectual Product|SIMPLE_SEGMENT|5833,5837|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|poor
Event|Event|SIMPLE_SEGMENT|5839,5843|false|false|false|||flow
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|5839,5843|false|false|false|C0806140|Flow|flow
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5850,5853|false|false|false|C2987138|Methylcytosine Dioxygenase TET1|LCx
Drug|Enzyme|SIMPLE_SEGMENT|5850,5853|false|false|false|C2987138|Methylcytosine Dioxygenase TET1|LCx
Finding|Gene or Genome|SIMPLE_SEGMENT|5850,5853|false|false|false|C1428863;C2987137|TET1 gene;TET1 wt Allele|LCx
Event|Event|SIMPLE_SEGMENT|5867,5875|false|false|false|||stenosis
Finding|Pathologic Function|SIMPLE_SEGMENT|5867,5875|false|false|false|C1261287|Stenosis|stenosis
Event|Event|SIMPLE_SEGMENT|5883,5889|false|false|false|||origin
Finding|Classification|SIMPLE_SEGMENT|5883,5889|false|false|false|C0079946;C1550512|National origin;Participation Type - origin|origin
Finding|Intellectual Product|SIMPLE_SEGMENT|5883,5889|false|false|false|C0079946;C1550512|National origin;Participation Type - origin|origin
Finding|Idea or Concept|SIMPLE_SEGMENT|5925,5933|false|false|false|C0750489|apparent|apparent
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5934,5941|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|5934,5941|false|false|false|||disease
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5947,5955|false|false|false|C0003842|Arteries|Arterial
Event|Event|SIMPLE_SEGMENT|5964,5975|false|false|false|||angiography
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5964,5975|false|false|false|C0002978|angiogram|angiography
Event|Event|SIMPLE_SEGMENT|5976,5988|false|false|false|||demonstrated
Anatomy|Tissue|SIMPLE_SEGMENT|5998,6003|false|false|false|C0332835|Transplanted tissue|graft
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5998,6003|false|false|false|C0181074;C1705210|Graft Dosage Form;Graft material|graft
Event|Event|SIMPLE_SEGMENT|5998,6003|false|false|false|||graft
Finding|Intellectual Product|SIMPLE_SEGMENT|5998,6003|false|false|false|C1546653|Graft - Specimen Source Codes|graft
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5998,6003|false|false|false|C1961139;C3683798|Graft Procedures on the Head;Grafting procedure|graft
Event|Event|SIMPLE_SEGMENT|6012,6018|false|false|false|||patent
Finding|Intellectual Product|SIMPLE_SEGMENT|6012,6018|false|false|false|C0030650|Legal patent|patent
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6024,6030|false|false|false|C0042449|Veins|Venous
Event|Event|SIMPLE_SEGMENT|6039,6050|false|false|false|||angiography
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6039,6050|false|false|false|C0002978|angiogram|angiography
Event|Event|SIMPLE_SEGMENT|6051,6063|false|false|false|||demonstrated
Finding|Intellectual Product|SIMPLE_SEGMENT|6066,6072|false|false|false|C0030650|Legal patent|patent
Event|Event|SIMPLE_SEGMENT|6073,6076|false|false|false|||SVG
Event|Event|SIMPLE_SEGMENT|6101,6109|false|false|false|||stenosis
Finding|Pathologic Function|SIMPLE_SEGMENT|6101,6109|false|false|false|C1261287|Stenosis|stenosis
Event|Event|SIMPLE_SEGMENT|6110,6119|false|false|false|||involving
Event|Event|SIMPLE_SEGMENT|6128,6138|false|false|false|||sub-branch
Event|Event|SIMPLE_SEGMENT|6170,6178|false|false|false|||diagonal
Event|Event|SIMPLE_SEGMENT|6183,6191|false|false|false|||presumed
Event|Event|SIMPLE_SEGMENT|6192,6200|false|false|false|||occluded
Finding|Finding|SIMPLE_SEGMENT|6192,6200|false|false|false|C0028778;C1947917|Obstruction;Occluded|occluded
Finding|Functional Concept|SIMPLE_SEGMENT|6192,6200|false|false|false|C0028778;C1947917|Obstruction;Occluded|occluded
Event|Event|SIMPLE_SEGMENT|6205,6211|false|false|false|||unable
Finding|Finding|SIMPLE_SEGMENT|6205,6211|false|false|false|C1299582|Unable|unable
Event|Event|SIMPLE_SEGMENT|6219,6229|false|false|false|||identified
Finding|Functional Concept|SIMPLE_SEGMENT|6235,6242|false|false|false|C0439801;C3542948|Limited (extensiveness);Limited component (foundation metadata concept)|Limited
Finding|Intellectual Product|SIMPLE_SEGMENT|6235,6242|false|false|false|C0439801;C3542948|Limited (extensiveness);Limited component (foundation metadata concept)|Limited
Event|Event|SIMPLE_SEGMENT|6251,6263|false|false|false|||hemodynamics
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|6251,6263|false|false|false|C0019010|Hemodynamics|hemodynamics
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6251,6263|false|false|false|C4281788|hemodynamics (procedure)|hemodynamics
Event|Event|SIMPLE_SEGMENT|6264,6272|false|false|false|||revealed
Finding|Functional Concept|SIMPLE_SEGMENT|6273,6281|false|false|false|C0205373;C5849094|Systemic;Systemic Route of Administration|systemic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6273,6294|false|false|false|C0020538|Hypertensive disease|systemic hypertension
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6282,6294|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|SIMPLE_SEGMENT|6282,6294|false|false|false|||hypertension
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6302,6308|false|false|false|C0003483|Aorta|aortic
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6302,6317|false|false|false|C0456180|Aortic Pressure|aortic pressure
Event|Event|SIMPLE_SEGMENT|6309,6317|false|false|false|||pressure
Finding|Finding|SIMPLE_SEGMENT|6309,6317|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|SIMPLE_SEGMENT|6309,6317|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|6309,6317|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|6309,6317|false|false|false|C0033095||pressure
Finding|Idea or Concept|SIMPLE_SEGMENT|6339,6344|false|false|false|C1546485|Diagnosis Type - Final|FINAL
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6345,6354|false|false|false|C0945731||DIAGNOSIS
Event|Event|SIMPLE_SEGMENT|6345,6354|false|false|false|||DIAGNOSIS
Finding|Classification|SIMPLE_SEGMENT|6345,6354|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|DIAGNOSIS
Finding|Functional Concept|SIMPLE_SEGMENT|6345,6354|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|DIAGNOSIS
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6345,6354|false|false|false|C0011900|Diagnosis|DIAGNOSIS
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6368,6374|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6368,6374|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6368,6383|false|false|false|C0010075|Coronary Vessels|vessel coronary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6375,6383|false|false|false|C0018787|Heart|coronary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6375,6390|false|false|false|C0205042|Coronary artery|coronary artery
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6375,6398|false|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|coronary artery disease
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6384,6390|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|SIMPLE_SEGMENT|6384,6390|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6384,6398|false|false|false|C0852949|Arteriopathic disease|artery disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6391,6398|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|6391,6398|false|false|false|||disease
Finding|Functional Concept|SIMPLE_SEGMENT|6406,6412|false|false|false|C0302891|Native (qualifier value)|native
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6413,6421|false|false|false|C0003842;C0226004|Arterial system;Arteries|arteries
Anatomy|Body System|SIMPLE_SEGMENT|6413,6421|false|false|false|C0003842;C0226004|Arterial system;Arteries|arteries
Procedure|Health Care Activity|SIMPLE_SEGMENT|6413,6421|false|false|false|C0397581|Procedure on artery|arteries
Finding|Intellectual Product|SIMPLE_SEGMENT|6426,6432|false|false|false|C0030650|Legal patent|Patent
Event|Event|SIMPLE_SEGMENT|6433,6437|false|false|false|||LIMA
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6441,6444|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6441,6444|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|SIMPLE_SEGMENT|6441,6444|false|false|false|||LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|6441,6444|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Finding|Intellectual Product|SIMPLE_SEGMENT|6446,6452|false|false|false|C0030650|Legal patent|patent
Event|Event|SIMPLE_SEGMENT|6453,6456|false|false|false|||SVG
Finding|Finding|SIMPLE_SEGMENT|6464,6472|false|false|false|C0028778;C1947917|Obstruction;Occluded|occluded
Finding|Functional Concept|SIMPLE_SEGMENT|6464,6472|false|false|false|C0028778;C1947917|Obstruction;Occluded|occluded
Event|Event|SIMPLE_SEGMENT|6473,6476|false|false|false|||SVG
Drug|Chemical Viewed Structurally|SIMPLE_SEGMENT|6497,6503|false|false|false|C1881507|Macromolecular Branch|branch
Event|Event|SIMPLE_SEGMENT|6497,6503|false|false|false|||branch
Finding|Intellectual Product|SIMPLE_SEGMENT|6509,6514|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|Brief
Finding|Idea or Concept|SIMPLE_SEGMENT|6515,6523|false|false|false|C1547192|Organization unit type - Hospital|Hospital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6515,6530|false|false|false|C0488549||Hospital Course
Finding|Finding|SIMPLE_SEGMENT|6515,6530|false|false|false|C0489547|Hospital course|Hospital Course
Finding|Idea or Concept|SIMPLE_SEGMENT|6536,6540|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|SIMPLE_SEGMENT|6536,6540|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Event|Event|SIMPLE_SEGMENT|6541,6544|false|false|false|||old
Event|Event|SIMPLE_SEGMENT|6559,6566|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|6559,6566|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|6559,6566|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|6559,6566|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|6559,6569|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6570,6573|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6570,6573|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|6570,6573|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|6570,6573|false|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|6570,6573|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6570,6573|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|6570,6573|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6570,6573|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6578,6581|false|false|false|C2713669|SERPINA5 protein, human|PCI
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6578,6581|false|false|false|C2713669|SERPINA5 protein, human|PCI
Event|Event|SIMPLE_SEGMENT|6578,6581|false|false|false|||PCI
Finding|Gene or Genome|SIMPLE_SEGMENT|6578,6581|false|false|false|C1418370;C1705930;C4049621|Peritoneal Cancer Index;SERPINA5 gene;SERPINA5 wt Allele|PCI
Finding|Intellectual Product|SIMPLE_SEGMENT|6578,6581|false|false|false|C1418370;C1705930;C4049621|Peritoneal Cancer Index;SERPINA5 gene;SERPINA5 wt Allele|PCI
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6578,6581|false|false|false|C1514496;C1532338;C4724254|Percutaneous Coronary Intervention;Prophylactic Cranial Irradiation;photochemical internalization|PCI
Event|Event|SIMPLE_SEGMENT|6582,6584|false|false|false|||x3
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6590,6594|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Event|Event|SIMPLE_SEGMENT|6595,6597|false|false|false|||x3
Event|Event|SIMPLE_SEGMENT|6606,6610|false|false|false|||type
Finding|Gene or Genome|SIMPLE_SEGMENT|6606,6610|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Finding|Intellectual Product|SIMPLE_SEGMENT|6606,6610|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Finding|Classification|SIMPLE_SEGMENT|6606,6612|false|false|false|C0441730|Type 2|type 2
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6619,6626|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|SIMPLE_SEGMENT|6619,6626|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6619,6626|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|SIMPLE_SEGMENT|6619,6626|false|false|false|||insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|6619,6626|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6619,6626|false|false|false|C0202098|Insulin measurement|insulin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6628,6631|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|SIMPLE_SEGMENT|6628,6631|false|false|false|||HTN
Event|Event|SIMPLE_SEGMENT|6637,6640|false|false|false|||HLD
Event|Event|SIMPLE_SEGMENT|6645,6654|false|false|false|||presented
Finding|Idea or Concept|SIMPLE_SEGMENT|6665,6668|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|6665,6668|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|6669,6676|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|6669,6676|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|6669,6676|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|6669,6676|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|6669,6679|false|false|false|C0262926|Medical History|history of
Finding|Functional Concept|SIMPLE_SEGMENT|6680,6684|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Finding|Sign or Symptom|SIMPLE_SEGMENT|6680,6701|false|false|false|C0541828|Left sided chest pain|left sided chest pain
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6691,6696|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|6691,6696|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6691,6701|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|6691,6701|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6697,6701|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|6697,6701|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|6697,6701|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|6697,6701|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|6706,6709|false|false|false|||SOB
Finding|Sign or Symptom|SIMPLE_SEGMENT|6706,6709|false|false|false|C0013404|Dyspnea|SOB
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6716,6721|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|SIMPLE_SEGMENT|6716,6721|false|false|false|C0741025|Chest problem|Chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6716,6726|false|false|false|C2926613||Chest Pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|6716,6726|false|false|false|C0008031|Chest Pain|Chest Pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6722,6726|false|false|false|C2598155||Pain
Event|Event|SIMPLE_SEGMENT|6722,6726|false|false|false|||Pain
Finding|Functional Concept|SIMPLE_SEGMENT|6722,6726|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|6722,6726|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Body Substance|SIMPLE_SEGMENT|6728,6735|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|6728,6735|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|6728,6735|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|6741,6752|false|false|false|C0750502|Significant|significant
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6753,6756|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6753,6756|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|6753,6756|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|6753,6756|false|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|6753,6756|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6753,6756|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|6753,6756|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6753,6756|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Event|Event|SIMPLE_SEGMENT|6757,6764|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|6757,6764|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|6757,6764|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|6757,6764|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Event|Event|SIMPLE_SEGMENT|6778,6782|false|false|false|||CABG
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6778,6782|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Event|Event|SIMPLE_SEGMENT|6784,6794|false|false|false|||presenting
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6800,6805|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|6800,6805|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6800,6810|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|6800,6810|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6806,6810|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|6806,6810|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|6806,6810|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|6806,6810|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6822,6831|false|false|false|C0041199|Troponin|troponins
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6822,6831|false|false|false|C0041199|Troponin|troponins
Event|Event|SIMPLE_SEGMENT|6822,6831|false|false|false|||troponins
Finding|Finding|SIMPLE_SEGMENT|6838,6841|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|6838,6841|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|6846,6857|false|false|false|C0011570|Mental Depression|depressions
Event|Event|SIMPLE_SEGMENT|6846,6857|false|false|false|||depressions
Event|Event|SIMPLE_SEGMENT|6879,6889|false|false|false|||consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|6879,6889|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|6879,6894|false|false|false|C0332290|Consistent with|consistent with
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6895,6901|false|false|false|C4255010||NSTEMI
Event|Event|SIMPLE_SEGMENT|6895,6901|false|false|false|||NSTEMI
Finding|Finding|SIMPLE_SEGMENT|6895,6901|false|false|false|C3537184||NSTEMI
Finding|Body Substance|SIMPLE_SEGMENT|6905,6912|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|6905,6912|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|6905,6912|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6915,6924|false|false|false|C0041199|Troponin|troponins
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6915,6924|false|false|false|C0041199|Troponin|troponins
Event|Event|SIMPLE_SEGMENT|6915,6924|false|false|false|||troponins
Event|Event|SIMPLE_SEGMENT|6925,6934|false|false|false|||plateaued
Event|Event|SIMPLE_SEGMENT|6953,6962|false|false|false|||initiated
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6969,6976|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Organic Chemical|SIMPLE_SEGMENT|6969,6976|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6969,6976|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Event|Event|SIMPLE_SEGMENT|6969,6976|false|false|false|||heparin
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6977,6980|false|false|false|C1135868|Gestational Trophoblastic Neoplasms|gtt
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6977,6980|false|false|false|C0991568|Drops - Drug Form|gtt
Event|Event|SIMPLE_SEGMENT|6977,6980|false|false|false|||gtt
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6977,6980|false|false|false|C0017741|Glucose tolerance test|gtt
Event|Event|SIMPLE_SEGMENT|7000,7005|false|false|false|||taken
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7009,7016|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|7009,7016|false|false|false|C1314974|Cardiac attachment|cardiac
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7009,7021|false|false|false|C0018795|Cardiac Catheterization Procedures|cardiac cath
Event|Event|SIMPLE_SEGMENT|7017,7021|false|false|false|||cath
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7017,7021|false|false|false|C0007430|Catheterization|cath
Event|Event|SIMPLE_SEGMENT|7047,7062|false|false|false|||Catheterization
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7047,7062|false|false|false|C0007430|Catheterization|Catheterization
Event|Event|SIMPLE_SEGMENT|7063,7069|false|false|false|||showed
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|7070,7079|false|false|false|C0001168|Complete obstruction|occlusion
Event|Event|SIMPLE_SEGMENT|7070,7079|false|false|false|||occlusion
Finding|Finding|SIMPLE_SEGMENT|7070,7079|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Functional Concept|SIMPLE_SEGMENT|7070,7079|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|7070,7079|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Pathologic Function|SIMPLE_SEGMENT|7070,7079|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Event|Event|SIMPLE_SEGMENT|7087,7090|false|false|false|||SVG
Finding|Finding|SIMPLE_SEGMENT|7109,7117|false|false|false|C0332149|Possible|possibly
Event|Event|SIMPLE_SEGMENT|7118,7125|false|false|false|||causing
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|7130,7137|false|false|false|C1705970|Electrical Current|current
Event|Event|SIMPLE_SEGMENT|7138,7146|false|false|false|||symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|7138,7146|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|7138,7146|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|SIMPLE_SEGMENT|7153,7165|false|false|false|||intervention
Procedure|Health Care Activity|SIMPLE_SEGMENT|7153,7165|false|false|false|C0184661;C0886296;C1273869|Intervention regimes;Interventional procedure;Nursing interventions|intervention
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7153,7165|false|false|false|C0184661;C0886296;C1273869|Intervention regimes;Interventional procedure;Nursing interventions|intervention
Finding|Body Substance|SIMPLE_SEGMENT|7182,7189|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|7182,7189|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|7182,7189|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|7204,7213|false|false|false|||optimized
Drug|Organic Chemical|SIMPLE_SEGMENT|7230,7240|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7230,7240|false|false|false|C0025859|metoprolol|metoprolol
Event|Event|SIMPLE_SEGMENT|7230,7240|false|false|false|||metoprolol
Event|Event|SIMPLE_SEGMENT|7242,7252|false|false|false|||initiation
Finding|Functional Concept|SIMPLE_SEGMENT|7242,7252|false|false|false|C0589507;C1158830;C1704686|Initiation;Transcription Initiation|initiation
Finding|Genetic Function|SIMPLE_SEGMENT|7242,7252|false|false|false|C0589507;C1158830;C1704686|Initiation;Transcription Initiation|initiation
Finding|Mental Process|SIMPLE_SEGMENT|7242,7252|false|false|false|C0589507;C1158830;C1704686|Initiation;Transcription Initiation|initiation
Drug|Organic Chemical|SIMPLE_SEGMENT|7256,7264|false|false|false|C0126174|losartan|losartan
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7256,7264|false|false|false|C0126174|losartan|losartan
Event|Event|SIMPLE_SEGMENT|7256,7264|false|false|false|||losartan
Event|Event|SIMPLE_SEGMENT|7271,7281|false|false|false|||initiation
Finding|Functional Concept|SIMPLE_SEGMENT|7271,7281|false|false|false|C0589507;C1158830;C1704686|Initiation;Transcription Initiation|initiation
Finding|Genetic Function|SIMPLE_SEGMENT|7271,7281|false|false|false|C0589507;C1158830;C1704686|Initiation;Transcription Initiation|initiation
Finding|Mental Process|SIMPLE_SEGMENT|7271,7281|false|false|false|C0589507;C1158830;C1704686|Initiation;Transcription Initiation|initiation
Drug|Organic Chemical|SIMPLE_SEGMENT|7285,7290|false|false|false|C0590690|Imdur|imdur
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7285,7290|false|false|false|C0590690|Imdur|imdur
Event|Event|SIMPLE_SEGMENT|7285,7290|false|false|false|||imdur
Event|Event|SIMPLE_SEGMENT|7309,7315|false|false|false|||causes
Finding|Functional Concept|SIMPLE_SEGMENT|7309,7315|false|false|false|C0015127;C1314792|Etiology;Etiology aspects|causes
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7323,7328|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|7323,7328|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7323,7333|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|7323,7333|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7329,7333|false|true|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|7329,7333|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|7329,7333|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|7329,7333|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|7340,7350|false|false|false|||considered
Finding|Classification|SIMPLE_SEGMENT|7380,7388|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|7380,7388|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|7380,7388|false|false|false|C5237010|Expression Negative|negative
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7389,7392|false|false|false|C3813556|Cancer/Testis Antigen|CTA
Event|Event|SIMPLE_SEGMENT|7389,7392|false|false|false|||CTA
Finding|Gene or Genome|SIMPLE_SEGMENT|7389,7392|false|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7389,7392|false|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7396,7408|false|false|false|C0031046|Pericarditis|pericarditis
Event|Event|SIMPLE_SEGMENT|7396,7408|false|false|false|||pericarditis
Event|Event|SIMPLE_SEGMENT|7410,7418|false|false|false|||symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|7410,7418|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|7410,7418|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|SIMPLE_SEGMENT|7419,7429|false|false|false|||consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|7419,7429|false|false|false|C0332290|Consistent with|consistent
Event|Event|SIMPLE_SEGMENT|7435,7439|false|false|false|||exam
Finding|Functional Concept|SIMPLE_SEGMENT|7435,7439|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|7435,7439|false|false|false|C0582103|Medical Examination|exam
Event|Event|SIMPLE_SEGMENT|7444,7447|false|false|false|||EKG
Finding|Intellectual Product|SIMPLE_SEGMENT|7444,7447|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7444,7447|false|false|false|C1623258|Electrocardiography|EKG
Event|Event|SIMPLE_SEGMENT|7453,7463|false|false|false|||consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|7453,7463|false|false|false|C0332290|Consistent with|consistent
Finding|Body Substance|SIMPLE_SEGMENT|7470,7477|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|7470,7477|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|7470,7477|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|SIMPLE_SEGMENT|7470,7481|false|false|false|C0332310|Has patient|patient has
Event|Event|SIMPLE_SEGMENT|7499,7506|false|false|false|||treated
Finding|Idea or Concept|SIMPLE_SEGMENT|7531,7541|false|false|false|C0332290|Consistent with|consistent
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7542,7548|false|false|false|C0003211;C0358845|Analgesics and non-steroidal anti-inflammatory drugs;Anti-Inflammatory Agents, Non-Steroidal|NSAIDs
Event|Event|SIMPLE_SEGMENT|7542,7548|false|false|false|||NSAIDs
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7551,7566|false|false|false|C0040213;C5779793|Costal chondritis;Tietze's Syndrome|costochondritis
Event|Event|SIMPLE_SEGMENT|7551,7566|false|false|false|||costochondritis
Event|Event|SIMPLE_SEGMENT|7568,7576|false|false|false|||symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|7568,7576|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|7568,7576|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|SIMPLE_SEGMENT|7593,7605|false|false|false|||reproducible
Event|Event|SIMPLE_SEGMENT|7609,7613|false|false|false|||exam
Finding|Functional Concept|SIMPLE_SEGMENT|7609,7613|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|7609,7613|false|false|false|C0582103|Medical Examination|exam
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7619,7628|false|false|false|C0032231|Pleurisy|pleuritis
Event|Event|SIMPLE_SEGMENT|7619,7628|false|false|false|||pleuritis
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7629,7638|false|false|false|C0027627|Neoplasm Metastasis|secondary
Event|Event|SIMPLE_SEGMENT|7629,7638|false|false|false|||secondary
Finding|Functional Concept|SIMPLE_SEGMENT|7629,7638|false|false|false|C1522484|metastatic qualifier|secondary
Anatomy|Tissue|SIMPLE_SEGMENT|7643,7650|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7643,7650|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Body Substance|SIMPLE_SEGMENT|7643,7659|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Finding|Finding|SIMPLE_SEGMENT|7643,7659|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|7643,7659|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Event|Event|SIMPLE_SEGMENT|7651,7659|false|false|false|||effusion
Finding|Body Substance|SIMPLE_SEGMENT|7651,7659|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|SIMPLE_SEGMENT|7651,7659|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|7651,7659|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Event|Event|SIMPLE_SEGMENT|7672,7680|false|false|false|||effusion
Finding|Body Substance|SIMPLE_SEGMENT|7672,7680|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|SIMPLE_SEGMENT|7672,7680|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|7672,7680|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Event|Event|SIMPLE_SEGMENT|7682,7688|false|false|false|||stable
Finding|Intellectual Product|SIMPLE_SEGMENT|7682,7688|false|false|false|C1547311|Patient Condition Code - Stable|stable
Event|Event|SIMPLE_SEGMENT|7695,7699|false|false|false|||CABG
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7695,7699|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7710,7714|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|7710,7714|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|7710,7714|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|7710,7714|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|7715,7723|false|false|false|||persists
Finding|Body Substance|SIMPLE_SEGMENT|7725,7732|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|7725,7732|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|7725,7732|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|7737,7747|false|false|false|||instructed
Event|Event|SIMPLE_SEGMENT|7751,7756|false|false|false|||speak
Event|Event|SIMPLE_SEGMENT|7767,7779|false|false|false|||cardiologist
Drug|Organic Chemical|SIMPLE_SEGMENT|7797,7802|false|false|false|C0590690|Imdur|imdur
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7797,7802|false|false|false|C0590690|Imdur|imdur
Event|Event|SIMPLE_SEGMENT|7797,7802|false|false|false|||imdur
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7814,7819|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|7814,7819|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|7814,7819|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Finding|SIMPLE_SEGMENT|7814,7828|false|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|blood pressure
Finding|Organism Function|SIMPLE_SEGMENT|7814,7828|false|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|blood pressure
Procedure|Health Care Activity|SIMPLE_SEGMENT|7814,7828|false|false|false|C0005824|Blood pressure determination|blood pressure
Event|Event|SIMPLE_SEGMENT|7820,7828|false|false|false|||pressure
Finding|Finding|SIMPLE_SEGMENT|7820,7828|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|SIMPLE_SEGMENT|7820,7828|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|7820,7828|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|7820,7828|false|false|false|C0033095||pressure
Event|Event|SIMPLE_SEGMENT|7830,7838|false|false|false|||tolerate
Finding|Intellectual Product|SIMPLE_SEGMENT|7847,7852|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|Acute
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7847,7872|false|false|false|C0022660;C1565662|Acute Kidney Insufficiency;Kidney Failure, Acute|Acute renal insufficiency
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7853,7858|false|false|false|C0022646|Kidney|renal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7853,7858|false|false|false|C0042075|Urologic Diseases|renal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7853,7872|false|false|false|C0035078;C1565489|Kidney Failure;Renal Insufficiency|renal insufficiency
Event|Event|SIMPLE_SEGMENT|7859,7872|false|false|false|||insufficiency
Finding|Functional Concept|SIMPLE_SEGMENT|7859,7872|false|false|false|C0231179|Insufficiency|insufficiency
Event|Event|SIMPLE_SEGMENT|7877,7886|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|7877,7886|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7888,7898|false|false|false|C0010294|creatinine|creatinine
Drug|Organic Chemical|SIMPLE_SEGMENT|7888,7898|false|false|false|C0010294|creatinine|creatinine
Event|Event|SIMPLE_SEGMENT|7888,7898|false|false|false|||creatinine
Finding|Physiologic Function|SIMPLE_SEGMENT|7888,7898|false|false|false|C4551889|Creatinine metabolic function|creatinine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7888,7898|false|false|false|C0201975|Creatinine measurement|creatinine
Finding|Finding|SIMPLE_SEGMENT|7888,7907|false|false|false|C0151578|Creatinine increased|creatinine elevated
Event|Event|SIMPLE_SEGMENT|7899,7907|false|false|false|||elevated
Finding|Finding|SIMPLE_SEGMENT|7917,7923|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|7917,7923|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7931,7942|false|false|false|C0011175;C2062903|Dehydration;dehydration (Na, H2O)|dehydration
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|7931,7942|false|false|false|C0011175;C2062903|Dehydration;dehydration (Na, H2O)|dehydration
Event|Event|SIMPLE_SEGMENT|7931,7942|false|false|false|||dehydration
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7931,7942|false|false|false|C4284399|Dehydration procedure|dehydration
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7947,7957|false|false|false|C0010294|creatinine|creatinine
Drug|Organic Chemical|SIMPLE_SEGMENT|7947,7957|false|false|false|C0010294|creatinine|creatinine
Event|Event|SIMPLE_SEGMENT|7947,7957|false|false|false|||creatinine
Finding|Physiologic Function|SIMPLE_SEGMENT|7947,7957|false|false|false|C4551889|Creatinine metabolic function|creatinine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7947,7957|false|false|false|C0201975|Creatinine measurement|creatinine
Event|Event|SIMPLE_SEGMENT|7958,7966|false|false|false|||improved
Event|Event|SIMPLE_SEGMENT|7968,7977|false|false|false|||overnight
Drug|Organic Chemical|SIMPLE_SEGMENT|7983,7989|false|false|false|C0720654|Gentle|gentle
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7983,7989|false|false|false|C0720654|Gentle|gentle
Drug|Substance|SIMPLE_SEGMENT|7990,7996|false|false|false|C0302908|Liquid substance|fluids
Event|Event|SIMPLE_SEGMENT|7990,7996|false|false|false|||fluids
Finding|Body Substance|SIMPLE_SEGMENT|7990,7996|false|false|false|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7990,7996|false|false|false|C0016286|Fluid Therapy|fluids
Event|Event|SIMPLE_SEGMENT|8001,8009|false|false|false|||remained
Event|Event|SIMPLE_SEGMENT|8010,8016|false|false|false|||stable
Finding|Intellectual Product|SIMPLE_SEGMENT|8010,8016|false|false|false|C1547311|Patient Condition Code - Stable|stable
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8022,8026|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8022,8026|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|SIMPLE_SEGMENT|8022,8026|false|false|false|||COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|8022,8026|false|false|false|C1412502|ARCN1 gene|COPD
Event|Event|SIMPLE_SEGMENT|8028,8037|false|false|false|||Continued
Finding|Idea or Concept|SIMPLE_SEGMENT|8041,8045|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|8041,8045|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|8041,8045|false|false|false|C1553498|home health encounter|home
Event|Event|SIMPLE_SEGMENT|8046,8054|false|false|false|||inhalers
Drug|Organic Chemical|SIMPLE_SEGMENT|8056,8065|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8056,8065|false|false|false|C0001927|albuterol|albuterol
Event|Event|SIMPLE_SEGMENT|8056,8065|false|false|false|||albuterol
Drug|Organic Chemical|SIMPLE_SEGMENT|8067,8078|false|false|false|C0082607|fluticasone|fluticasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8067,8078|false|false|false|C0082607|fluticasone|fluticasone
Event|Event|SIMPLE_SEGMENT|8067,8078|false|false|false|||fluticasone
Event|Event|SIMPLE_SEGMENT|8087,8096|false|false|false|||Continued
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8102,8110|false|false|false|C0907402|insulin glargine|glargine
Drug|Hormone|SIMPLE_SEGMENT|8102,8110|false|false|false|C0907402|insulin glargine|glargine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8102,8110|false|false|false|C0907402|insulin glargine|glargine
Event|Event|SIMPLE_SEGMENT|8102,8110|false|false|false|||glargine
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|8127,8130|false|false|false|C1845118|SHORT STATURE, IDIOPATHIC, X-LINKED|ISS
Event|Event|SIMPLE_SEGMENT|8127,8130|false|false|false|||ISS
Event|Event|SIMPLE_SEGMENT|8141,8150|false|false|false|||Continued
Finding|Idea or Concept|SIMPLE_SEGMENT|8154,8158|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|8154,8158|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|8154,8158|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|8159,8171|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8159,8171|false|false|false|C0286651|atorvastatin|atorvastatin
Event|Event|SIMPLE_SEGMENT|8159,8171|false|false|false|||atorvastatin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8176,8180|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Event|Event|SIMPLE_SEGMENT|8176,8180|false|false|false|||GERD
Event|Event|SIMPLE_SEGMENT|8182,8191|false|false|false|||Continued
Finding|Idea or Concept|SIMPLE_SEGMENT|8195,8199|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|8195,8199|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|8195,8199|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|8200,8212|false|false|false|C0081876|pantoprazole|pantoprazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8200,8212|false|false|false|C0081876|pantoprazole|pantoprazole
Event|Event|SIMPLE_SEGMENT|8200,8212|false|false|false|||pantoprazole
Finding|Idea or Concept|SIMPLE_SEGMENT|8216,8228|false|false|false|C1548597|Marketing basis - Transitional|Transitional
Event|Event|SIMPLE_SEGMENT|8229,8235|false|false|false|||issues
Event|Event|SIMPLE_SEGMENT|8239,8242|false|false|false|||NEW
Finding|Finding|SIMPLE_SEGMENT|8239,8242|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|NEW
Finding|Idea or Concept|SIMPLE_SEGMENT|8239,8242|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|NEW
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8239,8254|false|false|false|C1718097|New medications|NEW MEDICATIONS
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8243,8254|false|false|false|C0802604;C2598133||MEDICATIONS
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8243,8254|false|false|false|C0013227|Pharmaceutical Preparations|MEDICATIONS
Event|Event|SIMPLE_SEGMENT|8243,8254|false|false|false|||MEDICATIONS
Finding|Intellectual Product|SIMPLE_SEGMENT|8243,8254|false|false|false|C4284232|Medications|MEDICATIONS
Drug|Organic Chemical|SIMPLE_SEGMENT|8256,8264|false|false|false|C0126174|losartan|losartan
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8256,8264|false|false|false|C0126174|losartan|losartan
Event|Event|SIMPLE_SEGMENT|8256,8264|false|false|false|||losartan
Drug|Organic Chemical|SIMPLE_SEGMENT|8269,8274|false|false|false|C0590690|Imdur|imdur
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8269,8274|false|false|false|C0590690|Imdur|imdur
Event|Event|SIMPLE_SEGMENT|8269,8274|false|false|false|||imdur
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8277,8287|false|false|false|C0013227|Pharmaceutical Preparations|MEDICATION
Event|Event|SIMPLE_SEGMENT|8277,8287|false|false|false|||MEDICATION
Finding|Intellectual Product|SIMPLE_SEGMENT|8277,8287|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|MEDICATION
Event|Event|SIMPLE_SEGMENT|8288,8295|false|false|false|||CHANGES
Finding|Functional Concept|SIMPLE_SEGMENT|8288,8295|false|false|false|C0392747|Changing|CHANGES
Drug|Organic Chemical|SIMPLE_SEGMENT|8297,8307|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8297,8307|false|false|false|C0025859|metoprolol|metoprolol
Event|Event|SIMPLE_SEGMENT|8297,8307|false|false|false|||metoprolol
Event|Event|SIMPLE_SEGMENT|8308,8317|false|false|false|||increased
Event|Event|SIMPLE_SEGMENT|8329,8332|false|false|false|||TID
Event|Event|SIMPLE_SEGMENT|8353,8360|false|false|false|||ongoing
Finding|Idea or Concept|SIMPLE_SEGMENT|8353,8360|false|false|false|C0549178|Continuous|ongoing
Anatomy|Body Location or Region|SIMPLE_SEGMENT|8361,8366|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|8361,8366|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8361,8371|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|8361,8371|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8367,8371|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|8367,8371|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|8367,8371|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|8367,8371|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|8373,8381|false|false|false|||consider
Event|Event|SIMPLE_SEGMENT|8382,8391|false|false|false|||titrating
Drug|Organic Chemical|SIMPLE_SEGMENT|8398,8403|false|false|false|C0590690|Imdur|imdur
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8398,8403|false|false|false|C0590690|Imdur|imdur
Event|Event|SIMPLE_SEGMENT|8398,8403|false|false|false|||imdur
Finding|Sign or Symptom|SIMPLE_SEGMENT|8412,8424|false|false|false|C0002962|Angina Pectoris|anginal pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8420,8424|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|8420,8424|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|8420,8424|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|8420,8424|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|8437,8445|false|false|false|||consider
Event|Event|SIMPLE_SEGMENT|8446,8454|false|false|false|||treating
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8459,8474|false|false|false|C0040213;C5779793|Costal chondritis;Tietze's Syndrome|costochondritis
Event|Event|SIMPLE_SEGMENT|8459,8474|false|false|false|||costochondritis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8480,8492|false|false|false|C0031046|Pericarditis|pericarditis
Event|Event|SIMPLE_SEGMENT|8480,8492|false|false|false|||pericarditis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8495,8506|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8495,8506|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|8495,8506|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|8495,8506|false|false|false|C4284232|Medications|Medications
Finding|Finding|SIMPLE_SEGMENT|8495,8519|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|SIMPLE_SEGMENT|8510,8519|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|8510,8519|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8538,8548|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|8538,8548|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|8538,8553|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|SIMPLE_SEGMENT|8549,8553|false|false|false|||list
Finding|Intellectual Product|SIMPLE_SEGMENT|8549,8553|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|SIMPLE_SEGMENT|8557,8565|false|false|false|||accurate
Drug|Organic Chemical|SIMPLE_SEGMENT|8570,8578|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8570,8578|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|SIMPLE_SEGMENT|8570,8578|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|SIMPLE_SEGMENT|8570,8578|false|false|false|||complete
Finding|Functional Concept|SIMPLE_SEGMENT|8570,8578|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|SIMPLE_SEGMENT|8570,8578|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Organic Chemical|SIMPLE_SEGMENT|8583,8592|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8583,8592|false|false|false|C0001927|albuterol|Albuterol
Finding|Functional Concept|SIMPLE_SEGMENT|8593,8600|false|false|false|C4319647|Inhaler (unit of presentation)|Inhaler
Finding|Gene or Genome|SIMPLE_SEGMENT|8615,8618|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|SIMPLE_SEGMENT|8619,8622|false|false|false|||SOB
Finding|Sign or Symptom|SIMPLE_SEGMENT|8619,8622|false|false|false|C0013404|Dyspnea|SOB
Drug|Organic Chemical|SIMPLE_SEGMENT|8627,8639|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8627,8639|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|SIMPLE_SEGMENT|8659,8670|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8659,8670|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Organic Chemical|SIMPLE_SEGMENT|8690,8701|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8690,8701|false|false|false|C0082607|fluticasone|Fluticasone
Event|Event|SIMPLE_SEGMENT|8690,8701|false|false|false|||Fluticasone
Drug|Organic Chemical|SIMPLE_SEGMENT|8690,8712|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8690,8712|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Organic Chemical|SIMPLE_SEGMENT|8702,8712|false|false|false|C0033474;C0392214|Propionates;propionate|Propionate
Event|Event|SIMPLE_SEGMENT|8722,8726|false|false|false|||PUFF
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|8730,8733|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8730,8733|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8730,8733|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|8730,8733|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|8730,8733|false|false|false|C1332410|BID gene|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8738,8746|false|false|false|C0907402|insulin glargine|Glargine
Drug|Hormone|SIMPLE_SEGMENT|8738,8746|false|false|false|C0907402|insulin glargine|Glargine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8738,8746|false|false|false|C0907402|insulin glargine|Glargine
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8764,8771|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Hormone|SIMPLE_SEGMENT|8764,8771|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8764,8771|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Event|Event|SIMPLE_SEGMENT|8764,8771|false|false|false|||Insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|8764,8771|false|false|false|C1337112|INS gene|Insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8764,8771|false|false|false|C0202098|Insulin measurement|Insulin
Event|Event|SIMPLE_SEGMENT|8775,8782|false|false|false|||Sliding
Finding|Functional Concept|SIMPLE_SEGMENT|8775,8782|false|false|false|C0332246|Sliding|Sliding
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8775,8788|false|false|false|C2937251|sliding scale|Sliding Scale
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8783,8788|false|false|false|C0222045|Integumentary scale|Scale
Event|Activity|SIMPLE_SEGMENT|8783,8788|false|false|false|C1947916|Scaling|Scale
Finding|Conceptual Entity|SIMPLE_SEGMENT|8783,8788|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|Scale
Finding|Intellectual Product|SIMPLE_SEGMENT|8783,8788|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|Scale
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8799,8806|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Hormone|SIMPLE_SEGMENT|8799,8806|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8799,8806|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Event|Event|SIMPLE_SEGMENT|8799,8806|false|false|false|||Insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|8799,8806|false|false|false|C1337112|INS gene|Insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8799,8806|false|false|false|C0202098|Insulin measurement|Insulin
Drug|Organic Chemical|SIMPLE_SEGMENT|8810,8820|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8810,8820|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Organic Chemical|SIMPLE_SEGMENT|8810,8829|false|false|false|C0700548|metoprolol tartrate|Metoprolol Tartrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8810,8829|false|false|false|C0700548|metoprolol tartrate|Metoprolol Tartrate
Drug|Organic Chemical|SIMPLE_SEGMENT|8821,8829|false|false|false|C0039328;C0144544|Tartrates;tartrate|Tartrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8821,8829|false|false|false|C0039328;C0144544|Tartrates;tartrate|Tartrate
Event|Event|SIMPLE_SEGMENT|8821,8829|false|false|false|||Tartrate
Event|Event|SIMPLE_SEGMENT|8839,8842|false|false|false|||TID
Event|Activity|SIMPLE_SEGMENT|8844,8848|false|false|false|C1948035|Hold (action)|Hold
Event|Event|SIMPLE_SEGMENT|8844,8848|false|false|false|||Hold
Finding|Functional Concept|SIMPLE_SEGMENT|8844,8848|false|false|false|C1553387;C3853841|Hold - dosing instruction fragment;hold - Data Operation|Hold
Finding|Intellectual Product|SIMPLE_SEGMENT|8844,8848|false|false|false|C1553387;C3853841|Hold - dosing instruction fragment;hold - Data Operation|Hold
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8853,8856|false|false|false|C0871470|Systolic Pressure|SBP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8853,8856|false|false|false|C0085805|Androgen Binding Protein|SBP
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8853,8856|false|false|false|C0085805|Androgen Binding Protein|SBP
Event|Event|SIMPLE_SEGMENT|8853,8856|false|false|false|||SBP
Finding|Gene or Genome|SIMPLE_SEGMENT|8853,8856|false|false|false|C1705296;C3274833|CCHCR1 wt Allele;SHBG wt Allele|SBP
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8853,8856|false|false|false|C1306620|Systolic blood pressure measurement|SBP
Drug|Organic Chemical|SIMPLE_SEGMENT|8873,8881|false|false|false|C0699681|MetroGel|Metrogel
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8873,8881|false|false|false|C0699681|MetroGel|Metrogel
Event|Event|SIMPLE_SEGMENT|8873,8881|false|false|false|||Metrogel
Drug|Organic Chemical|SIMPLE_SEGMENT|8888,8901|false|false|false|C0025872|metronidazole|metroNIDAZOLE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8888,8901|false|false|false|C0025872|metronidazole|metroNIDAZOLE
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8910,8917|false|false|false|C1710439|Topical Dosage Form|Topical
Finding|Functional Concept|SIMPLE_SEGMENT|8910,8917|false|false|false|C1522168|Topical Route of Administration|Topical
Drug|Organic Chemical|SIMPLE_SEGMENT|8928,8937|false|false|false|C0030049|oxycodone|Oxycodone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8928,8937|false|false|false|C0030049|oxycodone|Oxycodone
Event|Event|SIMPLE_SEGMENT|8928,8937|false|false|false|||Oxycodone
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8928,8937|false|false|false|C0524222|Oxycodone measurement|Oxycodone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8928,8951|false|false|false|C0717368|acetaminophen / oxycodone|Oxycodone-Acetaminophen
Drug|Organic Chemical|SIMPLE_SEGMENT|8938,8951|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8938,8951|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|SIMPLE_SEGMENT|8938,8951|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8938,8951|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8966,8969|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|SIMPLE_SEGMENT|8966,8969|false|false|false|||TAB
Finding|Gene or Genome|SIMPLE_SEGMENT|8977,8980|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|SIMPLE_SEGMENT|8981,8987|false|false|false|||severe
Finding|Finding|SIMPLE_SEGMENT|8981,8987|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|SIMPLE_SEGMENT|8981,8987|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8989,8993|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|8989,8993|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|8989,8993|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|8989,8993|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|SIMPLE_SEGMENT|8998,9010|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8998,9010|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Organic Chemical|SIMPLE_SEGMENT|9030,9040|false|false|false|C0244821|ropinirole|Ropinirole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9030,9040|false|false|false|C0244821|ropinirole|Ropinirole
Event|Event|SIMPLE_SEGMENT|9052,9055|false|false|false|||QPM
Drug|Organic Chemical|SIMPLE_SEGMENT|9061,9068|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9061,9068|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|SIMPLE_SEGMENT|9090,9097|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9090,9097|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|SIMPLE_SEGMENT|9090,9097|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|SIMPLE_SEGMENT|9090,9099|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|SIMPLE_SEGMENT|9090,9099|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9090,9099|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|SIMPLE_SEGMENT|9090,9099|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Event|Event|SIMPLE_SEGMENT|9090,9099|false|false|false|||Vitamin D
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9090,9099|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Event|Event|SIMPLE_SEGMENT|9110,9112|false|false|false|||PO
Drug|Organic Chemical|SIMPLE_SEGMENT|9124,9133|false|false|false|C0020740|ibuprofen|Ibuprofen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9124,9133|false|false|false|C0020740|ibuprofen|Ibuprofen
Finding|Gene or Genome|SIMPLE_SEGMENT|9148,9151|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9152,9156|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|9152,9156|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|9152,9156|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|9152,9156|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|9161,9170|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|9161,9170|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|9161,9170|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|9161,9170|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|9161,9170|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|9161,9182|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9171,9182|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9171,9182|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|9171,9182|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|9171,9182|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|SIMPLE_SEGMENT|9187,9196|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9187,9196|false|false|false|C0001927|albuterol|Albuterol
Finding|Functional Concept|SIMPLE_SEGMENT|9197,9204|false|false|false|C4319647|Inhaler (unit of presentation)|Inhaler
Finding|Gene or Genome|SIMPLE_SEGMENT|9219,9222|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|SIMPLE_SEGMENT|9223,9226|false|false|false|||SOB
Finding|Sign or Symptom|SIMPLE_SEGMENT|9223,9226|false|false|false|C0013404|Dyspnea|SOB
Drug|Organic Chemical|SIMPLE_SEGMENT|9231,9238|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9231,9238|false|false|false|C0004057|aspirin|Aspirin
Event|Event|SIMPLE_SEGMENT|9255,9257|false|false|false|||RX
Drug|Organic Chemical|SIMPLE_SEGMENT|9259,9266|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9259,9266|false|false|false|C0004057|aspirin|aspirin
Event|Event|SIMPLE_SEGMENT|9259,9266|false|false|false|||aspirin
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9275,9281|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|SIMPLE_SEGMENT|9285,9293|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9288,9293|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|9288,9293|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9310,9316|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|9310,9316|false|false|false|||Tablet
Event|Event|SIMPLE_SEGMENT|9318,9325|false|false|false|||Refills
Finding|Idea or Concept|SIMPLE_SEGMENT|9318,9325|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|9332,9344|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9332,9344|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|SIMPLE_SEGMENT|9365,9377|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9365,9377|false|false|false|C0286651|atorvastatin|atorvastatin
Event|Event|SIMPLE_SEGMENT|9365,9377|false|false|false|||atorvastatin
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9386,9392|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|SIMPLE_SEGMENT|9396,9404|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9399,9404|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|9399,9404|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9422,9428|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|9429,9436|false|false|false|||Refills
Finding|Idea or Concept|SIMPLE_SEGMENT|9429,9436|false|false|false|C0807726|refill|Refills
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9443,9451|false|false|false|C0907402|insulin glargine|Glargine
Drug|Hormone|SIMPLE_SEGMENT|9443,9451|false|false|false|C0907402|insulin glargine|Glargine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9443,9451|false|false|false|C0907402|insulin glargine|Glargine
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9469,9476|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Hormone|SIMPLE_SEGMENT|9469,9476|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9469,9476|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Event|Event|SIMPLE_SEGMENT|9469,9476|false|false|false|||Insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|9469,9476|false|false|false|C1337112|INS gene|Insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9469,9476|false|false|false|C0202098|Insulin measurement|Insulin
Event|Event|SIMPLE_SEGMENT|9480,9487|false|false|false|||Sliding
Finding|Functional Concept|SIMPLE_SEGMENT|9480,9487|false|false|false|C0332246|Sliding|Sliding
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9480,9493|false|false|false|C2937251|sliding scale|Sliding Scale
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9488,9493|false|false|false|C0222045|Integumentary scale|Scale
Event|Activity|SIMPLE_SEGMENT|9488,9493|false|false|false|C1947916|Scaling|Scale
Finding|Conceptual Entity|SIMPLE_SEGMENT|9488,9493|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|Scale
Finding|Intellectual Product|SIMPLE_SEGMENT|9488,9493|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|Scale
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9504,9511|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Hormone|SIMPLE_SEGMENT|9504,9511|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9504,9511|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Event|Event|SIMPLE_SEGMENT|9504,9511|false|false|false|||Insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|9504,9511|false|false|false|C1337112|INS gene|Insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9504,9511|false|false|false|C0202098|Insulin measurement|Insulin
Drug|Organic Chemical|SIMPLE_SEGMENT|9515,9525|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9515,9525|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Organic Chemical|SIMPLE_SEGMENT|9515,9534|false|false|false|C0700548|metoprolol tartrate|Metoprolol Tartrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9515,9534|false|false|false|C0700548|metoprolol tartrate|Metoprolol Tartrate
Drug|Organic Chemical|SIMPLE_SEGMENT|9526,9534|false|false|false|C0039328;C0144544|Tartrates;tartrate|Tartrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9526,9534|false|false|false|C0039328;C0144544|Tartrates;tartrate|Tartrate
Event|Event|SIMPLE_SEGMENT|9526,9534|false|false|false|||Tartrate
Event|Event|SIMPLE_SEGMENT|9544,9547|false|false|false|||TID
Drug|Organic Chemical|SIMPLE_SEGMENT|9553,9563|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9553,9563|false|false|false|C0025859|metoprolol|metoprolol
Drug|Organic Chemical|SIMPLE_SEGMENT|9553,9572|false|false|false|C0700548|metoprolol tartrate|metoprolol tartrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9553,9572|false|false|false|C0700548|metoprolol tartrate|metoprolol tartrate
Drug|Organic Chemical|SIMPLE_SEGMENT|9564,9572|false|false|false|C0039328;C0144544|Tartrates;tartrate|tartrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9564,9572|false|false|false|C0039328;C0144544|Tartrates;tartrate|tartrate
Event|Event|SIMPLE_SEGMENT|9564,9572|false|false|false|||tartrate
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9581,9587|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|SIMPLE_SEGMENT|9591,9599|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9594,9599|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|9594,9599|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9606,9611|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|SIMPLE_SEGMENT|9615,9618|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|9615,9618|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9629,9635|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|9636,9643|false|false|false|||Refills
Finding|Idea or Concept|SIMPLE_SEGMENT|9636,9643|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|9650,9662|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9650,9662|false|false|false|C0081876|pantoprazole|Pantoprazole
Event|Event|SIMPLE_SEGMENT|9678,9680|false|false|false|||RX
Drug|Organic Chemical|SIMPLE_SEGMENT|9682,9694|false|false|false|C0081876|pantoprazole|pantoprazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9682,9694|false|false|false|C0081876|pantoprazole|pantoprazole
Event|Event|SIMPLE_SEGMENT|9682,9694|false|false|false|||pantoprazole
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9703,9709|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|SIMPLE_SEGMENT|9713,9721|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9716,9721|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|9716,9721|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9739,9745|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|9746,9753|false|false|false|||Refills
Finding|Idea or Concept|SIMPLE_SEGMENT|9746,9753|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|9760,9770|false|false|false|C0244821|ropinirole|Ropinirole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9760,9770|false|false|false|C0244821|ropinirole|Ropinirole
Event|Event|SIMPLE_SEGMENT|9782,9785|false|false|false|||QPM
Drug|Organic Chemical|SIMPLE_SEGMENT|9790,9797|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9790,9797|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|SIMPLE_SEGMENT|9790,9797|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|SIMPLE_SEGMENT|9790,9799|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|SIMPLE_SEGMENT|9790,9799|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9790,9799|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|SIMPLE_SEGMENT|9790,9799|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9790,9799|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Event|Event|SIMPLE_SEGMENT|9798,9799|false|false|false|||D
Event|Event|SIMPLE_SEGMENT|9805,9809|false|false|false|||UNIT
Drug|Organic Chemical|SIMPLE_SEGMENT|9823,9833|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9823,9833|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Organic Chemical|SIMPLE_SEGMENT|9823,9845|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9823,9845|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Event|Event|SIMPLE_SEGMENT|9834,9845|false|false|false|||Mononitrate
Finding|Finding|SIMPLE_SEGMENT|9847,9855|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|SIMPLE_SEGMENT|9847,9855|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|SIMPLE_SEGMENT|9856,9863|false|false|false|||Release
Finding|Functional Concept|SIMPLE_SEGMENT|9856,9863|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|9856,9863|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9856,9863|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|SIMPLE_SEGMENT|9885,9895|false|false|false|C0022251|isosorbide|isosorbide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9885,9895|false|false|false|C0022251|isosorbide|isosorbide
Drug|Organic Chemical|SIMPLE_SEGMENT|9885,9907|false|false|false|C0064079|isosorbide mononitrate|isosorbide mononitrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9885,9907|false|false|false|C0064079|isosorbide mononitrate|isosorbide mononitrate
Event|Event|SIMPLE_SEGMENT|9896,9907|false|false|false|||mononitrate
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9916,9922|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|SIMPLE_SEGMENT|9926,9934|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9929,9934|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|9929,9934|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Event|Activity|SIMPLE_SEGMENT|9941,9945|false|false|false|C1880359|Dispense (activity)|Disp
Finding|Gene or Genome|SIMPLE_SEGMENT|9941,9945|false|false|false|C2828567|PRSS30P gene|Disp
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9952,9958|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|9959,9966|false|false|false|||Refills
Finding|Idea or Concept|SIMPLE_SEGMENT|9959,9966|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|9974,9982|false|false|false|C0699681|MetroGel|Metrogel
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9974,9982|false|false|false|C0699681|MetroGel|Metrogel
Event|Event|SIMPLE_SEGMENT|9974,9982|false|false|false|||Metrogel
Drug|Organic Chemical|SIMPLE_SEGMENT|9989,10002|false|false|false|C0025872|metronidazole|metroNIDAZOLE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9989,10002|false|false|false|C0025872|metronidazole|metroNIDAZOLE
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10011,10018|false|false|false|C1710439|Topical Dosage Form|Topical
Finding|Functional Concept|SIMPLE_SEGMENT|10011,10018|false|false|false|C1522168|Topical Route of Administration|Topical
Drug|Organic Chemical|SIMPLE_SEGMENT|10030,10039|false|false|false|C0030049|oxycodone|Oxycodone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10030,10039|false|false|false|C0030049|oxycodone|Oxycodone
Event|Event|SIMPLE_SEGMENT|10030,10039|false|false|false|||Oxycodone
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10030,10039|false|false|false|C0524222|Oxycodone measurement|Oxycodone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10030,10053|false|false|false|C0717368|acetaminophen / oxycodone|Oxycodone-Acetaminophen
Drug|Organic Chemical|SIMPLE_SEGMENT|10040,10053|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10040,10053|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|SIMPLE_SEGMENT|10040,10053|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10040,10053|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10068,10071|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|SIMPLE_SEGMENT|10068,10071|false|false|false|||TAB
Finding|Gene or Genome|SIMPLE_SEGMENT|10079,10082|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|SIMPLE_SEGMENT|10083,10089|false|false|false|||severe
Finding|Finding|SIMPLE_SEGMENT|10083,10089|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|SIMPLE_SEGMENT|10083,10089|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10091,10095|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|10091,10095|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|10091,10095|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|10091,10095|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|SIMPLE_SEGMENT|10101,10109|false|false|false|C0126174|losartan|Losartan
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10101,10109|false|false|false|C0126174|losartan|Losartan
Event|Event|SIMPLE_SEGMENT|10101,10109|false|false|false|||Losartan
Drug|Organic Chemical|SIMPLE_SEGMENT|10101,10119|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10101,10119|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|10110,10119|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|10110,10119|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Food|SIMPLE_SEGMENT|10110,10119|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|10110,10119|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10110,10119|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Event|Event|SIMPLE_SEGMENT|10110,10119|false|false|false|||Potassium
Finding|Physiologic Function|SIMPLE_SEGMENT|10110,10119|false|false|false|C4553027|Potassium metabolic function|Potassium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10110,10119|false|false|false|C0202194|Potassium measurement|Potassium
Drug|Organic Chemical|SIMPLE_SEGMENT|10140,10148|false|false|false|C0126174|losartan|losartan
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10140,10148|false|false|false|C0126174|losartan|losartan
Event|Event|SIMPLE_SEGMENT|10140,10148|false|false|false|||losartan
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10157,10163|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|SIMPLE_SEGMENT|10167,10175|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|10170,10175|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|10170,10175|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10192,10198|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|10192,10198|false|false|false|||Tablet
Event|Event|SIMPLE_SEGMENT|10200,10207|false|false|false|||Refills
Finding|Idea or Concept|SIMPLE_SEGMENT|10200,10207|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|10215,10226|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10215,10226|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Organic Chemical|SIMPLE_SEGMENT|10247,10258|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10247,10258|false|false|false|C0082607|fluticasone|Fluticasone
Event|Event|SIMPLE_SEGMENT|10247,10258|false|false|false|||Fluticasone
Drug|Organic Chemical|SIMPLE_SEGMENT|10247,10269|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10247,10269|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Organic Chemical|SIMPLE_SEGMENT|10259,10269|false|false|false|C0033474;C0392214|Propionates;propionate|Propionate
Event|Event|SIMPLE_SEGMENT|10279,10283|false|false|false|||PUFF
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|10287,10290|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10287,10290|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|10287,10290|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|10287,10290|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|10287,10290|false|false|false|C1332410|BID gene|BID
Event|Event|SIMPLE_SEGMENT|10295,10304|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|10295,10304|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|10295,10304|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|10295,10304|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|10295,10304|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10295,10316|false|false|false|C4019243||Discharge Disposition
Finding|Finding|SIMPLE_SEGMENT|10295,10316|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10305,10316|false|false|false|C2926604||Disposition
Event|Event|SIMPLE_SEGMENT|10305,10316|false|false|false|||Disposition
Procedure|Health Care Activity|SIMPLE_SEGMENT|10305,10316|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|SIMPLE_SEGMENT|10318,10322|false|false|false|||Home
Finding|Idea or Concept|SIMPLE_SEGMENT|10318,10322|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|SIMPLE_SEGMENT|10318,10322|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|SIMPLE_SEGMENT|10318,10322|false|false|false|C1553498|home health encounter|Home
Event|Event|SIMPLE_SEGMENT|10325,10334|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|10325,10334|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|10325,10334|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|10325,10334|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|10325,10334|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|10325,10344|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10335,10344|false|false|false|C0945731||Diagnosis
Event|Event|SIMPLE_SEGMENT|10335,10344|false|false|false|||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|10335,10344|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|10335,10344|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10335,10344|false|false|false|C0011900|Diagnosis|Diagnosis
Event|Event|SIMPLE_SEGMENT|10362,10371|false|false|false|||elevation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10362,10371|false|false|false|C0439775|Elevation procedure|elevation
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10375,10383|false|false|false|C0018787|Heart|coronary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10375,10390|false|false|false|C0205042|Coronary artery|coronary artery
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10375,10398|false|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|coronary artery disease
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10384,10390|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|SIMPLE_SEGMENT|10384,10390|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10384,10398|false|false|false|C0852949|Arteriopathic disease|artery disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10391,10398|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|10391,10398|false|false|false|||disease
Disorder|Neoplastic Process|SIMPLE_SEGMENT|10400,10409|false|false|false|C0027627|Neoplasm Metastasis|Secondary
Event|Event|SIMPLE_SEGMENT|10400,10409|false|false|false|||Secondary
Finding|Functional Concept|SIMPLE_SEGMENT|10400,10409|false|false|false|C1522484|metastatic qualifier|Secondary
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10411,10419|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|diabetes
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10411,10428|false|false|false|C0011849|Diabetes Mellitus|diabetes mellitus
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10411,10435|false|false|false|C0011860|Diabetes Mellitus, Non-Insulin-Dependent|diabetes mellitus type 2
Event|Event|SIMPLE_SEGMENT|10429,10433|false|false|false|||type
Finding|Gene or Genome|SIMPLE_SEGMENT|10429,10433|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Finding|Intellectual Product|SIMPLE_SEGMENT|10429,10433|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Finding|Classification|SIMPLE_SEGMENT|10429,10435|false|false|false|C0441730|Type 2|type 2
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10436,10448|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|SIMPLE_SEGMENT|10436,10448|false|false|false|||hypertension
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10449,10463|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|hyperlipidemia
Event|Event|SIMPLE_SEGMENT|10449,10463|false|false|false|||hyperlipidemia
Finding|Finding|SIMPLE_SEGMENT|10449,10463|false|false|false|C0428465|Serum lipids high (finding)|hyperlipidemia
Event|Event|SIMPLE_SEGMENT|10467,10476|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|10467,10476|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|10467,10476|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|10467,10476|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|10467,10476|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10477,10486|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10477,10486|false|false|false|C0012634|Disease|Condition
Event|Event|SIMPLE_SEGMENT|10477,10486|false|false|false|||Condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|10477,10486|false|false|false|C1705253|Logical Condition|Condition
Finding|Mental Process|SIMPLE_SEGMENT|10488,10494|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10488,10501|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|SIMPLE_SEGMENT|10488,10501|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10495,10501|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|10495,10501|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|10503,10508|false|false|false|||Clear
Finding|Idea or Concept|SIMPLE_SEGMENT|10503,10508|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|SIMPLE_SEGMENT|10513,10521|false|false|false|||coherent
Finding|Finding|SIMPLE_SEGMENT|10513,10521|false|false|false|C4068804|Coherent|coherent
Event|Event|SIMPLE_SEGMENT|10523,10528|false|false|false|||Level
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10523,10545|false|false|false|C4050479||Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|10523,10545|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|SIMPLE_SEGMENT|10532,10545|false|false|false|||Consciousness
Finding|Finding|SIMPLE_SEGMENT|10532,10545|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|SIMPLE_SEGMENT|10532,10545|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10547,10552|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|10547,10552|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10547,10552|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|SIMPLE_SEGMENT|10547,10552|false|false|false|||Alert
Finding|Finding|SIMPLE_SEGMENT|10547,10552|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|10547,10552|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|10547,10552|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|SIMPLE_SEGMENT|10557,10568|false|false|false|||interactive
Finding|Functional Concept|SIMPLE_SEGMENT|10557,10568|false|false|false|C1704675|Interaction|interactive
Event|Activity|SIMPLE_SEGMENT|10570,10578|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|10570,10578|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|SIMPLE_SEGMENT|10570,10578|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10579,10585|false|false|false|C5889824||Status
Event|Event|SIMPLE_SEGMENT|10579,10585|false|false|false|||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|10579,10585|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|10587,10597|false|false|false|||Ambulatory
Finding|Functional Concept|SIMPLE_SEGMENT|10587,10597|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|SIMPLE_SEGMENT|10587,10597|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|SIMPLE_SEGMENT|10587,10597|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|SIMPLE_SEGMENT|10587,10597|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|SIMPLE_SEGMENT|10600,10611|false|false|false|||Independent
Finding|Finding|SIMPLE_SEGMENT|10600,10611|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|SIMPLE_SEGMENT|10600,10611|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Event|Event|SIMPLE_SEGMENT|10616,10625|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|10616,10625|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|10616,10625|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|10616,10625|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|10616,10625|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10616,10638|false|false|false|C3669312||Discharge Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|10616,10638|false|false|false|C4282220|Discharge instructions|Discharge Instructions
Procedure|Health Care Activity|SIMPLE_SEGMENT|10616,10638|false|false|false|C2266673|hospital discharge instructions (treatment)|Discharge Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10626,10638|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|10626,10638|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|10626,10638|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Event|Event|SIMPLE_SEGMENT|10649,10657|false|false|false|||pleasure
Finding|Intellectual Product|SIMPLE_SEGMENT|10649,10657|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|SIMPLE_SEGMENT|10649,10657|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|SIMPLE_SEGMENT|10665,10669|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|10665,10669|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|10665,10669|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|10665,10669|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|10665,10672|false|false|false|C1555558|care of - AddressPartType|care of
Event|Event|SIMPLE_SEGMENT|10697,10706|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|10697,10706|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|SIMPLE_SEGMENT|10725,10733|false|false|false|||admitted
Anatomy|Body Location or Region|SIMPLE_SEGMENT|10739,10744|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|10739,10744|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10739,10749|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|10739,10749|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10745,10749|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|10745,10749|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|10745,10749|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|10745,10749|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|SIMPLE_SEGMENT|10750,10758|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|SIMPLE_SEGMENT|10750,10758|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|10750,10758|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|10750,10758|false|false|false|C0033095||pressure
Event|Event|SIMPLE_SEGMENT|10759,10769|false|false|false|||concerning
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10777,10782|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|10777,10782|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|10777,10782|false|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10777,10789|false|false|false|C0027051|Myocardial Infarction|heart attack
Event|Event|SIMPLE_SEGMENT|10783,10789|false|false|false|||attack
Finding|Finding|SIMPLE_SEGMENT|10783,10789|false|false|false|C1261512;C1304680|Attack (finding);Attack behavior|attack
Finding|Social Behavior|SIMPLE_SEGMENT|10783,10789|false|false|false|C1261512;C1304680|Attack (finding);Attack behavior|attack
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10794,10801|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|10794,10801|false|false|false|C1314974|Cardiac attachment|cardiac
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|10794,10817|false|false|false|C0261588|Cardiac catheterisation as the cause of abnormal reaction of the patient, or of later complication, without mention of misadventure at the time of the procedure|cardiac catheterization
Finding|Intellectual Product|SIMPLE_SEGMENT|10794,10817|false|false|false|C1547981|Diagnostic Service Section ID - Cardiac Catheterization|cardiac catheterization
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10794,10817|false|false|false|C0018795;C1548828|Cardiac Catheterization Procedures;Consent Type - Cardiac Catheterization|cardiac catheterization
Procedure|Health Care Activity|SIMPLE_SEGMENT|10794,10817|false|false|false|C0018795;C1548828|Cardiac Catheterization Procedures;Consent Type - Cardiac Catheterization|cardiac catheterization
Event|Event|SIMPLE_SEGMENT|10802,10817|false|false|false|||catheterization
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10802,10817|false|false|false|C0007430|Catheterization|catheterization
Event|Event|SIMPLE_SEGMENT|10818,10824|false|false|false|||showed
Anatomy|Tissue|SIMPLE_SEGMENT|10843,10849|false|false|false|C0332835|Transplanted tissue|grafts
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10843,10849|false|false|false|C0181074|Graft material|grafts
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10867,10874|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|10867,10874|false|false|false|C1314974|Cardiac attachment|cardiac
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10875,10881|false|false|false|C0813207|Creation of shunt|bypass
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10875,10889|false|false|false|C1536078|Bypass surgery|bypass surgery
Event|Event|SIMPLE_SEGMENT|10882,10889|false|false|false|||surgery
Finding|Finding|SIMPLE_SEGMENT|10882,10889|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|SIMPLE_SEGMENT|10882,10889|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|SIMPLE_SEGMENT|10882,10889|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10882,10889|false|false|false|C0543467|Operative Surgical Procedures|surgery
Event|Event|SIMPLE_SEGMENT|10916,10923|false|false|false|||working
Event|Occupational Activity|SIMPLE_SEGMENT|10916,10923|false|false|false|C0043227|Work|working
Finding|Idea or Concept|SIMPLE_SEGMENT|10916,10923|false|false|false|C1563351|Diagnosis Type - Working|working
Event|Event|SIMPLE_SEGMENT|10937,10944|false|false|false|||causing
Event|Event|SIMPLE_SEGMENT|10950,10958|false|false|false|||symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|10950,10958|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|10950,10958|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|SIMPLE_SEGMENT|10971,10980|false|false|false|||increased
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10991,11002|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10991,11002|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|10991,11002|false|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|10991,11002|false|false|false|C4284232|Medications|medications
Event|Event|SIMPLE_SEGMENT|11006,11013|false|false|false|||control
Event|Event|SIMPLE_SEGMENT|11020,11028|false|false|false|||symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|11020,11028|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|11020,11028|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|SIMPLE_SEGMENT|11035,11042|false|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|11035,11042|false|false|false|C0392747|Changing|changes
Drug|Food|SIMPLE_SEGMENT|11054,11059|false|false|false|C0452588|Start brand of breakfast cereal|START
Event|Event|SIMPLE_SEGMENT|11054,11059|false|false|false|||START
Finding|Intellectual Product|SIMPLE_SEGMENT|11054,11059|false|false|false|C1552850|start - HtmlLinkType|START
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11054,11059|false|false|false|C5447432|Collagen Tile Brachytherapy|START
Drug|Organic Chemical|SIMPLE_SEGMENT|11060,11068|false|false|false|C0126174|losartan|losartan
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11060,11068|false|false|false|C0126174|losartan|losartan
Event|Event|SIMPLE_SEGMENT|11060,11068|false|false|false|||losartan
Drug|Food|SIMPLE_SEGMENT|11069,11074|false|false|false|C0452588|Start brand of breakfast cereal|START
Event|Event|SIMPLE_SEGMENT|11069,11074|false|false|false|||START
Finding|Intellectual Product|SIMPLE_SEGMENT|11069,11074|false|false|false|C1552850|start - HtmlLinkType|START
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11069,11074|false|false|false|C5447432|Collagen Tile Brachytherapy|START
Drug|Organic Chemical|SIMPLE_SEGMENT|11075,11085|false|false|false|C0022251|isosorbide|isosorbide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11075,11085|false|false|false|C0022251|isosorbide|isosorbide
Drug|Organic Chemical|SIMPLE_SEGMENT|11075,11097|false|false|false|C0064079|isosorbide mononitrate|isosorbide mononitrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11075,11097|false|false|false|C0064079|isosorbide mononitrate|isosorbide mononitrate
Event|Event|SIMPLE_SEGMENT|11086,11097|false|false|false|||mononitrate
Finding|Functional Concept|SIMPLE_SEGMENT|11098,11106|false|false|false|C0442805|Increase|INCREASE
Drug|Organic Chemical|SIMPLE_SEGMENT|11107,11119|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11107,11119|false|false|false|C0286651|atorvastatin|atorvastatin
Event|Event|SIMPLE_SEGMENT|11107,11119|false|false|false|||atorvastatin
Finding|Functional Concept|SIMPLE_SEGMENT|11120,11128|false|false|false|C0442805|Increase|INCREASE
Drug|Organic Chemical|SIMPLE_SEGMENT|11129,11139|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11129,11139|false|false|false|C0025859|metoprolol|metoprolol
Event|Event|SIMPLE_SEGMENT|11129,11139|false|false|false|||metoprolol
Finding|Finding|SIMPLE_SEGMENT|11140,11148|false|false|false|C0392756|Reduced|DECREASE
Drug|Organic Chemical|SIMPLE_SEGMENT|11149,11156|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11149,11156|false|false|false|C0004057|aspirin|aspirin
Event|Event|SIMPLE_SEGMENT|11149,11156|false|false|false|||aspirin
Finding|Finding|SIMPLE_SEGMENT|11157,11165|false|false|false|C0392756|Reduced|DECREASE
Drug|Organic Chemical|SIMPLE_SEGMENT|11166,11178|false|false|false|C0081876|pantoprazole|pantoprazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11166,11178|false|false|false|C0081876|pantoprazole|pantoprazole
Event|Event|SIMPLE_SEGMENT|11166,11178|false|false|false|||pantoprazole
Drug|Inorganic Chemical|SIMPLE_SEGMENT|11179,11183|false|false|false|C0723457|Stop brand of fluoride|STOP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11179,11183|false|false|false|C0723457|Stop brand of fluoride|STOP
Event|Activity|SIMPLE_SEGMENT|11179,11183|false|false|false|C1947925|Stop (Instruction Imperative)|STOP
Event|Event|SIMPLE_SEGMENT|11179,11183|false|false|false|||STOP
Finding|Gene or Genome|SIMPLE_SEGMENT|11179,11183|false|false|false|C1417022|MAP6 gene|STOP
Drug|Organic Chemical|SIMPLE_SEGMENT|11184,11193|false|false|false|C0020740|ibuprofen|ibuprofen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11184,11193|false|false|false|C0020740|ibuprofen|ibuprofen
Event|Event|SIMPLE_SEGMENT|11184,11193|false|false|false|||ibuprofen
Event|Event|SIMPLE_SEGMENT|11204,11210|false|false|false|||taking
Finding|Finding|SIMPLE_SEGMENT|11211,11219|false|false|false|C3843660|Too much|too much
Event|Event|SIMPLE_SEGMENT|11215,11219|false|false|false|||much
Finding|Finding|SIMPLE_SEGMENT|11215,11219|false|false|false|C4281574|Much|much
Drug|Organic Chemical|SIMPLE_SEGMENT|11226,11233|false|false|false|C0699142|Tylenol|tylenol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11226,11233|false|false|false|C0699142|Tylenol|tylenol
Event|Event|SIMPLE_SEGMENT|11226,11233|false|false|false|||tylenol
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11243,11247|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|11243,11247|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|11243,11247|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|11243,11247|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|11259,11264|false|false|false|||leave
Finding|Idea or Concept|SIMPLE_SEGMENT|11269,11277|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|SIMPLE_SEGMENT|11282,11291|false|false|false|||recommend
Event|Event|SIMPLE_SEGMENT|11300,11306|false|false|false|||workup
Drug|Substance|SIMPLE_SEGMENT|11313,11318|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|11313,11318|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|11313,11318|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|11319,11329|false|false|false|||collection
Finding|Conceptual Entity|SIMPLE_SEGMENT|11319,11329|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|SIMPLE_SEGMENT|11319,11329|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|SIMPLE_SEGMENT|11319,11329|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|SIMPLE_SEGMENT|11319,11329|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Event|Event|SIMPLE_SEGMENT|11330,11334|false|false|false|||seen
Finding|Functional Concept|SIMPLE_SEGMENT|11347,11351|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11347,11356|false|false|false|C0225730|Left lung|left lung
Anatomy|Body Location or Region|SIMPLE_SEGMENT|11352,11356|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11352,11356|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11352,11356|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|SIMPLE_SEGMENT|11352,11356|false|false|false|C0740941|Lung Problem|lung
Event|Event|SIMPLE_SEGMENT|11361,11367|false|false|false|||better
Finding|Idea or Concept|SIMPLE_SEGMENT|11361,11367|false|false|false|C1550462|Observation Interpretation - better|better
Event|Event|SIMPLE_SEGMENT|11369,11379|false|false|false|||management
Event|Occupational Activity|SIMPLE_SEGMENT|11369,11379|false|false|false|C0001554;C1273870|Administration occupational activities;Management procedure|management
Procedure|Health Care Activity|SIMPLE_SEGMENT|11369,11379|false|false|false|C0376636|Disease Management|management
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11388,11396|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|diabetes
Event|Event|SIMPLE_SEGMENT|11388,11396|false|false|false|||diabetes
Event|Event|SIMPLE_SEGMENT|11406,11410|false|false|false|||help
Finding|Intellectual Product|SIMPLE_SEGMENT|11406,11410|false|false|false|C1552861|Help document|help
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11419,11422|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|11419,11422|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|11419,11422|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|11419,11422|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|SIMPLE_SEGMENT|11419,11422|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|11419,11422|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|SIMPLE_SEGMENT|11419,11422|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11419,11422|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|SIMPLE_SEGMENT|11419,11422|false|false|false|||PCP
Finding|Gene or Genome|SIMPLE_SEGMENT|11419,11422|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|SIMPLE_SEGMENT|11419,11422|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Procedure|Health Care Activity|SIMPLE_SEGMENT|11426,11434|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11435,11447|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|11435,11447|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|11435,11447|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

