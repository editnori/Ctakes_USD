 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|42,51|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|42,51|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|42,56|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|76,85|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|76,85|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|76,85|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|76,85|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|76,85|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|76,90|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|108,113|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|108,113|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|108,113|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|132,135|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|143,150|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|143,150|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|152,160|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|SIMPLE_SEGMENT|163,172|false|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|163,172|false|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|163,172|false|false|false|C0020517|Hypersensitivity|Allergies
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|178,181|false|false|false|C0013343|Dyes|Dye
Event|Event|SIMPLE_SEGMENT|178,181|false|false|false|||Dye
Drug|Biologically Active Substance|SIMPLE_SEGMENT|183,189|false|false|false|C0021968;C0885449|Iodine, Homeopathic preparation;iodine|Iodine
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|183,189|false|false|false|C0021968;C0885449|Iodine, Homeopathic preparation;iodine|Iodine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|183,189|false|false|false|C0021968;C0885449|Iodine, Homeopathic preparation;iodine|Iodine
Event|Activity|SIMPLE_SEGMENT|190,200|false|false|false|C2700400|Contain (action)|Containing
Finding|Functional Concept|SIMPLE_SEGMENT|190,200|false|false|false|C0332256|Containing (qualifier value)|Containing
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|201,209|false|false|false|C0009924|Contrast Media|Contrast
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|201,215|false|false|false|C0009924|Contrast Media|Contrast Media
Anatomy|Tissue|SIMPLE_SEGMENT|210,215|false|false|false|C0162867;C1254021|Media layer;Tunica Media|Media
Finding|Intellectual Product|SIMPLE_SEGMENT|210,215|false|false|false|C0009458;C0677540|Communications Media;PAMS Media|Media
Drug|Organic Chemical|SIMPLE_SEGMENT|218,227|false|false|false|C0030049|oxycodone|Oxycodone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|218,227|false|false|false|C0030049|oxycodone|Oxycodone
Event|Event|SIMPLE_SEGMENT|218,227|false|false|false|||Oxycodone
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|218,227|false|false|false|C0524222|Oxycodone measurement|Oxycodone
Drug|Organic Chemical|SIMPLE_SEGMENT|231,241|false|false|false|C0055729|cilostazol|cilostazol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|231,241|false|false|false|C0055729|cilostazol|cilostazol
Event|Event|SIMPLE_SEGMENT|231,241|false|false|false|||cilostazol
Drug|Organic Chemical|SIMPLE_SEGMENT|244,255|false|false|false|C1569608|varenicline|Varenicline
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|244,255|false|false|false|C1569608|varenicline|Varenicline
Event|Event|SIMPLE_SEGMENT|244,255|false|false|false|||Varenicline
Event|Event|SIMPLE_SEGMENT|258,267|false|false|false|||Attending
Finding|Functional Concept|SIMPLE_SEGMENT|258,267|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|SIMPLE_SEGMENT|275,290|false|false|false|C0277786|Chief complaint (finding)|Chief Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|281,290|false|false|false|C3864418||Complaint
Event|Event|SIMPLE_SEGMENT|281,290|false|false|false|||Complaint
Finding|Finding|SIMPLE_SEGMENT|281,290|false|false|false|C5441521|Complaint (finding)|Complaint
Finding|Finding|SIMPLE_SEGMENT|292,299|false|false|false|C0013404;C2024878|Dyspnea|Dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|292,299|false|false|false|C0013404;C2024878|Dyspnea|Dyspnea
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|301,307|false|false|false|C0018792|Heart Atrium|Atrial
Attribute|Clinical Attribute|SIMPLE_SEGMENT|301,320|false|false|false|C2926591||Atrial Fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|301,320|false|false|false|C0004238|Atrial Fibrillation|Atrial Fibrillation
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|301,320|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Atrial Fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|308,320|false|false|false|C0232197|Fibrillation|Fibrillation
Event|Event|SIMPLE_SEGMENT|308,320|false|false|false|||Fibrillation
Finding|Classification|SIMPLE_SEGMENT|323,328|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|SIMPLE_SEGMENT|329,337|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|329,337|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|341,359|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|350,359|false|false|false|C0945766||Procedure
Event|Event|SIMPLE_SEGMENT|350,359|false|false|false|||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|350,359|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|350,359|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|350,359|false|false|false|C0184661|Interventional procedure|Procedure
Event|Event|SIMPLE_SEGMENT|369,376|true|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|369,376|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|369,376|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|369,376|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|369,379|true|false|false|C0262926|Medical History|History of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|369,395|true|false|false|C0488508||History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|369,395|true|false|false|C0262512|History of present illness (finding)|History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|380,387|true|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Idea or Concept|SIMPLE_SEGMENT|380,387|true|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Finding|SIMPLE_SEGMENT|380,395|true|false|false|C4264312|Present illness|Present Illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|388,395|true|false|false|C0221423|Illness (finding)|Illness
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|416,420|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|416,420|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|SIMPLE_SEGMENT|416,420|false|false|false|||COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|416,420|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|437,440|false|false|false|C0020538|Hypertensive disease|htn
Event|Event|SIMPLE_SEGMENT|437,440|false|false|false|||htn
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|442,446|false|false|false|C0004238|Atrial Fibrillation|afib
Event|Event|SIMPLE_SEGMENT|442,446|false|false|false|||afib
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|442,446|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|afib
Event|Event|SIMPLE_SEGMENT|451,459|false|false|false|||presents
Event|Event|SIMPLE_SEGMENT|466,473|false|false|false|||dyspnea
Finding|Finding|SIMPLE_SEGMENT|466,473|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|466,473|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Event|Event|SIMPLE_SEGMENT|491,498|false|false|false|||treated
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|503,507|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|503,507|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|SIMPLE_SEGMENT|503,507|false|false|false|||COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|503,507|false|false|false|C1412502|ARCN1 gene|COPD
Event|Event|SIMPLE_SEGMENT|512,520|false|false|false|||admitted
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|526,530|false|false|false|C0004238|Atrial Fibrillation|Afib
Event|Event|SIMPLE_SEGMENT|526,530|false|false|false|||Afib
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|526,530|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Afib
Event|Event|SIMPLE_SEGMENT|536,539|false|false|false|||RVR
Finding|Finding|SIMPLE_SEGMENT|536,539|false|false|false|C1417822;C3540498;C4050414|NR1D2 gene;NR1D2 wt Allele;Rapid Virologic Response|RVR
Finding|Gene or Genome|SIMPLE_SEGMENT|536,539|false|false|false|C1417822;C3540498;C4050414|NR1D2 gene;NR1D2 wt Allele;Rapid Virologic Response|RVR
Finding|Body Substance|SIMPLE_SEGMENT|548,555|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|548,555|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|548,555|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|586,595|false|false|false|||diagnosed
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|604,608|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|604,608|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|SIMPLE_SEGMENT|604,608|false|false|false|||COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|604,608|false|false|false|C1412502|ARCN1 gene|COPD
Event|Event|SIMPLE_SEGMENT|609,614|false|false|false|||flare
Finding|Finding|SIMPLE_SEGMENT|609,614|false|false|false|C1517205;C3540542|Exacerbation of cGVHD;Flare|flare
Finding|Sign or Symptom|SIMPLE_SEGMENT|609,614|false|false|false|C1517205;C3540542|Exacerbation of cGVHD;Flare|flare
Event|Event|SIMPLE_SEGMENT|624,634|false|false|false|||discharged
Drug|Hormone|SIMPLE_SEGMENT|642,652|false|false|false|C0032952|prednisone|prednisone
Drug|Organic Chemical|SIMPLE_SEGMENT|642,652|false|false|false|C0032952|prednisone|prednisone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|642,652|false|false|false|C0032952|prednisone|prednisone
Event|Event|SIMPLE_SEGMENT|653,658|false|false|false|||taper
Procedure|Health Care Activity|SIMPLE_SEGMENT|653,658|false|false|false|C0441640||taper
Drug|Antibiotic|SIMPLE_SEGMENT|684,696|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Clinical Drug|SIMPLE_SEGMENT|684,696|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Organic Chemical|SIMPLE_SEGMENT|684,696|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Event|Event|SIMPLE_SEGMENT|684,696|false|false|false|||azithromycin
Event|Event|SIMPLE_SEGMENT|720,724|false|false|false|||felt
Finding|Finding|SIMPLE_SEGMENT|726,730|false|false|false|C5575035|Well (answer to question)|well
Finding|Intellectual Product|SIMPLE_SEGMENT|732,736|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|SIMPLE_SEGMENT|737,746|false|false|false|||developed
Event|Event|SIMPLE_SEGMENT|747,754|false|false|false|||dyspnea
Finding|Finding|SIMPLE_SEGMENT|747,754|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|747,754|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Finding|SIMPLE_SEGMENT|747,762|false|false|false|C0743330|Rest Dyspnea|dyspnea at rest
Finding|Functional Concept|SIMPLE_SEGMENT|755,762|false|false|false|C0443144|At rest (qualifier value)|at rest
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|758,762|false|false|false|C1742913|REST protein, human|rest
Drug|Biologically Active Substance|SIMPLE_SEGMENT|758,762|false|false|false|C1742913|REST protein, human|rest
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|758,762|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Gene or Genome|SIMPLE_SEGMENT|758,762|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Molecular Function|SIMPLE_SEGMENT|758,762|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Event|Event|SIMPLE_SEGMENT|764,773|false|false|false|||worsening
Event|Event|SIMPLE_SEGMENT|779,787|false|false|false|||exertion
Finding|Organism Function|SIMPLE_SEGMENT|779,787|false|false|false|C0015264|Exertion|exertion
Event|Event|SIMPLE_SEGMENT|794,802|false|false|false|||inhalers
Event|Event|SIMPLE_SEGMENT|803,811|false|false|false|||improved
Event|Event|SIMPLE_SEGMENT|816,819|false|false|false|||SOB
Finding|Sign or Symptom|SIMPLE_SEGMENT|816,819|false|false|false|C0013404|Dyspnea|SOB
Event|Event|SIMPLE_SEGMENT|825,829|false|false|false|||felt
Event|Event|SIMPLE_SEGMENT|841,849|false|false|false|||symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|841,849|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|841,849|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|SIMPLE_SEGMENT|856,866|false|false|false|||consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|856,866|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|856,871|false|false|false|C0332290|Consistent with|consistent with
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|876,880|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|876,880|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|SIMPLE_SEGMENT|876,880|false|false|false|||COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|876,880|false|false|false|C1412502|ARCN1 gene|COPD
Event|Event|SIMPLE_SEGMENT|886,889|false|false|false|||saw
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|894,897|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|894,897|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|894,897|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|894,897|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|SIMPLE_SEGMENT|894,897|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|894,897|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|SIMPLE_SEGMENT|894,897|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|894,897|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|SIMPLE_SEGMENT|894,897|false|false|false|||PCP
Finding|Gene or Genome|SIMPLE_SEGMENT|894,897|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|SIMPLE_SEGMENT|894,897|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Event|SIMPLE_SEGMENT|933,938|false|false|false|||found
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|948,952|false|false|false|C0004238|Atrial Fibrillation|Afib
Event|Event|SIMPLE_SEGMENT|948,952|false|false|false|||Afib
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|948,952|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Afib
Event|Event|SIMPLE_SEGMENT|956,959|false|false|false|||RVR
Finding|Finding|SIMPLE_SEGMENT|956,959|false|false|false|C1417822;C3540498;C4050414|NR1D2 gene;NR1D2 wt Allele;Rapid Virologic Response|RVR
Finding|Gene or Genome|SIMPLE_SEGMENT|956,959|false|false|false|C1417822;C3540498;C4050414|NR1D2 gene;NR1D2 wt Allele;Rapid Virologic Response|RVR
Event|Activity|SIMPLE_SEGMENT|961,965|false|false|false|C0871208|Rating (action)|rate
Event|Event|SIMPLE_SEGMENT|961,965|false|false|false|||rate
Finding|Idea or Concept|SIMPLE_SEGMENT|961,965|false|false|false|C1549480|Amount type - Rate|rate
Event|Event|SIMPLE_SEGMENT|993,1000|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|993,1000|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|993,1000|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|993,1000|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|993,1003|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1004,1008|false|false|false|C0004238|Atrial Fibrillation|afib
Event|Event|SIMPLE_SEGMENT|1004,1008|false|false|false|||afib
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1004,1008|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|afib
Event|Event|SIMPLE_SEGMENT|1013,1021|false|false|false|||referred
Event|Event|SIMPLE_SEGMENT|1052,1055|false|false|false|||SOB
Finding|Sign or Symptom|SIMPLE_SEGMENT|1052,1055|false|false|false|C0013404|Dyspnea|SOB
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1060,1064|false|false|false|C0004238|Atrial Fibrillation|afib
Event|Event|SIMPLE_SEGMENT|1060,1064|false|false|false|||afib
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1060,1064|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|afib
Event|Event|SIMPLE_SEGMENT|1070,1073|false|false|false|||RVR
Finding|Finding|SIMPLE_SEGMENT|1070,1073|false|false|false|C1417822;C3540498;C4050414|NR1D2 gene;NR1D2 wt Allele;Rapid Virologic Response|RVR
Finding|Gene or Genome|SIMPLE_SEGMENT|1070,1073|false|false|false|C1417822;C3540498;C4050414|NR1D2 gene;NR1D2 wt Allele;Rapid Virologic Response|RVR
Event|Event|SIMPLE_SEGMENT|1079,1085|false|false|false|||states
Event|Event|SIMPLE_SEGMENT|1096,1105|false|false|false|||compliant
Finding|Individual Behavior|SIMPLE_SEGMENT|1096,1105|false|false|false|C1321605|Compliance behavior|compliant
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|1111,1115|false|false|false|C1300458|Nebulizer solution|nebs
Event|Event|SIMPLE_SEGMENT|1111,1115|false|false|false|||nebs
Drug|Organic Chemical|SIMPLE_SEGMENT|1120,1127|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1120,1127|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Event|Event|SIMPLE_SEGMENT|1120,1127|false|false|false|||steroid
Event|Event|SIMPLE_SEGMENT|1136,1143|false|false|false|||regimen
Finding|Intellectual Product|SIMPLE_SEGMENT|1136,1143|false|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1136,1143|false|false|false|C0040808|Treatment Protocols|regimen
Event|Event|SIMPLE_SEGMENT|1149,1155|true|false|false|||denies
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1165,1170|true|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|1165,1170|true|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|1165,1170|true|false|false|C0013604|Edema|edema
Event|Event|SIMPLE_SEGMENT|1172,1181|true|false|false|||orthopnea
Finding|Finding|SIMPLE_SEGMENT|1172,1181|true|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|1172,1181|true|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Event|Event|SIMPLE_SEGMENT|1187,1193|false|false|false|||denies
Event|Event|SIMPLE_SEGMENT|1201,1207|true|false|false|||travel
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|1201,1207|true|false|false|C0040802|travel|travel
Procedure|Health Care Activity|SIMPLE_SEGMENT|1201,1207|true|false|false|C1555670|travel charge|travel
Event|Event|SIMPLE_SEGMENT|1209,1218|true|false|false|||surgeries
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1209,1218|true|false|false|C0543467|Operative Surgical Procedures|surgeries
Event|Event|SIMPLE_SEGMENT|1232,1239|false|false|false|||episode
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1243,1248|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|1243,1248|false|false|false|C0741025|Chest problem|chest
Finding|Sign or Symptom|SIMPLE_SEGMENT|1243,1258|false|false|false|C0232292|Chest tightness|chest tightness
Event|Event|SIMPLE_SEGMENT|1249,1258|false|false|false|||tightness
Event|Event|SIMPLE_SEGMENT|1272,1276|false|false|false|||felt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1287,1291|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1287,1291|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|SIMPLE_SEGMENT|1287,1291|false|false|false|||COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|1287,1291|false|false|false|C1412502|ARCN1 gene|COPD
Event|Event|SIMPLE_SEGMENT|1292,1298|false|false|false|||flares
Event|Event|SIMPLE_SEGMENT|1300,1306|false|false|false|||Denies
Event|Event|SIMPLE_SEGMENT|1307,1313|true|false|false|||fevers
Finding|Sign or Symptom|SIMPLE_SEGMENT|1307,1313|true|false|false|C0015967|Fever|fevers
Event|Event|SIMPLE_SEGMENT|1317,1325|true|false|false|||coughing
Finding|Sign or Symptom|SIMPLE_SEGMENT|1317,1325|true|false|false|C0010200|Coughing|coughing
Event|Event|SIMPLE_SEGMENT|1329,1339|true|false|false|||production
Event|Occupational Activity|SIMPLE_SEGMENT|1329,1339|true|false|false|C0033268|production|production
Finding|Intellectual Product|SIMPLE_SEGMENT|1329,1339|true|false|false|C1548180|Production Processing ID|production
Event|Event|SIMPLE_SEGMENT|1343,1349|true|false|false|||sputum
Finding|Body Substance|SIMPLE_SEGMENT|1343,1349|true|false|false|C0038056;C1546789;C1576419|Specimen Type - Sputum;Sputum|sputum
Finding|Intellectual Product|SIMPLE_SEGMENT|1343,1349|true|false|false|C0038056;C1546789;C1576419|Specimen Type - Sputum;Sputum|sputum
Event|Event|SIMPLE_SEGMENT|1352,1363|false|false|false|||hemomptysis
Finding|Finding|SIMPLE_SEGMENT|1369,1389|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Event|Event|SIMPLE_SEGMENT|1374,1381|false|false|false|||Medical
Finding|Functional Concept|SIMPLE_SEGMENT|1374,1381|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|1374,1381|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|1374,1381|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|1374,1381|false|false|false|C0199168|Medical service|Medical
Finding|Finding|SIMPLE_SEGMENT|1374,1389|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1382,1389|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1382,1389|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|1382,1389|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1391,1397|false|false|false|C0004096|Asthma|ASTHMA
Event|Event|SIMPLE_SEGMENT|1391,1397|false|false|false|||ASTHMA
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1398,1402|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1398,1402|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|SIMPLE_SEGMENT|1398,1402|false|false|false|||COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|1398,1402|false|false|false|C1412502|ARCN1 gene|COPD
Finding|Finding|SIMPLE_SEGMENT|1406,1414|false|false|false|C0741302|atypia morphology|ATYPICAL
Finding|Sign or Symptom|SIMPLE_SEGMENT|1406,1425|false|false|false|C0262384|Atypical chest pain|ATYPICAL CHEST PAIN
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1415,1420|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|CHEST
Finding|Finding|SIMPLE_SEGMENT|1415,1420|false|false|false|C0741025|Chest problem|CHEST
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1415,1425|false|false|false|C2926613||CHEST PAIN
Finding|Sign or Symptom|SIMPLE_SEGMENT|1415,1425|false|false|false|C0008031|Chest Pain|CHEST PAIN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1421,1425|false|true|false|C2598155||PAIN
Event|Event|SIMPLE_SEGMENT|1421,1425|false|false|false|||PAIN
Finding|Functional Concept|SIMPLE_SEGMENT|1421,1425|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|PAIN
Finding|Sign or Symptom|SIMPLE_SEGMENT|1421,1425|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|PAIN
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1429,1437|false|false|false|C0027530|Neck|CERVICAL
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1429,1449|false|false|false|C0263884|Cervical radiculitis|CERVICAL RADICULITIS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1438,1449|false|false|false|C0034544|Radiculitis|RADICULITIS
Event|Event|SIMPLE_SEGMENT|1438,1449|false|false|false|||RADICULITIS
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1453,1461|false|false|false|C0027530|Neck|CERVICAL
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1453,1473|false|false|false|C0158241;C1384641|Cervical spondylosis;Cervical spondylosis without myelopathy|CERVICAL SPONDYLOSIS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1462,1473|false|false|false|C0038019|Spondylosis|SPONDYLOSIS
Event|Event|SIMPLE_SEGMENT|1462,1473|false|false|false|||SPONDYLOSIS
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1477,1485|false|false|false|C0018787|Heart|CORONARY
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1477,1492|false|false|false|C0205042|Coronary artery|CORONARY ARTERY
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1477,1500|false|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|CORONARY ARTERY DISEASE
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1486,1492|false|false|false|C0003842;C0226004|Arterial system;Arteries|ARTERY
Anatomy|Body System|SIMPLE_SEGMENT|1486,1492|false|false|false|C0003842;C0226004|Arterial system;Arteries|ARTERY
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1486,1500|false|false|false|C0852949|Arteriopathic disease|ARTERY DISEASE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1493,1500|false|false|false|C0012634|Disease|DISEASE
Event|Event|SIMPLE_SEGMENT|1493,1500|false|false|false|||DISEASE
Finding|Sign or Symptom|SIMPLE_SEGMENT|1504,1512|false|false|false|C0018681|Headache|HEADACHE
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1516,1519|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|HIP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1516,1519|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|HIP
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1516,1519|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|HIP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1516,1519|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|HIP
Event|Event|SIMPLE_SEGMENT|1516,1519|false|false|false|||HIP
Finding|Gene or Genome|SIMPLE_SEGMENT|1516,1519|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|HIP
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1516,1519|false|false|false|C1292890|Procedure on hip|HIP
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1516,1531|false|false|false|C0392806|Prosthetic arthroplasty of hip (procedure)|HIP REPLACEMENT
Event|Event|SIMPLE_SEGMENT|1520,1531|false|false|false|||REPLACEMENT
Finding|Functional Concept|SIMPLE_SEGMENT|1520,1531|false|false|false|C0559956|Replacement|REPLACEMENT
Procedure|Health Care Activity|SIMPLE_SEGMENT|1520,1531|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|REPLACEMENT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1520,1531|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|REPLACEMENT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1535,1549|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|HYPERLIPIDEMIA
Event|Event|SIMPLE_SEGMENT|1535,1549|false|false|false|||HYPERLIPIDEMIA
Finding|Finding|SIMPLE_SEGMENT|1535,1549|false|false|false|C0428465|Serum lipids high (finding)|HYPERLIPIDEMIA
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1553,1565|false|false|false|C0020538|Hypertensive disease|HYPERTENSION
Event|Event|SIMPLE_SEGMENT|1553,1565|false|false|false|||HYPERTENSION
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1569,1583|false|false|false|C0029408|Degenerative polyarthritis|OSTEOARTHRITIS
Event|Event|SIMPLE_SEGMENT|1569,1583|false|false|false|||OSTEOARTHRITIS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1587,1593|false|false|false|C0019340;C0854331|Herpes simplex dermatitis|HERPES
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1587,1600|false|false|false|C0019360;C0042338|Herpes zoster (disorder);herpesvirus 3, human|HERPES ZOSTER
Disorder|Virus|SIMPLE_SEGMENT|1587,1600|false|false|false|C0019360;C0042338|Herpes zoster (disorder);herpesvirus 3, human|HERPES ZOSTER
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1594,1600|false|false|false|C0019360|Herpes zoster (disorder)|ZOSTER
Event|Event|SIMPLE_SEGMENT|1594,1600|false|false|false|||ZOSTER
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1604,1610|false|false|false|C0018792|Heart Atrium|ATRIAL
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1604,1623|false|false|false|C2926591||ATRIAL FIBRILLATION
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1604,1623|false|false|false|C0004238|Atrial Fibrillation|ATRIAL FIBRILLATION
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1604,1623|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|ATRIAL FIBRILLATION
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1611,1623|false|false|false|C0232197|Fibrillation|FIBRILLATION
Event|Event|SIMPLE_SEGMENT|1611,1623|false|false|false|||FIBRILLATION
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|1627,1634|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|ANXIETY
Event|Event|SIMPLE_SEGMENT|1627,1634|false|false|false|||ANXIETY
Finding|Sign or Symptom|SIMPLE_SEGMENT|1627,1634|false|false|false|C0860603|Anxiety symptoms|ANXIETY
Finding|Intellectual Product|SIMPLE_SEGMENT|1638,1654|false|false|false|C1314977|Gastrointestinal attachment|GASTROINTESTINAL
Finding|Pathologic Function|SIMPLE_SEGMENT|1638,1663|false|false|false|C0017181|Gastrointestinal Hemorrhage|GASTROINTESTINAL BLEEDING
Finding|Pathologic Function|SIMPLE_SEGMENT|1655,1663|false|false|false|C0019080|Hemorrhage|BLEEDING
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1667,1681|false|false|false|C0029408|Degenerative polyarthritis|OSTEOARTHRITIS
Event|Event|SIMPLE_SEGMENT|1667,1681|false|false|false|||OSTEOARTHRITIS
Finding|Functional Concept|SIMPLE_SEGMENT|1685,1700|false|false|false|C0333482|atherosclerotic|ATHEROSCLEROTIC
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1685,1723|false|false|false|C0004153|Atherosclerosis|ATHEROSCLEROTIC CARDIOVASCULAR DISEASE
Anatomy|Body System|SIMPLE_SEGMENT|1701,1715|false|false|false|C0007226;C3887460|Cardiovascular;Cardiovascular system|CARDIOVASCULAR
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1701,1723|false|false|false|C0007222|Cardiovascular Diseases|CARDIOVASCULAR DISEASE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1716,1723|false|false|false|C0012634|Disease|DISEASE
Event|Event|SIMPLE_SEGMENT|1716,1723|false|false|false|||DISEASE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1727,1754|false|false|false|C0085096|Peripheral Vascular Diseases|PERIPHERAL VASCULAR DISEASE
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1738,1746|false|false|false|C0005847|Blood Vessel|VASCULAR
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1738,1754|false|false|false|C0042373|Vascular Diseases|VASCULAR DISEASE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1747,1754|false|false|false|C0012634|Disease|DISEASE
Event|Event|SIMPLE_SEGMENT|1747,1754|false|false|false|||DISEASE
Finding|Functional Concept|SIMPLE_SEGMENT|1757,1763|false|false|false|C0728831|Social|Social
Finding|Finding|SIMPLE_SEGMENT|1757,1771|false|false|false|C0424945;C3714536|Social History;Social and personal history|Social History
Event|Event|SIMPLE_SEGMENT|1764,1771|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1764,1771|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1764,1771|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|1764,1771|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Classification|SIMPLE_SEGMENT|1777,1783|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|SIMPLE_SEGMENT|1777,1783|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|SIMPLE_SEGMENT|1777,1783|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|SIMPLE_SEGMENT|1777,1783|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Finding|SIMPLE_SEGMENT|1777,1791|false|false|false|C0241889|Family Medical History|Family History
Event|Event|SIMPLE_SEGMENT|1784,1791|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1784,1791|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1784,1791|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|1784,1791|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Idea or Concept|SIMPLE_SEGMENT|1793,1799|false|false|false|C1546508|Relationship - Mother|Mother
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1806,1809|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|SIMPLE_SEGMENT|1806,1809|false|false|false|||HTN
Finding|Conceptual Entity|SIMPLE_SEGMENT|1812,1818|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Idea or Concept|SIMPLE_SEGMENT|1812,1818|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Event|Event|SIMPLE_SEGMENT|1829,1836|false|false|false|||Brother
Finding|Conceptual Entity|SIMPLE_SEGMENT|1829,1836|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Finding|Idea or Concept|SIMPLE_SEGMENT|1829,1836|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Event|Event|SIMPLE_SEGMENT|1844,1851|false|false|false|||Brother
Finding|Conceptual Entity|SIMPLE_SEGMENT|1844,1851|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Finding|Idea or Concept|SIMPLE_SEGMENT|1844,1851|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Event|Event|SIMPLE_SEGMENT|1860,1868|false|false|false|||Physical
Finding|Finding|SIMPLE_SEGMENT|1860,1868|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|1860,1868|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|1860,1868|false|false|false|C0031809|Physical Examination|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|1874,1883|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|SIMPLE_SEGMENT|1884,1892|false|false|false|||PHYSICAL
Finding|Finding|SIMPLE_SEGMENT|1884,1892|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|SIMPLE_SEGMENT|1884,1892|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|1884,1892|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|SIMPLE_SEGMENT|1884,1897|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAM
Procedure|Health Care Activity|SIMPLE_SEGMENT|1884,1897|false|false|false|C0031809|Physical Examination|PHYSICAL EXAM
Event|Event|SIMPLE_SEGMENT|1893,1897|false|false|false|||EXAM
Finding|Functional Concept|SIMPLE_SEGMENT|1893,1897|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|SIMPLE_SEGMENT|1893,1897|false|false|false|C0582103|Medical Examination|EXAM
Event|Event|SIMPLE_SEGMENT|1932,1939|false|false|false|||GENERAL
Finding|Classification|SIMPLE_SEGMENT|1932,1939|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|1932,1939|false|false|false|C3812897|General medical service|GENERAL
Finding|Finding|SIMPLE_SEGMENT|1941,1945|true|false|false|C5575035|Well (answer to question)|Well
Event|Event|SIMPLE_SEGMENT|1946,1955|true|false|false|||appearing
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1957,1960|true|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1957,1960|true|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1957,1960|true|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|1957,1960|true|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1957,1960|true|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|SIMPLE_SEGMENT|1957,1960|true|false|false|||NAD
Finding|Finding|SIMPLE_SEGMENT|1957,1960|true|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|1965,1981|true|false|false|C0158784|Accessory skeletal muscle|accessory muscle
Finding|Finding|SIMPLE_SEGMENT|1965,1985|true|false|false|C1821466|Use of accessory muscles|accessory muscle use
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1975,1981|true|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Anatomy|Tissue|SIMPLE_SEGMENT|1975,1981|true|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Event|Event|SIMPLE_SEGMENT|1982,1985|true|false|false|||use
Finding|Functional Concept|SIMPLE_SEGMENT|1982,1985|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|SIMPLE_SEGMENT|1982,1985|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1990,1995|false|false|false|C1512338|HEENT|HEENT
Event|Event|SIMPLE_SEGMENT|1997,2001|false|false|false|||NCAT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2003,2009|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2003,2009|false|false|false|C0036412|Scleral Diseases|Sclera
Event|Event|SIMPLE_SEGMENT|2003,2009|false|false|false|||Sclera
Procedure|Health Care Activity|SIMPLE_SEGMENT|2003,2009|false|false|false|C2228481|examination of sclera|Sclera
Event|Event|SIMPLE_SEGMENT|2010,2019|false|false|false|||anicteric
Finding|Finding|SIMPLE_SEGMENT|2010,2019|false|false|false|C0205180|Anicteric|anicteric
Event|Event|SIMPLE_SEGMENT|2021,2026|false|false|false|||PERRL
Finding|Finding|SIMPLE_SEGMENT|2021,2026|false|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Event|Event|SIMPLE_SEGMENT|2028,2032|false|false|false|||EOMI
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2037,2041|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|SIMPLE_SEGMENT|2037,2041|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|SIMPLE_SEGMENT|2037,2041|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Event|Event|SIMPLE_SEGMENT|2046,2049|true|false|false|||JVD
Finding|Finding|SIMPLE_SEGMENT|2046,2049|true|false|false|C0425687|Jugular venous engorgement|JVD
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2053,2060|true|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|SIMPLE_SEGMENT|2053,2060|true|false|false|C1314974|Cardiac attachment|CARDIAC
Event|Event|SIMPLE_SEGMENT|2072,2078|false|false|false|||rhythm
Finding|Finding|SIMPLE_SEGMENT|2072,2078|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|SIMPLE_SEGMENT|2072,2078|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Event|Activity|SIMPLE_SEGMENT|2087,2091|false|false|false|C0871208|Rating (action)|rate
Event|Event|SIMPLE_SEGMENT|2087,2091|false|false|false|||rate
Finding|Idea or Concept|SIMPLE_SEGMENT|2087,2091|false|false|false|C1549480|Amount type - Rate|rate
Event|Event|SIMPLE_SEGMENT|2112,2119|true|false|false|||murmurs
Finding|Finding|SIMPLE_SEGMENT|2112,2119|true|false|false|C0018808|Heart murmur|murmurs
Event|Event|SIMPLE_SEGMENT|2120,2124|true|false|false|||rubs
Finding|Finding|SIMPLE_SEGMENT|2120,2124|true|false|false|C0232267|Pericardial friction rub|rubs
Event|Event|SIMPLE_SEGMENT|2125,2132|true|false|false|||gallops
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2137,2142|false|false|false|C0024109|Lung|LUNGS
Drug|Inorganic Chemical|SIMPLE_SEGMENT|2151,2154|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2151,2154|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|SIMPLE_SEGMENT|2151,2154|false|false|false|C0001861;C3536832|Air (substance);air|air
Finding|Finding|SIMPLE_SEGMENT|2151,2154|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|SIMPLE_SEGMENT|2151,2154|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|SIMPLE_SEGMENT|2151,2154|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Event|Event|SIMPLE_SEGMENT|2155,2159|false|false|false|||well
Finding|Finding|SIMPLE_SEGMENT|2155,2159|false|false|false|C5575035|Well (answer to question)|well
Finding|Functional Concept|SIMPLE_SEGMENT|2173,2178|false|false|false|C1883002|Sequence Chromatogram|Trace
Finding|Organism Function|SIMPLE_SEGMENT|2179,2190|false|false|false|C0004048|Inspiration (function)|inspiratory
Finding|Sign or Symptom|SIMPLE_SEGMENT|2179,2199|false|false|false|C0231874|Inspiratory wheezing|inspiratory wheezing
Event|Event|SIMPLE_SEGMENT|2191,2199|false|false|false|||wheezing
Finding|Sign or Symptom|SIMPLE_SEGMENT|2191,2199|false|false|false|C0043144|Wheezing|wheezing
Finding|Organism Function|SIMPLE_SEGMENT|2212,2222|false|false|false|C0231800|Expiration, Respiratory|expiratory
Finding|Sign or Symptom|SIMPLE_SEGMENT|2212,2231|false|false|false|C0231875|Expiratory wheezing|expiratory wheezing
Event|Event|SIMPLE_SEGMENT|2223,2231|false|false|false|||wheezing
Finding|Sign or Symptom|SIMPLE_SEGMENT|2223,2231|false|false|false|C0043144|Wheezing|wheezing
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2239,2243|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2239,2243|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2239,2243|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|SIMPLE_SEGMENT|2239,2243|false|false|false|C0740941|Lung Problem|lung
Event|Event|SIMPLE_SEGMENT|2244,2250|false|false|false|||fields
Event|Event|SIMPLE_SEGMENT|2256,2264|true|false|false|||crackles
Finding|Finding|SIMPLE_SEGMENT|2256,2264|true|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Event|Event|SIMPLE_SEGMENT|2265,2272|true|false|false|||rhonchi
Finding|Finding|SIMPLE_SEGMENT|2265,2272|true|false|false|C0035508|Rhonchi|rhonchi
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2277,2284|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2277,2284|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Event|Event|SIMPLE_SEGMENT|2277,2284|false|false|false|||ABDOMEN
Finding|Finding|SIMPLE_SEGMENT|2277,2284|false|false|false|C0941288|Abdomen problem|ABDOMEN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2286,2290|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Event|Event|SIMPLE_SEGMENT|2286,2290|false|false|false|||Soft
Event|Event|SIMPLE_SEGMENT|2292,2296|false|false|false|||NTND
Event|Event|SIMPLE_SEGMENT|2301,2304|true|false|false|||HSM
Finding|Gene or Genome|SIMPLE_SEGMENT|2301,2304|true|false|false|C1537594|LRRC4B gene|HSM
Event|Event|SIMPLE_SEGMENT|2308,2318|true|false|false|||tenderness
Finding|Mental Process|SIMPLE_SEGMENT|2308,2318|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|SIMPLE_SEGMENT|2308,2318|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2323,2334|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2349,2356|true|false|false|C0015811|Femur|femoral
Event|Event|SIMPLE_SEGMENT|2357,2363|true|false|false|||bruits
Finding|Finding|SIMPLE_SEGMENT|2357,2363|true|false|false|C0006318|Bruit|bruits
Finding|Body Substance|SIMPLE_SEGMENT|2368,2377|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|2368,2377|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|2368,2377|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|2368,2377|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|SIMPLE_SEGMENT|2378,2386|false|false|false|||PHYSICAL
Finding|Finding|SIMPLE_SEGMENT|2378,2386|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|SIMPLE_SEGMENT|2378,2386|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|2378,2386|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|SIMPLE_SEGMENT|2378,2391|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAM
Procedure|Health Care Activity|SIMPLE_SEGMENT|2378,2391|false|false|false|C0031809|Physical Examination|PHYSICAL EXAM
Event|Event|SIMPLE_SEGMENT|2387,2391|false|false|false|||EXAM
Finding|Functional Concept|SIMPLE_SEGMENT|2387,2391|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|SIMPLE_SEGMENT|2387,2391|false|false|false|C0582103|Medical Examination|EXAM
Event|Event|SIMPLE_SEGMENT|2420,2427|false|false|false|||GENERAL
Finding|Classification|SIMPLE_SEGMENT|2420,2427|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|2420,2427|false|false|false|C3812897|General medical service|GENERAL
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2429,2432|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2429,2432|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2429,2432|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|2429,2432|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2429,2432|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|SIMPLE_SEGMENT|2429,2432|false|false|false|||NAD
Finding|Finding|SIMPLE_SEGMENT|2429,2432|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2433,2438|false|false|false|C1512338|HEENT|HEENT
Event|Event|SIMPLE_SEGMENT|2440,2444|false|false|false|||NCAT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2446,2452|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2446,2452|false|false|false|C0036412|Scleral Diseases|Sclera
Event|Event|SIMPLE_SEGMENT|2446,2452|false|false|false|||Sclera
Procedure|Health Care Activity|SIMPLE_SEGMENT|2446,2452|false|false|false|C2228481|examination of sclera|Sclera
Event|Event|SIMPLE_SEGMENT|2453,2462|false|false|false|||anicteric
Finding|Finding|SIMPLE_SEGMENT|2453,2462|false|false|false|C0205180|Anicteric|anicteric
Event|Event|SIMPLE_SEGMENT|2477,2488|false|false|false|||noninjected
Event|Event|SIMPLE_SEGMENT|2494,2499|false|false|false|||clear
Finding|Idea or Concept|SIMPLE_SEGMENT|2494,2499|false|false|false|C1550016|Remote control command - Clear|clear
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2501,2505|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|SIMPLE_SEGMENT|2501,2505|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|SIMPLE_SEGMENT|2501,2505|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Event|Event|SIMPLE_SEGMENT|2510,2513|true|false|false|||JVD
Finding|Finding|SIMPLE_SEGMENT|2510,2513|true|false|false|C0425687|Jugular venous engorgement|JVD
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2516,2523|true|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|SIMPLE_SEGMENT|2516,2523|true|false|false|C1314974|Cardiac attachment|CARDIAC
Event|Event|SIMPLE_SEGMENT|2525,2528|false|false|false|||RRR
Event|Event|SIMPLE_SEGMENT|2548,2555|true|false|false|||murmurs
Finding|Finding|SIMPLE_SEGMENT|2548,2555|true|false|false|C0018808|Heart murmur|murmurs
Finding|Finding|SIMPLE_SEGMENT|2556,2560|true|false|false|C0232267|Pericardial friction rub|rubs
Event|Event|SIMPLE_SEGMENT|2561,2568|true|false|false|||gallops
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2572,2577|false|false|false|C0024109|Lung|LUNGS
Event|Event|SIMPLE_SEGMENT|2586,2593|false|false|false|||reduced
Drug|Inorganic Chemical|SIMPLE_SEGMENT|2594,2597|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2594,2597|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|SIMPLE_SEGMENT|2594,2597|false|false|false|C0001861;C3536832|Air (substance);air|air
Finding|Finding|SIMPLE_SEGMENT|2594,2597|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|SIMPLE_SEGMENT|2594,2597|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|SIMPLE_SEGMENT|2594,2597|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|2594,2606|false|false|false|C0001868|Air Movements|air movement
Event|Event|SIMPLE_SEGMENT|2598,2606|false|false|false|||movement
Finding|Organism Function|SIMPLE_SEGMENT|2598,2606|false|false|false|C0026649|Movement|movement
Finding|Idea or Concept|SIMPLE_SEGMENT|2608,2619|false|false|false|C0750502|Significant|significant
Event|Event|SIMPLE_SEGMENT|2620,2628|true|false|false|||wheezing
Finding|Sign or Symptom|SIMPLE_SEGMENT|2620,2628|true|false|false|C0043144|Wheezing|wheezing
Event|Event|SIMPLE_SEGMENT|2644,2651|true|false|false|||rhonchi
Finding|Finding|SIMPLE_SEGMENT|2644,2651|true|false|false|C0035508|Rhonchi|rhonchi
Event|Event|SIMPLE_SEGMENT|2656,2664|true|false|false|||crackles
Finding|Finding|SIMPLE_SEGMENT|2656,2664|true|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2667,2674|true|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2667,2674|true|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Event|Event|SIMPLE_SEGMENT|2667,2674|true|false|false|||ABDOMEN
Finding|Finding|SIMPLE_SEGMENT|2667,2674|true|false|false|C0941288|Abdomen problem|ABDOMEN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2676,2680|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Event|Event|SIMPLE_SEGMENT|2676,2680|false|false|false|||Soft
Event|Event|SIMPLE_SEGMENT|2682,2686|false|false|false|||NTND
Event|Event|SIMPLE_SEGMENT|2691,2694|true|false|false|||HSM
Finding|Gene or Genome|SIMPLE_SEGMENT|2691,2694|true|false|false|C1537594|LRRC4B gene|HSM
Event|Event|SIMPLE_SEGMENT|2698,2708|true|false|false|||tenderness
Finding|Mental Process|SIMPLE_SEGMENT|2698,2708|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|SIMPLE_SEGMENT|2698,2708|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2712,2723|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Procedure|Health Care Activity|SIMPLE_SEGMENT|2757,2766|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|SIMPLE_SEGMENT|2767,2771|false|false|false|||LABS
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2767,2771|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2785,2790|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|2785,2790|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|2785,2790|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|2791,2794|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|2799,2802|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2799,2802|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2799,2802|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2808,2811|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2808,2811|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|2808,2811|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2808,2811|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2817,2820|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2817,2820|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|2828,2831|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|2828,2831|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2828,2831|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2828,2831|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2828,2831|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|2836,2839|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2836,2839|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|2836,2839|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|2836,2839|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|2836,2839|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2836,2839|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2846,2850|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2879,2882|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2899,2904|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|2899,2904|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|2899,2904|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|2917,2923|false|false|false|C0024202|Lymph|Lymphs
Drug|Antibiotic|SIMPLE_SEGMENT|2929,2934|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|2929,2934|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|SIMPLE_SEGMENT|2929,2934|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2941,2944|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|Eos
Event|Event|SIMPLE_SEGMENT|2941,2944|false|false|false|||Eos
Finding|Gene or Genome|SIMPLE_SEGMENT|2941,2944|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|Eos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3049,3054|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3049,3054|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3049,3054|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3059,3062|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|SIMPLE_SEGMENT|3059,3062|false|false|false|||PTT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3059,3062|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3084,3089|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3084,3089|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3084,3089|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|3084,3097|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3084,3097|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3084,3097|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3090,3097|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|3090,3097|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3090,3097|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|3090,3097|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3090,3097|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3090,3097|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|SIMPLE_SEGMENT|3143,3147|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3143,3147|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3143,3147|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3172,3177|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3172,3177|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3172,3177|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3172,3185|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3178,3185|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|3178,3185|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|3178,3185|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3178,3185|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|3178,3185|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|SIMPLE_SEGMENT|3178,3185|false|false|false|||Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|3178,3185|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3178,3185|false|false|false|C0201925|Calcium measurement|Calcium
Event|Event|SIMPLE_SEGMENT|3217,3221|false|false|false|||LABS
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3217,3221|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3235,3240|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3235,3240|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3235,3240|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3267,3272|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3267,3272|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3267,3272|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3273,3278|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|SIMPLE_SEGMENT|3273,3278|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|SIMPLE_SEGMENT|3273,3278|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3273,3278|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3307,3312|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3307,3312|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3307,3312|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3336,3339|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3336,3339|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Drug|Hormone|SIMPLE_SEGMENT|3336,3339|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3336,3339|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Event|Event|SIMPLE_SEGMENT|3336,3339|false|false|false|||TRF
Finding|Gene or Genome|SIMPLE_SEGMENT|3336,3339|false|false|false|C1334121;C1336604;C1705002|IL5 gene;TERF1 gene;TERF1 wt Allele|TRF
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3356,3361|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3356,3361|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3356,3361|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3362,3365|false|false|false|C2708739||TSH
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3362,3365|false|false|false|C0040160|thyrotropin|TSH
Drug|Hormone|SIMPLE_SEGMENT|3362,3365|false|false|false|C0040160|thyrotropin|TSH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3362,3365|false|false|false|C0040160|thyrotropin|TSH
Event|Event|SIMPLE_SEGMENT|3362,3365|false|false|false|||TSH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3362,3365|false|false|false|C0202230|Thyroid stimulating hormone measurement|TSH
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3383,3388|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3383,3388|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3383,3388|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Event|Event|SIMPLE_SEGMENT|3393,3396|false|false|false|||pO2
Finding|Classification|SIMPLE_SEGMENT|3393,3396|false|false|false|C0391840;C4521535|Partial pressure of Oxygen;US Military enlisted E5|pO2
Finding|Molecular Function|SIMPLE_SEGMENT|3393,3396|false|false|false|C0391840;C4521535|Partial pressure of Oxygen;US Military enlisted E5|pO2
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3393,3396|false|false|false|C1283004|PO2 measurement|pO2
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3401,3405|false|false|false|C0391839|Carbon dioxide, partial pressure|pCO2
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3401,3405|false|false|false|C0201931|Carbon dioxide measurement, partial pressure|pCO2
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3431,3435|false|false|false|C2987514|Anatomical base|Base
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3431,3435|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|Base
Drug|Chemical Viewed Functionally|SIMPLE_SEGMENT|3431,3435|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|Base
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|3431,3435|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|Base
Finding|Gene or Genome|SIMPLE_SEGMENT|3431,3435|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|Base
Finding|Idea or Concept|SIMPLE_SEGMENT|3431,3435|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|Base
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3458,3463|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3458,3463|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3458,3463|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Event|Event|SIMPLE_SEGMENT|3468,3472|false|false|false|||FREE
Finding|Functional Concept|SIMPLE_SEGMENT|3468,3472|false|false|false|C0332296|Free of (attribute)|FREE
Finding|Intellectual Product|SIMPLE_SEGMENT|3474,3480|false|false|false|C1552596;C3244286|Direct - PostalAddressUse;direct address|DIRECT
Event|Event|SIMPLE_SEGMENT|3481,3489|false|false|false|||DIALYSIS
Finding|Functional Concept|SIMPLE_SEGMENT|3481,3489|false|false|false|C4723631|Dialysis Method of Administration|DIALYSIS
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3481,3489|false|false|false|C0011945|Physical Dialysis|DIALYSIS
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3481,3489|false|false|false|C0011946;C4551529|Dialysis procedure;Renal Dialysis|DIALYSIS
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3490,3494|false|false|false|C4318744|Test - temporal region|Test
Event|Event|SIMPLE_SEGMENT|3490,3494|false|false|false|||Test
Finding|Functional Concept|SIMPLE_SEGMENT|3490,3494|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|Test
Finding|Intellectual Product|SIMPLE_SEGMENT|3490,3494|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|Test
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3490,3494|false|false|false|C0456984|Test Result|Test
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3490,3494|false|false|false|C0022885|Laboratory Procedures|Test
Finding|Body Substance|SIMPLE_SEGMENT|3498,3507|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|3498,3507|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|3498,3507|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|3498,3507|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|SIMPLE_SEGMENT|3508,3512|false|false|false|||LABS
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3508,3512|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3530,3535|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3530,3535|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3530,3535|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|3536,3539|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|3546,3549|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3546,3549|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3546,3549|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3555,3558|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3555,3558|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|3555,3558|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3555,3558|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3564,3567|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3564,3567|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|3575,3578|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|3575,3578|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3575,3578|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3575,3578|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3575,3578|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|3583,3586|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3583,3586|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|3583,3586|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|3583,3586|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|3583,3586|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3583,3586|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3593,3597|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3626,3629|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3646,3651|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3646,3651|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3646,3651|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|3646,3659|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3646,3659|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3646,3659|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3652,3659|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|3652,3659|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3652,3659|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|3652,3659|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3652,3659|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3652,3659|false|false|false|C0337438|Glucose measurement|Glucose
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3733,3738|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3733,3738|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3733,3738|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3733,3746|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3739,3746|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|3739,3746|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|3739,3746|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3739,3746|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|3739,3746|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|SIMPLE_SEGMENT|3739,3746|false|false|false|||Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|3739,3746|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3739,3746|false|false|false|C0201925|Calcium measurement|Calcium
Event|Event|SIMPLE_SEGMENT|3768,3775|false|false|false|||IMAGING
Finding|Finding|SIMPLE_SEGMENT|3768,3775|false|false|false|C0740845|Imaging problem|IMAGING
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3768,3775|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|IMAGING
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3781,3786|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|SIMPLE_SEGMENT|3781,3786|false|false|false|C0741025|Chest problem|Chest
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3781,3792|false|false|false|C0039985|Plain chest X-ray|Chest X ray
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3787,3792|false|false|false|C0043309|Roentgen Rays|X ray
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3787,3792|false|false|false|C1306645;C1962945|Plain x-ray;Radiographic imaging procedure|X ray
Event|Event|SIMPLE_SEGMENT|3789,3792|false|false|false|||ray
Finding|Gene or Genome|SIMPLE_SEGMENT|3789,3792|false|false|false|C1428870;C5444437|RAB35 wt Allele;SH3YL1 gene|ray
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3789,3792|false|false|false|C0851346|Radiation|ray
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3794,3802|false|false|false|C3172260||Relative
Finding|Idea or Concept|SIMPLE_SEGMENT|3794,3802|false|false|false|C1546849|Living Arrangement - Relative|Relative
Event|Event|SIMPLE_SEGMENT|3803,3811|false|false|false|||increase
Finding|Functional Concept|SIMPLE_SEGMENT|3803,3811|false|false|false|C0442805|Increase|increase
Event|Event|SIMPLE_SEGMENT|3815,3822|false|false|false|||opacity
Finding|Finding|SIMPLE_SEGMENT|3815,3822|false|false|false|C0029053;C1265876|Abnormally opaque structure (morphologic abnormality);Decreased translucency|opacity
Finding|Pathologic Function|SIMPLE_SEGMENT|3815,3822|false|false|false|C0029053;C1265876|Abnormally opaque structure (morphologic abnormality);Decreased translucency|opacity
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3832,3836|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3832,3836|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3832,3836|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|SIMPLE_SEGMENT|3832,3836|false|false|false|C0740941|Lung Problem|lung
Drug|Chemical Viewed Functionally|SIMPLE_SEGMENT|3838,3843|false|false|false|C0178499|Base|bases
Event|Event|SIMPLE_SEGMENT|3838,3843|false|false|false|||bases
Event|Event|SIMPLE_SEGMENT|3856,3860|false|false|false|||felt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3878,3882|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3878,3889|false|false|false|C0225317;C4532079|Neck+Chest>Soft tissue;soft tissue|soft tissue
Anatomy|Tissue|SIMPLE_SEGMENT|3878,3889|false|false|false|C0225317;C4532079|Neck+Chest>Soft tissue;soft tissue|soft tissue
Anatomy|Tissue|SIMPLE_SEGMENT|3883,3889|false|false|false|C0040300|Body tissue|tissue
Finding|Intellectual Product|SIMPLE_SEGMENT|3883,3889|false|true|false|C1547928|Tissue Specimen Code|tissue
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3903,3916|false|false|false|C0521530|Lung consolidation|consolidation
Event|Event|SIMPLE_SEGMENT|3903,3916|false|false|false|||consolidation
Event|Event|SIMPLE_SEGMENT|3939,3946|false|false|false|||helpful
Event|Event|SIMPLE_SEGMENT|3951,3963|false|false|false|||confirmation
Finding|Finding|SIMPLE_SEGMENT|3951,3963|false|false|false|C0750484;C1611825|Confirmation;confirmation - ResponseLevel|confirmation
Finding|Intellectual Product|SIMPLE_SEGMENT|3951,3963|false|false|false|C0750484;C1611825|Confirmation;confirmation - ResponseLevel|confirmation
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3970,3975|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|SIMPLE_SEGMENT|3970,3975|false|false|false|C0741025|Chest problem|Chest
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3970,3981|false|false|false|C0039985|Plain chest X-ray|Chest X ray
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3976,3981|false|false|false|C0043309|Roentgen Rays|X ray
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3976,3981|false|false|false|C1306645;C1962945|Plain x-ray;Radiographic imaging procedure|X ray
Event|Event|SIMPLE_SEGMENT|3978,3981|false|false|false|||ray
Finding|Gene or Genome|SIMPLE_SEGMENT|3978,3981|false|false|false|C1428870;C5444437|RAB35 wt Allele;SH3YL1 gene|ray
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3978,3981|false|false|false|C0851346|Radiation|ray
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|3992,4006|false|false|false|C0020449|Hyperdistention|hyperinflation
Event|Event|SIMPLE_SEGMENT|3992,4006|false|false|false|||hyperinflation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4022,4034|true|false|false|C0032326|Pneumothorax|pneumothorax
Event|Event|SIMPLE_SEGMENT|4022,4034|true|false|false|||pneumothorax
Event|Event|SIMPLE_SEGMENT|4036,4044|true|false|false|||effusion
Finding|Body Substance|SIMPLE_SEGMENT|4036,4044|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|SIMPLE_SEGMENT|4036,4044|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|4036,4044|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4046,4059|true|false|false|C0521530|Lung consolidation|consolidation
Event|Event|SIMPLE_SEGMENT|4046,4059|true|false|false|||consolidation
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4063,4066|false|false|false|C0262212|Choroidal fissure|CHF
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4063,4066|false|false|false|C0018802|Congestive heart failure|CHF
Event|Event|SIMPLE_SEGMENT|4063,4066|false|false|false|||CHF
Event|Event|SIMPLE_SEGMENT|4078,4086|false|false|false|||probable
Finding|Finding|SIMPLE_SEGMENT|4078,4086|false|false|false|C0332148|Probable diagnosis|probable
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4088,4098|false|false|false|C0029453|Osteopenia|osteopenia
Event|Event|SIMPLE_SEGMENT|4088,4098|false|false|false|||osteopenia
Finding|Intellectual Product|SIMPLE_SEGMENT|4102,4107|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|Brief
Finding|Idea or Concept|SIMPLE_SEGMENT|4108,4116|false|false|false|C1547192|Organization unit type - Hospital|Hospital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4108,4123|false|false|false|C0488549||Hospital Course
Finding|Finding|SIMPLE_SEGMENT|4108,4123|false|false|false|C0489547|Hospital course|Hospital Course
Event|Event|SIMPLE_SEGMENT|4145,4152|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|4145,4152|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|4145,4152|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|4145,4152|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|4145,4155|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4156,4159|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4156,4159|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|4156,4159|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|4156,4159|false|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|4156,4159|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4156,4159|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|4156,4159|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4156,4159|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4161,4164|false|false|false|C0085096|Peripheral Vascular Diseases|PVD
Event|Event|SIMPLE_SEGMENT|4161,4164|false|false|false|||PVD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4161,4164|false|false|false|C4521226|Pomalidomide/Bortezomib/Dexamethasone Regimen|PVD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4171,4175|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4171,4175|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|SIMPLE_SEGMENT|4171,4175|false|false|false|||COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|4171,4175|false|false|false|C1412502|ARCN1 gene|COPD
Event|Event|SIMPLE_SEGMENT|4180,4187|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|4180,4187|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|4180,4187|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|4180,4187|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|4180,4190|false|false|false|C0262926|Medical History|history of
Event|Event|SIMPLE_SEGMENT|4191,4200|false|false|false|||recurrent
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4201,4206|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|4201,4206|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4201,4211|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|4201,4211|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4207,4211|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|4207,4211|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|4207,4211|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|4207,4211|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|4216,4225|false|false|false|||presented
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4231,4235|false|false|false|C0004238|Atrial Fibrillation|afib
Event|Event|SIMPLE_SEGMENT|4231,4235|false|false|false|||afib
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4231,4235|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|afib
Event|Event|SIMPLE_SEGMENT|4242,4245|false|false|false|||RVR
Finding|Finding|SIMPLE_SEGMENT|4242,4245|false|false|false|C1417822;C3540498;C4050414|NR1D2 gene;NR1D2 wt Allele;Rapid Virologic Response|RVR
Finding|Gene or Genome|SIMPLE_SEGMENT|4242,4245|false|false|false|C1417822;C3540498;C4050414|NR1D2 gene;NR1D2 wt Allele;Rapid Virologic Response|RVR
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4250,4254|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4250,4254|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|SIMPLE_SEGMENT|4250,4254|false|false|false|||COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|4250,4254|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4250,4267|false|false|false|C0740304|COPD exacerbation|COPD exacerbation
Event|Event|SIMPLE_SEGMENT|4255,4267|false|false|false|||exacerbation
Finding|Finding|SIMPLE_SEGMENT|4255,4267|false|false|false|C4086268|Exacerbation|exacerbation
Finding|Intellectual Product|SIMPLE_SEGMENT|4273,4278|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|ACUTE
Event|Event|SIMPLE_SEGMENT|4279,4287|false|false|false|||PROBLEMS
Finding|Idea or Concept|SIMPLE_SEGMENT|4279,4287|false|false|false|C1546466|Problems - What subject filter|PROBLEMS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4291,4295|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4291,4295|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|SIMPLE_SEGMENT|4291,4295|false|false|false|||COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|4291,4295|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4291,4308|false|false|false|C0740304|COPD exacerbation|COPD exacerbation
Event|Event|SIMPLE_SEGMENT|4296,4308|false|false|false|||exacerbation
Finding|Finding|SIMPLE_SEGMENT|4296,4308|false|false|false|C4086268|Exacerbation|exacerbation
Event|Event|SIMPLE_SEGMENT|4340,4346|false|false|false|||visits
Finding|Social Behavior|SIMPLE_SEGMENT|4340,4346|false|false|false|C0545082|Visit|visits
Procedure|Health Care Activity|SIMPLE_SEGMENT|4340,4346|false|false|false|C1512346|Patient Visit|visits
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4352,4356|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4352,4356|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|SIMPLE_SEGMENT|4352,4356|false|false|false|||COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|4352,4356|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4352,4369|false|false|false|C0740304|COPD exacerbation|COPD exacerbation
Event|Event|SIMPLE_SEGMENT|4357,4369|false|false|false|||exacerbation
Finding|Finding|SIMPLE_SEGMENT|4357,4369|false|false|false|C4086268|Exacerbation|exacerbation
Event|Event|SIMPLE_SEGMENT|4402,4409|false|false|false|||started
Drug|Hormone|SIMPLE_SEGMENT|4414,4424|false|false|false|C0032952|prednisone|prednisone
Drug|Organic Chemical|SIMPLE_SEGMENT|4414,4424|false|false|false|C0032952|prednisone|prednisone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4414,4424|false|false|false|C0032952|prednisone|prednisone
Event|Event|SIMPLE_SEGMENT|4436,4445|false|false|false|||presented
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4453,4456|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|4453,4456|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4453,4456|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4453,4456|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|SIMPLE_SEGMENT|4453,4456|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|4453,4456|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|SIMPLE_SEGMENT|4453,4456|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4453,4456|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|SIMPLE_SEGMENT|4453,4456|false|false|false|||PCP
Finding|Gene or Genome|SIMPLE_SEGMENT|4453,4456|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|SIMPLE_SEGMENT|4453,4456|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Event|SIMPLE_SEGMENT|4459,4465|false|false|false|||office
Finding|Idea or Concept|SIMPLE_SEGMENT|4459,4465|false|false|false|C1549636|Address type - Office|office
Event|Event|SIMPLE_SEGMENT|4482,4489|false|false|false|||dyspnea
Finding|Finding|SIMPLE_SEGMENT|4482,4489|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|4482,4489|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Event|Event|SIMPLE_SEGMENT|4503,4510|false|false|false|||therapy
Finding|Finding|SIMPLE_SEGMENT|4503,4510|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|SIMPLE_SEGMENT|4503,4510|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4503,4510|false|false|false|C0087111|Therapeutic procedure|therapy
Event|Event|SIMPLE_SEGMENT|4524,4535|false|false|false|||complaining
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4540,4545|false|false|false|C0028429||nasal
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4540,4545|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Organic Chemical|SIMPLE_SEGMENT|4540,4545|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4540,4545|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Finding|Finding|SIMPLE_SEGMENT|4540,4545|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Functional Concept|SIMPLE_SEGMENT|4540,4545|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Sign or Symptom|SIMPLE_SEGMENT|4540,4556|false|false|false|C0027424|Nasal congestion (finding)|nasal congestion
Event|Event|SIMPLE_SEGMENT|4546,4556|false|false|false|||congestion
Finding|Pathologic Function|SIMPLE_SEGMENT|4546,4556|false|false|false|C0700148|Congestion|congestion
Event|Event|SIMPLE_SEGMENT|4558,4568|false|false|false|||suggesting
Finding|Functional Concept|SIMPLE_SEGMENT|4571,4576|false|false|false|C0521026|Viral|viral
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4577,4580|false|false|false|C0041912|Upper Respiratory Infections|URI
Event|Event|SIMPLE_SEGMENT|4577,4580|false|false|false|||URI
Finding|Gene or Genome|SIMPLE_SEGMENT|4577,4580|false|false|false|C1421895;C1548524;C3272713|URI1 gene;URI1 wt Allele;Uniform Resource Identifier|URI
Finding|Intellectual Product|SIMPLE_SEGMENT|4577,4580|false|false|false|C1421895;C1548524;C3272713|URI1 gene;URI1 wt Allele;Uniform Resource Identifier|URI
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4581,4588|false|false|false|C0032930|Precipitating Factors|trigger
Event|Event|SIMPLE_SEGMENT|4581,4588|false|false|false|||trigger
Event|Event|SIMPLE_SEGMENT|4614,4619|false|false|false|||noted
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4629,4633|false|false|false|C0004238|Atrial Fibrillation|afib
Event|Event|SIMPLE_SEGMENT|4629,4633|false|false|false|||afib
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4629,4633|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|afib
Event|Event|SIMPLE_SEGMENT|4639,4642|false|false|false|||RVR
Finding|Finding|SIMPLE_SEGMENT|4639,4642|false|false|false|C1417822;C3540498;C4050414|NR1D2 gene;NR1D2 wt Allele;Rapid Virologic Response|RVR
Finding|Gene or Genome|SIMPLE_SEGMENT|4639,4642|false|false|false|C1417822;C3540498;C4050414|NR1D2 gene;NR1D2 wt Allele;Rapid Virologic Response|RVR
Event|Event|SIMPLE_SEGMENT|4650,4658|false|false|false|||referred
Event|Event|SIMPLE_SEGMENT|4667,4669|false|false|false|||ED
Event|Event|SIMPLE_SEGMENT|4684,4692|false|false|false|||admitted
Drug|Organic Chemical|SIMPLE_SEGMENT|4699,4706|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4699,4706|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Substance|SIMPLE_SEGMENT|4699,4706|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Event|Event|SIMPLE_SEGMENT|4699,4706|false|false|false|||control
Finding|Conceptual Entity|SIMPLE_SEGMENT|4699,4706|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Functional Concept|SIMPLE_SEGMENT|4699,4706|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Idea or Concept|SIMPLE_SEGMENT|4699,4706|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4714,4719|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4714,4719|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|4714,4719|false|false|false|C0795691|HEART PROBLEM|heart
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4714,4724|false|false|false|C0018810;C0488794|heart rate|heart rate
Finding|Finding|SIMPLE_SEGMENT|4714,4724|false|false|false|C2041121||heart rate
Procedure|Health Care Activity|SIMPLE_SEGMENT|4714,4724|false|false|false|C2197023|examination of heart rate|heart rate
Event|Activity|SIMPLE_SEGMENT|4720,4724|false|false|false|C0871208|Rating (action)|rate
Event|Event|SIMPLE_SEGMENT|4720,4724|false|false|false|||rate
Finding|Idea or Concept|SIMPLE_SEGMENT|4720,4724|false|false|false|C1549480|Amount type - Rate|rate
Event|Event|SIMPLE_SEGMENT|4726,4729|false|false|false|||see
Event|Event|SIMPLE_SEGMENT|4742,4751|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|4742,4751|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|4759,4764|false|false|false|C3714591|Floor (anatomic)|floor
Event|Event|SIMPLE_SEGMENT|4774,4779|false|false|false|||noted
Event|Event|SIMPLE_SEGMENT|4789,4797|false|false|false|||wheezing
Finding|Sign or Symptom|SIMPLE_SEGMENT|4789,4797|false|false|false|C0043144|Wheezing|wheezing
Event|Event|SIMPLE_SEGMENT|4799,4808|false|false|false|||increased
Finding|Finding|SIMPLE_SEGMENT|4799,4808|false|false|false|C0442805;C5236002|Increase;Increased (finding)|increased
Finding|Functional Concept|SIMPLE_SEGMENT|4799,4808|false|false|false|C0442805;C5236002|Increase;Increased (finding)|increased
Finding|Sign or Symptom|SIMPLE_SEGMENT|4799,4826|false|false|false|C0859927|Increased work of breathing|increased work of breathing
Event|Event|SIMPLE_SEGMENT|4809,4813|false|false|false|||work
Event|Occupational Activity|SIMPLE_SEGMENT|4809,4813|false|false|false|C0043227|Work|work
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|4809,4826|false|false|false|C0043229|Work of Breathing|work of breathing
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4817,4826|false|false|false|C5885990||breathing
Event|Event|SIMPLE_SEGMENT|4817,4826|false|false|false|||breathing
Finding|Finding|SIMPLE_SEGMENT|4817,4826|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|SIMPLE_SEGMENT|4817,4826|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|SIMPLE_SEGMENT|4817,4826|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|SIMPLE_SEGMENT|4817,4826|false|false|false|C1160636|respiratory system process|breathing
Finding|Intellectual Product|SIMPLE_SEGMENT|4832,4836|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|poor
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4837,4840|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4837,4840|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|SIMPLE_SEGMENT|4837,4840|false|false|false|C0001861;C3536832|Air (substance);air|air
Finding|Finding|SIMPLE_SEGMENT|4837,4840|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|SIMPLE_SEGMENT|4837,4840|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|SIMPLE_SEGMENT|4837,4840|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|4837,4849|false|false|false|C0001868|Air Movements|air movement
Event|Event|SIMPLE_SEGMENT|4841,4849|false|false|false|||movement
Finding|Organism Function|SIMPLE_SEGMENT|4841,4849|false|false|false|C0026649|Movement|movement
Event|Event|SIMPLE_SEGMENT|4860,4867|false|false|false|||treated
Drug|Organic Chemical|SIMPLE_SEGMENT|4880,4890|false|false|false|C0701466|Solu-Medrol|solumedrol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4880,4890|false|false|false|C0701466|Solu-Medrol|solumedrol
Event|Event|SIMPLE_SEGMENT|4880,4890|false|false|false|||solumedrol
Event|Event|SIMPLE_SEGMENT|4895,4905|false|false|false|||maintained
Drug|Hormone|SIMPLE_SEGMENT|4919,4929|false|false|false|C0032952|prednisone|prednisone
Drug|Organic Chemical|SIMPLE_SEGMENT|4919,4929|false|false|false|C0032952|prednisone|prednisone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4919,4929|false|false|false|C0032952|prednisone|prednisone
Event|Event|SIMPLE_SEGMENT|4919,4929|false|false|false|||prednisone
Finding|Idea or Concept|SIMPLE_SEGMENT|4941,4945|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|4941,4945|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|4941,4945|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|4946,4958|false|false|false|C0039771|theophylline|theophylline
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4946,4958|false|false|false|C0039771|theophylline|theophylline
Event|Event|SIMPLE_SEGMENT|4946,4958|false|false|false|||theophylline
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4946,4958|false|false|false|C0039773|Assay of theophylline|theophylline
Event|Event|SIMPLE_SEGMENT|4963,4972|false|false|false|||decreased
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|4986,4989|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4986,4989|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4986,4989|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|4986,4989|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|4986,4989|false|false|false|C1332410|BID gene|BID
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|5000,5003|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5000,5003|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5000,5003|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|5000,5003|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|5000,5003|false|false|false|C1332410|BID gene|BID
Event|Event|SIMPLE_SEGMENT|5011,5019|false|false|false|||concerns
Event|Event|SIMPLE_SEGMENT|5027,5039|false|false|false|||contributing
Event|Event|SIMPLE_SEGMENT|5048,5063|false|false|false|||tachyarrhythmia
Finding|Finding|SIMPLE_SEGMENT|5048,5063|false|false|false|C0080203|Tachyarrhythmia|tachyarrhythmia
Event|Event|SIMPLE_SEGMENT|5073,5079|false|false|false|||placed
Drug|Organic Chemical|SIMPLE_SEGMENT|5083,5094|false|false|false|C0027235|ipratropium|ipratropium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5083,5094|false|false|false|C0027235|ipratropium|ipratropium
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5095,5099|false|false|false|C1300458|Nebulizer solution|nebs
Event|Event|SIMPLE_SEGMENT|5100,5103|false|false|false|||q6h
Drug|Organic Chemical|SIMPLE_SEGMENT|5106,5115|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5106,5115|false|false|false|C0001927|albuterol|albuterol
Event|Event|SIMPLE_SEGMENT|5106,5115|false|false|false|||albuterol
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5116,5120|false|false|false|C1300458|Nebulizer solution|nebs
Event|Event|SIMPLE_SEGMENT|5121,5124|false|false|false|||q2h
Drug|Organic Chemical|SIMPLE_SEGMENT|5130,5141|false|false|false|C0082607|fluticasone|fluticasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5130,5141|false|false|false|C0082607|fluticasone|fluticasone
Event|Event|SIMPLE_SEGMENT|5130,5141|false|false|false|||fluticasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5130,5152|false|false|false|C0939232|fluticasone / salmeterol|fluticasone-salmeterol
Drug|Organic Chemical|SIMPLE_SEGMENT|5142,5152|false|false|false|C0073992|salmeterol|salmeterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5142,5152|false|false|false|C0073992|salmeterol|salmeterol
Event|Event|SIMPLE_SEGMENT|5142,5152|false|false|false|||salmeterol
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5154,5163|false|false|false|C0024109|Lung|Pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5154,5163|false|false|false|C2707265||Pulmonary
Finding|Finding|SIMPLE_SEGMENT|5154,5163|false|false|false|C4522268|Pulmonary (intended site)|Pulmonary
Event|Event|SIMPLE_SEGMENT|5169,5178|false|false|false|||consulted
Event|Event|SIMPLE_SEGMENT|5183,5194|false|false|false|||recommended
Event|Event|SIMPLE_SEGMENT|5197,5202|false|false|false|||trial
Procedure|Research Activity|SIMPLE_SEGMENT|5197,5202|false|false|false|C0008976|Clinical Trials|trial
Event|Event|SIMPLE_SEGMENT|5206,5214|false|false|false|||diuresis
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|5206,5214|false|false|false|C0012797|Diuresis|diuresis
Drug|Organic Chemical|SIMPLE_SEGMENT|5241,5246|false|false|false|C0699992|Lasix|Lasix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5241,5246|false|false|false|C0699992|Lasix|Lasix
Event|Event|SIMPLE_SEGMENT|5241,5246|false|false|false|||Lasix
Finding|Finding|SIMPLE_SEGMENT|5250,5254|false|false|false|C5575035|Well (answer to question)|well
Drug|Antibiotic|SIMPLE_SEGMENT|5256,5268|true|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|Azithromycin
Drug|Clinical Drug|SIMPLE_SEGMENT|5256,5268|true|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|Azithromycin
Drug|Organic Chemical|SIMPLE_SEGMENT|5256,5268|true|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|Azithromycin
Event|Event|SIMPLE_SEGMENT|5256,5268|true|false|false|||Azithromycin
Event|Event|SIMPLE_SEGMENT|5277,5282|true|false|false|||given
Event|Event|SIMPLE_SEGMENT|5290,5298|true|false|false|||concerns
Event|Event|SIMPLE_SEGMENT|5307,5319|false|false|false|||prolongation
Drug|Organic Chemical|SIMPLE_SEGMENT|5325,5337|false|false|false|C0039771|theophylline|theophylline
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5325,5337|false|false|false|C0039771|theophylline|theophylline
Event|Event|SIMPLE_SEGMENT|5325,5337|false|false|false|||theophylline
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5325,5337|false|false|false|C0039773|Assay of theophylline|theophylline
Drug|Organic Chemical|SIMPLE_SEGMENT|5342,5352|false|false|false|C0002598|amiodarone|amiodarone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5342,5352|false|false|false|C0002598|amiodarone|amiodarone
Event|Event|SIMPLE_SEGMENT|5342,5352|false|false|false|||amiodarone
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5342,5352|false|false|false|C5399868|Drug assay amiodarone|amiodarone
Event|Event|SIMPLE_SEGMENT|5377,5384|false|false|false|||started
Finding|Idea or Concept|SIMPLE_SEGMENT|5392,5395|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|5392,5395|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|5396,5402|false|false|false|||course
Drug|Antibiotic|SIMPLE_SEGMENT|5406,5417|false|false|false|C0007561|ceftriaxone|ceftriaxone
Drug|Organic Chemical|SIMPLE_SEGMENT|5406,5417|false|false|false|C0007561|ceftriaxone|ceftriaxone
Event|Event|SIMPLE_SEGMENT|5406,5417|false|false|false|||ceftriaxone
Event|Event|SIMPLE_SEGMENT|5432,5442|false|false|false|||discharged
Event|Event|SIMPLE_SEGMENT|5446,5452|false|false|false|||finish
Event|Event|SIMPLE_SEGMENT|5457,5463|false|false|false|||course
Drug|Antibiotic|SIMPLE_SEGMENT|5469,5480|false|false|false|C0055011|cefpodoxime|cefpodoxime
Drug|Organic Chemical|SIMPLE_SEGMENT|5469,5480|false|false|false|C0055011|cefpodoxime|cefpodoxime
Event|Event|SIMPLE_SEGMENT|5469,5480|false|false|false|||cefpodoxime
Event|Event|SIMPLE_SEGMENT|5491,5501|false|false|false|||discharged
Drug|Hormone|SIMPLE_SEGMENT|5509,5519|false|false|false|C0032952|prednisone|prednisone
Drug|Organic Chemical|SIMPLE_SEGMENT|5509,5519|false|false|false|C0032952|prednisone|prednisone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5509,5519|false|false|false|C0032952|prednisone|prednisone
Event|Event|SIMPLE_SEGMENT|5520,5525|false|false|false|||taper
Procedure|Health Care Activity|SIMPLE_SEGMENT|5520,5525|false|false|false|C0441640||taper
Event|Event|SIMPLE_SEGMENT|5533,5541|false|false|false|||decrease
Finding|Intellectual Product|SIMPLE_SEGMENT|5563,5567|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|SIMPLE_SEGMENT|5568,5572|false|false|false|||stay
Procedure|Health Care Activity|SIMPLE_SEGMENT|5588,5592|false|false|false|C1315068|Pulmonary ventilator management|pulm
Event|Event|SIMPLE_SEGMENT|5593,5599|false|false|false|||follow
Finding|Functional Concept|SIMPLE_SEGMENT|5593,5599|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|SIMPLE_SEGMENT|5593,5599|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|SIMPLE_SEGMENT|5593,5602|false|false|false|C0589120|Follow-up status|follow up
Procedure|Health Care Activity|SIMPLE_SEGMENT|5593,5602|false|false|false|C1522577|follow-up|follow up
Finding|Finding|SIMPLE_SEGMENT|5607,5611|false|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|5616,5622|false|false|false|||follow
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5631,5640|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5631,5640|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|5631,5640|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Event|Event|SIMPLE_SEGMENT|5641,5646|false|false|false|||rehab
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5641,5646|false|false|false|C0034991|Rehabilitation therapy|rehab
Event|Event|SIMPLE_SEGMENT|5720,5730|false|false|false|||discharged
Event|Event|SIMPLE_SEGMENT|5735,5737|false|false|false|||2L
Event|Event|SIMPLE_SEGMENT|5738,5750|false|false|false|||supplemental
Finding|Functional Concept|SIMPLE_SEGMENT|5738,5750|false|false|false|C2348609|Supplement|supplemental
Event|Event|SIMPLE_SEGMENT|5760,5764|false|false|false|||worn
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5772,5777|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5782,5788|false|false|false|C0018792|Heart Atrium|Atrial
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5782,5801|false|false|false|C2926591||Atrial fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5782,5801|false|false|false|C0004238|Atrial Fibrillation|Atrial fibrillation
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5782,5801|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Atrial fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5789,5801|false|false|false|C0232197|Fibrillation|fibrillation
Event|Event|SIMPLE_SEGMENT|5789,5801|false|false|false|||fibrillation
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5821,5827|false|false|false|C0018792|Heart Atrium|atrial
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5829,5841|false|false|false|C0232197|Fibrillation|fibrillation
Event|Event|SIMPLE_SEGMENT|5829,5841|false|false|false|||fibrillation
Drug|Organic Chemical|SIMPLE_SEGMENT|5863,5873|false|false|false|C0002598|amiodarone|amiodarone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5863,5873|false|false|false|C0002598|amiodarone|amiodarone
Event|Event|SIMPLE_SEGMENT|5863,5873|false|false|false|||amiodarone
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5863,5873|false|false|false|C5399868|Drug assay amiodarone|amiodarone
Drug|Organic Chemical|SIMPLE_SEGMENT|5878,5886|false|false|false|C1831808|apixaban|apixaban
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5878,5886|false|false|false|C1831808|apixaban|apixaban
Event|Event|SIMPLE_SEGMENT|5878,5886|false|false|false|||apixaban
Event|Event|SIMPLE_SEGMENT|5896,5901|false|false|false|||found
Event|Event|SIMPLE_SEGMENT|5910,5912|false|false|false|||HR
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5932,5935|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|5932,5935|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5932,5935|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5932,5935|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|SIMPLE_SEGMENT|5932,5935|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|5932,5935|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|SIMPLE_SEGMENT|5932,5935|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5932,5935|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|SIMPLE_SEGMENT|5932,5935|false|false|false|||PCP
Finding|Gene or Genome|SIMPLE_SEGMENT|5932,5935|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|SIMPLE_SEGMENT|5932,5935|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Event|SIMPLE_SEGMENT|5938,5944|false|false|false|||office
Finding|Idea or Concept|SIMPLE_SEGMENT|5938,5944|false|false|false|C1549636|Address type - Office|office
Event|Event|SIMPLE_SEGMENT|5946,5955|false|false|false|||prompting
Finding|Functional Concept|SIMPLE_SEGMENT|5946,5955|false|false|false|C0871157|Prompting|prompting
Event|Event|SIMPLE_SEGMENT|5961,5969|false|false|false|||referral
Procedure|Health Care Activity|SIMPLE_SEGMENT|5961,5969|false|false|false|C0034927|Patient referral|referral
Procedure|Health Care Activity|SIMPLE_SEGMENT|5961,5972|false|false|false|C2585021|Referral to|referral to
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5985,5989|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5985,5989|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|SIMPLE_SEGMENT|5985,5989|false|false|false|||COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|5985,5989|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5985,6002|false|false|false|C0740304|COPD exacerbation|COPD exacerbation
Event|Event|SIMPLE_SEGMENT|5990,6002|false|false|false|||exacerbation
Finding|Finding|SIMPLE_SEGMENT|5990,6002|false|false|false|C4086268|Exacerbation|exacerbation
Event|Event|SIMPLE_SEGMENT|6011,6017|false|false|false|||likely
Finding|Finding|SIMPLE_SEGMENT|6011,6017|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|6011,6017|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6037,6048|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6037,6048|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|6037,6048|false|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|6037,6048|false|false|false|C4284232|Medications|medications
Finding|Finding|SIMPLE_SEGMENT|6054,6062|false|false|false|C0332149|Possible|possibly
Event|Event|SIMPLE_SEGMENT|6063,6075|false|false|false|||contributing
Drug|Organic Chemical|SIMPLE_SEGMENT|6091,6103|false|false|false|C0039771|theophylline|theophylline
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6091,6103|false|false|false|C0039771|theophylline|theophylline
Event|Event|SIMPLE_SEGMENT|6091,6103|false|false|false|||theophylline
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6091,6103|false|false|false|C0039773|Assay of theophylline|theophylline
Event|Event|SIMPLE_SEGMENT|6113,6120|false|false|false|||started
Drug|Organic Chemical|SIMPLE_SEGMENT|6126,6135|false|false|false|C0012373|diltiazem|diltiazem
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6126,6135|false|false|false|C0012373|diltiazem|diltiazem
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6136,6139|false|false|false|C1135868|Gestational Trophoblastic Neoplasms|gtt
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6136,6139|false|false|false|C0991568|Drops - Drug Form|gtt
Event|Event|SIMPLE_SEGMENT|6136,6139|false|false|false|||gtt
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6136,6139|false|false|false|C0017741|Glucose tolerance test|gtt
Event|Event|SIMPLE_SEGMENT|6154,6161|false|false|false|||control
Event|Event|SIMPLE_SEGMENT|6166,6171|false|false|false|||rates
Event|Event|SIMPLE_SEGMENT|6177,6189|false|false|false|||transitioned
Drug|Organic Chemical|SIMPLE_SEGMENT|6193,6202|false|false|false|C0012373|diltiazem|diltiazem
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6193,6202|false|false|false|C0012373|diltiazem|diltiazem
Event|Event|SIMPLE_SEGMENT|6193,6202|false|false|false|||diltiazem
Event|Event|SIMPLE_SEGMENT|6210,6213|false|false|false|||q6h
Event|Activity|SIMPLE_SEGMENT|6221,6228|false|false|false|C1706079||arrival
Event|Event|SIMPLE_SEGMENT|6221,6228|false|false|false|||arrival
Finding|Functional Concept|SIMPLE_SEGMENT|6221,6228|false|false|false|C1555577|arrival - ActRelationshipType|arrival
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|6236,6241|false|false|false|C3714591|Floor (anatomic)|floor
Event|Event|SIMPLE_SEGMENT|6253,6261|false|false|false|||remained
Event|Event|SIMPLE_SEGMENT|6262,6272|false|false|false|||controlled
Drug|Organic Chemical|SIMPLE_SEGMENT|6279,6289|false|false|false|C0002598|amiodarone|amiodarone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6279,6289|false|false|false|C0002598|amiodarone|amiodarone
Event|Event|SIMPLE_SEGMENT|6279,6289|false|false|false|||amiodarone
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6279,6289|false|false|false|C5399868|Drug assay amiodarone|amiodarone
Drug|Organic Chemical|SIMPLE_SEGMENT|6294,6302|false|false|false|C1831808|apixaban|apixaban
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6294,6302|false|false|false|C1831808|apixaban|apixaban
Event|Event|SIMPLE_SEGMENT|6294,6302|false|false|false|||apixaban
Event|Event|SIMPLE_SEGMENT|6308,6317|false|false|false|||continued
Drug|Organic Chemical|SIMPLE_SEGMENT|6323,6335|false|false|false|C0039771|theophylline|theophylline
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6323,6335|false|false|false|C0039771|theophylline|theophylline
Event|Event|SIMPLE_SEGMENT|6323,6335|false|false|false|||theophylline
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6323,6335|false|false|false|C0039773|Assay of theophylline|theophylline
Event|Event|SIMPLE_SEGMENT|6341,6350|false|false|false|||decreased
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|6361,6364|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6361,6364|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6361,6364|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|6361,6364|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|6361,6364|false|false|false|C1332410|BID gene|BID
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|6377,6380|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6377,6380|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6377,6380|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|6377,6380|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|6377,6380|false|false|false|C1332410|BID gene|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6384,6388|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|6384,6388|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6384,6388|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6384,6388|false|false|false|C0337439|Iron measurement|Iron
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6384,6399|false|false|false|C0162316;C0240066|Iron deficiency;Iron deficiency anemia|Iron deficiency
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6384,6406|false|false|false|C0162316|Iron deficiency anemia|Iron deficiency anemia
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6389,6399|false|false|false|C0162429|Malnutrition|deficiency
Event|Event|SIMPLE_SEGMENT|6389,6399|false|false|false|||deficiency
Finding|Functional Concept|SIMPLE_SEGMENT|6389,6399|false|false|false|C0011155|Deficiency|deficiency
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6389,6406|false|false|false|C0041782|Deficiency anemias|deficiency anemia
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6400,6406|false|false|false|C0002871|Anemia|anemia
Event|Event|SIMPLE_SEGMENT|6400,6406|false|false|false|||anemia
Finding|Body Substance|SIMPLE_SEGMENT|6408,6415|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|6408,6415|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|6408,6415|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|6420,6425|false|false|false|||found
Event|Event|SIMPLE_SEGMENT|6434,6444|false|false|false|||microcytic
Finding|Finding|SIMPLE_SEGMENT|6434,6444|false|false|false|C0302870|microcytic|microcytic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6446,6452|false|false|false|C0002871|Anemia|anemia
Event|Event|SIMPLE_SEGMENT|6446,6452|false|false|false|||anemia
Finding|Finding|SIMPLE_SEGMENT|6458,6461|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|SIMPLE_SEGMENT|6458,6461|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Finding|SIMPLE_SEGMENT|6458,6466|false|false|false|C0860975|Iron low|low iron
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6462,6466|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|6462,6466|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6462,6466|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Event|Event|SIMPLE_SEGMENT|6462,6466|false|false|false|||iron
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6462,6466|false|false|false|C0337439|Iron measurement|iron
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6471,6479|false|false|false|C0015879|Ferritin|ferritin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6471,6479|false|false|false|C0015879|Ferritin|ferritin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6471,6479|false|false|false|C0015879|Ferritin|ferritin
Event|Event|SIMPLE_SEGMENT|6471,6479|false|false|false|||ferritin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6471,6479|false|false|false|C0373607|Ferritin measurement|ferritin
Event|Event|SIMPLE_SEGMENT|6489,6496|false|false|false|||started
Finding|Finding|SIMPLE_SEGMENT|6497,6502|false|false|false|C3714655|On IV|on IV
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|6500,6507|false|false|false|C0082568|ferryl iron|IV iron
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6503,6507|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|6503,6507|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6503,6507|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Event|Event|SIMPLE_SEGMENT|6503,6507|false|false|false|||iron
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6503,6507|false|false|false|C0337439|Iron measurement|iron
Drug|Inorganic Chemical|SIMPLE_SEGMENT|6516,6522|false|false|false|C3848561|ferric cation|ferric
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6516,6522|false|false|false|C3848561|ferric cation|ferric
Drug|Organic Chemical|SIMPLE_SEGMENT|6516,6532|false|false|false|C0060235|ferric gluconate|ferric gluconate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6516,6532|false|false|false|C0060235|ferric gluconate|ferric gluconate
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6523,6532|false|false|false|C0017714;C0220836|Gluconates;gluconate|gluconate
Drug|Organic Chemical|SIMPLE_SEGMENT|6523,6532|false|false|false|C0017714;C0220836|Gluconates;gluconate|gluconate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6523,6532|false|false|false|C0017714;C0220836|Gluconates;gluconate|gluconate
Event|Event|SIMPLE_SEGMENT|6523,6532|false|false|false|||gluconate
Event|Event|SIMPLE_SEGMENT|6536,6541|false|false|false|||doses
Event|Event|SIMPLE_SEGMENT|6546,6559|false|false|false|||wasdischarged
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6566,6570|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|6566,6570|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6566,6570|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Event|Event|SIMPLE_SEGMENT|6566,6570|false|false|false|||iron
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6566,6570|false|false|false|C0337439|Iron measurement|iron
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6579,6584|false|false|false|C0021853|Intestines|bowel
Procedure|Health Care Activity|SIMPLE_SEGMENT|6579,6592|false|false|false|C5979615|Bowel Regimen|bowel regimen
Event|Event|SIMPLE_SEGMENT|6585,6592|false|false|false|||regimen
Finding|Intellectual Product|SIMPLE_SEGMENT|6585,6592|false|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6585,6592|false|false|false|C0040808|Treatment Protocols|regimen
Event|Event|SIMPLE_SEGMENT|6606,6612|false|false|false|||stable
Finding|Intellectual Product|SIMPLE_SEGMENT|6606,6612|false|false|false|C1547311|Patient Condition Code - Stable|stable
Event|Event|SIMPLE_SEGMENT|6629,6641|false|false|false|||hospitalized
Event|Event|SIMPLE_SEGMENT|6656,6664|true|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|6656,6664|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|6656,6667|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Event|Event|SIMPLE_SEGMENT|6668,6676|true|false|false|||bleeding
Finding|Pathologic Function|SIMPLE_SEGMENT|6668,6676|true|false|false|C0019080|Hemorrhage|bleeding
Finding|Idea or Concept|SIMPLE_SEGMENT|6679,6691|false|false|false|C1548597|Marketing basis - Transitional|Transitional
Event|Event|SIMPLE_SEGMENT|6692,6698|false|false|false|||issues
Finding|Body Substance|SIMPLE_SEGMENT|6702,6709|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|6702,6709|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|6702,6709|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|6710,6720|false|false|false|||discharged
Drug|Hormone|SIMPLE_SEGMENT|6724,6734|false|false|false|C0032952|prednisone|prednisone
Drug|Organic Chemical|SIMPLE_SEGMENT|6724,6734|false|false|false|C0032952|prednisone|prednisone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6724,6734|false|false|false|C0032952|prednisone|prednisone
Event|Event|SIMPLE_SEGMENT|6735,6740|false|false|false|||taper
Procedure|Health Care Activity|SIMPLE_SEGMENT|6735,6740|false|false|false|C0441640||taper
Event|Event|SIMPLE_SEGMENT|6742,6750|false|false|false|||decrease
Finding|Finding|SIMPLE_SEGMENT|6742,6750|false|false|false|C0392756|Reduced|decrease
Finding|Intellectual Product|SIMPLE_SEGMENT|6790,6794|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|SIMPLE_SEGMENT|6795,6799|false|false|false|||keep
Finding|Body Substance|SIMPLE_SEGMENT|6838,6845|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|6838,6845|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|6838,6845|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|6846,6856|false|false|false|||discharged
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6862,6866|false|false|false|C0270724|Infantile Neuroaxonal Dystrophy|plan
Event|Event|SIMPLE_SEGMENT|6862,6866|false|false|false|||plan
Finding|Functional Concept|SIMPLE_SEGMENT|6862,6866|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Intellectual Product|SIMPLE_SEGMENT|6862,6866|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Mental Process|SIMPLE_SEGMENT|6862,6866|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Event|Event|SIMPLE_SEGMENT|6870,6876|false|false|false|||follow
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6902,6911|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6902,6911|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|6902,6911|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Event|Event|SIMPLE_SEGMENT|6912,6917|false|false|false|||rehab
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6912,6917|false|false|false|C0034991|Rehabilitation therapy|rehab
Event|Event|SIMPLE_SEGMENT|6923,6927|false|false|false|||call
Event|Event|SIMPLE_SEGMENT|6935,6943|false|false|false|||schedule
Event|Activity|SIMPLE_SEGMENT|6944,6955|false|false|false|C0003629|Appointments|appointment
Event|Event|SIMPLE_SEGMENT|6944,6955|false|false|false|||appointment
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6962,6971|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6962,6971|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|6962,6971|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Event|Event|SIMPLE_SEGMENT|6972,6977|false|false|false|||rehab
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6972,6977|false|false|false|C0034991|Rehabilitation therapy|rehab
Finding|Body Substance|SIMPLE_SEGMENT|6981,6988|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|6981,6988|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|6981,6988|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|6989,6999|false|false|false|||discharged
Drug|Antibiotic|SIMPLE_SEGMENT|7018,7029|false|false|false|C0055011|cefpodoxime|cefpodoxime
Drug|Organic Chemical|SIMPLE_SEGMENT|7018,7029|false|false|false|C0055011|cefpodoxime|cefpodoxime
Event|Event|SIMPLE_SEGMENT|7018,7029|false|false|false|||cefpodoxime
Drug|Organic Chemical|SIMPLE_SEGMENT|7033,7041|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7033,7041|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|SIMPLE_SEGMENT|7033,7041|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|SIMPLE_SEGMENT|7033,7041|false|false|false|||complete
Finding|Functional Concept|SIMPLE_SEGMENT|7033,7041|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|SIMPLE_SEGMENT|7033,7041|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|SIMPLE_SEGMENT|7045,7048|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|7045,7048|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|7049,7055|false|false|false|||course
Drug|Antibiotic|SIMPLE_SEGMENT|7059,7070|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|SIMPLE_SEGMENT|7059,7070|false|false|false|||antibiotics
Finding|Finding|SIMPLE_SEGMENT|7075,7081|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|SIMPLE_SEGMENT|7075,7081|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7082,7086|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7082,7086|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|SIMPLE_SEGMENT|7082,7086|false|false|false|||COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|7082,7086|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7082,7099|false|false|false|C0740304|COPD exacerbation|COPD exacerbation
Event|Event|SIMPLE_SEGMENT|7087,7099|false|false|false|||exacerbation
Finding|Finding|SIMPLE_SEGMENT|7087,7099|false|false|false|C4086268|Exacerbation|exacerbation
Finding|Body Substance|SIMPLE_SEGMENT|7102,7109|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|7102,7109|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|7102,7109|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|7110,7120|false|false|false|||discharged
Event|Event|SIMPLE_SEGMENT|7129,7141|false|false|false|||concentrator
Finding|Idea or Concept|SIMPLE_SEGMENT|7146,7156|false|false|false|C0549178|Continuous|continuous
Event|Event|SIMPLE_SEGMENT|7157,7161|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|7157,7161|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|7157,7161|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|7157,7161|false|false|false|C1553498|home health encounter|home
Finding|Body Substance|SIMPLE_SEGMENT|7167,7174|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|7167,7174|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|7167,7174|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Organic Chemical|SIMPLE_SEGMENT|7177,7189|false|false|false|C0039771|theophylline|theophylline
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7177,7189|false|false|false|C0039771|theophylline|theophylline
Event|Event|SIMPLE_SEGMENT|7177,7189|false|false|false|||theophylline
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7177,7189|false|false|false|C0039773|Assay of theophylline|theophylline
Event|Event|SIMPLE_SEGMENT|7190,7199|false|false|false|||decreased
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|7212,7215|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7212,7215|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7212,7215|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|7212,7215|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|7212,7215|false|false|false|C1332410|BID gene|BID
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|7226,7229|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7226,7229|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7226,7229|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|7226,7229|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|7226,7229|false|false|false|C1332410|BID gene|BID
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7242,7246|false|false|false|C0004238|Atrial Fibrillation|afib
Event|Event|SIMPLE_SEGMENT|7242,7246|false|false|false|||afib
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|7242,7246|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|afib
Event|Event|SIMPLE_SEGMENT|7252,7255|false|false|false|||RVR
Finding|Finding|SIMPLE_SEGMENT|7252,7255|false|false|false|C1417822;C3540498;C4050414|NR1D2 gene;NR1D2 wt Allele;Rapid Virologic Response|RVR
Finding|Gene or Genome|SIMPLE_SEGMENT|7252,7255|false|false|false|C1417822;C3540498;C4050414|NR1D2 gene;NR1D2 wt Allele;Rapid Virologic Response|RVR
Event|Event|SIMPLE_SEGMENT|7261,7265|false|false|false|||want
Event|Event|SIMPLE_SEGMENT|7269,7277|false|false|false|||consider
Drug|Organic Chemical|SIMPLE_SEGMENT|7287,7299|false|false|false|C0039771|theophylline|theophylline
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7287,7299|false|false|false|C0039771|theophylline|theophylline
Event|Event|SIMPLE_SEGMENT|7287,7299|false|false|false|||theophylline
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7287,7299|false|false|false|C0039773|Assay of theophylline|theophylline
Event|Event|SIMPLE_SEGMENT|7300,7304|false|false|false|||wean
Finding|Finding|SIMPLE_SEGMENT|7300,7304|false|false|false|C0043084|Weaning|wean
Event|Event|SIMPLE_SEGMENT|7310,7318|false|false|false|||addition
Finding|Functional Concept|SIMPLE_SEGMENT|7310,7318|false|false|false|C0332287;C1883712|Add - instruction imperative;In addition to|addition
Drug|Antibiotic|SIMPLE_SEGMENT|7322,7334|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Clinical Drug|SIMPLE_SEGMENT|7322,7334|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Organic Chemical|SIMPLE_SEGMENT|7322,7334|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Event|Event|SIMPLE_SEGMENT|7322,7334|false|false|false|||azithromycin
Event|Event|SIMPLE_SEGMENT|7347,7356|false|false|false|||decreased
Finding|Body Substance|SIMPLE_SEGMENT|7360,7367|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|7360,7367|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|7360,7367|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Organic Chemical|SIMPLE_SEGMENT|7376,7386|false|false|false|C0002598|amiodarone|amiodarone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7376,7386|false|false|false|C0002598|amiodarone|amiodarone
Event|Event|SIMPLE_SEGMENT|7376,7386|false|false|false|||amiodarone
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7376,7386|false|false|false|C5399868|Drug assay amiodarone|amiodarone
Drug|Organic Chemical|SIMPLE_SEGMENT|7396,7407|false|false|false|C0965618|roflumilast|roflumilast
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7396,7407|false|false|false|C0965618|roflumilast|roflumilast
Event|Event|SIMPLE_SEGMENT|7396,7407|false|false|false|||roflumilast
Event|Event|SIMPLE_SEGMENT|7409,7416|false|false|false|||therapy
Finding|Finding|SIMPLE_SEGMENT|7409,7416|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|SIMPLE_SEGMENT|7409,7416|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7409,7416|false|false|false|C0087111|Therapeutic procedure|therapy
Finding|Body Substance|SIMPLE_SEGMENT|7419,7426|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|7419,7426|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|7419,7426|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|7427,7432|false|false|false|||found
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7439,7443|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|7439,7443|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7439,7443|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Event|Event|SIMPLE_SEGMENT|7439,7443|false|false|false|||iron
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7439,7443|false|false|false|C0337439|Iron measurement|iron
Event|Event|SIMPLE_SEGMENT|7444,7453|false|false|false|||deficient
Finding|Functional Concept|SIMPLE_SEGMENT|7444,7453|false|false|false|C0011155|Deficiency|deficient
Event|Event|SIMPLE_SEGMENT|7455,7462|false|false|false|||started
Finding|Finding|SIMPLE_SEGMENT|7463,7468|false|false|false|C3714655|On IV|on IV
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|7466,7473|false|false|false|C0082568|ferryl iron|IV iron
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7469,7473|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|7469,7473|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7469,7473|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Event|Event|SIMPLE_SEGMENT|7469,7473|false|false|false|||iron
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7469,7473|false|false|false|C0337439|Iron measurement|iron
Event|Event|SIMPLE_SEGMENT|7475,7484|false|false|false|||repletion
Event|Event|SIMPLE_SEGMENT|7486,7496|false|false|false|||discharged
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7503,7507|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|7503,7507|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7503,7507|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Event|Event|SIMPLE_SEGMENT|7503,7507|false|false|false|||iron
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7503,7507|false|false|false|C0337439|Iron measurement|iron
Finding|Body Substance|SIMPLE_SEGMENT|7510,7517|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|7510,7517|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|7510,7517|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|7518,7523|false|false|false|||found
Finding|Finding|SIMPLE_SEGMENT|7532,7544|false|false|false|C0586553|Raised TSH level|elevated TSH
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7541,7544|false|false|false|C2708739||TSH
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7541,7544|false|false|false|C0040160|thyrotropin|TSH
Drug|Hormone|SIMPLE_SEGMENT|7541,7544|false|false|false|C0040160|thyrotropin|TSH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7541,7544|false|false|false|C0040160|thyrotropin|TSH
Event|Event|SIMPLE_SEGMENT|7541,7544|false|false|false|||TSH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7541,7544|false|false|false|C0202230|Thyroid stimulating hormone measurement|TSH
Event|Event|SIMPLE_SEGMENT|7546,7552|false|false|false|||please
Event|Event|SIMPLE_SEGMENT|7553,7559|false|false|false|||follow
Finding|Functional Concept|SIMPLE_SEGMENT|7563,7567|false|false|false|C0332296|Free of (attribute)|free
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7563,7570|false|false|false|C0202225|T4 free measurement|free T4
Event|Event|SIMPLE_SEGMENT|7582,7589|false|false|false|||pending
Finding|Idea or Concept|SIMPLE_SEGMENT|7582,7589|false|false|false|C1691786;C1704475|Pending - Allergy Clinical Status;Pending - referral status|pending
Event|Event|SIMPLE_SEGMENT|7593,7602|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|7593,7602|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|7593,7602|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|7593,7602|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|7593,7602|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|SIMPLE_SEGMENT|7605,7609|false|false|false|||Code
Event|Occupational Activity|SIMPLE_SEGMENT|7605,7609|false|false|false|C0009219|Coding|Code
Finding|Intellectual Product|SIMPLE_SEGMENT|7605,7609|false|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|Code
Event|Event|SIMPLE_SEGMENT|7618,7627|false|false|false|||Emergency
Finding|Finding|SIMPLE_SEGMENT|7618,7627|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Finding|Idea or Concept|SIMPLE_SEGMENT|7618,7627|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Finding|Intellectual Product|SIMPLE_SEGMENT|7618,7627|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Finding|Pathologic Function|SIMPLE_SEGMENT|7618,7627|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|7618,7627|false|false|false|C0013956|Emergency Situation|Emergency
Procedure|Health Care Activity|SIMPLE_SEGMENT|7618,7627|false|false|false|C1553500|emergency encounter|Emergency
Finding|Functional Concept|SIMPLE_SEGMENT|7618,7635|false|false|false|C1552023|emergency contact|Emergency Contact
Event|Activity|SIMPLE_SEGMENT|7628,7635|false|false|false|C3812666|Personal Contact|Contact
Finding|Functional Concept|SIMPLE_SEGMENT|7628,7635|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|Contact
Finding|Idea or Concept|SIMPLE_SEGMENT|7628,7635|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|Contact
Finding|Intellectual Product|SIMPLE_SEGMENT|7628,7635|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|Contact
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|7628,7635|false|false|false|C0392367|Physical contact|Contact
Procedure|Health Care Activity|SIMPLE_SEGMENT|7683,7692|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7711,7721|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|7711,7721|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|7711,7726|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|SIMPLE_SEGMENT|7722,7726|false|false|false|||list
Finding|Intellectual Product|SIMPLE_SEGMENT|7722,7726|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|SIMPLE_SEGMENT|7730,7738|false|false|false|||accurate
Drug|Organic Chemical|SIMPLE_SEGMENT|7743,7751|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7743,7751|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|SIMPLE_SEGMENT|7743,7751|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|SIMPLE_SEGMENT|7743,7751|false|false|false|||complete
Finding|Functional Concept|SIMPLE_SEGMENT|7743,7751|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|SIMPLE_SEGMENT|7743,7751|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Organic Chemical|SIMPLE_SEGMENT|7756,7769|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7756,7769|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|SIMPLE_SEGMENT|7756,7769|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7756,7769|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|SIMPLE_SEGMENT|7784,7787|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7788,7792|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|7788,7792|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|7788,7792|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|7788,7792|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|SIMPLE_SEGMENT|7797,7805|false|false|false|C1831808|apixaban|Apixaban
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7797,7805|false|false|false|C1831808|apixaban|Apixaban
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|7814,7817|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7814,7817|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7814,7817|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|7814,7817|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|7814,7817|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|7822,7831|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7822,7831|false|false|false|C0001927|albuterol|Albuterol
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7839,7842|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7839,7842|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7839,7842|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Finding|Cell Function|SIMPLE_SEGMENT|7839,7842|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Finding|Gene or Genome|SIMPLE_SEGMENT|7839,7842|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7850,7853|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7850,7853|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7850,7853|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Event|Event|SIMPLE_SEGMENT|7850,7853|false|false|false|||NEB
Finding|Cell Function|SIMPLE_SEGMENT|7850,7853|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|SIMPLE_SEGMENT|7850,7853|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|SIMPLE_SEGMENT|7861,7864|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|SIMPLE_SEGMENT|7865,7874|false|false|false|||shortness
Finding|Body Substance|SIMPLE_SEGMENT|7879,7885|false|false|false|C0225386|Breath|breath
Drug|Organic Chemical|SIMPLE_SEGMENT|7890,7900|false|false|false|C0002598|amiodarone|Amiodarone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7890,7900|false|false|false|C0002598|amiodarone|Amiodarone
Event|Event|SIMPLE_SEGMENT|7890,7900|false|false|false|||Amiodarone
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7890,7900|false|false|false|C5399868|Drug assay amiodarone|Amiodarone
Drug|Organic Chemical|SIMPLE_SEGMENT|7921,7933|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7921,7933|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7951,7967|false|false|false|C0003921;C2608262;C3853661|Artificial Tears;Lubricant Eye Drops;artificial tears (medication)|Artificial Tears
Finding|Body Substance|SIMPLE_SEGMENT|7962,7967|false|false|false|C0039409;C1547924;C1611838|Tears (substance);Tears specimen|Tears
Finding|Intellectual Product|SIMPLE_SEGMENT|7962,7967|false|false|false|C0039409;C1547924;C1611838|Tears (substance);Tears specimen|Tears
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7972,7976|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|SIMPLE_SEGMENT|7972,7976|false|false|false|C1705648|Dropping|DROP
Event|Event|SIMPLE_SEGMENT|7972,7976|false|false|false|||DROP
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7977,7986|false|false|false|C0229118|Structure of both eyes|BOTH EYES
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7982,7986|false|false|false|C0015392|Eye|EYES
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7982,7986|false|false|false|C5848506||EYES
Finding|Gene or Genome|SIMPLE_SEGMENT|7987,7990|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|SIMPLE_SEGMENT|7991,8001|false|false|false|||irritation
Finding|Intellectual Product|SIMPLE_SEGMENT|7991,8001|false|false|false|C1706307;C2700617;C5575347|Have Vulvar Irritation question;Irritability - emotion;Irritation (finding)|irritation
Finding|Mental Process|SIMPLE_SEGMENT|7991,8001|false|false|false|C1706307;C2700617;C5575347|Have Vulvar Irritation question;Irritability - emotion;Irritation (finding)|irritation
Finding|Pathologic Function|SIMPLE_SEGMENT|7991,8001|false|false|false|C1706307;C2700617;C5575347|Have Vulvar Irritation question;Irritability - emotion;Irritation (finding)|irritation
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|7991,8001|false|false|false|C0441723|Irritation|irritation
Drug|Organic Chemical|SIMPLE_SEGMENT|8006,8017|false|false|false|C0090306|latanoprost|Latanoprost
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8006,8017|false|false|false|C0090306|latanoprost|Latanoprost
Finding|Functional Concept|SIMPLE_SEGMENT|8025,8030|false|false|false|C1522230|Ophthalmic Route of Administration|Ophth
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8040,8044|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|SIMPLE_SEGMENT|8040,8044|false|false|false|C1705648|Dropping|DROP
Event|Event|SIMPLE_SEGMENT|8045,8049|false|false|false|||LEFT
Finding|Functional Concept|SIMPLE_SEGMENT|8045,8049|false|false|false|C1552822|Table Cell Horizontal Align - left|LEFT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8045,8053|false|false|false|C0229090|Left eye structure|LEFT EYE
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8045,8053|false|false|false|C2141124|examination of left eye|LEFT EYE
Anatomy|Body Location or Region|SIMPLE_SEGMENT|8050,8053|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|EYE
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8050,8053|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|EYE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8050,8053|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|EYE
Disorder|Neoplastic Process|SIMPLE_SEGMENT|8050,8053|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|EYE
Event|Event|SIMPLE_SEGMENT|8050,8053|false|false|false|||EYE
Finding|Body Substance|SIMPLE_SEGMENT|8050,8053|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|EYE
Finding|Finding|SIMPLE_SEGMENT|8050,8053|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|EYE
Finding|Intellectual Product|SIMPLE_SEGMENT|8050,8053|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|EYE
Event|Event|SIMPLE_SEGMENT|8054,8057|false|false|false|||QHS
Drug|Organic Chemical|SIMPLE_SEGMENT|8062,8071|false|false|false|C0012373|diltiazem|Diltiazem
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8062,8071|false|false|false|C0012373|diltiazem|Diltiazem
Finding|Finding|SIMPLE_SEGMENT|8072,8080|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|SIMPLE_SEGMENT|8072,8080|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|SIMPLE_SEGMENT|8081,8088|false|false|false|||Release
Finding|Functional Concept|SIMPLE_SEGMENT|8081,8088|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|8081,8088|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8081,8088|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|8099,8102|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8099,8102|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8099,8102|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|8099,8102|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|8099,8102|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|8107,8118|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8107,8118|false|false|false|C0082607|fluticasone|Fluticasone
Event|Event|SIMPLE_SEGMENT|8107,8118|false|false|false|||Fluticasone
Drug|Organic Chemical|SIMPLE_SEGMENT|8107,8129|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8107,8129|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Organic Chemical|SIMPLE_SEGMENT|8119,8129|false|false|false|C0033474;C0392214|Propionates;propionate|Propionate
Event|Event|SIMPLE_SEGMENT|8119,8129|false|false|false|||Propionate
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8130,8135|false|false|false|C0028429||NASAL
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8130,8135|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Drug|Organic Chemical|SIMPLE_SEGMENT|8130,8135|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8130,8135|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Finding|Finding|SIMPLE_SEGMENT|8130,8135|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|NASAL
Finding|Functional Concept|SIMPLE_SEGMENT|8130,8135|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|NASAL
Event|Event|SIMPLE_SEGMENT|8138,8142|false|false|false|||SPRY
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|8146,8149|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8146,8149|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8146,8149|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|8146,8149|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|8146,8149|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|8155,8166|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8155,8166|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8155,8177|false|false|false|C0939232|fluticasone / salmeterol|Fluticasone-Salmeterol
Drug|Organic Chemical|SIMPLE_SEGMENT|8155,8184|false|false|false|C4762496|Fluticasone-Salmeterol Diskus|Fluticasone-Salmeterol Diskus
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8155,8184|false|false|false|C4762496|Fluticasone-Salmeterol Diskus|Fluticasone-Salmeterol Diskus
Drug|Organic Chemical|SIMPLE_SEGMENT|8167,8177|false|false|false|C0073992|salmeterol|Salmeterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8167,8177|false|false|false|C0073992|salmeterol|Salmeterol
Event|Event|SIMPLE_SEGMENT|8178,8184|false|false|false|||Diskus
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8197,8200|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Organic Chemical|SIMPLE_SEGMENT|8197,8200|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8197,8200|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Event|Event|SIMPLE_SEGMENT|8197,8200|false|false|false|||INH
Finding|Functional Concept|SIMPLE_SEGMENT|8197,8200|false|false|false|C0205535|Inhalation Route of Administration|INH
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|8204,8207|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8204,8207|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8204,8207|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|8204,8207|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|8204,8207|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|8213,8232|false|false|false|C0020261|hydrochlorothiazide|Hydrochlorothiazide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8213,8232|false|false|false|C0020261|hydrochlorothiazide|Hydrochlorothiazide
Drug|Organic Chemical|SIMPLE_SEGMENT|8253,8263|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8253,8263|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Organic Chemical|SIMPLE_SEGMENT|8253,8275|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8253,8275|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Event|Event|SIMPLE_SEGMENT|8264,8275|false|false|false|||Mononitrate
Finding|Finding|SIMPLE_SEGMENT|8277,8285|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|SIMPLE_SEGMENT|8277,8285|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|SIMPLE_SEGMENT|8286,8293|false|false|false|||Release
Finding|Functional Concept|SIMPLE_SEGMENT|8286,8293|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|8286,8293|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8286,8293|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|SIMPLE_SEGMENT|8316,8325|false|false|false|C0024002|lorazepam|Lorazepam
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8316,8325|false|false|false|C0024002|lorazepam|Lorazepam
Event|Event|SIMPLE_SEGMENT|8336,8339|false|false|false|||QHS
Finding|Gene or Genome|SIMPLE_SEGMENT|8340,8343|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8344,8352|false|false|false|C1950154|Insomnia homeopathic medication|insomnia
Event|Event|SIMPLE_SEGMENT|8344,8352|false|false|false|||insomnia
Finding|Sign or Symptom|SIMPLE_SEGMENT|8344,8352|false|false|false|C0917801|Sleeplessness|insomnia
Drug|Organic Chemical|SIMPLE_SEGMENT|8358,8370|false|false|false|C0039771|theophylline|Theophylline
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8358,8370|false|false|false|C0039771|theophylline|Theophylline
Event|Event|SIMPLE_SEGMENT|8358,8370|false|false|false|||Theophylline
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8358,8370|false|false|false|C0039773|Assay of theophylline|Theophylline
Drug|Organic Chemical|SIMPLE_SEGMENT|8358,8373|false|false|false|C2241157|Theophylline ER|Theophylline ER
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8358,8373|false|false|false|C2241157|Theophylline ER|Theophylline ER
Event|Event|SIMPLE_SEGMENT|8371,8373|false|false|false|||ER
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|8384,8387|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8384,8387|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8384,8387|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|8384,8387|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|8384,8387|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|8393,8403|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8393,8403|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Organic Chemical|SIMPLE_SEGMENT|8425,8435|false|false|false|C0213771|tiotropium|Tiotropium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8425,8435|false|false|false|C0213771|tiotropium|Tiotropium
Event|Event|SIMPLE_SEGMENT|8425,8435|false|false|false|||Tiotropium
Drug|Organic Chemical|SIMPLE_SEGMENT|8425,8443|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8425,8443|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Inorganic Chemical|SIMPLE_SEGMENT|8436,8443|false|false|false|C0006222|Bromides|Bromide
Event|Event|SIMPLE_SEGMENT|8436,8443|false|false|false|||Bromide
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8436,8443|false|false|false|C0202341|Bromides measurement|Bromide
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|8446,8449|false|false|false|C1855179|CATARACT, ANTERIOR POLAR|CAP
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8446,8449|false|false|false|C0006935|capsule (pharmacologic)|CAP
Event|Event|SIMPLE_SEGMENT|8446,8449|false|false|false|||CAP
Finding|Gene or Genome|SIMPLE_SEGMENT|8446,8449|false|false|false|C1416891;C1418551;C1419093;C1422073;C1422760;C2985259;C4522312|BRD4 gene;BRD4 wt Allele;CAP1 gene;HACD1 gene;LNPEP gene;SERPINB6 gene;SORBS1 gene|CAP
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8446,8449|false|false|false|C0278651;C0280547;C1879916|CAP Regimen;cisplatin/cyclophosphamide/doxorubicin protocol;cyclophosphamide/doxorubicin/prednisone protocol|CAP
Drug|Organic Chemical|SIMPLE_SEGMENT|8464,8477|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8464,8477|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|SIMPLE_SEGMENT|8464,8477|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Event|Event|SIMPLE_SEGMENT|8464,8477|false|false|false|||Multivitamins
Drug|Inorganic Chemical|SIMPLE_SEGMENT|8480,8488|false|false|false|C0026162|Minerals|minerals
Event|Event|SIMPLE_SEGMENT|8480,8488|false|false|false|||minerals
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8491,8494|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|SIMPLE_SEGMENT|8491,8494|false|false|false|||TAB
Drug|Organic Chemical|SIMPLE_SEGMENT|8509,8516|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8509,8516|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|SIMPLE_SEGMENT|8537,8548|false|false|false|C0165590|dorzolamide|Dorzolamide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8537,8548|false|false|false|C0165590|dorzolamide|Dorzolamide
Finding|Functional Concept|SIMPLE_SEGMENT|8552,8557|false|false|false|C1522230|Ophthalmic Route of Administration|Ophth
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8567,8571|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|SIMPLE_SEGMENT|8567,8571|false|false|false|C1705648|Dropping|DROP
Event|Event|SIMPLE_SEGMENT|8567,8571|false|false|false|||DROP
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8572,8581|false|false|false|C0229118|Structure of both eyes|BOTH EYES
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8577,8581|false|false|false|C0015392|Eye|EYES
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8577,8581|false|false|false|C5848506||EYES
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|8582,8585|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8582,8585|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8582,8585|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|8582,8585|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|8582,8585|false|false|false|C1332410|BID gene|BID
Event|Event|SIMPLE_SEGMENT|8590,8599|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|8590,8599|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|8590,8599|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|8590,8599|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|8590,8599|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|8590,8611|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8600,8611|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8600,8611|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|8600,8611|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|8600,8611|false|false|false|C4284232|Medications|Medications
Event|Event|SIMPLE_SEGMENT|8616,8620|false|false|false|||Home
Finding|Idea or Concept|SIMPLE_SEGMENT|8616,8620|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|SIMPLE_SEGMENT|8616,8620|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|SIMPLE_SEGMENT|8616,8620|false|false|false|C1553498|home health encounter|Home
Event|Event|SIMPLE_SEGMENT|8633,8643|false|false|false|||continuous
Finding|Idea or Concept|SIMPLE_SEGMENT|8633,8643|false|false|false|C0549178|Continuous|continuous
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8644,8649|false|false|false|C0028429||nasal
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8644,8649|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Organic Chemical|SIMPLE_SEGMENT|8644,8649|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8644,8649|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Finding|Finding|SIMPLE_SEGMENT|8644,8649|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Functional Concept|SIMPLE_SEGMENT|8644,8649|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8650,8657|false|false|false|C1550232|Body Parts - Cannula|cannula
Event|Event|SIMPLE_SEGMENT|8650,8657|false|false|false|||cannula
Finding|Body Substance|SIMPLE_SEGMENT|8650,8657|false|false|false|C1546577;C1550622|Specimen Type - Cannula|cannula
Finding|Intellectual Product|SIMPLE_SEGMENT|8650,8657|false|false|false|C1546577;C1550622|Specimen Type - Cannula|cannula
Event|Event|SIMPLE_SEGMENT|8663,8671|false|false|false|||exertion
Finding|Organism Function|SIMPLE_SEGMENT|8663,8671|false|false|false|C0015264|Exertion|exertion
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8672,8681|false|false|false|C0945731||Diagnosis
Event|Event|SIMPLE_SEGMENT|8672,8681|false|false|false|||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|8672,8681|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|8672,8681|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8672,8681|false|false|false|C0011900|Diagnosis|Diagnosis
Event|Event|SIMPLE_SEGMENT|8683,8690|false|false|false|||chronic
Finding|Intellectual Product|SIMPLE_SEGMENT|8683,8690|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|8683,8690|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8683,8720|false|false|false|C0024117|Chronic Obstructive Airway Disease|chronic obstructive pulmonary disease
Finding|Functional Concept|SIMPLE_SEGMENT|8691,8702|false|false|false|C0549186|Obstructed|obstructive
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8691,8720|false|false|false|C0600260|Lung Diseases, Obstructive|obstructive pulmonary disease
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8703,8712|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8703,8712|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|8703,8712|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8703,8720|false|false|false|C0024115|Lung diseases|pulmonary disease
Finding|Finding|SIMPLE_SEGMENT|8703,8720|false|false|false|C0455540|History of - respiratory disease|pulmonary disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8713,8720|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|8713,8720|false|false|false|||disease
Event|Event|SIMPLE_SEGMENT|8729,8735|false|false|false|||Length
Event|Event|SIMPLE_SEGMENT|8739,8744|false|false|false|||Needs
Finding|Functional Concept|SIMPLE_SEGMENT|8739,8744|false|false|false|C0686904|Patient need for (contextual qualifier)|Needs
Event|Event|SIMPLE_SEGMENT|8746,8753|false|false|false|||ongoing
Finding|Idea or Concept|SIMPLE_SEGMENT|8746,8753|false|false|false|C0549178|Continuous|ongoing
Drug|Organic Chemical|SIMPLE_SEGMENT|8765,8778|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8765,8778|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|SIMPLE_SEGMENT|8765,8778|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8765,8778|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|SIMPLE_SEGMENT|8793,8796|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8797,8801|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|8797,8801|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|8797,8801|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|8797,8801|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|SIMPLE_SEGMENT|8806,8816|false|false|false|C0002598|amiodarone|Amiodarone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8806,8816|false|false|false|C0002598|amiodarone|Amiodarone
Event|Event|SIMPLE_SEGMENT|8806,8816|false|false|false|||Amiodarone
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8806,8816|false|false|false|C5399868|Drug assay amiodarone|Amiodarone
Drug|Organic Chemical|SIMPLE_SEGMENT|8837,8845|false|false|false|C1831808|apixaban|Apixaban
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8837,8845|false|false|false|C1831808|apixaban|Apixaban
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|8854,8857|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8854,8857|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8854,8857|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|8854,8857|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|8854,8857|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|8862,8871|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8862,8871|false|false|false|C0001927|albuterol|Albuterol
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8879,8882|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8879,8882|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8879,8882|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Finding|Cell Function|SIMPLE_SEGMENT|8879,8882|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Finding|Gene or Genome|SIMPLE_SEGMENT|8879,8882|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8890,8893|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8890,8893|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8890,8893|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Event|Event|SIMPLE_SEGMENT|8890,8893|false|false|false|||NEB
Finding|Cell Function|SIMPLE_SEGMENT|8890,8893|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|SIMPLE_SEGMENT|8890,8893|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|SIMPLE_SEGMENT|8901,8904|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|SIMPLE_SEGMENT|8905,8914|false|false|false|||shortness
Finding|Body Substance|SIMPLE_SEGMENT|8919,8925|false|false|false|C0225386|Breath|breath
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8930,8946|false|false|false|C0003921;C2608262;C3853661|Artificial Tears;Lubricant Eye Drops;artificial tears (medication)|Artificial Tears
Finding|Body Substance|SIMPLE_SEGMENT|8941,8946|false|false|false|C0039409;C1547924;C1611838|Tears (substance);Tears specimen|Tears
Finding|Intellectual Product|SIMPLE_SEGMENT|8941,8946|false|false|false|C0039409;C1547924;C1611838|Tears (substance);Tears specimen|Tears
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8951,8955|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|SIMPLE_SEGMENT|8951,8955|false|false|false|C1705648|Dropping|DROP
Event|Event|SIMPLE_SEGMENT|8951,8955|false|false|false|||DROP
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8956,8965|false|false|false|C0229118|Structure of both eyes|BOTH EYES
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8961,8965|false|false|false|C0015392|Eye|EYES
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8961,8965|false|false|false|C5848506||EYES
Finding|Gene or Genome|SIMPLE_SEGMENT|8966,8969|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|SIMPLE_SEGMENT|8970,8980|false|false|false|||irritation
Finding|Intellectual Product|SIMPLE_SEGMENT|8970,8980|false|false|false|C1706307;C2700617;C5575347|Have Vulvar Irritation question;Irritability - emotion;Irritation (finding)|irritation
Finding|Mental Process|SIMPLE_SEGMENT|8970,8980|false|false|false|C1706307;C2700617;C5575347|Have Vulvar Irritation question;Irritability - emotion;Irritation (finding)|irritation
Finding|Pathologic Function|SIMPLE_SEGMENT|8970,8980|false|false|false|C1706307;C2700617;C5575347|Have Vulvar Irritation question;Irritability - emotion;Irritation (finding)|irritation
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|8970,8980|false|false|false|C0441723|Irritation|irritation
Drug|Organic Chemical|SIMPLE_SEGMENT|8985,8992|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8985,8992|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|SIMPLE_SEGMENT|9012,9024|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9012,9024|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|SIMPLE_SEGMENT|9042,9051|false|false|false|C0012373|diltiazem|Diltiazem
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9042,9051|false|false|false|C0012373|diltiazem|Diltiazem
Finding|Finding|SIMPLE_SEGMENT|9052,9060|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|SIMPLE_SEGMENT|9052,9060|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|SIMPLE_SEGMENT|9061,9068|false|false|false|||Release
Finding|Functional Concept|SIMPLE_SEGMENT|9061,9068|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|9061,9068|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9061,9068|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|9079,9082|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9079,9082|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9079,9082|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|9079,9082|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|9079,9082|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|9088,9099|false|false|false|C0165590|dorzolamide|Dorzolamide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9088,9099|false|false|false|C0165590|dorzolamide|Dorzolamide
Finding|Functional Concept|SIMPLE_SEGMENT|9103,9108|false|false|false|C1522230|Ophthalmic Route of Administration|Ophth
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9118,9122|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|SIMPLE_SEGMENT|9118,9122|false|false|false|C1705648|Dropping|DROP
Event|Event|SIMPLE_SEGMENT|9118,9122|false|false|false|||DROP
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9123,9132|false|false|false|C0229118|Structure of both eyes|BOTH EYES
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9128,9132|false|false|false|C0015392|Eye|EYES
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9128,9132|false|false|false|C5848506||EYES
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|9133,9136|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9133,9136|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9133,9136|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|9133,9136|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|9133,9136|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|9142,9153|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9142,9153|false|false|false|C0082607|fluticasone|Fluticasone
Event|Event|SIMPLE_SEGMENT|9142,9153|false|false|false|||Fluticasone
Drug|Organic Chemical|SIMPLE_SEGMENT|9142,9164|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9142,9164|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Organic Chemical|SIMPLE_SEGMENT|9154,9164|false|false|false|C0033474;C0392214|Propionates;propionate|Propionate
Event|Event|SIMPLE_SEGMENT|9154,9164|false|false|false|||Propionate
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9165,9170|false|false|false|C0028429||NASAL
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9165,9170|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Drug|Organic Chemical|SIMPLE_SEGMENT|9165,9170|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9165,9170|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Finding|Finding|SIMPLE_SEGMENT|9165,9170|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|NASAL
Finding|Functional Concept|SIMPLE_SEGMENT|9165,9170|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|NASAL
Event|Event|SIMPLE_SEGMENT|9173,9177|false|false|false|||SPRY
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|9181,9184|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9181,9184|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9181,9184|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|9181,9184|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|9181,9184|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|9190,9201|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9190,9201|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9190,9212|false|false|false|C0939232|fluticasone / salmeterol|Fluticasone-Salmeterol
Drug|Organic Chemical|SIMPLE_SEGMENT|9190,9219|false|false|false|C4762496|Fluticasone-Salmeterol Diskus|Fluticasone-Salmeterol Diskus
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9190,9219|false|false|false|C4762496|Fluticasone-Salmeterol Diskus|Fluticasone-Salmeterol Diskus
Drug|Organic Chemical|SIMPLE_SEGMENT|9202,9212|false|false|false|C0073992|salmeterol|Salmeterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9202,9212|false|false|false|C0073992|salmeterol|Salmeterol
Event|Event|SIMPLE_SEGMENT|9213,9219|false|false|false|||Diskus
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9232,9235|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Organic Chemical|SIMPLE_SEGMENT|9232,9235|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9232,9235|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Event|Event|SIMPLE_SEGMENT|9232,9235|false|false|false|||INH
Finding|Functional Concept|SIMPLE_SEGMENT|9232,9235|false|false|false|C0205535|Inhalation Route of Administration|INH
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|9239,9242|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9239,9242|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9239,9242|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|9239,9242|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|9239,9242|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|9248,9267|false|false|false|C0020261|hydrochlorothiazide|Hydrochlorothiazide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9248,9267|false|false|false|C0020261|hydrochlorothiazide|Hydrochlorothiazide
Drug|Organic Chemical|SIMPLE_SEGMENT|9288,9298|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9288,9298|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Organic Chemical|SIMPLE_SEGMENT|9288,9310|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9288,9310|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Event|Event|SIMPLE_SEGMENT|9299,9310|false|false|false|||Mononitrate
Finding|Finding|SIMPLE_SEGMENT|9312,9320|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|SIMPLE_SEGMENT|9312,9320|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|SIMPLE_SEGMENT|9321,9328|false|false|false|||Release
Finding|Functional Concept|SIMPLE_SEGMENT|9321,9328|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|9321,9328|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9321,9328|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|SIMPLE_SEGMENT|9351,9362|false|false|false|C0090306|latanoprost|Latanoprost
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9351,9362|false|false|false|C0090306|latanoprost|Latanoprost
Finding|Functional Concept|SIMPLE_SEGMENT|9370,9375|false|false|false|C1522230|Ophthalmic Route of Administration|Ophth
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9385,9389|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|SIMPLE_SEGMENT|9385,9389|false|false|false|C1705648|Dropping|DROP
Event|Event|SIMPLE_SEGMENT|9390,9394|false|false|false|||LEFT
Finding|Functional Concept|SIMPLE_SEGMENT|9390,9394|false|false|false|C1552822|Table Cell Horizontal Align - left|LEFT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9390,9398|false|false|false|C0229090|Left eye structure|LEFT EYE
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|9390,9398|false|false|false|C2141124|examination of left eye|LEFT EYE
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9395,9398|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|EYE
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9395,9398|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|EYE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9395,9398|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|EYE
Disorder|Neoplastic Process|SIMPLE_SEGMENT|9395,9398|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|EYE
Event|Event|SIMPLE_SEGMENT|9395,9398|false|false|false|||EYE
Finding|Body Substance|SIMPLE_SEGMENT|9395,9398|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|EYE
Finding|Finding|SIMPLE_SEGMENT|9395,9398|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|EYE
Finding|Intellectual Product|SIMPLE_SEGMENT|9395,9398|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|EYE
Event|Event|SIMPLE_SEGMENT|9399,9402|false|false|false|||QHS
Drug|Organic Chemical|SIMPLE_SEGMENT|9408,9417|false|false|false|C0024002|lorazepam|Lorazepam
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9408,9417|false|false|false|C0024002|lorazepam|Lorazepam
Event|Event|SIMPLE_SEGMENT|9428,9431|false|false|false|||QHS
Finding|Gene or Genome|SIMPLE_SEGMENT|9432,9435|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9436,9444|false|false|false|C1950154|Insomnia homeopathic medication|insomnia
Event|Event|SIMPLE_SEGMENT|9436,9444|false|false|false|||insomnia
Finding|Sign or Symptom|SIMPLE_SEGMENT|9436,9444|false|false|false|C0917801|Sleeplessness|insomnia
Drug|Organic Chemical|SIMPLE_SEGMENT|9450,9463|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9450,9463|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|SIMPLE_SEGMENT|9450,9463|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Event|Event|SIMPLE_SEGMENT|9450,9463|false|false|false|||Multivitamins
Drug|Inorganic Chemical|SIMPLE_SEGMENT|9466,9474|false|false|false|C0026162|Minerals|minerals
Event|Event|SIMPLE_SEGMENT|9466,9474|false|false|false|||minerals
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9477,9480|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|SIMPLE_SEGMENT|9477,9480|false|false|false|||TAB
Drug|Organic Chemical|SIMPLE_SEGMENT|9495,9505|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9495,9505|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Organic Chemical|SIMPLE_SEGMENT|9527,9537|false|false|false|C0213771|tiotropium|Tiotropium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9527,9537|false|false|false|C0213771|tiotropium|Tiotropium
Event|Event|SIMPLE_SEGMENT|9527,9537|false|false|false|||Tiotropium
Drug|Organic Chemical|SIMPLE_SEGMENT|9527,9545|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9527,9545|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Inorganic Chemical|SIMPLE_SEGMENT|9538,9545|false|false|false|C0006222|Bromides|Bromide
Event|Event|SIMPLE_SEGMENT|9538,9545|false|false|false|||Bromide
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9538,9545|false|false|false|C0202341|Bromides measurement|Bromide
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|9548,9551|false|false|false|C1855179|CATARACT, ANTERIOR POLAR|CAP
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9548,9551|false|false|false|C0006935|capsule (pharmacologic)|CAP
Event|Event|SIMPLE_SEGMENT|9548,9551|false|false|false|||CAP
Finding|Gene or Genome|SIMPLE_SEGMENT|9548,9551|false|false|false|C1416891;C1418551;C1419093;C1422073;C1422760;C2985259;C4522312|BRD4 gene;BRD4 wt Allele;CAP1 gene;HACD1 gene;LNPEP gene;SERPINB6 gene;SORBS1 gene|CAP
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9548,9551|false|false|false|C0278651;C0280547;C1879916|CAP Regimen;cisplatin/cyclophosphamide/doxorubicin protocol;cyclophosphamide/doxorubicin/prednisone protocol|CAP
Drug|Organic Chemical|SIMPLE_SEGMENT|9566,9578|false|false|false|C0039771|theophylline|Theophylline
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9566,9578|false|false|false|C0039771|theophylline|Theophylline
Event|Event|SIMPLE_SEGMENT|9566,9578|false|false|false|||Theophylline
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9566,9578|false|false|false|C0039773|Assay of theophylline|Theophylline
Drug|Organic Chemical|SIMPLE_SEGMENT|9566,9581|false|false|false|C0939729|Theophylline SR|Theophylline SR
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9566,9581|false|false|false|C0939729|Theophylline SR|Theophylline SR
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|9592,9595|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9592,9595|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9592,9595|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|9592,9595|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|9592,9595|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|9601,9613|false|false|false|C0039771|theophylline|theophylline
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9601,9613|false|false|false|C0039771|theophylline|theophylline
Event|Event|SIMPLE_SEGMENT|9601,9613|false|false|false|||theophylline
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9601,9613|false|false|false|C0039773|Assay of theophylline|theophylline
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9623,9629|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|SIMPLE_SEGMENT|9633,9641|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9636,9641|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|9636,9641|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Idea or Concept|SIMPLE_SEGMENT|9650,9653|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|9650,9653|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Activity|SIMPLE_SEGMENT|9654,9658|false|false|false|C1880359|Dispense (activity)|Disp
Finding|Gene or Genome|SIMPLE_SEGMENT|9654,9658|false|false|false|C2828567|PRSS30P gene|Disp
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9665,9671|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|9672,9679|false|false|false|||Refills
Finding|Idea or Concept|SIMPLE_SEGMENT|9672,9679|false|false|false|C0807726|refill|Refills
Drug|Antibiotic|SIMPLE_SEGMENT|9687,9698|false|false|false|C0055011|cefpodoxime|Cefpodoxime
Drug|Organic Chemical|SIMPLE_SEGMENT|9687,9698|false|false|false|C0055011|cefpodoxime|Cefpodoxime
Drug|Antibiotic|SIMPLE_SEGMENT|9687,9707|false|false|false|C0108938|cefpodoxime proxetil|Cefpodoxime Proxetil
Drug|Organic Chemical|SIMPLE_SEGMENT|9687,9707|false|false|false|C0108938|cefpodoxime proxetil|Cefpodoxime Proxetil
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9723,9731|false|false|false|C0720099|Duration brand of oxymetazoline|Duration
Event|Event|SIMPLE_SEGMENT|9723,9731|false|false|false|||Duration
Event|Event|SIMPLE_SEGMENT|9735,9739|false|false|false|||Days
Drug|Antibiotic|SIMPLE_SEGMENT|9745,9756|false|false|false|C0055011|cefpodoxime|cefpodoxime
Drug|Organic Chemical|SIMPLE_SEGMENT|9745,9756|false|false|false|C0055011|cefpodoxime|cefpodoxime
Event|Event|SIMPLE_SEGMENT|9745,9756|false|false|false|||cefpodoxime
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9766,9772|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|SIMPLE_SEGMENT|9776,9784|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9779,9784|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|9779,9784|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Idea or Concept|SIMPLE_SEGMENT|9793,9796|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|9793,9796|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9807,9813|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|9814,9821|false|false|false|||Refills
Finding|Idea or Concept|SIMPLE_SEGMENT|9814,9821|false|false|false|C0807726|refill|Refills
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|9829,9836|false|false|false|C2346592|Ferrous|Ferrous
Drug|Inorganic Chemical|SIMPLE_SEGMENT|9829,9844|false|false|false|C0060282|ferrous sulfate|Ferrous Sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9829,9844|false|false|false|C0060282|ferrous sulfate|Ferrous Sulfate
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|9837,9844|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Inorganic Chemical|SIMPLE_SEGMENT|9837,9844|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9837,9844|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Event|Event|SIMPLE_SEGMENT|9837,9844|false|false|false|||Sulfate
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|9866,9873|false|false|false|C2346592|Ferrous|ferrous
Drug|Inorganic Chemical|SIMPLE_SEGMENT|9866,9881|false|false|false|C0060282|ferrous sulfate|ferrous sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9866,9881|false|false|false|C0060282|ferrous sulfate|ferrous sulfate
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|9874,9881|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Inorganic Chemical|SIMPLE_SEGMENT|9874,9881|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9874,9881|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Event|Event|SIMPLE_SEGMENT|9874,9881|false|false|false|||sulfate
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9896,9900|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|9896,9900|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9896,9900|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Event|Event|SIMPLE_SEGMENT|9896,9900|false|false|false|||iron
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9896,9900|false|false|false|C0337439|Iron measurement|iron
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9904,9910|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|SIMPLE_SEGMENT|9914,9922|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9917,9922|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|9917,9922|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9940,9946|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|9947,9954|false|false|false|||Refills
Finding|Idea or Concept|SIMPLE_SEGMENT|9947,9954|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|9962,9970|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9962,9970|false|false|false|C1692318|docusate|Docusate
Drug|Organic Chemical|SIMPLE_SEGMENT|9962,9977|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9962,9977|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9971,9977|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|9971,9977|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9971,9977|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|SIMPLE_SEGMENT|9971,9977|false|false|false|||Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|9971,9977|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9971,9977|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|9988,9991|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9988,9991|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9988,9991|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|9988,9991|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|9988,9991|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|9997,10005|false|false|false|C1692318|docusate|docusate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9997,10005|false|false|false|C1692318|docusate|docusate
Drug|Organic Chemical|SIMPLE_SEGMENT|9997,10012|false|false|false|C0243237|docusate sodium|docusate sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9997,10012|false|false|false|C0243237|docusate sodium|docusate sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|10006,10012|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|10006,10012|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10006,10012|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Event|Event|SIMPLE_SEGMENT|10006,10012|false|false|false|||sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|10006,10012|false|false|false|C4553025|Sodium metabolic function|sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10006,10012|false|false|false|C0337443|Sodium measurement|sodium
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10022,10029|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Anatomy|Cell Component|SIMPLE_SEGMENT|10022,10029|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10022,10029|false|false|false|C0006935|capsule (pharmacologic)|capsule
Finding|Functional Concept|SIMPLE_SEGMENT|10033,10041|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|10036,10041|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|10036,10041|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Idea or Concept|SIMPLE_SEGMENT|10050,10053|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|10050,10053|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10065,10072|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|SIMPLE_SEGMENT|10065,10072|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10065,10072|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Event|Event|SIMPLE_SEGMENT|10073,10080|false|false|false|||Refills
Finding|Idea or Concept|SIMPLE_SEGMENT|10073,10080|false|false|false|C0807726|refill|Refills
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10088,10100|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|Polyethylene
Drug|Organic Chemical|SIMPLE_SEGMENT|10088,10100|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|Polyethylene
Event|Event|SIMPLE_SEGMENT|10088,10100|false|false|false|||Polyethylene
Drug|Organic Chemical|SIMPLE_SEGMENT|10088,10107|false|false|false|C0032483|polyethylene glycols|Polyethylene Glycol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10088,10107|false|false|false|C0032483|polyethylene glycols|Polyethylene Glycol
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|10101,10107|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|Glycol
Drug|Organic Chemical|SIMPLE_SEGMENT|10101,10107|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|Glycol
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10127,10139|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|polyethylene
Drug|Organic Chemical|SIMPLE_SEGMENT|10127,10139|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|polyethylene
Drug|Organic Chemical|SIMPLE_SEGMENT|10127,10146|false|false|false|C0032483|polyethylene glycols|polyethylene glycol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10127,10146|false|false|false|C0032483|polyethylene glycols|polyethylene glycol
Drug|Organic Chemical|SIMPLE_SEGMENT|10127,10151|false|false|false|C0724672|polyethylene glycol 3350|polyethylene glycol 3350
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10127,10151|false|false|false|C0724672|polyethylene glycol 3350|polyethylene glycol 3350
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|10140,10146|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|glycol
Drug|Organic Chemical|SIMPLE_SEGMENT|10140,10146|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|glycol
Event|Event|SIMPLE_SEGMENT|10140,10146|false|false|false|||glycol
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10167,10173|false|false|false|C0032861;C1382110|Powder dose form;powder physical state|powder
Drug|Substance|SIMPLE_SEGMENT|10167,10173|false|false|false|C0032861;C1382110|Powder dose form;powder physical state|powder
Event|Event|SIMPLE_SEGMENT|10167,10173|false|false|false|||powder
Finding|Functional Concept|SIMPLE_SEGMENT|10177,10185|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|10180,10185|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|10180,10185|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Event|Event|SIMPLE_SEGMENT|10193,10200|false|false|false|||Refills
Finding|Idea or Concept|SIMPLE_SEGMENT|10193,10200|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|10208,10219|false|false|false|C0027235|ipratropium|Ipratropium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10208,10219|false|false|false|C0027235|ipratropium|Ipratropium
Event|Event|SIMPLE_SEGMENT|10208,10219|false|false|false|||Ipratropium
Drug|Organic Chemical|SIMPLE_SEGMENT|10208,10227|false|false|false|C0700580|ipratropium bromide|Ipratropium Bromide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10208,10227|false|false|false|C0700580|ipratropium bromide|Ipratropium Bromide
Drug|Inorganic Chemical|SIMPLE_SEGMENT|10220,10227|false|false|false|C0006222|Bromides|Bromide
Event|Event|SIMPLE_SEGMENT|10220,10227|false|false|false|||Bromide
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10220,10227|false|false|false|C0202341|Bromides measurement|Bromide
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10228,10231|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|10228,10231|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10228,10231|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Event|Event|SIMPLE_SEGMENT|10228,10231|false|false|false|||Neb
Finding|Cell Function|SIMPLE_SEGMENT|10228,10231|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Finding|Gene or Genome|SIMPLE_SEGMENT|10228,10231|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10234,10237|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biologically Active Substance|SIMPLE_SEGMENT|10234,10237|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10234,10237|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Event|Event|SIMPLE_SEGMENT|10234,10237|false|false|false|||NEB
Finding|Cell Function|SIMPLE_SEGMENT|10234,10237|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|SIMPLE_SEGMENT|10234,10237|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Event|Event|SIMPLE_SEGMENT|10241,10244|false|false|false|||Q6H
Finding|Gene or Genome|SIMPLE_SEGMENT|10245,10248|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|SIMPLE_SEGMENT|10249,10256|false|false|false|||dyspnea
Finding|Finding|SIMPLE_SEGMENT|10249,10256|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|10249,10256|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Event|Event|SIMPLE_SEGMENT|10258,10266|false|false|false|||wheezing
Finding|Sign or Symptom|SIMPLE_SEGMENT|10258,10266|false|false|false|C0043144|Wheezing|wheezing
Drug|Organic Chemical|SIMPLE_SEGMENT|10272,10283|false|false|false|C0027235|ipratropium|ipratropium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10272,10283|false|false|false|C0027235|ipratropium|ipratropium
Drug|Organic Chemical|SIMPLE_SEGMENT|10272,10291|false|false|false|C0700580|ipratropium bromide|ipratropium bromide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10272,10291|false|false|false|C0700580|ipratropium bromide|ipratropium bromide
Drug|Inorganic Chemical|SIMPLE_SEGMENT|10284,10291|false|false|false|C0006222|Bromides|bromide
Event|Event|SIMPLE_SEGMENT|10284,10291|false|false|false|||bromide
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10284,10291|false|false|false|C0202341|Bromides measurement|bromide
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10314,10317|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|neb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|10314,10317|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|neb
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10314,10317|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|neb
Finding|Cell Function|SIMPLE_SEGMENT|10314,10317|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|neb
Finding|Gene or Genome|SIMPLE_SEGMENT|10314,10317|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|neb
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10318,10321|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Organic Chemical|SIMPLE_SEGMENT|10318,10321|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10318,10321|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Event|Event|SIMPLE_SEGMENT|10318,10321|false|false|false|||INH
Finding|Functional Concept|SIMPLE_SEGMENT|10318,10321|false|false|false|C0205535|Inhalation Route of Administration|INH
Finding|Intellectual Product|SIMPLE_SEGMENT|10322,10327|false|false|false|C1720374|Every - dosing instruction fragment|Every
Event|Event|SIMPLE_SEGMENT|10356,10363|false|false|false|||Refills
Finding|Idea or Concept|SIMPLE_SEGMENT|10356,10363|false|false|false|C0807726|refill|Refills
Drug|Hormone|SIMPLE_SEGMENT|10371,10381|false|false|false|C0032952|prednisone|PredniSONE
Drug|Organic Chemical|SIMPLE_SEGMENT|10371,10381|false|false|false|C0032952|prednisone|PredniSONE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10371,10381|false|false|false|C0032952|prednisone|PredniSONE
Finding|Intellectual Product|SIMPLE_SEGMENT|10409,10413|false|false|false|C1720594|Then - dosing instruction fragment|then
Finding|Intellectual Product|SIMPLE_SEGMENT|10426,10430|false|false|false|C1720594|Then - dosing instruction fragment|then
Finding|Intellectual Product|SIMPLE_SEGMENT|10442,10446|false|false|false|C1720594|Then - dosing instruction fragment|then
Finding|Intellectual Product|SIMPLE_SEGMENT|10458,10462|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|SIMPLE_SEGMENT|10469,10476|false|false|false|||ongoing
Finding|Idea or Concept|SIMPLE_SEGMENT|10469,10476|false|false|false|C0549178|Continuous|ongoing
Procedure|Health Care Activity|SIMPLE_SEGMENT|10478,10485|false|false|false|C0441640||Tapered
Event|Event|SIMPLE_SEGMENT|10493,10497|false|false|false|||DOWN
Drug|Hormone|SIMPLE_SEGMENT|10503,10513|false|false|false|C0032952|prednisone|prednisone
Drug|Organic Chemical|SIMPLE_SEGMENT|10503,10513|false|false|false|C0032952|prednisone|prednisone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10503,10513|false|false|false|C0032952|prednisone|prednisone
Event|Event|SIMPLE_SEGMENT|10503,10513|false|false|false|||prednisone
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10527,10533|false|false|false|C0039225|Tablet Dosage Form|tablet
Event|Event|SIMPLE_SEGMENT|10527,10533|false|false|false|||tablet
Finding|Functional Concept|SIMPLE_SEGMENT|10537,10545|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|10540,10545|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|10540,10545|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Event|Event|SIMPLE_SEGMENT|10558,10562|false|false|false|||Disp
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10569,10575|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|10576,10583|false|false|false|||Refills
Finding|Idea or Concept|SIMPLE_SEGMENT|10576,10583|false|false|false|C0807726|refill|Refills
Event|Event|SIMPLE_SEGMENT|10590,10599|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|10590,10599|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|10590,10599|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|10590,10599|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|10590,10599|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10590,10611|false|false|false|C4019243||Discharge Disposition
Finding|Finding|SIMPLE_SEGMENT|10590,10611|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10600,10611|false|false|false|C2926604||Disposition
Event|Event|SIMPLE_SEGMENT|10600,10611|false|false|false|||Disposition
Procedure|Health Care Activity|SIMPLE_SEGMENT|10600,10611|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|SIMPLE_SEGMENT|10613,10617|false|false|false|||Home
Finding|Idea or Concept|SIMPLE_SEGMENT|10613,10617|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|SIMPLE_SEGMENT|10613,10617|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|SIMPLE_SEGMENT|10613,10617|false|false|false|C1553498|home health encounter|Home
Event|Occupational Activity|SIMPLE_SEGMENT|10623,10630|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|10623,10630|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Event|Event|SIMPLE_SEGMENT|10633,10641|false|false|false|||Facility
Finding|Intellectual Product|SIMPLE_SEGMENT|10633,10641|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|SIMPLE_SEGMENT|10649,10658|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|10649,10658|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|10649,10658|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|10649,10658|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|10649,10658|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|10649,10668|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10659,10668|false|false|false|C0945731||Diagnosis
Event|Event|SIMPLE_SEGMENT|10659,10668|false|false|false|||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|10659,10668|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|10659,10668|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10659,10668|false|false|false|C0011900|Diagnosis|Diagnosis
Event|Event|SIMPLE_SEGMENT|10678,10687|false|false|false|||diagnoses
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10678,10687|false|false|false|C0011900|Diagnosis|diagnoses
Event|Event|SIMPLE_SEGMENT|10689,10696|false|false|false|||Chronic
Finding|Intellectual Product|SIMPLE_SEGMENT|10689,10696|false|false|false|C1547296|Chronic - Admission Level of Care Code|Chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|10689,10696|false|false|false|C1555457|Provision of recurring care for chronic illness|Chronic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10689,10726|false|false|false|C0024117|Chronic Obstructive Airway Disease|Chronic obstructive pulmonary disease
Finding|Functional Concept|SIMPLE_SEGMENT|10697,10708|false|false|false|C0549186|Obstructed|obstructive
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10697,10726|false|false|false|C0600260|Lung Diseases, Obstructive|obstructive pulmonary disease
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10709,10718|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10709,10718|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|10709,10718|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10709,10726|false|false|false|C0024115|Lung diseases|pulmonary disease
Finding|Finding|SIMPLE_SEGMENT|10709,10726|false|false|false|C0455540|History of - respiratory disease|pulmonary disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10719,10726|false|true|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|10719,10726|false|false|false|||disease
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10727,10733|false|false|false|C0018792|Heart Atrium|Atrial
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10727,10746|false|false|false|C2926591||Atrial fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10727,10746|false|false|false|C0004238|Atrial Fibrillation|Atrial fibrillation
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|10727,10746|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Atrial fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10727,10778|false|false|false|C1142306|Atrial fibrillation with rapid ventricular response|Atrial fibrillation with rapid ventricular response
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10727,10778|false|false|false|C3853730|continuous electrocardiogram monitoring atrial fibrillation with rapid ventricular response|Atrial fibrillation with rapid ventricular response
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10734,10746|false|false|false|C0232197|Fibrillation|fibrillation
Event|Event|SIMPLE_SEGMENT|10734,10746|false|false|false|||fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10752,10778|false|false|false|C0748243|rapid ventricular response|rapid ventricular response
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10758,10769|false|false|false|C0018827|Heart Ventricle|ventricular
Event|Event|SIMPLE_SEGMENT|10770,10778|false|false|false|||response
Finding|Finding|SIMPLE_SEGMENT|10770,10778|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Intellectual Product|SIMPLE_SEGMENT|10770,10778|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Mental Process|SIMPLE_SEGMENT|10770,10778|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Disorder|Neoplastic Process|SIMPLE_SEGMENT|10780,10789|false|false|false|C0027627|Neoplasm Metastasis|Secondary
Event|Event|SIMPLE_SEGMENT|10780,10789|false|false|false|||Secondary
Finding|Functional Concept|SIMPLE_SEGMENT|10780,10789|false|false|false|C1522484|metastatic qualifier|Secondary
Event|Event|SIMPLE_SEGMENT|10790,10799|false|false|false|||diagnoses
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10790,10799|false|false|false|C0011900|Diagnosis|diagnoses
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10801,10813|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|SIMPLE_SEGMENT|10801,10813|false|false|false|||Hypertension
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10814,10822|false|false|false|C0018787|Heart|Coronary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10814,10829|false|false|false|C0205042|Coronary artery|Coronary artery
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10814,10837|false|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|Coronary artery disease
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10823,10829|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|SIMPLE_SEGMENT|10823,10829|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10823,10837|false|false|false|C0852949|Arteriopathic disease|artery disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10830,10837|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|10830,10837|false|false|false|||disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10838,10865|false|false|false|C0085096|Peripheral Vascular Diseases|Peripheral vascular disease
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10849,10857|false|false|false|C0005847|Blood Vessel|vascular
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10849,10865|false|false|false|C0042373|Vascular Diseases|vascular disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10858,10865|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|10858,10865|false|false|false|||disease
Event|Event|SIMPLE_SEGMENT|10869,10878|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|10869,10878|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|10869,10878|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|10869,10878|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|10869,10878|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10879,10888|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10879,10888|false|false|false|C0012634|Disease|Condition
Event|Event|SIMPLE_SEGMENT|10879,10888|false|false|false|||Condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|10879,10888|false|false|false|C1705253|Logical Condition|Condition
Finding|Mental Process|SIMPLE_SEGMENT|10890,10896|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10890,10903|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|SIMPLE_SEGMENT|10890,10903|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10897,10903|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|10897,10903|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|10905,10910|false|false|false|||Clear
Finding|Idea or Concept|SIMPLE_SEGMENT|10905,10910|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|SIMPLE_SEGMENT|10915,10923|false|false|false|||coherent
Finding|Finding|SIMPLE_SEGMENT|10915,10923|false|false|false|C4068804|Coherent|coherent
Event|Event|SIMPLE_SEGMENT|10925,10930|false|false|false|||Level
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10925,10947|false|false|false|C4050479||Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|10925,10947|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|SIMPLE_SEGMENT|10934,10947|false|false|false|||Consciousness
Finding|Finding|SIMPLE_SEGMENT|10934,10947|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|SIMPLE_SEGMENT|10934,10947|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10949,10954|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|10949,10954|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10949,10954|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|SIMPLE_SEGMENT|10949,10954|false|false|false|||Alert
Finding|Finding|SIMPLE_SEGMENT|10949,10954|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|10949,10954|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|10949,10954|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|SIMPLE_SEGMENT|10959,10970|false|false|false|||interactive
Finding|Functional Concept|SIMPLE_SEGMENT|10959,10970|false|false|false|C1704675|Interaction|interactive
Event|Activity|SIMPLE_SEGMENT|10972,10980|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|10972,10980|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|SIMPLE_SEGMENT|10972,10980|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10981,10987|false|false|false|C5889824||Status
Event|Event|SIMPLE_SEGMENT|10981,10987|false|false|false|||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|10981,10987|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|10989,10999|false|false|false|||Ambulatory
Finding|Functional Concept|SIMPLE_SEGMENT|10989,10999|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|SIMPLE_SEGMENT|10989,10999|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|SIMPLE_SEGMENT|10989,10999|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|SIMPLE_SEGMENT|10989,10999|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|SIMPLE_SEGMENT|11002,11013|false|false|false|||Independent
Finding|Finding|SIMPLE_SEGMENT|11002,11013|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|SIMPLE_SEGMENT|11002,11013|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Event|Event|SIMPLE_SEGMENT|11018,11027|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|11018,11027|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|11018,11027|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|11018,11027|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|11018,11027|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11018,11040|false|false|false|C3669312||Discharge Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|11018,11040|false|false|false|C4282220|Discharge instructions|Discharge Instructions
Procedure|Health Care Activity|SIMPLE_SEGMENT|11018,11040|false|false|false|C2266673|hospital discharge instructions (treatment)|Discharge Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11028,11040|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|11028,11040|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|11028,11040|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Finding|Gene or Genome|SIMPLE_SEGMENT|11042,11046|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Event|Event|SIMPLE_SEGMENT|11066,11078|false|false|false|||hospitalized
Event|Event|SIMPLE_SEGMENT|11111,11121|false|false|false|||difficulty
Finding|Finding|SIMPLE_SEGMENT|11111,11121|false|false|false|C1299586|Has difficulty doing (qualifier value)|difficulty
Finding|Sign or Symptom|SIMPLE_SEGMENT|11111,11131|false|false|false|C0013404;C0476273|Dyspnea;Respiratory distress|difficulty breathing
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11122,11131|false|false|false|C5885990||breathing
Event|Event|SIMPLE_SEGMENT|11122,11131|false|false|false|||breathing
Finding|Finding|SIMPLE_SEGMENT|11122,11131|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|SIMPLE_SEGMENT|11122,11131|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|SIMPLE_SEGMENT|11122,11131|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|SIMPLE_SEGMENT|11122,11131|false|false|false|C1160636|respiratory system process|breathing
Event|Event|SIMPLE_SEGMENT|11141,11146|false|false|false|||found
Finding|Finding|SIMPLE_SEGMENT|11168,11172|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|fast
Finding|Gene or Genome|SIMPLE_SEGMENT|11168,11172|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|fast
Finding|Molecular Function|SIMPLE_SEGMENT|11168,11172|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|fast
Finding|Finding|SIMPLE_SEGMENT|11168,11183|false|false|false|C0039231|Tachycardia|fast heart rate
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11173,11178|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|11173,11178|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|11173,11178|false|false|false|C0795691|HEART PROBLEM|heart
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11173,11183|false|false|false|C0018810;C0488794|heart rate|heart rate
Finding|Finding|SIMPLE_SEGMENT|11173,11183|false|false|false|C2041121||heart rate
Procedure|Health Care Activity|SIMPLE_SEGMENT|11173,11183|false|false|false|C2197023|examination of heart rate|heart rate
Event|Activity|SIMPLE_SEGMENT|11179,11183|false|false|false|C0871208|Rating (action)|rate
Event|Event|SIMPLE_SEGMENT|11179,11183|false|false|false|||rate
Finding|Idea or Concept|SIMPLE_SEGMENT|11179,11183|false|false|false|C1549480|Amount type - Rate|rate
Event|Event|SIMPLE_SEGMENT|11190,11200|false|false|false|||difficulty
Finding|Finding|SIMPLE_SEGMENT|11190,11200|false|false|false|C1299586|Has difficulty doing (qualifier value)|difficulty
Finding|Sign or Symptom|SIMPLE_SEGMENT|11190,11210|false|false|false|C0013404;C0476273|Dyspnea;Respiratory distress|difficulty breathing
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11201,11210|false|false|false|C5885990||breathing
Event|Event|SIMPLE_SEGMENT|11201,11210|false|false|false|||breathing
Finding|Finding|SIMPLE_SEGMENT|11201,11210|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|SIMPLE_SEGMENT|11201,11210|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|SIMPLE_SEGMENT|11201,11210|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|SIMPLE_SEGMENT|11201,11210|false|false|false|C1160636|respiratory system process|breathing
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11228,11232|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11228,11232|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|SIMPLE_SEGMENT|11228,11232|false|false|false|||COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|11228,11232|false|false|false|C1412502|ARCN1 gene|COPD
Event|Event|SIMPLE_SEGMENT|11233,11240|false|false|false|||flaring
Finding|Finding|SIMPLE_SEGMENT|11247,11251|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|fast
Finding|Gene or Genome|SIMPLE_SEGMENT|11247,11251|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|fast
Finding|Molecular Function|SIMPLE_SEGMENT|11247,11251|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|fast
Finding|Finding|SIMPLE_SEGMENT|11247,11262|false|false|false|C0039231|Tachycardia|fast heart rate
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11252,11257|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|11252,11257|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|11252,11257|false|false|false|C0795691|HEART PROBLEM|heart
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11252,11262|false|false|false|C0018810;C0488794|heart rate|heart rate
Finding|Finding|SIMPLE_SEGMENT|11252,11262|false|false|false|C2041121||heart rate
Procedure|Health Care Activity|SIMPLE_SEGMENT|11252,11262|false|false|false|C2197023|examination of heart rate|heart rate
Event|Activity|SIMPLE_SEGMENT|11258,11262|false|false|false|C0871208|Rating (action)|rate
Event|Event|SIMPLE_SEGMENT|11258,11262|false|false|false|||rate
Finding|Idea or Concept|SIMPLE_SEGMENT|11258,11262|false|false|false|C1549480|Amount type - Rate|rate
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11280,11286|false|false|false|C0018792|Heart Atrium|atrial
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11280,11299|false|false|false|C2926591||atrial fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11280,11299|false|false|false|C0004238|Atrial Fibrillation|atrial fibrillation
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|11280,11299|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|atrial fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11287,11299|false|false|false|C0232197|Fibrillation|fibrillation
Event|Event|SIMPLE_SEGMENT|11287,11299|false|false|false|||fibrillation
Finding|Finding|SIMPLE_SEGMENT|11313,11333|false|false|false|C0237314|Irregular heart beat|irregular heart rate
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11323,11328|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|11323,11328|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|11323,11328|false|false|false|C0795691|HEART PROBLEM|heart
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11323,11333|false|false|false|C0018810;C0488794|heart rate|heart rate
Finding|Finding|SIMPLE_SEGMENT|11323,11333|false|false|false|C2041121||heart rate
Procedure|Health Care Activity|SIMPLE_SEGMENT|11323,11333|false|false|false|C2197023|examination of heart rate|heart rate
Event|Activity|SIMPLE_SEGMENT|11329,11333|false|false|false|C0871208|Rating (action)|rate
Event|Event|SIMPLE_SEGMENT|11329,11333|false|false|false|||rate
Finding|Idea or Concept|SIMPLE_SEGMENT|11329,11333|false|false|false|C1549480|Amount type - Rate|rate
Event|Event|SIMPLE_SEGMENT|11354,11359|false|false|false|||cause
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11364,11369|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|11364,11369|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Event|Event|SIMPLE_SEGMENT|11364,11369|false|false|false|||heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|11364,11369|false|false|false|C0795691|HEART PROBLEM|heart
Event|Event|SIMPLE_SEGMENT|11373,11377|false|false|false|||beat
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11392,11403|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11392,11403|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|11392,11403|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|11392,11403|false|false|false|C4284232|Medications|Medications
Event|Event|SIMPLE_SEGMENT|11419,11425|false|false|false|||taking
Drug|Organic Chemical|SIMPLE_SEGMENT|11435,11447|false|false|false|C0039771|theophylline|theophylline
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11435,11447|false|false|false|C0039771|theophylline|theophylline
Event|Event|SIMPLE_SEGMENT|11435,11447|false|false|false|||theophylline
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|11435,11447|false|false|false|C0039773|Assay of theophylline|theophylline
Finding|Finding|SIMPLE_SEGMENT|11454,11460|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|11454,11460|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|SIMPLE_SEGMENT|11461,11473|false|false|false|||contributing
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11481,11486|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|11481,11486|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|11481,11486|false|false|false|C0795691|HEART PROBLEM|heart
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11481,11491|false|false|false|C0018810;C0488794|heart rate|heart rate
Finding|Finding|SIMPLE_SEGMENT|11481,11491|false|false|false|C2041121||heart rate
Procedure|Health Care Activity|SIMPLE_SEGMENT|11481,11491|false|false|false|C2197023|examination of heart rate|heart rate
Event|Activity|SIMPLE_SEGMENT|11487,11491|false|false|false|C0871208|Rating (action)|rate
Event|Event|SIMPLE_SEGMENT|11487,11491|false|false|false|||rate
Finding|Idea or Concept|SIMPLE_SEGMENT|11487,11491|false|false|false|C1549480|Amount type - Rate|rate
Event|Event|SIMPLE_SEGMENT|11496,11503|false|false|false|||lowered
Event|Event|SIMPLE_SEGMENT|11504,11509|false|false|false|||using
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11519,11529|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|11519,11529|false|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|11519,11529|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|SIMPLE_SEGMENT|11540,11544|false|false|false|||take
Finding|Finding|SIMPLE_SEGMENT|11545,11552|false|false|false|C4534363|At home|at home
Event|Event|SIMPLE_SEGMENT|11548,11552|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|11548,11552|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|11548,11552|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|11548,11552|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|11554,11563|false|false|false|C0012373|diltiazem|diltiazem
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11554,11563|false|false|false|C0012373|diltiazem|diltiazem
Event|Event|SIMPLE_SEGMENT|11554,11563|false|false|false|||diltiazem
Event|Event|SIMPLE_SEGMENT|11565,11570|false|false|false|||given
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11595,11599|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11595,11599|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|SIMPLE_SEGMENT|11595,11599|false|false|false|||COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|11595,11599|false|false|false|C1412502|ARCN1 gene|COPD
Finding|Finding|SIMPLE_SEGMENT|11604,11610|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|11604,11610|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|SIMPLE_SEGMENT|11611,11619|false|false|false|||worsened
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11633,11637|false|false|false|C0009443;C0024117|Chronic Obstructive Airway Disease;Common Cold|cold
Drug|Organic Chemical|SIMPLE_SEGMENT|11633,11637|false|false|false|C0719425|Cold brand of chlorpheniramine-phenylpropanolamine|cold
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11633,11637|false|false|false|C0719425|Cold brand of chlorpheniramine-phenylpropanolamine|cold
Event|Event|SIMPLE_SEGMENT|11633,11637|false|false|false|||cold
Finding|Organism Function|SIMPLE_SEGMENT|11633,11637|false|false|false|C0234192|Cold Sensation|cold
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|11633,11637|false|false|false|C0009264|Cold Temperature|cold
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11633,11637|false|false|false|C0010412|Cold Therapy|cold
Event|Event|SIMPLE_SEGMENT|11654,11659|false|false|false|||flare
Finding|Finding|SIMPLE_SEGMENT|11654,11659|false|false|false|C1517205;C3540542|Exacerbation of cGVHD;Flare|flare
Finding|Sign or Symptom|SIMPLE_SEGMENT|11654,11659|false|false|false|C1517205;C3540542|Exacerbation of cGVHD;Flare|flare
Event|Event|SIMPLE_SEGMENT|11669,11676|false|false|false|||serious
Finding|Finding|SIMPLE_SEGMENT|11669,11676|false|false|false|C1551395;C1552745;C1561576|Alert level - Serious;Device Alert Level - Serious;Equipment Alert Level - Serious|serious
Finding|Idea or Concept|SIMPLE_SEGMENT|11669,11676|false|false|false|C1551395;C1552745;C1561576|Alert level - Serious;Device Alert Level - Serious;Equipment Alert Level - Serious|serious
Event|Event|SIMPLE_SEGMENT|11677,11686|false|false|false|||requiring
Drug|Organic Chemical|SIMPLE_SEGMENT|11690,11698|false|false|false|C0038317|Steroids|steroids
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11690,11698|false|false|false|C0038317|Steroids|steroids
Event|Event|SIMPLE_SEGMENT|11690,11698|false|false|false|||steroids
Finding|Organism Function|SIMPLE_SEGMENT|11708,11715|false|false|false|C0004048|Inspiration (function)|inhaled
Event|Event|SIMPLE_SEGMENT|11717,11727|false|false|false|||treatments
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11717,11727|false|false|false|C0087111|Therapeutic procedure|treatments
Event|Event|SIMPLE_SEGMENT|11740,11746|false|false|false|||follow
Anatomy|Body Location or Region|SIMPLE_SEGMENT|11759,11763|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11759,11763|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11759,11763|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|SIMPLE_SEGMENT|11759,11763|false|false|false|C0740941|Lung Problem|lung
Event|Event|SIMPLE_SEGMENT|11764,11771|false|false|false|||doctors
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11788,11797|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11788,11797|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|11788,11797|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Event|Event|SIMPLE_SEGMENT|11798,11803|false|false|false|||rehab
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11798,11803|false|false|false|C0034991|Rehabilitation therapy|rehab
Event|Event|SIMPLE_SEGMENT|11812,11816|false|false|false|||sure
Finding|Intellectual Product|SIMPLE_SEGMENT|11812,11816|false|false|false|C4724437|SURE Test|sure
Anatomy|Body Location or Region|SIMPLE_SEGMENT|11822,11826|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11822,11826|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11822,11826|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|SIMPLE_SEGMENT|11822,11826|false|false|false|C0740941|Lung Problem|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11822,11834|false|false|false|C0024115|Lung diseases|lung disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11827,11834|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|11827,11834|false|false|false|||disease
Event|Event|SIMPLE_SEGMENT|11838,11843|false|false|false|||being
Event|Event|SIMPLE_SEGMENT|11845,11852|false|false|false|||treated
Event|Event|SIMPLE_SEGMENT|11856,11860|false|false|false|||well
Finding|Finding|SIMPLE_SEGMENT|11856,11860|false|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|11864,11872|false|false|false|||possible
Finding|Finding|SIMPLE_SEGMENT|11864,11872|false|false|false|C0332149|Possible|possible
Event|Event|SIMPLE_SEGMENT|11876,11883|false|false|false|||prevent
Event|Event|SIMPLE_SEGMENT|11893,11899|false|false|false|||coming
Event|Event|SIMPLE_SEGMENT|11910,11918|false|false|false|||hospital
Finding|Idea or Concept|SIMPLE_SEGMENT|11910,11918|false|false|false|C1547192|Organization unit type - Hospital|hospital
Finding|Intellectual Product|SIMPLE_SEGMENT|11922,11927|false|false|false|C4050225|Often - answer to question|often
Event|Event|SIMPLE_SEGMENT|11936,11940|false|false|false|||call
Event|Event|SIMPLE_SEGMENT|11948,11956|false|false|false|||schedule
Event|Activity|SIMPLE_SEGMENT|11961,11972|false|false|false|C0003629|Appointments|appointment
Event|Event|SIMPLE_SEGMENT|11961,11972|false|false|false|||appointment
Event|Event|SIMPLE_SEGMENT|11994,12002|false|false|false|||pleasure
Finding|Intellectual Product|SIMPLE_SEGMENT|11994,12002|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|SIMPLE_SEGMENT|11994,12002|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Event|SIMPLE_SEGMENT|12003,12016|false|false|false|||participating
Event|Activity|SIMPLE_SEGMENT|12025,12029|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|12025,12029|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|12025,12029|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|12025,12029|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Event|Event|SIMPLE_SEGMENT|12034,12038|false|false|false|||wish
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12052,12056|false|false|false|C0339510|Vitelliform Macular Dystrophy|best
Event|Event|SIMPLE_SEGMENT|12052,12056|false|false|false|||best
Finding|Gene or Genome|SIMPLE_SEGMENT|12052,12056|false|false|false|C1826421;C5781213|BEST1 gene;BEST1 wt Allele|best
Procedure|Health Care Activity|SIMPLE_SEGMENT|12101,12109|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12110,12122|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|12110,12122|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|12110,12122|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

