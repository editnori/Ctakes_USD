 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|29,33
No|34,36
:|36,37
_|40,41
_|41,42
_|42,43
<EOL>|43,44
<EOL>|45,46
Admission|46,55
Date|56,60
:|60,61
_|63,64
_|64,65
_|65,66
Discharge|80,89
Date|90,94
:|94,95
_|98,99
_|99,100
_|100,101
<EOL>|101,102
<EOL>|103,104
Date|104,108
of|109,111
Birth|112,117
:|117,118
_|120,121
_|121,122
_|122,123
Sex|136,139
:|139,140
F|143,144
<EOL>|144,145
<EOL>|146,147
Service|147,154
:|154,155
ORTHOPAEDICS|156,168
<EOL>|168,169
<EOL>|170,171
Allergies|171,180
:|180,181
<EOL>|182,183
omeprazole|183,193
/|194,195
Iodine|196,202
and|203,206
Iodide|207,213
Containing|214,224
Products|225,233
/|234,235
<EOL>|236,237
hallucinogens|237,250
<EOL>|250,251
<EOL>|252,253
Attending|253,262
:|262,263
_|264,265
_|265,266
_|266,267
.|267,268
<EOL>|268,269
<EOL>|270,271
Chief|271,276
Complaint|277,286
:|286,287
<EOL>|287,288
Left|288,292
hip|293,296
pain|297,301
<EOL>|302,303
<EOL>|304,305
Major|305,310
Surgical|311,319
or|320,322
Invasive|323,331
Procedure|332,341
:|341,342
<EOL>|342,343
Status|343,349
post|350,354
left|355,359
CRPP|360,364
_|365,366
_|366,367
_|367,368
,|368,369
_|370,371
_|371,372
_|372,373
<EOL>|373,374
<EOL>|374,375
<EOL>|376,377
History|377,384
of|385,387
Present|388,395
Illness|396,403
:|403,404
<EOL>|404,405
REASON|405,411
FOR|412,415
CONSULT|416,423
:|423,424
Femur|425,430
fracture|431,439
<EOL>|439,440
<EOL>|440,441
HPI|441,444
:|444,445
_|446,447
_|447,448
_|448,449
female|450,456
presents|457,465
with|466,470
the|471,474
above|475,480
fracture|481,489
s|490,491
/|491,492
p|492,493
mechanical|494,504
<EOL>|504,505
fall|505,509
.|509,510
This|511,515
morning|516,523
,|523,524
pt|525,527
was|528,531
walking|532,539
_|540,541
_|541,542
_|542,543
,|543,544
when|545,549
dog|550,553
<EOL>|553,554
pulled|554,560
on|561,563
leash|564,569
.|569,570
Pt|571,573
fell|574,578
on|579,581
L|582,583
hip.|584,588
Immediate|589,598
pain|599,603
.|603,604
_|605,606
_|606,607
_|607,608
_|609,610
_|610,611
_|611,612
with|613,617
movement|618,626
.|626,627
Denies|628,634
Head|635,639
strike|640,646
,|646,647
LOC|648,651
or|652,654
blood|655,660
thinners|661,669
.|669,670
<EOL>|670,671
Denies|671,677
numbness|678,686
or|687,689
weakness|690,698
in|699,701
the|702,705
extremities|706,717
.|717,718
<EOL>|719,720
<EOL>|721,722
Past|722,726
Medical|727,734
History|735,742
:|742,743
<EOL>|743,744
-|744,745
GERD|746,750
<EOL>|752,753
-|754,755
Hypercholesterolemia|756,776
<EOL>|778,779
-|780,781
Kidney|782,788
stones|789,795
<EOL>|797,798
-|799,800
Mitral|801,807
valve|808,813
prolapse|814,822
<EOL>|824,825
-|826,827
Uterine|828,835
fibroids|836,844
<EOL>|846,847
-|848,849
Osteoporosis|850,862
<EOL>|864,865
-|866,867
Migraine|868,876
headaches|877,886
<EOL>|887,888
<EOL>|889,890
Social|890,896
History|897,904
:|904,905
<EOL>|905,906
_|906,907
_|907,908
_|908,909
<EOL>|909,910
Family|910,916
History|917,924
:|924,925
<EOL>|925,926
+|926,927
HTN|928,931
-|932,933
father|934,940
<EOL>|942,943
+|943,944
Dementia|945,953
-|954,955
father|956,962
<EOL>|964,965
<EOL>|966,967
<EOL>|968,969
Physical|969,977
Exam|978,982
:|982,983
<EOL>|983,984
General|984,991
:|991,992
Well|993,997
-|997,998
appearing|998,1007
female|1008,1014
in|1015,1017
no|1018,1020
acute|1021,1026
distress|1027,1035
.|1035,1036
<EOL>|1036,1037
<EOL>|1037,1038
Left|1038,1042
Lower|1043,1048
extremity|1049,1058
:|1058,1059
<EOL>|1059,1060
-|1060,1061
Skin|1062,1066
intact|1067,1073
<EOL>|1073,1074
-|1074,1075
No|1076,1078
deformity|1079,1088
,|1088,1089
edema|1090,1095
,|1095,1096
ecchymosis|1097,1107
,|1107,1108
erythema|1109,1117
,|1117,1118
induration|1119,1129
<EOL>|1129,1130
-|1130,1131
Soft|1132,1136
,|1136,1137
non-tender|1138,1148
thigh|1149,1154
and|1155,1158
leg|1159,1162
<EOL>|1162,1163
-|1163,1164
Full|1165,1169
,|1169,1170
painless|1171,1179
ROM|1180,1183
knee|1184,1188
,|1188,1189
and|1190,1193
ankle|1194,1199
<EOL>|1199,1200
-|1200,1201
Fires|1202,1207
_|1208,1209
_|1209,1210
_|1210,1211
<EOL>|1211,1212
-|1212,1213
SILT|1214,1218
S|1219,1220
/|1220,1221
S|1221,1222
/|1222,1223
SP|1223,1225
/|1225,1226
DP|1226,1228
/|1228,1229
T|1229,1230
distributions|1231,1244
<EOL>|1244,1245
-|1245,1246
1|1247,1248
+|1248,1249
_|1250,1251
_|1251,1252
_|1252,1253
pulses|1254,1260
,|1260,1261
WWP|1262,1265
<EOL>|1265,1266
<EOL>|1267,1268
Brief|1268,1273
Hospital|1274,1282
Course|1283,1289
:|1289,1290
<EOL>|1290,1291
The|1291,1294
patient|1295,1302
presented|1303,1312
to|1313,1315
the|1316,1319
emergency|1320,1329
department|1330,1340
and|1341,1344
was|1345,1348
<EOL>|1349,1350
evaluated|1350,1359
by|1360,1362
the|1363,1366
orthopedic|1367,1377
surgery|1378,1385
team|1386,1390
.|1390,1391
The|1392,1395
patient|1396,1403
was|1404,1407
found|1408,1413
<EOL>|1414,1415
to|1415,1417
have|1418,1422
a|1423,1424
left|1425,1429
valgus|1430,1436
impacted|1437,1445
femoral|1446,1453
neck|1454,1458
fracture|1459,1467
and|1468,1471
was|1472,1475
<EOL>|1476,1477
admitted|1477,1485
to|1486,1488
the|1489,1492
orthopedic|1493,1503
surgery|1504,1511
service|1512,1519
.|1519,1520
The|1521,1524
patient|1525,1532
was|1533,1536
<EOL>|1537,1538
taken|1538,1543
to|1544,1546
the|1547,1550
operating|1551,1560
room|1561,1565
on|1566,1568
_|1569,1570
_|1570,1571
_|1571,1572
for|1573,1576
left|1577,1581
closed|1582,1588
reduction|1589,1598
<EOL>|1599,1600
and|1600,1603
percutaneous|1604,1616
pinning|1617,1624
of|1625,1627
hip|1628,1631
,|1631,1632
which|1633,1638
the|1639,1642
patient|1643,1650
tolerated|1651,1660
<EOL>|1661,1662
well|1662,1666
.|1666,1667
For|1668,1671
full|1672,1676
details|1677,1684
of|1685,1687
the|1688,1691
procedure|1692,1701
please|1702,1708
see|1709,1712
the|1713,1716
<EOL>|1717,1718
separately|1718,1728
dictated|1729,1737
operative|1738,1747
report|1748,1754
.|1754,1755
The|1756,1759
patient|1760,1767
was|1768,1771
taken|1772,1777
from|1778,1782
<EOL>|1783,1784
the|1784,1787
OR|1788,1790
to|1791,1793
the|1794,1797
PACU|1798,1802
in|1803,1805
stable|1806,1812
condition|1813,1822
and|1823,1826
after|1827,1832
satisfactory|1833,1845
<EOL>|1846,1847
recovery|1847,1855
from|1856,1860
anesthesia|1861,1871
was|1872,1875
transferred|1876,1887
to|1888,1890
the|1891,1894
floor|1895,1900
.|1900,1901
The|1902,1905
<EOL>|1906,1907
patient|1907,1914
was|1915,1918
initially|1919,1928
given|1929,1934
IV|1935,1937
fluids|1938,1944
and|1945,1948
IV|1949,1951
pain|1952,1956
medications|1957,1968
,|1968,1969
<EOL>|1970,1971
and|1971,1974
progressed|1975,1985
to|1986,1988
a|1989,1990
regular|1991,1998
diet|1999,2003
and|2004,2007
oral|2008,2012
medications|2013,2024
by|2025,2027
POD|2028,2031
#|2031,2032
1|2032,2033
.|2033,2034
<EOL>|2035,2036
The|2036,2039
patient|2040,2047
was|2048,2051
given|2052,2057
_|2058,2059
_|2059,2060
_|2060,2061
antibiotics|2062,2073
and|2074,2077
<EOL>|2078,2079
anticoagulation|2079,2094
per|2095,2098
routine|2099,2106
.|2106,2107
The|2108,2111
patient|2112,2119
's|2119,2121
home|2122,2126
medications|2127,2138
were|2139,2143
<EOL>|2144,2145
continued|2145,2154
throughout|2155,2165
this|2166,2170
hospitalization|2171,2186
.|2186,2187
The|2188,2191
patient|2192,2199
worked|2200,2206
<EOL>|2207,2208
with|2208,2212
_|2213,2214
_|2214,2215
_|2215,2216
who|2217,2220
determined|2221,2231
that|2232,2236
discharge|2237,2246
to|2247,2249
home|2250,2254
with|2255,2259
services|2260,2268
was|2269,2272
<EOL>|2273,2274
appropriate|2274,2285
.|2285,2286
The|2287,2290
_|2291,2292
_|2292,2293
_|2293,2294
hospital|2295,2303
course|2304,2310
was|2311,2314
otherwise|2315,2324
<EOL>|2325,2326
unremarkable|2326,2338
.|2338,2339
<EOL>|2339,2340
<EOL>|2340,2341
At|2341,2343
the|2344,2347
time|2348,2352
of|2353,2355
discharge|2356,2365
the|2366,2369
patient|2370,2377
's|2377,2379
pain|2380,2384
was|2385,2388
well|2389,2393
controlled|2394,2404
<EOL>|2405,2406
with|2406,2410
oral|2411,2415
medications|2416,2427
,|2427,2428
incisions|2429,2438
were|2439,2443
clean|2444,2449
/|2449,2450
dry|2450,2453
/|2453,2454
intact|2454,2460
,|2460,2461
and|2462,2465
the|2466,2469
<EOL>|2470,2471
patient|2471,2478
was|2479,2482
voiding|2483,2490
/|2490,2491
moving|2491,2497
bowels|2498,2504
spontaneously|2505,2518
.|2518,2519
The|2520,2523
patient|2524,2531
is|2532,2534
<EOL>|2536,2537
weightbearing|2537,2550
as|2551,2553
tolerated|2554,2563
in|2564,2566
the|2567,2570
left|2571,2575
lower|2576,2581
extremity|2582,2591
,|2591,2592
and|2593,2596
will|2597,2601
<EOL>|2602,2603
be|2603,2605
discharged|2606,2616
on|2617,2619
Lovenox|2620,2627
for|2628,2631
DVT|2632,2635
prophylaxis|2636,2647
.|2647,2648
The|2649,2652
patient|2653,2660
will|2661,2665
<EOL>|2666,2667
follow|2667,2673
up|2674,2676
with|2677,2681
Dr.|2682,2685
_|2686,2687
_|2687,2688
_|2688,2689
routine|2690,2697
.|2697,2698
A|2699,2700
thorough|2701,2709
discussion|2710,2720
<EOL>|2721,2722
was|2722,2725
had|2726,2729
with|2730,2734
the|2735,2738
patient|2739,2746
regarding|2747,2756
the|2757,2760
diagnosis|2761,2770
and|2771,2774
expected|2775,2783
<EOL>|2784,2785
post-discharge|2785,2799
course|2800,2806
including|2807,2816
reasons|2817,2824
to|2825,2827
call|2828,2832
the|2833,2836
office|2837,2843
or|2844,2846
<EOL>|2847,2848
return|2848,2854
to|2855,2857
the|2858,2861
hospital|2862,2870
,|2870,2871
and|2872,2875
all|2876,2879
questions|2880,2889
were|2890,2894
answered|2895,2903
.|2903,2904
The|2905,2908
<EOL>|2909,2910
patient|2910,2917
was|2918,2921
also|2922,2926
given|2927,2932
written|2933,2940
instructions|2941,2953
concerning|2954,2964
<EOL>|2965,2966
precautionary|2966,2979
instructions|2980,2992
and|2993,2996
the|2997,3000
appropriate|3001,3012
follow|3013,3019
-|3019,3020
up|3020,3022
care|3023,3027
.|3027,3028
<EOL>|3029,3030
The|3030,3033
patient|3034,3041
expressed|3042,3051
readiness|3052,3061
for|3062,3065
discharge|3066,3075
.|3075,3076
<EOL>|3076,3077
<EOL>|3077,3078
<EOL>|3079,3080
Medications|3080,3091
on|3092,3094
Admission|3095,3104
:|3104,3105
<EOL>|3105,3106
The|3106,3109
Preadmission|3110,3122
Medication|3123,3133
list|3134,3138
is|3139,3141
accurate|3142,3150
and|3151,3154
complete|3155,3163
.|3163,3164
<EOL>|3164,3165
1.|3165,3167
Lactaid|3168,3175
(|3176,3177
lactase|3177,3184
)|3184,3185
3,000|3186,3191
unit|3192,3196
oral|3197,3201
DAILY|3202,3207
:|3207,3208
PRN|3208,3211
<EOL>|3212,3213
2|3213,3214
.|3214,3215
Calcium|3216,3223
Citrate|3224,3231
+|3232,3233
D|3234,3235
(|3236,3237
calcium|3237,3244
citrate|3245,3252
-|3252,3253
vitamin|3253,3260
D3|3261,3263
)|3263,3264
315|3265,3268
-|3268,3269
200|3269,3272
<EOL>|3273,3274
mg|3274,3276
-|3276,3277
unit|3277,3281
oral|3282,3286
DAILY|3287,3292
<EOL>|3293,3294
<EOL>|3294,3295
<EOL>|3296,3297
Discharge|3297,3306
Medications|3307,3318
:|3318,3319
<EOL>|3319,3320
1.|3320,3322
Acetaminophen|3324,3337
1000|3338,3342
mg|3343,3345
PO|3346,3348
Q6H|3349,3352
:|3352,3353
PRN|3353,3356
Pain|3357,3361
-|3362,3363
Mild|3364,3368
/|3368,3369
Fever|3369,3374
<EOL>|3376,3377
2.|3377,3379
Bisacodyl|3381,3390
10|3391,3393
mg|3394,3396
PO|3397,3399
/|3399,3400
PR|3400,3402
DAILY|3403,3408
:|3408,3409
PRN|3409,3412
Constipation|3413,3425
<EOL>|3427,3428
3.|3428,3430
Docusate|3432,3440
Sodium|3441,3447
100|3448,3451
mg|3452,3454
PO|3455,3457
BID|3458,3461
<EOL>|3463,3464
4.|3464,3466
Enoxaparin|3468,3478
Sodium|3479,3485
40|3486,3488
mg|3489,3491
SC|3492,3494
QHS|3495,3498
<EOL>|3499,3500
RX|3500,3502
*|3503,3504
enoxaparin|3504,3514
40|3515,3517
mg|3518,3520
/|3520,3521
0.4|3521,3524
mL|3525,3527
40|3528,3530
mg|3531,3533
Subcutaneously|3534,3548
Nightly|3549,3556
Disp|3557,3561
<EOL>|3562,3563
#|3563,3564
*|3564,3565
30|3565,3567
Syringe|3568,3575
Refills|3576,3583
:|3583,3584
*|3584,3585
0|3585,3586
<EOL>|3587,3588
5.|3588,3590
OxyCODONE|3592,3601
(|3602,3603
Immediate|3603,3612
Release|3613,3620
)|3620,3621
_|3622,3623
_|3623,3624
_|3624,3625
mg|3626,3628
PO|3629,3631
Q4H|3632,3635
:|3635,3636
PRN|3636,3639
Pain|3640,3644
-|3645,3646
<EOL>|3647,3648
Moderate|3648,3656
<EOL>|3657,3658
RX|3658,3660
*|3661,3662
oxycodone|3662,3671
5|3672,3673
mg|3674,3676
1|3677,3678
tablet|3679,3685
(|3685,3686
s|3686,3687
)|3687,3688
by|3689,3691
mouth|3692,3697
q4|3698,3700
PRN|3701,3704
Disp|3705,3709
#|3710,3711
*|3711,3712
25|3712,3714
Tablet|3715,3721
<EOL>|3722,3723
Refills|3723,3730
:|3730,3731
*|3731,3732
0|3732,3733
<EOL>|3734,3735
6.|3735,3737
Senna|3739,3744
8.6|3745,3748
mg|3749,3751
PO|3752,3754
BID|3755,3758
<EOL>|3760,3761
7.|3761,3763
Calcium|3765,3772
Citrate|3773,3780
+|3781,3782
D|3783,3784
(|3785,3786
calcium|3786,3793
citrate|3794,3801
-|3801,3802
vitamin|3802,3809
D3|3810,3812
)|3812,3813
315|3814,3817
-|3817,3818
200|3818,3821
<EOL>|3822,3823
mg|3823,3825
-|3825,3826
unit|3826,3830
oral|3831,3835
DAILY|3836,3841
<EOL>|3843,3844
8.|3844,3846
Lactaid|3848,3855
(|3856,3857
lactase|3857,3864
)|3864,3865
3,000|3866,3871
unit|3872,3876
oral|3877,3881
DAILY|3882,3887
:|3887,3888
PRN|3888,3891
<EOL>|3893,3894
9.|3894,3896
Multivitamins|3898,3911
1|3912,3913
TAB|3914,3917
PO|3918,3920
DAILY|3921,3926
<EOL>|3928,3929
10|3929,3931
.|3931,3932
Vitamin|3934,3941
D|3942,3943
400|3944,3947
UNIT|3948,3952
PO|3953,3955
DAILY|3956,3961
<EOL>|3963,3964
<EOL>|3964,3965
<EOL>|3966,3967
Discharge|3967,3976
Disposition|3977,3988
:|3988,3989
<EOL>|3989,3990
Home|3990,3994
With|3995,3999
Service|4000,4007
<EOL>|4007,4008
<EOL>|4009,4010
Facility|4010,4018
:|4018,4019
<EOL>|4019,4020
_|4020,4021
_|4021,4022
_|4022,4023
<EOL>|4023,4024
<EOL>|4025,4026
Discharge|4026,4035
Diagnosis|4036,4045
:|4045,4046
<EOL>|4046,4047
Left|4047,4051
valgus|4052,4058
impacted|4059,4067
femoral|4068,4075
neck|4076,4080
fracture|4081,4089
<EOL>|4089,4090
<EOL>|4090,4091
<EOL>|4092,4093
Discharge|4093,4102
Condition|4103,4112
:|4112,4113
<EOL>|4113,4114
AVSS|4114,4118
<EOL>|4118,4119
NAD|4119,4122
,|4122,4123
A|4124,4125
&|4125,4126
Ox3|4126,4129
<EOL>|4129,4130
LLE|4130,4133
:|4133,4134
Incision|4135,4143
well|4144,4148
approximated|4149,4161
.|4161,4162
Dressing|4163,4171
clean|4172,4177
and|4178,4181
dry|4182,4185
.|4185,4186
Fires|4187,4192
<EOL>|4193,4194
FHL|4194,4197
,|4197,4198
_|4199,4200
_|4200,4201
_|4201,4202
,|4202,4203
TA|4204,4206
,|4206,4207
GCS|4208,4211
.|4211,4212
SILT|4213,4217
_|4218,4219
_|4219,4220
_|4220,4221
n|4222,4223
distributions|4224,4237
.|4237,4238
1|4239,4240
+|4240,4241
DP|4242,4244
<EOL>|4245,4246
pulse|4246,4251
,|4251,4252
wwp|4253,4256
distally|4257,4265
.|4265,4266
<EOL>|4266,4267
<EOL>|4267,4268
<EOL>|4269,4270
Discharge|4270,4279
Instructions|4280,4292
:|4292,4293
<EOL>|4293,4294
INSTRUCTIONS|4294,4306
AFTER|4307,4312
ORTHOPAEDIC|4313,4324
SURGERY|4325,4332
:|4332,4333
<EOL>|4333,4334
<EOL>|4334,4335
-|4335,4336
You|4337,4340
were|4341,4345
in|4346,4348
the|4349,4352
hospital|4353,4361
for|4362,4365
orthopedic|4366,4376
surgery|4377,4384
.|4384,4385
It|4386,4388
is|4389,4391
normal|4392,4398
<EOL>|4399,4400
to|4400,4402
feel|4403,4407
tired|4408,4413
or|4414,4416
"|4417,4418
washed|4418,4424
out|4425,4428
"|4428,4429
after|4430,4435
surgery|4436,4443
,|4443,4444
and|4445,4448
this|4449,4453
feeling|4454,4461
<EOL>|4462,4463
should|4463,4469
improve|4470,4477
over|4478,4482
the|4483,4486
first|4487,4492
few|4493,4496
days|4497,4501
to|4502,4504
week|4505,4509
.|4509,4510
<EOL>|4511,4512
-|4512,4513
Resume|4514,4520
your|4521,4525
regular|4526,4533
activities|4534,4544
as|4545,4547
tolerated|4548,4557
,|4557,4558
but|4559,4562
please|4563,4569
follow|4570,4576
<EOL>|4577,4578
your|4578,4582
weight|4583,4589
bearing|4590,4597
precautions|4598,4609
strictly|4610,4618
at|4619,4621
all|4622,4625
times|4626,4631
.|4631,4632
<EOL>|4632,4633
<EOL>|4633,4634
ACTIVITY|4634,4642
AND|4643,4646
WEIGHT|4647,4653
BEARING|4654,4661
:|4661,4662
<EOL>|4662,4663
-|4663,4664
Weightbearing|4665,4678
as|4679,4681
tolerated|4682,4691
left|4692,4696
lower|4697,4702
extremity|4703,4712
<EOL>|4712,4713
<EOL>|4713,4714
MEDICATIONS|4714,4725
:|4725,4726
<EOL>|4726,4727
1|4729,4730
)|4730,4731
Take|4733,4737
Tylenol|4738,4745
_|4746,4747
_|4747,4748
_|4748,4749
every|4750,4755
6|4756,4757
hours|4758,4763
around|4764,4770
the|4771,4774
clock|4775,4780
.|4780,4781
This|4782,4786
is|4787,4789
<EOL>|4790,4791
an|4791,4793
over|4794,4798
the|4799,4802
counter|4803,4810
medication|4811,4821
.|4821,4822
<EOL>|4822,4823
2|4825,4826
)|4826,4827
Add|4829,4832
oxycodone|4833,4842
as|4843,4845
needed|4846,4852
for|4853,4856
increased|4857,4866
pain|4867,4871
.|4871,4872
Aim|4873,4876
to|4877,4879
wean|4880,4884
<EOL>|4885,4886
off|4886,4889
this|4890,4894
medication|4895,4905
in|4906,4908
1|4909,4910
week|4911,4915
or|4916,4918
sooner|4919,4925
.|4925,4926
This|4928,4932
is|4933,4935
an|4936,4938
example|4939,4946
on|4947,4949
<EOL>|4950,4951
how|4951,4954
to|4955,4957
wean|4958,4962
down|4963,4967
:|4967,4968
<EOL>|4968,4969
Take|4969,4973
1|4974,4975
tablet|4976,4982
every|4983,4988
3|4989,4990
hours|4991,4996
as|4997,4999
needed|5000,5006
x|5007,5008
1|5009,5010
day|5011,5014
,|5014,5015
<EOL>|5015,5016
then|5016,5020
1|5021,5022
tablet|5023,5029
every|5030,5035
4|5036,5037
hours|5038,5043
as|5044,5046
needed|5047,5053
x|5054,5055
1|5056,5057
day|5058,5061
,|5061,5062
<EOL>|5062,5063
then|5063,5067
1|5068,5069
tablet|5070,5076
every|5077,5082
6|5083,5084
hours|5085,5090
as|5091,5093
needed|5094,5100
x|5101,5102
1|5103,5104
day|5105,5108
,|5108,5109
<EOL>|5109,5110
then|5110,5114
1|5115,5116
tablet|5117,5123
every|5124,5129
8|5130,5131
hours|5132,5137
as|5138,5140
needed|5141,5147
x|5148,5149
2|5150,5151
days|5152,5156
,|5156,5157
<EOL>|5158,5159
then|5159,5163
1|5164,5165
tablet|5166,5172
every|5173,5178
12|5179,5181
hours|5182,5187
as|5188,5190
needed|5191,5197
x|5198,5199
1|5200,5201
day|5202,5205
,|5205,5206
<EOL>|5206,5207
then|5207,5211
1|5212,5213
tablet|5214,5220
every|5221,5226
before|5227,5233
bedtime|5234,5241
as|5242,5244
needed|5245,5251
x|5252,5253
1|5254,5255
day|5256,5259
.|5259,5260
<EOL>|5262,5263
Then|5263,5267
continue|5268,5276
with|5277,5281
Tylenol|5282,5289
for|5290,5293
pain|5294,5298
.|5298,5299
<EOL>|5299,5300
3|5302,5303
)|5303,5304
Do|5306,5308
not|5309,5312
stop|5313,5317
the|5318,5321
Tylenol|5322,5329
until|5330,5335
you|5336,5339
are|5340,5343
off|5344,5347
of|5348,5350
the|5351,5354
narcotic|5355,5363
<EOL>|5364,5365
medication|5365,5375
.|5375,5376
<EOL>|5376,5377
4|5379,5380
)|5380,5381
Per|5383,5386
state|5387,5392
regulations|5393,5404
,|5404,5405
we|5406,5408
are|5409,5412
limited|5413,5420
in|5421,5423
the|5424,5427
amount|5428,5434
of|5435,5437
<EOL>|5438,5439
narcotics|5439,5448
we|5449,5451
can|5452,5455
prescribe|5456,5465
.|5465,5466
If|5467,5469
you|5470,5473
require|5474,5481
more|5482,5486
,|5486,5487
you|5488,5491
must|5492,5496
<EOL>|5497,5498
contact|5498,5505
the|5506,5509
office|5510,5516
to|5517,5519
set|5520,5523
up|5524,5526
an|5527,5529
appointment|5530,5541
because|5542,5549
we|5550,5552
can|5553,5556
not|5556,5559
<EOL>|5560,5561
refill|5561,5567
this|5568,5572
type|5573,5577
of|5578,5580
pain|5581,5585
medication|5586,5596
over|5597,5601
the|5602,5605
phone|5606,5611
.|5611,5612
<EOL>|5613,5614
5|5616,5617
)|5617,5618
Narcotic|5620,5628
pain|5629,5633
relievers|5634,5643
can|5644,5647
cause|5648,5653
constipation|5654,5666
,|5666,5667
so|5668,5670
you|5671,5674
<EOL>|5675,5676
should|5676,5682
drink|5683,5688
eight|5689,5694
8oz|5695,5698
glasses|5699,5706
of|5707,5709
water|5710,5715
daily|5716,5721
and|5722,5725
continue|5726,5734
<EOL>|5735,5736
following|5736,5745
the|5746,5749
bowel|5750,5755
regimen|5756,5763
as|5764,5766
stated|5767,5773
on|5774,5776
your|5777,5781
medication|5782,5792
<EOL>|5793,5794
prescription|5794,5806
list|5807,5811
.|5811,5812
These|5813,5818
meds|5819,5823
(|5824,5825
senna|5825,5830
,|5830,5831
colace|5832,5838
,|5838,5839
miralax|5840,5847
)|5847,5848
are|5849,5852
over|5853,5857
<EOL>|5858,5859
the|5859,5862
counter|5863,5870
and|5871,5874
may|5875,5878
be|5879,5881
obtained|5882,5890
at|5891,5893
any|5894,5897
pharmacy|5898,5906
.|5906,5907
<EOL>|5907,5908
6|5910,5911
)|5911,5912
Do|5914,5916
not|5917,5920
drink|5921,5926
alcohol|5927,5934
,|5934,5935
drive|5936,5941
a|5942,5943
motor|5944,5949
vehicle|5950,5957
,|5957,5958
or|5959,5961
operate|5962,5969
<EOL>|5970,5971
machinery|5971,5980
while|5981,5986
taking|5987,5993
narcotic|5994,6002
pain|6003,6007
relievers|6008,6017
.|6017,6018
<EOL>|6018,6019
7|6021,6022
)|6022,6023
Please|6025,6031
take|6032,6036
all|6037,6040
medications|6041,6052
as|6053,6055
prescribed|6056,6066
by|6067,6069
your|6070,6074
<EOL>|6075,6076
physicians|6076,6086
at|6087,6089
discharge|6090,6099
.|6099,6100
<EOL>|6100,6101
8|6103,6104
)|6104,6105
Continue|6107,6115
all|6116,6119
home|6120,6124
medications|6125,6136
unless|6137,6143
specifically|6144,6156
<EOL>|6157,6158
instructed|6158,6168
to|6169,6171
stop|6172,6176
by|6177,6179
your|6180,6184
surgeon|6185,6192
.|6192,6193
<EOL>|6193,6194
<EOL>|6200,6201
ANTICOAGULATION|6201,6216
:|6216,6217
<EOL>|6217,6218
-|6218,6219
Please|6220,6226
take|6227,6231
Lovenox|6233,6240
daily|6241,6246
for|6247,6250
4|6251,6252
weeks|6253,6258
<EOL>|6258,6259
<EOL>|6260,6261
Followup|6261,6269
Instructions|6270,6282
:|6282,6283
<EOL>|6283,6284
_|6284,6285
_|6285,6286
_|6286,6287
<EOL>|6287,6288

