 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|33,37
No|38,40
:|40,41
_|44,45
_|45,46
_|46,47
<EOL>|47,48
<EOL>|49,50
Admission|50,59
Date|60,64
:|64,65
_|67,68
_|68,69
_|69,70
Discharge|84,93
Date|94,98
:|98,99
_|102,103
_|103,104
_|104,105
<EOL>|105,106
<EOL>|107,108
Date|108,112
of|113,115
Birth|116,121
:|121,122
_|124,125
_|125,126
_|126,127
Sex|140,143
:|143,144
F|147,148
<EOL>|148,149
<EOL>|150,151
Service|151,158
:|158,159
UROLOGY|160,167
<EOL>|167,168
<EOL>|169,170
Patient|182,189
recorded|190,198
as|199,201
having|202,208
No|209,211
Known|212,217
Allergies|218,227
to|228,230
Drugs|231,236
<EOL>|236,237
<EOL>|238,239
Attending|239,248
:|248,249
_|250,251
_|251,252
_|252,253
.|253,254
<EOL>|254,255
<EOL>|256,257
renal|274,279
mass|280,284
<EOL>|284,285
<EOL>|286,287
Major|287,292
Surgical|293,301
or|302,304
Invasive|305,313
Procedure|314,323
:|323,324
<EOL>|324,325
right|325,330
laparascopic|331,343
radical|344,351
nephrectomy|352,363
-|363,364
Dr.|365,368
_|369,370
_|370,371
_|371,372
,|372,373
Dr|374,376
.|376,377
<EOL>|378,379
_|379,380
_|380,381
_|381,382
_|383,384
_|384,385
_|385,386
<EOL>|386,387
<EOL>|387,388
<EOL>|389,390
_|418,419
_|419,420
_|420,421
y|422,423
/|423,424
o|424,425
healthy|426,433
female|434,440
with|441,445
incidental|446,456
finding|457,464
of|465,467
right|468,473
renal|474,479
<EOL>|480,481
mass|481,485
suspicious|486,496
for|497,500
RCC|501,504
following|505,514
MRI|515,518
on|519,521
_|522,523
_|523,524
_|524,525
.|525,526
<EOL>|527,528
<EOL>|529,530
PMH|552,555
:|555,556
nonspecific|557,568
right|569,574
axis|575,579
deviation|580,589
<EOL>|591,592
<EOL>|592,593
PSH|593,596
-|596,597
cesarean|598,606
section|607,614
<EOL>|614,615
<EOL>|615,616
ALL|616,619
-|619,620
NKDA|620,624
<EOL>|624,625
<EOL>|626,627
:|641,642
<EOL>|642,643
_|643,644
_|644,645
_|645,646
<EOL>|646,647
:|661,662
<EOL>|662,663
no|663,665
history|666,673
of|674,676
RCC|677,680
<EOL>|680,681
<EOL>|682,683
Pertinent|683,692
Results|693,700
:|700,701
<EOL>|701,702
_|702,703
_|703,704
_|704,705
07|706,708
:|708,709
15AM|709,713
BLOOD|714,719
WBC|720,723
-|723,724
7.6|724,727
RBC|728,731
-|731,732
3|732,733
.|733,734
82|734,736
*|736,737
Hgb|738,741
-|741,742
11|742,744
.|744,745
9|745,746
*|746,747
Hct|748,751
-|751,752
33|752,754
.|754,755
8|755,756
*|756,757
<EOL>|758,759
MCV|759,762
-|762,763
89|763,765
MCH|766,769
-|769,770
31.2|770,774
MCHC|775,779
-|779,780
35|780,782
.|782,783
2|783,784
*|784,785
RDW|786,789
-|789,790
12.8|790,794
Plt|795,798
_|799,800
_|800,801
_|801,802
<EOL>|802,803
_|803,804
_|804,805
_|805,806
07|807,809
:|809,810
15AM|810,814
BLOOD|815,820
Glucose|821,828
-|828,829
150|829,832
*|832,833
UreaN|834,839
-|839,840
10|840,842
Creat|843,848
-|848,849
0.9|849,852
Na|853,855
-|855,856
138|856,859
<EOL>|860,861
K|861,862
-|862,863
3.8|863,866
Cl|867,869
-|869,870
104|870,873
HCO3|874,878
-|878,879
27|879,881
AnGap|882,887
-|887,888
11|888,890
<EOL>|890,891
<EOL>|892,893
Patient|916,923
was|924,927
admitted|928,936
to|937,939
Urology|940,947
after|948,953
undergoing|954,964
laparoscopic|965,977
<EOL>|978,979
right|979,984
radical|985,992
nephrectomy|993,1004
.|1004,1005
No|1006,1008
concerning|1009,1019
intraoperative|1020,1034
events|1035,1041
<EOL>|1042,1043
occurred|1043,1051
;|1051,1052
please|1053,1059
see|1060,1063
dictated|1064,1072
operative|1073,1082
note|1083,1087
for|1088,1091
details|1092,1099
.|1099,1100
The|1101,1104
<EOL>|1105,1106
patient|1106,1113
received|1114,1122
perioperative|1123,1136
antibiotic|1137,1147
prophylaxis|1148,1159
.|1159,1160
The|1161,1164
<EOL>|1165,1166
patient|1166,1173
was|1174,1177
transferred|1178,1189
to|1190,1192
the|1193,1196
floor|1197,1202
from|1203,1207
the|1208,1211
PACU|1212,1216
in|1217,1219
stable|1220,1226
<EOL>|1227,1228
condition|1228,1237
.|1237,1238
On|1240,1242
POD0|1243,1247
,|1247,1248
pain|1249,1253
was|1254,1257
well|1258,1262
controlled|1263,1273
on|1274,1276
PCA|1277,1280
,|1280,1281
hydrated|1282,1290
<EOL>|1291,1292
for|1292,1295
urine|1296,1301
output|1302,1308
>|1309,1310
30cc|1310,1314
/|1314,1315
hour|1315,1319
,|1319,1320
provided|1321,1329
with|1330,1334
pneumoboots|1335,1346
and|1347,1350
<EOL>|1351,1352
incentive|1352,1361
spirometry|1362,1372
for|1373,1376
prophylaxis|1377,1388
,|1388,1389
and|1390,1393
ambulated|1394,1403
once|1404,1408
.|1408,1409
On|1410,1412
<EOL>|1413,1414
POD1|1414,1418
,|1418,1419
foley|1419,1424
was|1425,1428
removed|1429,1436
without|1437,1444
difficulty|1445,1455
,|1455,1456
basic|1457,1462
metabolic|1463,1472
panel|1473,1478
<EOL>|1479,1480
and|1480,1483
complete|1484,1492
blood|1493,1498
count|1499,1504
were|1505,1509
checked|1510,1517
,|1517,1518
pain|1519,1523
control|1524,1531
was|1532,1535
<EOL>|1536,1537
transitioned|1537,1549
from|1550,1554
PCA|1555,1558
to|1559,1561
oral|1562,1566
analgesics|1567,1577
,|1577,1578
diet|1579,1583
was|1584,1587
advanced|1588,1596
to|1597,1599
a|1600,1601
<EOL>|1602,1603
clears|1603,1609
/|1609,1610
toast|1610,1615
and|1616,1619
crackers|1620,1628
diet|1629,1633
.|1633,1634
On|1635,1637
POD2|1638,1642
,|1642,1643
diet|1644,1648
was|1649,1652
advanced|1653,1661
as|1662,1664
<EOL>|1665,1666
tolerated|1666,1675
.|1675,1676
The|1677,1680
remainder|1681,1690
of|1691,1693
the|1694,1697
hospital|1698,1706
course|1707,1713
was|1714,1717
relatively|1718,1728
<EOL>|1729,1730
unremarkable|1730,1742
.|1742,1743
The|1744,1747
patient|1748,1755
was|1756,1759
discharged|1760,1770
in|1771,1773
stable|1774,1780
condition|1781,1790
,|1790,1791
<EOL>|1792,1793
eating|1793,1799
well|1800,1804
,|1804,1805
ambulating|1806,1816
independently|1817,1830
,|1830,1831
voiding|1832,1839
without|1840,1847
<EOL>|1848,1849
difficulty|1849,1859
,|1859,1860
and|1861,1864
with|1865,1869
pain|1870,1874
control|1875,1882
on|1883,1885
oral|1886,1890
analgesics|1891,1901
.|1901,1902
On|1903,1905
exam|1906,1910
,|1910,1911
<EOL>|1912,1913
incision|1913,1921
was|1922,1925
clean|1926,1931
,|1931,1932
dry|1933,1936
,|1936,1937
and|1938,1941
intact|1942,1948
,|1948,1949
with|1950,1954
no|1955,1957
evidence|1958,1966
of|1967,1969
<EOL>|1970,1971
hematoma|1971,1979
collection|1980,1990
or|1991,1993
infection|1994,2003
.|2003,2004
The|2005,2008
patient|2009,2016
was|2017,2020
given|2021,2026
explicit|2027,2035
<EOL>|2036,2037
instructions|2037,2049
to|2050,2052
follow|2053,2059
-|2059,2060
up|2060,2062
in|2063,2065
clinic|2066,2072
with|2073,2077
_|2078,2079
_|2079,2080
_|2080,2081
in|2082,2084
3|2085,2086
weeks|2087,2092
.|2092,2093
<EOL>|2093,2094
<EOL>|2094,2095
<EOL>|2096,2097
Medications|2097,2108
on|2109,2111
Admission|2112,2121
:|2121,2122
<EOL>|2122,2123
none|2123,2127
<EOL>|2127,2128
<EOL>|2129,2130
Discharge|2130,2139
Medications|2140,2151
:|2151,2152
<EOL>|2152,2153
1.|2153,2155
Hydrocodone|2156,2167
-|2167,2168
Acetaminophen|2168,2181
_|2182,2183
_|2183,2184
_|2184,2185
mg|2186,2188
Tablet|2189,2195
Sig|2196,2199
:|2199,2200
_|2201,2202
_|2202,2203
_|2203,2204
Tablets|2205,2212
PO|2213,2215
<EOL>|2216,2217
Q6H|2217,2220
(|2221,2222
every|2222,2227
6|2228,2229
hours|2230,2235
)|2235,2236
as|2237,2239
needed|2240,2246
for|2247,2250
break|2251,2256
through|2257,2264
pain|2265,2269
only|2270,2274
(|2275,2276
score|2276,2281
<EOL>|2282,2283
>|2283,2284
4|2284,2285
)|2285,2286
.|2287,2288
<EOL>|2288,2289
Disp|2289,2293
:|2293,2294
*|2294,2295
60|2295,2297
Tablet|2298,2304
(|2304,2305
s|2305,2306
)|2306,2307
*|2307,2308
Refills|2309,2316
:|2316,2317
*|2317,2318
0|2318,2319
*|2319,2320
<EOL>|2320,2321
2.|2321,2323
Docusate|2324,2332
Sodium|2333,2339
100|2340,2343
mg|2344,2346
Capsule|2347,2354
Sig|2355,2358
:|2358,2359
One|2360,2363
(|2364,2365
1|2365,2366
)|2366,2367
Capsule|2368,2375
PO|2376,2378
BID|2379,2382
(|2383,2384
2|2384,2385
<EOL>|2386,2387
times|2387,2392
a|2393,2394
day|2395,2398
)|2398,2399
.|2399,2400
<EOL>|2400,2401
Disp|2401,2405
:|2405,2406
*|2406,2407
60|2407,2409
Capsule|2410,2417
(|2417,2418
s|2418,2419
)|2419,2420
*|2420,2421
Refills|2422,2429
:|2429,2430
*|2430,2431
2|2431,2432
*|2432,2433
<EOL>|2433,2434
<EOL>|2434,2435
<EOL>|2436,2437
Discharge|2437,2446
Disposition|2447,2458
:|2458,2459
<EOL>|2459,2460
Home|2460,2464
<EOL>|2464,2465
<EOL>|2466,2467
Discharge|2467,2476
Diagnosis|2477,2486
:|2486,2487
<EOL>|2487,2488
renal|2488,2493
cell|2494,2498
carcinoma|2499,2508
<EOL>|2508,2509
<EOL>|2509,2510
<EOL>|2511,2512
stable|2533,2539
<EOL>|2539,2540
<EOL>|2540,2541
<EOL>|2542,2543
-|2567,2568
You|2568,2571
may|2572,2575
shower|2576,2582
but|2583,2586
do|2587,2589
not|2590,2593
bathe|2594,2599
,|2599,2600
swim|2601,2605
or|2606,2608
immerse|2609,2616
your|2617,2621
incision|2622,2630
.|2630,2631
<EOL>|2631,2632
<EOL>|2632,2633
-|2633,2634
Do|2634,2636
not|2637,2640
eat|2641,2644
constipating|2645,2657
foods|2658,2663
for|2664,2667
_|2668,2669
_|2669,2670
_|2670,2671
weeks|2672,2677
,|2677,2678
drink|2679,2684
plenty|2685,2691
of|2692,2694
<EOL>|2695,2696
fluids|2696,2702
<EOL>|2702,2703
<EOL>|2703,2704
-|2704,2705
Do|2705,2707
not|2708,2711
lift|2712,2716
anything|2717,2725
heavier|2726,2733
than|2734,2738
a|2739,2740
phone|2741,2746
book|2747,2751
(|2752,2753
10|2753,2755
pounds|2756,2762
)|2762,2763
or|2764,2766
<EOL>|2767,2768
drive|2768,2773
until|2774,2779
you|2780,2783
are|2784,2787
seen|2788,2792
by|2793,2795
your|2796,2800
Urologist|2801,2810
in|2811,2813
follow|2814,2820
-|2820,2821
up|2821,2823
<EOL>|2823,2824
<EOL>|2824,2825
-|2825,2826
Tylenol|2826,2833
should|2834,2840
be|2841,2843
used|2844,2848
as|2849,2851
your|2852,2856
first|2857,2862
line|2863,2867
pain|2868,2872
medication|2873,2883
.|2883,2884
If|2885,2887
<EOL>|2888,2889
your|2889,2893
pain|2894,2898
is|2899,2901
not|2902,2905
well|2906,2910
controlled|2911,2921
on|2922,2924
Tylenol|2925,2932
you|2933,2936
have|2937,2941
been|2942,2946
<EOL>|2947,2948
prescribed|2948,2958
a|2959,2960
narcotic|2961,2969
pain|2970,2974
medication|2975,2985
.|2985,2986
Use|2987,2990
in|2991,2993
place|2994,2999
of|3000,3002
Tylenol|3003,3010
.|3010,3011
<EOL>|3012,3013
Do|3013,3015
not|3016,3019
exceed|3020,3026
4|3027,3028
gms|3029,3032
of|3033,3035
Tylenol|3036,3043
in|3044,3046
total|3047,3052
daily|3053,3058
<EOL>|3058,3059
<EOL>|3059,3060
-|3060,3061
Do|3061,3063
not|3064,3067
drive|3068,3073
or|3074,3076
drink|3077,3082
alcohol|3083,3090
while|3091,3096
taking|3097,3103
narcotics|3104,3113
<EOL>|3113,3114
<EOL>|3114,3115
-|3115,3116
Resume|3116,3122
all|3123,3126
of|3127,3129
your|3130,3134
home|3135,3139
medications|3140,3151
,|3151,3152
except|3153,3159
hold|3160,3164
NSAID|3165,3170
<EOL>|3171,3172
(|3172,3173
aspirin|3173,3180
,|3180,3181
advil|3182,3187
,|3187,3188
motrin|3189,3195
,|3195,3196
ibuprofen|3197,3206
)|3206,3207
until|3208,3213
you|3214,3217
see|3218,3221
your|3222,3226
urologist|3227,3236
<EOL>|3237,3238
in|3238,3240
follow|3241,3247
-|3247,3248
up|3248,3250
<EOL>|3250,3251
<EOL>|3251,3252
-|3252,3253
If|3253,3255
you|3256,3259
have|3260,3264
fevers|3265,3271
>|3272,3273
101.5|3274,3279
F|3280,3281
,|3281,3282
vomiting|3283,3291
,|3291,3292
or|3293,3295
increased|3296,3305
redness|3306,3313
,|3313,3314
<EOL>|3315,3316
swelling|3316,3324
,|3324,3325
or|3326,3328
discharge|3329,3338
from|3339,3343
your|3344,3348
incision|3349,3357
,|3357,3358
call|3359,3363
your|3364,3368
doctor|3369,3375
or|3376,3378
<EOL>|3379,3380
go|3380,3382
to|3383,3385
the|3386,3389
nearest|3390,3397
ER|3398,3400
<EOL>|3400,3401
<EOL>|3401,3402
-|3402,3403
Call|3403,3407
Dr.|3408,3411
_|3412,3413
_|3413,3414
_|3414,3415
to|3416,3418
set|3419,3422
up|3423,3425
follow|3426,3432
-|3432,3433
up|3433,3435
appointment|3436,3447
and|3448,3451
if|3452,3454
<EOL>|3455,3456
you|3456,3459
have|3460,3464
any|3465,3468
urological|3469,3479
questions|3480,3489
.|3489,3490
_|3491,3492
_|3492,3493
_|3493,3494
<EOL>|3494,3495
<EOL>|3495,3496
<EOL>|3497,3498
Followup|3498,3506
Instructions|3507,3519
:|3519,3520
<EOL>|3520,3521
_|3521,3522
_|3522,3523
_|3523,3524
<EOL>|3524,3525

