 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|33,37
No|38,40
:|40,41
_|44,45
_|45,46
_|46,47
<EOL>|47,48
<EOL>|49,50
Admission|50,59
Date|60,64
:|64,65
_|67,68
_|68,69
_|69,70
Discharge|84,93
Date|94,98
:|98,99
_|102,103
_|103,104
_|104,105
<EOL>|105,106
<EOL>|107,108
Date|108,112
of|113,115
Birth|116,121
:|121,122
_|124,125
_|125,126
_|126,127
Sex|140,143
:|143,144
F|147,148
<EOL>|148,149
<EOL>|150,151
Service|151,158
:|158,159
MEDICINE|160,168
<EOL>|168,169
<EOL>|170,171
Allergies|171,180
:|180,181
<EOL>|182,183
No|183,185
Known|186,191
Allergies|192,201
/|202,203
Adverse|204,211
Drug|212,216
Reactions|217,226
<EOL>|226,227
<EOL>|228,229
Attending|229,238
:|238,239
_|240,241
_|241,242
_|242,243
<EOL>|243,244
<EOL>|245,246
Chief|246,251
Complaint|252,261
:|261,262
<EOL>|262,263
Worsening|263,272
ABD|273,276
distension|277,287
and|288,291
pain|292,296
<EOL>|297,298
<EOL>|299,300
Major|300,305
Surgical|306,314
or|315,317
Invasive|318,326
Procedure|327,336
:|336,337
<EOL>|337,338
Paracentesis|338,350
<EOL>|350,351
<EOL>|351,352
<EOL>|353,354
History|354,361
of|362,364
Present|365,372
Illness|373,380
:|380,381
<EOL>|381,382
_|382,383
_|383,384
_|384,385
HCV|386,389
cirrhosis|390,399
c|400,401
/|401,402
b|402,403
ascites|404,411
,|411,412
hiv|413,416
on|417,419
ART|420,423
,|423,424
h|425,426
/|426,427
o|427,428
IVDU|429,433
,|433,434
COPD|435,439
,|439,440
<EOL>|441,442
bioplar|442,449
,|449,450
PTSD|451,455
,|455,456
presented|457,466
from|467,471
OSH|472,475
ED|476,478
with|479,483
worsening|484,493
abd|494,497
<EOL>|498,499
distension|499,509
over|510,514
past|515,519
week|520,524
.|524,525
<EOL>|527,528
Pt|528,530
reports|531,538
self|539,543
-|543,544
discontinuing|544,557
lasix|558,563
and|564,567
spirnolactone|568,581
_|582,583
_|583,584
_|584,585
weeks|586,591
<EOL>|592,593
ago|593,596
,|596,597
because|598,605
she|606,609
feels|610,615
like|616,620
"|621,622
they|622,626
do|627,629
n't|629,632
do|633,635
anything|636,644
"|644,645
and|646,649
that|650,654
<EOL>|655,656
she|656,659
"|660,661
does|661,665
n't|665,668
want|669,673
to|674,676
put|677,680
more|681,685
chemicals|686,695
in|696,698
her|699,702
.|702,703
"|703,704
She|705,708
does|709,713
not|714,717
<EOL>|718,719
follow|719,725
Na|726,728
-|728,729
restricted|729,739
diets|740,745
.|745,746
In|747,749
the|750,753
past|754,758
week|759,763
,|763,764
she|765,768
notes|769,774
that|775,779
she|780,783
<EOL>|784,785
has|785,788
been|789,793
having|794,800
worsening|801,810
abd|811,814
distension|815,825
and|826,829
discomfort|830,840
.|840,841
She|842,845
<EOL>|846,847
denies|847,853
_|854,855
_|855,856
_|856,857
edema|858,863
,|863,864
or|865,867
SOB|868,871
,|871,872
or|873,875
orthopnea|876,885
.|885,886
She|887,890
denies|891,897
f|898,899
/|899,900
c|900,901
/|901,902
n|902,903
/|903,904
v|904,905
,|905,906
d|907,908
/|908,909
c|909,910
,|910,911
<EOL>|912,913
dysuria|913,920
.|920,921
She|922,925
had|926,929
food|930,934
poisoning|935,944
a|945,946
week|947,951
ago|952,955
from|956,960
eating|961,967
stale|968,973
<EOL>|974,975
cake|975,979
(|980,981
n|981,982
/|982,983
v|983,984
20|985,987
min|988,991
after|992,997
food|998,1002
ingestion|1003,1012
)|1012,1013
,|1013,1014
which|1015,1020
resolved|1021,1029
the|1030,1033
same|1034,1038
<EOL>|1039,1040
day|1040,1043
.|1043,1044
She|1045,1048
denies|1049,1055
other|1056,1061
recent|1062,1068
illness|1069,1076
or|1077,1079
sick|1080,1084
contacts|1085,1093
.|1093,1094
She|1095,1098
notes|1099,1104
<EOL>|1105,1106
that|1106,1110
she|1111,1114
has|1115,1118
been|1119,1123
noticing|1124,1132
gum|1133,1136
bleeding|1137,1145
while|1146,1151
brushing|1152,1160
her|1161,1164
teeth|1165,1170
<EOL>|1171,1172
in|1172,1174
recent|1175,1181
weeks|1182,1187
.|1187,1188
she|1189,1192
denies|1193,1199
easy|1200,1204
bruising|1205,1213
,|1213,1214
melena|1215,1221
,|1221,1222
BRBPR|1223,1228
,|1228,1229
<EOL>|1230,1231
hemetesis|1231,1240
,|1240,1241
hemoptysis|1242,1252
,|1252,1253
or|1254,1256
hematuria|1257,1266
.|1266,1267
<EOL>|1269,1270
Because|1270,1277
of|1278,1280
her|1281,1284
abd|1285,1288
pain|1289,1293
,|1293,1294
she|1295,1298
went|1299,1303
to|1304,1306
OSH|1307,1310
ED|1311,1313
and|1314,1317
was|1318,1321
transferred|1322,1333
<EOL>|1334,1335
to|1335,1337
_|1338,1339
_|1339,1340
_|1340,1341
for|1342,1345
further|1346,1353
care|1354,1358
.|1358,1359
Per|1360,1363
ED|1364,1366
report|1367,1373
,|1373,1374
pt|1375,1377
has|1378,1381
brief|1382,1387
period|1388,1394
of|1395,1397
<EOL>|1398,1399
confusion|1399,1408
-|1409,1410
she|1411,1414
did|1415,1418
not|1419,1422
recall|1423,1429
the|1430,1433
ultrasound|1434,1444
or|1445,1447
bloodwork|1448,1457
at|1458,1460
<EOL>|1461,1462
osh|1462,1465
.|1465,1466
She|1467,1470
denies|1471,1477
recent|1478,1484
drug|1485,1489
use|1490,1493
or|1494,1496
alcohol|1497,1504
use.|1505,1509
She|1510,1513
denies|1514,1520
<EOL>|1521,1522
feeling|1522,1529
confused|1530,1538
,|1538,1539
but|1540,1543
reports|1544,1551
that|1552,1556
she|1557,1560
is|1561,1563
forgetful|1564,1573
at|1574,1576
times|1577,1582
.|1582,1583
<EOL>|1585,1586
In|1586,1588
the|1589,1592
ED|1593,1595
,|1595,1596
initial|1597,1604
vitals|1605,1611
were|1612,1616
98.4|1617,1621
70|1622,1624
106|1625,1628
/|1628,1629
63|1629,1631
16|1632,1634
97|1635,1637
%|1637,1638
RA|1638,1640
<EOL>|1642,1643
Labs|1643,1647
notable|1648,1655
for|1656,1659
ALT|1660,1663
/|1663,1664
AST|1664,1667
/|1667,1668
AP|1668,1670
_|1671,1672
_|1672,1673
_|1673,1674
_|1675,1676
_|1676,1677
_|1677,1678
:|1678,1679
_|1680,1681
_|1681,1682
_|1682,1683
,|1683,1684
<EOL>|1685,1686
Tbili1|1686,1692
.|1692,1693
6|1693,1694
,|1694,1695
WBC|1696,1699
5K|1700,1702
,|1702,1703
platelet|1704,1712
77|1713,1715
,|1715,1716
INR|1717,1720
1.6|1721,1724
<EOL>|1726,1727
<EOL>|1727,1728
<EOL>|1729,1730
Past|1730,1734
Medical|1735,1742
History|1743,1750
:|1750,1751
<EOL>|1751,1752
1.|1752,1754
HCV|1755,1758
Cirrhosis|1759,1768
<EOL>|1770,1771
2.|1771,1773
No|1774,1776
history|1777,1784
of|1785,1787
abnormal|1788,1796
Pap|1797,1800
smears|1801,1807
.|1807,1808
<EOL>|1810,1811
3.|1811,1813
She|1814,1817
had|1818,1821
calcification|1822,1835
in|1836,1838
her|1839,1842
breast|1843,1849
,|1849,1850
which|1851,1856
was|1857,1860
removed|1861,1868
<EOL>|1870,1871
previously|1871,1881
and|1882,1885
per|1886,1889
patient|1890,1897
not|1898,1901
,|1901,1902
it|1903,1905
was|1906,1909
benign|1910,1916
.|1916,1917
<EOL>|1919,1920
4|1920,1921
.|1921,1922
For|1923,1926
HIV|1927,1930
disease|1931,1938
,|1938,1939
she|1940,1943
is|1944,1946
being|1947,1952
followed|1953,1961
by|1962,1964
Dr.|1965,1968
_|1969,1970
_|1970,1971
_|1971,1972
Dr|1973,1975
.|1975,1976
<EOL>|1978,1979
_|1979,1980
_|1980,1981
_|1981,1982
.|1982,1983
<EOL>|1985,1986
5.|1986,1988
COPD|1989,1993
<EOL>|1995,1996
6.|1996,1998
Past|1999,2003
history|2004,2011
of|2012,2014
smoking|2015,2022
.|2022,2023
<EOL>|2025,2026
7.|2026,2028
She|2029,2032
also|2033,2037
had|2038,2041
a|2042,2043
skin|2044,2048
lesion|2049,2055
,|2055,2056
which|2057,2062
was|2063,2066
biopsied|2067,2075
and|2076,2079
showed|2080,2086
<EOL>|2088,2089
skin|2089,2093
cancer|2094,2100
per|2101,2104
patient|2105,2112
report|2113,2119
and|2120,2123
is|2124,2126
scheduled|2127,2136
for|2137,2140
a|2141,2142
complete|2143,2151
<EOL>|2153,2154
removal|2154,2161
of|2162,2164
the|2165,2168
skin|2169,2173
lesion|2174,2180
in|2181,2183
_|2184,2185
_|2185,2186
_|2186,2187
of|2188,2190
this|2191,2195
year|2196,2200
.|2200,2201
<EOL>|2203,2204
8.|2204,2206
She|2207,2210
also|2211,2215
had|2216,2219
another|2220,2227
lesion|2228,2234
in|2235,2237
her|2238,2241
forehead|2242,2250
with|2251,2255
purple|2256,2262
<EOL>|2264,2265
discoloration|2265,2278
.|2278,2279
It|2280,2282
was|2283,2286
biopsied|2287,2295
to|2296,2298
exclude|2299,2306
the|2307,2310
possibility|2311,2322
of|2323,2325
<EOL>|2327,2328
_|2328,2329
_|2329,2330
_|2330,2331
'|2331,2332
s|2332,2333
sarcoma|2334,2341
,|2341,2342
the|2343,2346
results|2347,2354
is|2355,2357
pending|2358,2365
.|2365,2366
<EOL>|2368,2369
9|2369,2370
.|2370,2371
A|2372,2373
15|2374,2376
mm|2377,2379
hypoechoic|2380,2390
lesion|2391,2397
on|2398,2400
her|2401,2404
ultrasound|2405,2415
on|2416,2418
_|2419,2420
_|2420,2421
_|2421,2422
<EOL>|2424,2425
and|2425,2428
is|2429,2431
being|2432,2437
monitored|2438,2447
by|2448,2450
an|2451,2453
MRI|2454,2457
.|2457,2458
<EOL>|2460,2461
10|2461,2463
.|2463,2464
History|2465,2472
of|2473,2475
dysplasia|2476,2485
of|2486,2488
anus|2489,2493
in|2494,2496
_|2497,2498
_|2498,2499
_|2499,2500
.|2500,2501
<EOL>|2503,2504
11|2504,2506
.|2506,2507
Bipolar|2508,2515
affective|2516,2525
disorder|2526,2534
,|2534,2535
currently|2536,2545
manic|2546,2551
,|2551,2552
mild|2553,2557
,|2557,2558
and|2559,2562
PTSD|2563,2567
.|2567,2568
<EOL>|2569,2570
<EOL>|2571,2572
12.|2572,2575
History|2576,2583
of|2584,2586
cocaine|2587,2594
and|2595,2598
heroin|2599,2605
use|2606,2609
.|2609,2610
<EOL>|2612,2613
<EOL>|2613,2614
<EOL>|2615,2616
Social|2616,2622
History|2623,2630
:|2630,2631
<EOL>|2631,2632
_|2632,2633
_|2633,2634
_|2634,2635
<EOL>|2635,2636
Family|2636,2642
History|2643,2650
:|2650,2651
<EOL>|2651,2652
She|2652,2655
a|2656,2657
total|2658,2663
of|2664,2666
five|2667,2671
siblings|2672,2680
,|2680,2681
but|2682,2685
she|2686,2689
is|2690,2692
not|2693,2696
<EOL>|2698,2699
talking|2699,2706
to|2707,2709
most|2710,2714
of|2715,2717
them|2718,2722
.|2722,2723
She|2724,2727
only|2728,2732
has|2733,2736
one|2737,2740
brother|2741,2748
that|2749,2753
she|2754,2757
is|2758,2760
in|2761,2763
<EOL>|2764,2765
<EOL>|2766,2767
touch|2767,2772
with|2773,2777
and|2778,2781
lives|2782,2787
in|2788,2790
_|2791,2792
_|2792,2793
_|2793,2794
.|2794,2795
She|2796,2799
is|2800,2802
not|2803,2806
aware|2807,2812
of|2813,2815
any|2816,2819
<EOL>|2821,2822
known|2822,2827
GI|2828,2830
or|2831,2833
liver|2834,2839
disease|2840,2847
in|2848,2850
her|2851,2854
family|2855,2861
.|2861,2862
<EOL>|2864,2865
Her|2865,2868
last|2869,2873
alcohol|2874,2881
consumption|2882,2893
was|2894,2897
one|2898,2901
drink|2902,2907
two|2908,2911
months|2912,2918
ago|2919,2922
.|2922,2923
No|2924,2926
<EOL>|2928,2929
regular|2929,2936
alcohol|2937,2944
consumption|2945,2956
.|2956,2957
Last|2958,2962
drug|2963,2967
use|2968,2971
_|2972,2973
_|2973,2974
_|2974,2975
years|2976,2981
ago|2982,2985
.|2985,2986
She|2987,2990
<EOL>|2992,2993
quit|2993,2997
smoking|2998,3005
a|3006,3007
couple|3008,3014
of|3015,3017
years|3018,3023
ago|3024,3027
.|3027,3028
<EOL>|3030,3031
<EOL>|3031,3032
<EOL>|3033,3034
Physical|3034,3042
Exam|3043,3047
:|3047,3048
<EOL>|3048,3049
VS|3049,3051
:|3051,3052
98.1|3053,3057
107|3058,3061
/|3061,3062
61|3062,3064
78|3065,3067
18|3068,3070
97RA|3071,3075
<EOL>|3077,3078
General|3078,3085
:|3085,3086
in|3087,3089
NAD|3090,3093
<EOL>|3095,3096
HEENT|3096,3101
:|3101,3102
CTAB|3103,3107
,|3107,3108
anicteric|3109,3118
sclera|3119,3125
,|3125,3126
OP|3127,3129
clear|3130,3135
<EOL>|3137,3138
Neck|3138,3142
:|3142,3143
supple|3144,3150
,|3150,3151
no|3152,3154
LAD|3155,3158
<EOL>|3160,3161
CV|3161,3163
:|3163,3164
RRR|3165,3168
,|3168,3169
S1S2|3169,3173
,|3173,3174
no|3175,3177
m|3178,3179
/|3179,3180
r|3180,3181
/|3181,3182
g|3182,3183
<EOL>|3185,3186
Lungs|3186,3191
:|3191,3192
CTAb|3193,3197
,|3197,3198
prolonged|3199,3208
expiratory|3209,3219
phase|3220,3225
,|3225,3226
no|3227,3229
w|3230,3231
/|3231,3232
r|3232,3233
/|3233,3234
r|3234,3235
<EOL>|3237,3238
Abdomen|3238,3245
:|3245,3246
distended|3247,3256
,|3256,3257
mild|3258,3262
diffuse|3263,3270
tenderness|3271,3281
,|3281,3282
+|3283,3284
flank|3284,3289
dullness|3290,3298
,|3298,3299
<EOL>|3300,3301
can|3301,3304
not|3304,3307
percuss|3308,3315
liver|3316,3321
/|3321,3322
spleen|3322,3328
edge|3329,3333
_|3334,3335
_|3335,3336
_|3336,3337
distension|3338,3348
<EOL>|3350,3351
GU|3351,3353
:|3353,3354
no|3355,3357
foley|3358,3363
<EOL>|3365,3366
Ext|3366,3369
:|3369,3370
wwp|3371,3374
,|3374,3375
no|3376,3378
c|3379,3380
/|3380,3381
e|3381,3382
/|3382,3383
e|3383,3384
,|3384,3385
+|3386,3387
clubbing|3388,3396
<EOL>|3398,3399
Neuro|3399,3404
:|3404,3405
AAO3|3406,3410
,|3410,3411
converse|3412,3420
normally|3421,3429
,|3429,3430
able|3431,3435
to|3436,3438
recall|3439,3445
3|3446,3447
times|3448,3453
after|3454,3459
5|3460,3461
<EOL>|3462,3463
minutes|3463,3470
,|3470,3471
CN|3472,3474
II|3475,3477
-|3477,3478
XII|3478,3481
intact|3482,3488
<EOL>|3490,3491
<EOL>|3491,3492
Discharge|3492,3501
:|3501,3502
<EOL>|3502,3503
<EOL>|3503,3504
PHYSICAL|3504,3512
EXAMINATION|3513,3524
:|3524,3525
<EOL>|3527,3528
VS|3528,3530
:|3530,3531
98|3532,3534
105|3535,3538
/|3538,3539
70|3539,3541
95|3542,3544
<EOL>|3544,3545
General|3545,3552
:|3552,3553
in|3554,3556
NAD|3557,3560
<EOL>|3562,3563
HEENT|3563,3568
:|3568,3569
anicteric|3570,3579
sclera|3580,3586
,|3586,3587
OP|3588,3590
clear|3591,3596
<EOL>|3598,3599
Neck|3599,3603
:|3603,3604
supple|3605,3611
,|3611,3612
no|3613,3615
LAD|3616,3619
<EOL>|3621,3622
CV|3622,3624
:|3624,3625
RRR|3626,3629
,|3629,3630
S1S2|3630,3634
,|3634,3635
no|3636,3638
m|3639,3640
/|3640,3641
r|3641,3642
/|3642,3643
g|3643,3644
<EOL>|3646,3647
Lungs|3647,3652
:|3652,3653
CTAb|3654,3658
,|3658,3659
prolonged|3660,3669
expiratory|3670,3680
phase|3681,3686
,|3686,3687
no|3688,3690
w|3691,3692
/|3692,3693
r|3693,3694
/|3694,3695
r|3695,3696
<EOL>|3698,3699
Abdomen|3699,3706
:|3706,3707
distended|3708,3717
but|3718,3721
improved|3722,3730
,|3730,3731
TTP|3732,3735
in|3736,3738
RUQ|3739,3742
,|3742,3743
<EOL>|3744,3745
GU|3745,3747
:|3747,3748
no|3749,3751
foley|3752,3757
<EOL>|3759,3760
Ext|3760,3763
:|3763,3764
wwp|3765,3768
,|3768,3769
no|3770,3772
c|3773,3774
/|3774,3775
e|3775,3776
/|3776,3777
e|3777,3778
,|3778,3779
+|3780,3781
clubbing|3782,3790
<EOL>|3792,3793
Neuro|3793,3798
:|3798,3799
AAO3|3800,3804
,|3804,3805
CN|3807,3809
II|3810,3812
-|3812,3813
XII|3813,3816
intact|3817,3823
<EOL>|3825,3826
<EOL>|3826,3827
<EOL>|3828,3829
Pertinent|3829,3838
Results|3839,3846
:|3846,3847
<EOL>|3847,3848
_|3848,3849
_|3849,3850
_|3850,3851
10|3852,3854
:|3854,3855
25PM|3855,3859
GLUCOSE|3862,3869
-|3869,3870
109|3870,3873
*|3873,3874
UREA|3875,3879
N|3880,3881
-|3881,3882
25|3882,3884
*|3884,3885
CREAT|3886,3891
-|3891,3892
0|3892,3893
.|3893,3894
3|3894,3895
*|3895,3896
SODIUM|3897,3903
-|3903,3904
138|3904,3907
<EOL>|3908,3909
POTASSIUM|3909,3918
-|3918,3919
3.4|3919,3922
CHLORIDE|3923,3931
-|3931,3932
105|3932,3935
TOTAL|3936,3941
CO2|3942,3945
-|3945,3946
27|3946,3948
ANION|3949,3954
GAP|3955,3958
-|3958,3959
9|3959,3960
<EOL>|3960,3961
_|3961,3962
_|3962,3963
_|3963,3964
10|3965,3967
:|3967,3968
25PM|3968,3972
estGFR|3975,3981
-|3981,3982
Using|3982,3987
this|3988,3992
<EOL>|3992,3993
_|3993,3994
_|3994,3995
_|3995,3996
10|3997,3999
:|3999,4000
25PM|4000,4004
ALT|4007,4010
(|4010,4011
SGPT|4011,4015
)|4015,4016
-|4016,4017
100|4017,4020
*|4020,4021
AST|4022,4025
(|4025,4026
SGOT|4026,4030
)|4030,4031
-|4031,4032
114|4032,4035
*|4035,4036
ALK|4037,4040
PHOS|4041,4045
-|4045,4046
114|4046,4049
*|4049,4050
<EOL>|4051,4052
TOT|4052,4055
BILI|4056,4060
-|4060,4061
1|4061,4062
.|4062,4063
6|4063,4064
*|4064,4065
<EOL>|4065,4066
_|4066,4067
_|4067,4068
_|4068,4069
10|4070,4072
:|4072,4073
25PM|4073,4077
LIPASE|4080,4086
-|4086,4087
77|4087,4089
*|4089,4090
<EOL>|4090,4091
_|4091,4092
_|4092,4093
_|4093,4094
10|4095,4097
:|4097,4098
25PM|4098,4102
ALBUMIN|4105,4112
-|4112,4113
3|4113,4114
.|4114,4115
3|4115,4116
*|4116,4117
<EOL>|4117,4118
_|4118,4119
_|4119,4120
_|4120,4121
10|4122,4124
:|4124,4125
25PM|4125,4129
WBC|4132,4135
-|4135,4136
5|4136,4137
.|4137,4138
0|4138,4139
#|4139,4140
RBC|4141,4144
-|4144,4145
4.29|4145,4149
HGB|4150,4153
-|4153,4154
14.3|4154,4158
HCT|4159,4162
-|4162,4163
42.6|4163,4167
MCV|4168,4171
-|4171,4172
99|4172,4174
*|4174,4175
<EOL>|4176,4177
MCH|4177,4180
-|4180,4181
33|4181,4183
.|4183,4184
3|4184,4185
*|4185,4186
MCHC|4187,4191
-|4191,4192
33.5|4192,4196
RDW|4197,4200
-|4200,4201
15|4201,4203
.|4203,4204
7|4204,4205
*|4205,4206
<EOL>|4206,4207
_|4207,4208
_|4208,4209
_|4209,4210
10|4211,4213
:|4213,4214
25PM|4214,4218
NEUTS|4221,4226
-|4226,4227
70|4227,4229
.|4229,4230
3|4230,4231
*|4231,4232
LYMPHS|4233,4239
-|4239,4240
16|4240,4242
.|4242,4243
5|4243,4244
*|4244,4245
MONOS|4246,4251
-|4251,4252
8.1|4252,4255
EOS|4256,4259
-|4259,4260
4|4260,4261
.|4261,4262
2|4262,4263
*|4263,4264
<EOL>|4265,4266
BASOS|4266,4271
-|4271,4272
0.8|4272,4275
<EOL>|4275,4276
_|4276,4277
_|4277,4278
_|4278,4279
10|4280,4282
:|4282,4283
25PM|4283,4287
PLT|4290,4293
COUNT|4294,4299
-|4299,4300
71|4300,4302
*|4302,4303
<EOL>|4303,4304
_|4304,4305
_|4305,4306
_|4306,4307
10|4308,4310
:|4310,4311
25PM|4311,4315
_|4318,4319
_|4319,4320
_|4320,4321
PTT|4322,4325
-|4325,4326
30.9|4326,4330
_|4331,4332
_|4332,4333
_|4333,4334
<EOL>|4334,4335
_|4335,4336
_|4336,4337
_|4337,4338
10|4339,4341
:|4341,4342
25PM|4342,4346
_|4349,4350
_|4350,4351
_|4351,4352
<EOL>|4352,4353
.|4353,4354
<EOL>|4354,4355
<EOL>|4355,4356
CXR|4356,4359
:|4359,4360
No|4361,4363
acute|4364,4369
cardiopulmonary|4370,4385
process|4386,4393
.|4393,4394
<EOL>|4396,4397
U|4397,4398
/|4398,4399
S|4399,4400
:|4400,4401
<EOL>|4403,4404
1.|4404,4406
Nodular|4407,4414
appearance|4415,4425
of|4426,4428
the|4429,4432
liver|4433,4438
compatible|4439,4449
with|4450,4454
cirrhosis|4455,4464
.|4464,4465
<EOL>|4466,4467
Signs|4467,4472
of|4473,4475
portal|4476,4482
<EOL>|4484,4485
hypertension|4485,4497
including|4498,4507
small|4508,4513
amount|4514,4520
of|4521,4523
ascites|4524,4531
and|4532,4535
splenomegaly|4536,4548
.|4548,4549
<EOL>|4550,4551
<EOL>|4552,4553
2.|4553,4555
Cholelithiasis|4556,4570
.|4570,4571
<EOL>|4573,4574
3.|4574,4576
Patent|4577,4583
portal|4584,4590
veins|4591,4596
with|4597,4601
normal|4602,4608
hepatopetal|4609,4620
flow|4621,4625
.|4625,4626
<EOL>|4628,4629
Diagnostic|4629,4639
para|4640,4644
attempted|4645,4654
in|4655,4657
the|4658,4661
ED|4662,4664
,|4664,4665
unsuccessful|4666,4678
.|4678,4679
<EOL>|4681,4682
On|4682,4684
the|4685,4688
floor|4689,4694
,|4694,4695
pt|4696,4698
c|4699,4700
/|4700,4701
o|4701,4702
abd|4703,4706
distension|4707,4717
and|4718,4721
discomfort|4722,4732
.|4732,4733
<EOL>|4733,4734
<EOL>|4735,4736
Brief|4736,4741
Hospital|4742,4750
Course|4751,4757
:|4757,4758
<EOL>|4758,4759
_|4759,4760
_|4760,4761
_|4761,4762
HCV|4763,4766
cirrhosis|4767,4776
c|4777,4778
/|4778,4779
b|4779,4780
ascites|4781,4788
,|4788,4789
hiv|4790,4793
on|4794,4796
ART|4797,4800
,|4800,4801
h|4802,4803
/|4803,4804
o|4804,4805
IVDU|4806,4810
,|4810,4811
COPD|4812,4816
,|4816,4817
<EOL>|4818,4819
bioplar|4819,4826
,|4826,4827
PTSD|4828,4832
,|4832,4833
presented|4834,4843
from|4844,4848
OSH|4849,4852
ED|4853,4855
with|4856,4860
worsening|4861,4870
abd|4871,4874
<EOL>|4875,4876
distension|4876,4886
over|4887,4891
past|4892,4896
week|4897,4901
and|4902,4905
confusion|4906,4915
.|4915,4916
<EOL>|4918,4919
<EOL>|4919,4920
#|4920,4921
Ascites|4922,4929
-|4930,4931
p|4932,4933
/|4933,4934
w|4934,4935
worsening|4936,4945
abd|4946,4949
distension|4950,4960
and|4961,4964
discomfort|4965,4975
for|4976,4979
last|4980,4984
<EOL>|4985,4986
week|4986,4990
.|4990,4991
likely|4992,4998
_|4999,5000
_|5000,5001
_|5001,5002
portal|5003,5009
HTN|5010,5013
given|5014,5019
underlying|5020,5030
liver|5031,5036
disease|5037,5044
,|5044,5045
<EOL>|5046,5047
though|5047,5053
no|5054,5056
ascitic|5057,5064
fluid|5065,5070
available|5071,5080
on|5081,5083
night|5084,5089
of|5090,5092
admission|5093,5102
.|5102,5103
No|5104,5106
<EOL>|5107,5108
signs|5108,5113
of|5114,5116
heart|5117,5122
failure|5123,5130
noted|5131,5136
on|5137,5139
exam|5140,5144
.|5144,5145
This|5146,5150
was|5151,5154
_|5155,5156
_|5156,5157
_|5157,5158
to|5159,5161
med|5162,5165
<EOL>|5166,5167
non-compliance|5167,5181
and|5182,5185
lack|5186,5190
of|5191,5193
diet|5194,5198
restriction|5199,5210
.|5210,5211
SBP|5212,5215
negative|5216,5224
<EOL>|5224,5225
diuretics|5225,5234
:|5234,5235
<EOL>|5237,5238
>|5238,5239
Furosemide|5240,5250
40|5251,5253
mg|5254,5256
PO|5257,5259
DAILY|5260,5265
<EOL>|5267,5268
>|5268,5269
Spironolactone|5270,5284
50|5285,5287
mg|5288,5290
PO|5291,5293
DAILY|5294,5299
,|5299,5300
chosen|5301,5307
over|5308,5312
the|5313,5316
usual|5317,5322
100mg|5323,5328
<EOL>|5329,5330
dose|5330,5334
d|5335,5336
/|5336,5337
t|5337,5338
K|5339,5340
+|5340,5341
of|5342,5344
4.5|5345,5348
.|5348,5349
<EOL>|5352,5353
CXR|5354,5357
was|5358,5361
wnl|5362,5365
,|5365,5366
UA|5367,5369
negative|5370,5378
,|5378,5379
Urine|5380,5385
culture|5386,5393
blood|5394,5399
culture|5400,5407
negative|5408,5416
.|5416,5417
<EOL>|5418,5419
<EOL>|5420,5421
Pt|5421,5423
was|5424,5427
losing|5428,5434
excess|5435,5441
fluid|5442,5447
appropriately|5448,5461
with|5462,5466
stable|5467,5473
lytes|5474,5479
on|5480,5482
<EOL>|5483,5484
the|5484,5487
above|5488,5493
regimen|5494,5501
.|5501,5502
Pt|5503,5505
was|5506,5509
scheduled|5510,5519
with|5520,5524
current|5525,5532
PCP|5533,5536
for|5537,5540
<EOL>|5541,5542
_|5542,5543
_|5543,5544
_|5544,5545
check|5546,5551
upon|5552,5556
discharge|5557,5566
.|5566,5567
<EOL>|5570,5571
Pt|5571,5573
was|5574,5577
scheduled|5578,5587
for|5588,5591
new|5592,5595
PCP|5596,5599
with|5600,5604
Dr.|5605,5608
_|5609,5610
_|5610,5611
_|5611,5612
at|5613,5615
_|5616,5617
_|5617,5618
_|5618,5619
and|5620,5623
<EOL>|5624,5625
follow|5625,5631
up|5632,5634
in|5635,5637
Liver|5638,5643
clinic|5644,5650
to|5651,5653
schedule|5654,5662
outpatient|5663,5673
screening|5674,5683
EGD|5684,5687
<EOL>|5688,5689
and|5689,5692
_|5693,5694
_|5694,5695
_|5695,5696
.|5696,5697
<EOL>|5700,5701
<EOL>|5702,5703
<EOL>|5703,5704
<EOL>|5705,5706
Medications|5706,5717
on|5718,5720
Admission|5721,5730
:|5730,5731
<EOL>|5731,5732
The|5732,5735
Preadmission|5736,5748
Medication|5749,5759
list|5760,5764
is|5765,5767
accurate|5768,5776
and|5777,5780
complete|5781,5789
.|5789,5790
<EOL>|5790,5791
1.|5791,5793
Furosemide|5794,5804
20|5805,5807
mg|5808,5810
PO|5811,5813
DAILY|5814,5819
<EOL>|5820,5821
2.|5821,5823
Spironolactone|5824,5838
50|5839,5841
mg|5842,5844
PO|5845,5847
DAILY|5848,5853
<EOL>|5854,5855
3.|5855,5857
Albuterol|5858,5867
Inhaler|5868,5875
2|5876,5877
PUFF|5878,5882
IH|5883,5885
Q4H|5886,5889
:|5889,5890
PRN|5890,5893
wheezing|5894,5902
,|5902,5903
SOB|5904,5907
<EOL>|5908,5909
4.|5909,5911
Raltegravir|5912,5923
400|5924,5927
mg|5928,5930
PO|5931,5933
BID|5934,5937
<EOL>|5938,5939
5.|5939,5941
Emtricitabine|5942,5955
-|5955,5956
Tenofovir|5956,5965
(|5966,5967
Truvada|5967,5974
)|5974,5975
1|5976,5977
TAB|5978,5981
PO|5982,5984
DAILY|5985,5990
<EOL>|5991,5992
6.|5992,5994
Nicotine|5995,6003
Patch|6004,6009
14|6010,6012
mg|6013,6015
TD|6016,6018
DAILY|6019,6024
<EOL>|6025,6026
7.|6026,6028
Ipratropium|6029,6040
Bromide|6041,6048
Neb|6049,6052
1|6053,6054
NEB|6055,6058
IH|6059,6061
Q6H|6062,6065
SOB|6066,6069
<EOL>|6070,6071
<EOL>|6071,6072
<EOL>|6073,6074
Discharge|6074,6083
Medications|6084,6095
:|6095,6096
<EOL>|6096,6097
1.|6097,6099
Albuterol|6100,6109
Inhaler|6110,6117
2|6118,6119
PUFF|6120,6124
IH|6125,6127
Q4H|6128,6131
:|6131,6132
PRN|6132,6135
wheezing|6136,6144
,|6144,6145
SOB|6146,6149
<EOL>|6150,6151
2.|6151,6153
Emtricitabine|6154,6167
-|6167,6168
Tenofovir|6168,6177
(|6178,6179
Truvada|6179,6186
)|6186,6187
1|6188,6189
TAB|6190,6193
PO|6194,6196
DAILY|6197,6202
<EOL>|6203,6204
3.|6204,6206
Furosemide|6207,6217
40|6218,6220
mg|6221,6223
PO|6224,6226
DAILY|6227,6232
<EOL>|6233,6234
RX|6234,6236
*|6237,6238
furosemide|6238,6248
40|6249,6251
mg|6252,6254
1|6255,6256
tablet|6257,6263
(|6263,6264
s|6264,6265
)|6265,6266
by|6267,6269
mouth|6270,6275
Daily|6276,6281
Disp|6282,6286
#|6287,6288
*|6288,6289
30|6289,6291
Tablet|6292,6298
<EOL>|6299,6300
Refills|6300,6307
:|6307,6308
*|6308,6309
3|6309,6310
<EOL>|6310,6311
4.|6311,6313
Ipratropium|6314,6325
Bromide|6326,6333
Neb|6334,6337
1|6338,6339
NEB|6340,6343
IH|6344,6346
Q6H|6347,6350
SOB|6351,6354
<EOL>|6355,6356
5.|6356,6358
Nicotine|6359,6367
Patch|6368,6373
14|6374,6376
mg|6377,6379
TD|6380,6382
DAILY|6383,6388
<EOL>|6389,6390
6.|6390,6392
Raltegravir|6393,6404
400|6405,6408
mg|6409,6411
PO|6412,6414
BID|6415,6418
<EOL>|6419,6420
7.|6420,6422
Spironolactone|6423,6437
50|6438,6440
mg|6441,6443
PO|6444,6446
DAILY|6447,6452
<EOL>|6453,6454
8.|6454,6456
Acetaminophen|6457,6470
500|6471,6474
mg|6475,6477
PO|6478,6480
Q6H|6481,6484
:|6484,6485
PRN|6485,6488
pain|6489,6493
<EOL>|6494,6495
<EOL>|6495,6496
<EOL>|6497,6498
Discharge|6498,6507
Disposition|6508,6519
:|6519,6520
<EOL>|6520,6521
Home|6521,6525
<EOL>|6525,6526
<EOL>|6527,6528
Discharge|6528,6537
Diagnosis|6538,6547
:|6547,6548
<EOL>|6548,6549
Ascites|6549,6556
from|6557,6561
Portal|6562,6568
HTN|6569,6572
<EOL>|6572,6573
<EOL>|6573,6574
<EOL>|6575,6576
Discharge|6576,6585
Condition|6586,6595
:|6595,6596
<EOL>|6596,6597
Mental|6597,6603
Status|6604,6610
:|6610,6611
Clear|6612,6617
and|6618,6621
coherent|6622,6630
.|6630,6631
<EOL>|6631,6632
Level|6632,6637
of|6638,6640
Consciousness|6641,6654
:|6654,6655
Alert|6656,6661
and|6662,6665
interactive|6666,6677
.|6677,6678
<EOL>|6678,6679
Activity|6679,6687
Status|6688,6694
:|6694,6695
Ambulatory|6696,6706
-|6707,6708
Independent|6709,6720
.|6720,6721
<EOL>|6721,6722
<EOL>|6722,6723
<EOL>|6724,6725
Discharge|6725,6734
Instructions|6735,6747
:|6747,6748
<EOL>|6748,6749
Dear|6749,6753
Ms.|6754,6757
_|6758,6759
_|6759,6760
_|6760,6761
,|6761,6762
<EOL>|6762,6763
It|6763,6765
was|6766,6769
a|6770,6771
pleasure|6772,6780
taking|6781,6787
care|6788,6792
of|6793,6795
you|6796,6799
!|6799,6800
You|6801,6804
came|6805,6809
to|6810,6812
us|6813,6815
with|6816,6820
<EOL>|6821,6822
stomach|6822,6829
pain|6830,6834
and|6835,6838
worsening|6839,6848
distension|6849,6859
.|6859,6860
While|6861,6866
you|6867,6870
were|6871,6875
here|6876,6880
we|6881,6883
<EOL>|6884,6885
did|6885,6888
a|6889,6890
paracentesis|6891,6903
to|6904,6906
remove|6907,6913
1.5|6914,6917
L|6917,6918
of|6919,6921
fluid|6922,6927
from|6928,6932
your|6933,6937
belly|6938,6943
.|6943,6944
We|6945,6947
<EOL>|6948,6949
also|6949,6953
placed|6954,6960
you|6961,6964
on|6965,6967
you|6968,6971
40|6972,6974
mg|6975,6977
of|6978,6980
Lasix|6981,6986
and|6987,6990
50|6991,6993
mg|6994,6996
of|6997,6999
Aldactone|7000,7009
to|7010,7012
<EOL>|7013,7014
help|7014,7018
you|7019,7022
urinate|7023,7030
the|7031,7034
excess|7035,7041
fluid|7042,7047
still|7048,7053
in|7054,7056
your|7057,7061
belly|7062,7067
.|7067,7068
As|7069,7071
we|7072,7074
<EOL>|7075,7076
discussed|7076,7085
,|7085,7086
everyone|7087,7095
has|7096,7099
a|7100,7101
different|7102,7111
dose|7112,7116
of|7117,7119
lasix|7120,7125
required|7126,7134
to|7135,7137
<EOL>|7138,7139
make|7139,7143
them|7144,7148
urinate|7149,7156
and|7157,7160
it|7161,7163
's|7163,7165
likely|7166,7172
that|7173,7177
you|7178,7181
were|7182,7186
n't|7186,7189
taking|7190,7196
a|7197,7198
high|7199,7203
<EOL>|7204,7205
enough|7205,7211
dose|7212,7216
.|7216,7217
Please|7218,7224
take|7225,7229
these|7230,7235
medications|7236,7247
daily|7248,7253
to|7254,7256
keep|7257,7261
excess|7262,7268
<EOL>|7269,7270
fluid|7270,7275
off|7276,7279
and|7280,7283
eat|7284,7287
a|7288,7289
low|7290,7293
salt|7294,7298
diet|7299,7303
.|7303,7304
You|7305,7308
will|7309,7313
follow|7314,7320
up|7321,7323
with|7324,7328
Dr|7329,7331
.|7331,7332
<EOL>|7333,7334
_|7334,7335
_|7335,7336
_|7336,7337
in|7338,7340
liver|7341,7346
clinic|7347,7353
and|7354,7357
from|7358,7362
there|7363,7368
have|7369,7373
your|7374,7378
colonoscopy|7379,7390
<EOL>|7391,7392
and|7392,7395
EGD|7396,7399
scheduled|7400,7409
.|7409,7410
Of|7411,7413
course|7414,7420
,|7420,7421
we|7422,7424
are|7425,7428
always|7429,7435
here|7436,7440
if|7441,7443
you|7444,7447
need|7448,7452
us|7453,7455
.|7455,7456
<EOL>|7457,7458
We|7458,7460
wish|7461,7465
you|7466,7469
all|7470,7473
the|7474,7477
best|7478,7482
!|7482,7483
<EOL>|7483,7484
Your|7484,7488
_|7489,7490
_|7490,7491
_|7491,7492
Team|7493,7497
.|7497,7498
<EOL>|7500,7501
<EOL>|7502,7503
Followup|7503,7511
Instructions|7512,7524
:|7524,7525
<EOL>|7525,7526
_|7526,7527
_|7527,7528
_|7528,7529
<EOL>|7529,7530

