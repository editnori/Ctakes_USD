CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Neurosurgical Procedures|Procedure|false|false||NEUROSURGERYnull|Science of neurosurgery|Title|false|false||NEUROSURGERYnull|penicillins|Drug|false|false||Penicillins
null|penicillins|Drug|false|false||Penicillinsnull|Poisoning by, adverse effect of and underdosing of penicillins|Disorder|false|false||Penicillins
null|Poisoning by penicillin|Disorder|false|false||Penicillinsnull|Adverse reaction to penicillins|Finding|false|false||Penicillinsnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Wound Infection|Finding|false|false||Wound Infectionnull|Traumatic Wound|Disorder|false|false||Wound
null|Wounds and Injuries|Disorder|false|false||Wound
null|Traumatic injury|Disorder|false|false||Woundnull|Route of Administration - Wound|Finding|false|false||Wound
null|null|Finding|false|false||Wound
null|Specimen Type - Wound|Finding|false|false||Woundnull|Communicable Diseases|Disorder|false|false||Infectionnull|Infection|Finding|false|false||Infectionnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Table Cell Horizontal Align - right|Finding|false|false||Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|Craniotomy|Procedure|false|false||Craniotomynull|Evacuation procedure|Procedure|false|false||Evacuationnull|Abscess|Disorder|false|false||Abscessnull|null|Finding|false|false||Abscessnull|Woman|Subject|false|false||woman
null|Human, Female adult|Subject|false|false||womannull|PMH - past medical history|Finding|false|false||past medical history
null|Medical History|Finding|false|false||past medical historynull|Medical History|Finding|false|false||medical historynull|Medical referral type|Finding|false|false||medical
null|Medical|Finding|false|false||medical
null|Medical school type|Finding|false|false||medicalnull|Medical service|Procedure|false|false||medicalnull|Medical History|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|History of present illness (finding)|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Parietal|Modifier|false|false||parietalnull|Brain Abscess|Disorder|false|false|C4266577;C0006104|brain abscess
null|Cerebral abscess|Disorder|false|false|C4266577;C0006104|brain abscessnull|Brain Diseases|Disorder|false|false|C4266577;C0006104|brainnull|Head>Brain|Anatomy|false|false|C1546533;C0006111;C0006105;C1510428;C0000833|brain
null|Brain|Anatomy|false|false|C1546533;C0006111;C0006105;C1510428;C0000833|brainnull|Abscess|Disorder|false|false|C4266577;C0006104|abscessnull|null|Finding|false|false|C4266577;C0006104|abscessnull|One month|Time|false|false||one monthnull|Transaction counts and value totals - month|Finding|false|false||month
null|Precision - month|Finding|false|false||monthnull|month|Time|false|false||month
null|Monthly (qualifier value)|Time|false|false||monthnull|FBXW7 wt Allele|Finding|false|false||ago
null|FBXW7 gene|Finding|false|false||agonull|Left upper arm structure|Anatomy|false|false|C1824218;C3715044;C3495676;C1522541;C5400986;C4761640|left arm
null|Left arm|Anatomy|false|false|C1824218;C3715044;C3495676;C1522541;C5400986;C4761640|left armnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Anorectal Malformations|Disorder|false|false|C0230347;C5779993;C0446516;C1140618;C1269078|armnull|AKR1A1 wt Allele|Finding|false|false|C0230347;C5779993;C0446516;C1140618;C1269078|arm
null|ARMC9 gene|Finding|false|false|C0230347;C5779993;C0446516;C1140618;C1269078|armnull|Protocol Treatment Arm|Procedure|false|false|C0446516;C1140618;C1269078;C0230347;C5779993|arm
null|Axillary Reverse Mapping|Procedure|false|false|C0446516;C1140618;C1269078;C0230347;C5779993|arm
null|Study Arm|Procedure|false|false|C0446516;C1140618;C1269078;C0230347;C5779993|armnull|Upper arm|Anatomy|false|false|C1522541;C5400986;C4761640;C3495676;C1824218;C3715044|arm
null|null|Anatomy|false|false|C1522541;C5400986;C4761640;C3495676;C1824218;C3715044|arm
null|Upper Extremity|Anatomy|false|false|C1522541;C5400986;C4761640;C3495676;C1824218;C3715044|armnull|Numbness of face|Finding|false|false|C0015450;C4266571|face numbnessnull|FANCONI ANEMIA, COMPLEMENTATION GROUP E|Disorder|false|false|C0015450;C4266571|facenull|FANCE wt Allele|Finding|false|false|C0015450;C4266571|face
null|FANCE gene|Finding|false|false|C0015450;C4266571|face
null|ELOVL6 gene|Finding|false|false|C0015450;C4266571|facenull|Head>Face|Anatomy|false|false|C3160739;C0239511;C1423759;C2828055;C1414531;C0028643;C0020580|face
null|Face|Anatomy|false|false|C3160739;C0239511;C1423759;C2828055;C1414531;C0028643;C0020580|facenull|Face (spatial concept)|Modifier|false|false||facenull|Numbness|Finding|false|false|C0015450;C4266571|numbness
null|Hypesthesia|Finding|false|false|C0015450;C4266571|numbnessnull|Abscess|Disorder|false|false||abscessnull|null|Finding|false|false||abscessnull|Initially|Time|false|false||initiallynull|Widening|Modifier|false|false||broadnull|Spectrum|Finding|false|false||spectrumnull|Electromagnetic Spectrum|LabModifier|false|false||spectrumnull|Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE|Drug|false|false||antibiotics
null|Antibiotics|Drug|false|false||antibiotics
null|Antibiotics, ophthalmologic|Drug|false|false||antibiotics
null|Antibiotics, Gynecological|Drug|false|false||antibiotics
null|antibiotics, intestinal|Drug|false|false||antibiotics
null|Antibiotic throat preparations|Drug|false|false||antibiotics
null|Antibiotics, Antitubercular|Drug|false|false||antibiotics
null|Antibiotics for systemic use|Drug|false|false||antibiotics
null|Antifungal Antibiotics, Topical|Drug|false|false||antibioticsnull|Culture Dose Form|Drug|false|false||culturenull|Culture (Anthropological)|Finding|false|false||culture
null|Cultural aspects|Finding|false|false||culturenull|Microbial culture (procedure)|Procedure|false|false||culture
null|Laboratory culture|Procedure|false|false||culturenull|Data|Finding|false|false||datanull|Data call receiving device|Device|false|false||datanull|Data <Amphipyrinae>|Entity|false|false||datanull|Genus Fusobacterium|Entity|false|false||fusobacteriumnull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|ceftriaxone|Drug|false|false||Ceftriaxone
null|ceftriaxone|Drug|false|false||Ceftriaxonenull|Every twelve hours|Time|false|false||q12hnull|Flagyl|Drug|false|false||flagyl
null|Flagyl|Drug|false|false||flagylnull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|Peripherally inserted central catheter (physical object)|Device|false|false||PICC linenull|Peripherally Inserted Central Catheter Line Insertion|Procedure|false|false||PICCnull|Peripherally inserted central catheter (physical object)|Device|false|false||PICCnull|Line Specimen|Drug|false|false||line
null|Long Interspersed Elements|Drug|false|false||line
null|Long Interspersed Elements|Drug|false|false||linenull|line source specimen code|Finding|false|false||linenull|Intravascular line|Device|false|false||linenull|Linear|Modifier|false|false||linenull|Line Unit of Length|LabModifier|false|false||linenull|Clinic|Device|false|false||clinic
null|Ambulatory Care Facilities|Device|false|false||clinicnull|Clinic|Entity|false|false||clinic
null|Ambulatory Care Facilities|Entity|false|false||clinicnull|Patient location type - Clinic|Modifier|false|false||clinic
null|Person location type - Clinic|Modifier|false|false||clinicnull|Repeat Object|Finding|false|false||repeat
null|Repeat|Finding|false|false||repeatnull|Repeat Pattern|Time|false|false||repeatnull|CYREN gene|Finding|false|false||MRInull|Magnetic resonance imaging service|Procedure|false|false||MRI
null|Magnetic Resonance Imaging|Procedure|false|false||MRInull|Maori Language|Entity|false|false||MRInull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Persistent|Time|false|false||persistentnull|Ring Dosage Form|Drug|false|false||ringnull|Ring device|Device|false|false||ringnull|Annular shape|Modifier|false|false||ringnull|Ring Dosing Unit|LabModifier|false|false||ringnull|Congenital Abnormality|Disorder|false|false|C1515974|abnormalitynull|Abnormality|Finding|false|false|C1515974|abnormalitynull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Parietal|Modifier|false|false||parietalnull|Operative site|Modifier|false|false||surgical sitenull|Operative Surgical Procedures|Procedure|false|false|C1515974|surgical
null|Surgical service|Procedure|false|false|C1515974|surgicalnull|null|Finding|false|false|C1515974|sitenull|Anatomic Site|Anatomy|false|false|C1546778;C1704258;C0000768;C0543467;C0587668|sitenull|Study Site|Modifier|false|false||site
null|Site|Modifier|false|false||sitenull|Continuous|Finding|false|false||ongoingnull|Abscess|Disorder|false|false||abscessnull|null|Finding|false|false||abscessnull|Repeat Object|Finding|false|false||repeat
null|Repeat|Finding|false|false||repeatnull|Repeat Pattern|Time|false|false||repeatnull|Body Substance Discharge|Finding|false|false||drainage
null|Body Fluid Discharge|Finding|false|false||drainagenull|Drainage procedure|Procedure|false|false||drainagenull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|Communicable Diseases|Disorder|false|false||infectious diseasenull|Infectious Disease Medicine|Title|false|false||infectious diseasenull|Communicable Diseases|Disorder|false|false||infectiousnull|infectious - Entity Risk|Modifier|false|false||infectiousnull|Disease|Disorder|false|false||diseasenull|Address type - Office|Finding|false|false||officenull|Office|Device|false|false||officenull|Organization unit type - Office|Entity|false|false||officenull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|One day|Time|false|false||one daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Early|Time|false|false||earlynull|Antibiotics|Drug|false|false||antibioticnull|GDC Regimen Terminology|Finding|false|false||regimennull|Treatment Protocols|Procedure|false|false||regimennull|null|Time|false|false||prior tonull|null|Time|false|false||priornull|Body Substance Discharge|Finding|false|false||drainage
null|Body Fluid Discharge|Finding|false|false||drainagenull|Drainage procedure|Procedure|false|false||drainagenull|Past 30 days|Time|false|false||past monthnull|Transaction counts and value totals - month|Finding|false|false||month
null|Precision - month|Finding|false|false||monthnull|month|Time|false|false||month
null|Monthly (qualifier value)|Time|false|false||monthnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Upper Extremity Paresis|Finding|false|false|C1140618;C0015385|upper extremity weaknessnull|Upper Extremity|Anatomy|false|false|C0751409;C0028643;C0020580;C0587246;C3714552;C0004093|upper extremitynull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|Muscle weakness of limb|Finding|false|false|C0015385;C1140618|extremity weaknessnull|Limb structure|Anatomy|false|false|C0028643;C0020580;C0587246;C0751409;C3714552;C0004093|extremitynull|Weakness|Finding|false|false|C0015385;C1140618|weakness
null|Asthenia|Finding|false|false|C0015385;C1140618|weaknessnull|Numbness|Finding|false|false|C1140618;C0015385|numbness
null|Hypesthesia|Finding|false|false|C1140618;C0015385|numbnessnull|Overall Publication Type|Finding|false|false||overallnull|Overall|Modifier|false|false||overallnull|Slightly (qualifier value)|Modifier|false|false||slightly
null|Slight (qualifier value)|Modifier|false|false||slightlynull|Fever|Finding|false|false||feversnull|Chills|Finding|true|false||chillsnull|Headache|Finding|true|false||headachesnull|Changing|Finding|true|false||changesnull|Changed status|LabModifier|false|false||changesnull|Vision|Finding|false|false||visionnull|null|Attribute|false|false||visionnull|Specialized Stand Alone Plan - Vision|Entity|false|false||visionnull|Leg|Anatomy|false|false||leg
null|Lower Extremity|Anatomy|false|false||legnull|Weakness|Finding|false|false||weakness
null|Asthenia|Finding|false|false||weaknessnull|Trouble with Coordination|Finding|false|false||trouble with coordinationnull|Coordination of Benefits - Coordination|Finding|false|false||coordination
null|Coordinated|Finding|false|false||coordination
null|Physiologic Coordination|Finding|false|false||coordinationnull|Balance (substance)|Drug|false|false||balance
null|Balance (substance)|Drug|false|false||balancenull|Ability to balance|Finding|false|false||balance
null|Equilibrium|Finding|false|false||balancenull|examination of balance|Procedure|false|false||balancenull|balance device|Device|false|false||balancenull|Balanced (qualifier value)|Modifier|false|false||balancenull|Dyspnea|Finding|true|false||shortness of breathnull|null|Attribute|true|false||shortness of breathnull|Breath|Finding|false|false||breathnull|Chest Pain|Finding|true|false|C1527391;C0817096|chest painnull|null|Attribute|true|false|C1527391;C0817096|chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0008031;C2926613;C1549543;C0030193;C0741025|chest
null|Anterior thoracic region|Anatomy|false|false|C0008031;C2926613;C1549543;C0030193;C0741025|chestnull|Abdominal Pain|Finding|false|false|C0000726|pain, abdominalnull|Administration Method - Pain|Finding|false|false|C1527391;C0817096|pain
null|Pain|Finding|false|false|C1527391;C0817096|painnull|null|Attribute|false|false||painnull|Abdominal Pain|Finding|true|false|C0000726|abdominal painnull|Abdomen|Anatomy|false|false|C0000737;C1549543;C0030193;C0000737|abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Administration Method - Pain|Finding|true|false|C0000726|pain
null|Pain|Finding|true|false|C0000726|painnull|null|Attribute|true|false||painnull|Multiple Sclerosis|Disorder|false|false||Multiple sclerosisnull|Numerous|LabModifier|false|false||Multiplenull|Sclerosis|Finding|false|false||sclerosisnull|Relationship - Mother|Finding|false|false||Mothernull|Mother (person)|Subject|false|false||Mothernull|Pancreatic carcinoma|Disorder|false|false|C0030274|pancreatic cancer
null|Malignant neoplasm of pancreas|Disorder|false|false|C0030274|pancreatic cancernull|Pancreatic Hormones|Drug|false|false||pancreatic
null|Pancreatic Hormones|Drug|false|false||pancreatic
null|Pancreatic Hormones|Drug|false|false||pancreaticnull|Pancreas|Anatomy|false|false|C0346647;C0235974|pancreaticnull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Brother - courtesy title|Finding|false|false||brother
null|Relationship - Brother|Finding|false|false||brothernull|Brothers|Subject|false|false||brothernull|Malignant neoplasm of lung|Disorder|false|false|C4037972;C0024109|lung cancer
null|Carcinoma of lung|Disorder|false|false|C4037972;C0024109|lung cancernull|Lung diseases|Disorder|false|false|C4037972;C0024109|lungnull|Lung Problem|Finding|false|false|C4037972;C0024109|lungnull|Chest>Lung|Anatomy|false|false|C0024115;C0242379;C0684249;C0740941|lung
null|Lung|Anatomy|false|false|C0024115;C0242379;C0684249;C0740941|lungnull|Malignant Neoplasms|Disorder|false|true||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|true||cancernull|Sister|Subject|false|false||sistersnull|Malignant neoplasm of brain|Disorder|false|false|C4266577;C0006104|brain cancer
null|Brain Neoplasms|Disorder|false|false|C4266577;C0006104|brain cancernull|Brain Diseases|Disorder|false|false|C4266577;C0006104|brainnull|Head>Brain|Anatomy|false|false|C0006826;C0006111;C0153633;C0006118|brain
null|Brain|Anatomy|false|false|C0006826;C0006111;C0153633;C0006118|brainnull|Malignant Neoplasms|Disorder|false|false|C4266577;C0006104|cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|physical examination (physical finding)|Finding|false|false||PHYSICAL EXAMINATIONnull|Physical Examination|Procedure|false|false||PHYSICAL EXAMINATIONnull|physical examination (physical finding)|Finding|false|false||PHYSICAL
null|Physical|Finding|false|false||PHYSICALnull|Physical Examination|Procedure|false|false||PHYSICALnull|Physical Examination|Procedure|false|false||EXAMINATION
null|Medical Examination|Procedure|false|false||EXAMINATIONnull|Examination|Event|false|false||EXAMINATIONnull|On admission|Time|false|false||ON ADMISSIONnull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||Generalnull|General medical service|Procedure|false|false||Generalnull|Generalized|Modifier|false|false||Generalnull|Feeling comfortable|Finding|false|false||comfortablenull|HEENT|Anatomy|false|false|C0026987|HEENTnull|Myelofibrosis|Disorder|false|false|C0694605;C1512338|MMMnull|Medial part of medial mammillary nucleus|Anatomy|false|false|C0026987|MMMnull|Scleral icterus|Finding|true|false|C0036410|scleral icterusnull|Sclera|Anatomy|false|false|C0240962|scleralnull|Icterus|Finding|true|false||icterusnull|Icterus <Icteridae>|Entity|true|false||icterusnull|null|LabModifier|false|false||icterusnull|Exophthalmos|Disorder|true|false||proptosisnull|Scleral Diseases|Disorder|true|false|C0036410|scleranull|examination of sclera|Procedure|true|false|C0036410|scleranull|Sclera|Anatomy|false|false|C0036412;C2228481|scleranull|Malignant neoplasm of conjunctiva|Disorder|false|false|C0229274;C0009758|conjunctiva
null|Benign neoplasm of conjunctiva|Disorder|false|false|C0229274;C0009758|conjunctiva
null|Conjunctival Diseases|Disorder|false|false|C0229274;C0009758|conjunctivanull|Specimen Type - Conjunctiva|Finding|false|false|C0229274;C0009758|conjunctiva
null|null|Finding|false|false|C0229274;C0009758|conjunctivanull|examination of conjunctiva|Procedure|false|false|C0229274;C0009758|conjunctiva
null|Procedure on conjunctiva|Procedure|false|false|C0229274;C0009758|conjunctivanull|Structure of palpebral conjunctiva|Anatomy|false|false|C0021485;C1533685;C1828121;C1550624;C1546576;C0872390;C2228431;C0153628;C0154025;C0009759;C1272883;C0013604|conjunctiva
null|conjunctiva|Anatomy|false|false|C0021485;C1533685;C1828121;C1550624;C1546576;C0872390;C2228431;C0153628;C0154025;C0009759;C1272883;C0013604|conjunctivanull|Edema|Finding|true|false|C0229274;C0009758|edemanull|null|Attribute|true|false||edemanull|Injection|Drug|true|false|C0229274;C0009758|injectionnull|Injection Route of Administration|Finding|true|false|C0229274;C0009758|injectionnull|Injection of therapeutic agent|Procedure|true|false|C0229274;C0009758|injection
null|Injection procedure|Procedure|true|false|C0229274;C0009758|injectionnull|Passive joint movement of neck (finding)|Finding|false|false|C0027530;C3159206|Neck
null|Neck problem|Finding|false|false|C0027530;C3159206|Necknull|dendritic spine neck|Anatomy|false|false|C0332254;C0812434;C0684335|Neck
null|Neck|Anatomy|false|false|C0332254;C0812434;C0684335|Necknull|Supple|Finding|false|false|C0027530;C3159206|supplenull|Heart murmur|Finding|true|false||murmursnull|Pericardial friction rub|Finding|true|false||rubsnull|Carotid bruit|Finding|true|false|C0007272|carotid bruitsnull|Carotid Arteries|Anatomy|false|false|C0007280;C0006318|carotidnull|Bruit|Finding|true|false|C0007272|bruitsnull|Pulmonary ventilator management|Procedure|false|false||Pulmnull|Cancer/Testis Antigen|Drug|false|false||CTAnull|PCYT1A wt Allele|Finding|false|false||CTA
null|CERNA3 gene|Finding|false|false||CTAnull|Cardiac Computerized Tomographic Angiography|Procedure|false|false||CTAnull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false|C0449202;C0000726|Abdnull|ABD (body structure)|Anatomy|false|false|C3811055|Abd
null|Abdomen|Anatomy|false|false|C3811055|Abdnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||softnull|Soft|Modifier|false|false||softnull|Bowel sounds|Finding|false|false|C0021853|bowel soundsnull|Intestines|Anatomy|false|false|C0232693|bowelnull|null|Device|false|false||soundsnull|null|Phenomenon|false|false||soundsnull|All extremities|Anatomy|false|false|C0013604;C0010520|Extremities
null|Limb structure|Anatomy|false|false|C0013604;C0010520|Extremitiesnull|Cyanosis|Finding|true|false|C0278454;C0015385|cyanosisnull|Edema|Finding|true|false|C0278454;C0015385|edemanull|null|Attribute|true|false||edemanull|Skin and subcutaneous tissue disorders|Disorder|false|false|C1123023;C4520765|Skin
null|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false|C1123023;C4520765|Skinnull|Skin Specimen Source Code|Finding|false|false|C1123023;C4520765|Skin
null|Skin Specimen|Finding|false|false|C1123023;C4520765|Skinnull|Skin, Human|Anatomy|false|false|C0687712;C0178298;C0496955;C0582051;C1546781;C0444099|Skin
null|Skin|Anatomy|false|false|C0687712;C0178298;C0496955;C0582051;C1546781;C0444099|Skinnull|Feels warm|Finding|false|false|C1123023;C4520765|warmnull|warming process|Phenomenon|false|false|C1123023;C4520765|warmnull|Pink color|Modifier|false|false||pinknull|Skin rash|Finding|true|false||rashes
null|Exanthema|Finding|true|false||rashesnull|Neurologic (qualifier value)|Modifier|false|false||Neurologicnull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|Mental state|Finding|false|false||MENTAL STATUSnull|null|Attribute|false|false||MENTAL STATUS
null|null|Attribute|false|false||MENTAL STATUSnull|Psyche structure|Finding|false|false||MENTALnull|What subject filter - Status|Finding|false|false||STATUSnull|null|Attribute|false|false||STATUSnull|Social status|Modifier|false|false||STATUS
null|Status|Modifier|false|false||STATUSnull|Alert brand of caffeine|Drug|false|false||alert
null|Alert brand of caffeine|Drug|false|false||alertnull|Mentally alert|Finding|false|false||alert
null|Consciousness clear|Finding|false|false||alert
null|Alert note|Finding|false|false||alert
null|Alert|Finding|false|false||alertnull|null|Attribute|false|false||alertnull|Oriented to place|Finding|false|false||orientednull|Orientation, Spatial|Modifier|false|false||orientednull|midline cell component|Anatomy|false|false||midlinenull|Midline (qualifier value)|Modifier|false|false||midlinenull|Recent|Time|false|false||recentnull|Distant Metastasis|Finding|false|false||distantnull|Distant|Modifier|false|false||distantnull|Event|Event|false|false||eventsnull|Visual neglect|Finding|true|false||visual neglectnull|Visual|Finding|false|false||visualnull|Victim of neglect (finding)|Finding|true|false||neglectnull|Neglect (event)|Event|true|false||neglectnull|physical examination (physical finding)|Finding|false|false||PHYSICAL EXAMINATIONnull|Physical Examination|Procedure|false|false||PHYSICAL EXAMINATIONnull|physical examination (physical finding)|Finding|false|false||PHYSICAL
null|Physical|Finding|false|false||PHYSICALnull|Physical Examination|Procedure|false|false||PHYSICALnull|Physical Examination|Procedure|false|false||EXAMINATION
null|Medical Examination|Procedure|false|false||EXAMINATIONnull|Examination|Event|false|false||EXAMINATIONnull|On discharge|Time|false|false||ON DISCHARGEnull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|Nuclear magnetic resonance imaging brain|Procedure|false|false|C4266577;C0006104|MRI Brainnull|CYREN gene|Finding|false|false|C4266577;C0006104|MRInull|Magnetic resonance imaging service|Procedure|false|false|C4266577;C0006104|MRI
null|Magnetic Resonance Imaging|Procedure|false|false|C4266577;C0006104|MRInull|Maori Language|Entity|false|false||MRInull|Brain Diseases|Disorder|false|false|C4266577;C0006104|Brainnull|Head>Brain|Anatomy|false|false|C0024485;C0587658;C0006111;C1824234;C4028269|Brain
null|Brain|Anatomy|false|false|C0024485;C0587658;C0006111;C1824234;C4028269|Brainnull|Operative|Time|false|false||Operativenull|null|Finding|false|false||Planning
null|Planned|Finding|false|false||Planningnull|Reduced|Finding|false|false|C0230003|Decreasenull|Decrease|LabModifier|false|false||Decreasenull|size|Modifier|false|false||sizenull|size - solid dosage form|LabModifier|false|false||sizenull|Known|Modifier|false|false||knownnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Coronal (qualifier value)|Modifier|false|false||frontalnull|Graph Node|Finding|false|false|C0230003|vertexnull|Vertex|Anatomy|false|false|C0392756;C1308727;C2697524;C5575294;C1419293;C1424873;C2347743|vertexnull|RBBP8 protein, human|Drug|false|false|C0230003|rim
null|RBBP8 protein, human|Drug|false|false|C0230003|rimnull|RIMS1 wt Allele|Finding|false|false|C0230003|rim
null|RBBP8 gene|Finding|false|false|C0230003|rim
null|RIMS1 gene|Finding|false|false|C0230003|rim
null|RBBP8 wt Allele|Finding|false|false|C0230003|rimnull|HL7 Reference Information Model|Device|false|false||rimnull|Rim|Modifier|false|false||rimnull|Lesion|Finding|false|false||lesion
null|null|Finding|false|false||lesionnull|null|Finding|false|false||unchangednull|About The Same|Modifier|false|false||unchangednull|Vasogenic Edema|Finding|false|false||vasogenic edemanull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Mass Effect|Finding|false|false||mass effectnull|Morphology, Attenuation, Size, and Structure Criteria|Finding|false|false||mass
null|null|Finding|false|false||mass
null|FBN1 wt Allele|Finding|false|false||mass
null|FBN1 gene|Finding|false|false||mass
null|Mass of body region|Finding|false|false||mass
null|Mass of body structure|Finding|false|false||massnull|Mass, a measure of quantity of matter|LabModifier|false|false||mass
null|Molecular Mass|LabModifier|false|false||massnull|Effect, Appearance|Modifier|false|false||effect
null|Effect|Modifier|false|false||effectnull|CAT scan of head|Procedure|false|false|C0018670;C0152336|Head CTnull|Problems with head|Disorder|false|false|C0018670;C0152336|Headnull|Procedure on head|Procedure|false|false|C0018670;C0152336|Headnull|Structure of head of caudate nucleus|Anatomy|false|false|C0202691;C0362076;C0876917|Head
null|Head|Anatomy|false|false|C0202691;C0362076;C0876917|Headnull|Head Device|Device|false|false||Headnull|Radionuclide Imaging|Procedure|false|false||SCAN
null|Scanning|Procedure|false|false||SCANnull|Status post|Time|false|false||Status post
null|Post|Time|false|false||Status postnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Revision|Time|false|false||redonull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Parietal|Modifier|false|false||parietalnull|Graph Node|Finding|false|false|C0230003|vertexnull|Vertex|Anatomy|false|false|C2697524;C0010280|vertexnull|Craniotomy|Procedure|false|false|C0230003|craniotomynull|Evidence of (contextual qualifier)|Finding|false|false||evidence ofnull|Evidence|Finding|false|false||evidencenull|Hemorrhage|Finding|false|false||hemorrhagenull|Patient Condition Code - Stable|Finding|false|false||Stablenull|Stable status|Modifier|false|false||Stablenull|Vasogenic Edema|Finding|false|false||vasogenic edemanull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Table Cell Horizontal Align - right|Finding|false|false|C0796494;C0030560;C0546003|rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Frontal and parietal lobes|Anatomy|false|false|C1552823|frontal and parietal lobesnull|Coronal (qualifier value)|Modifier|false|false||frontalnull|Parietal Lobe|Anatomy|false|false|C1552823|parietal lobesnull|Parietal|Modifier|false|false||parietalnull|lobe|Anatomy|false|false|C1552823|lobesnull|Neurosurgical Procedures|Procedure|false|false||neurosurgerynull|Science of neurosurgery|Title|false|false||neurosurgerynull|ActInformationPrivacyReason - service|Finding|false|false||servicenull|Software Service|Device|false|false||servicenull|Services|Event|false|false||servicenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Communicable Diseases|Disorder|false|false||Infectiousnull|infectious - Entity Risk|Modifier|false|false||Infectiousnull|Disease|Disorder|false|false|C4266577;C0006104|Diseasenull|Clinic|Device|false|false||Clinic
null|Ambulatory Care Facilities|Device|false|false||Clinicnull|Clinic|Entity|false|false||Clinic
null|Ambulatory Care Facilities|Entity|false|false||Clinicnull|Patient location type - Clinic|Modifier|false|false||Clinic
null|Person location type - Clinic|Modifier|false|false||Clinicnull|anticipation|Finding|false|false|C4266577;C0006104|anticipationnull|Evacuation procedure|Procedure|false|false|C4266577;C0006104|evacuationnull|Brain Diseases|Disorder|false|false|C4266577;C0006104|brainnull|Head>Brain|Anatomy|false|false|C0679106;C0012634;C1282573;C0006111|brain
null|Brain|Anatomy|false|false|C0679106;C0012634;C1282573;C0006111|brainnull|Abscess|Disorder|false|false||abscessnull|null|Finding|false|false||abscessnull|CYREN gene|Finding|false|false||MRInull|Magnetic resonance imaging service|Procedure|false|false||MRI
null|Magnetic Resonance Imaging|Procedure|false|false||MRInull|Maori Language|Entity|false|false||MRInull|History of surgery|Finding|false|false||prior surgerynull|null|Time|false|false||priornull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Operative|Time|false|false||operativenull|null|Finding|false|false||planning
null|Planned|Finding|false|false||planningnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Craniotomy|Procedure|false|false||craniotomynull|Evacuation procedure|Procedure|false|false||evacuationnull|Abscess|Disorder|false|false||abscessnull|null|Finding|false|false||abscessnull|Procedure (set of actions)|Finding|false|false||procedurenull|Interventional procedure|Procedure|false|false||procedurenull|null|Attribute|false|false||procedurenull|Act Class - procedure|Event|false|false||procedurenull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Operating Room|Device|false|false||operating roomnull|Operating Room|Entity|false|false||operating roomnull|Patient location type - Operating Room|Modifier|false|false||operating roomnull|Operating|Finding|false|false||operatingnull|Room - Patient location type|Modifier|false|false||room
null|Room|Modifier|false|false||roomnull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|Inventory of Callous-Unemotional Traits|Finding|false|false|C0228479|ICUnull|Structure of intraculminate fissure|Anatomy|false|false|C2004454;C0237820;C4554035|ICUnull|intensive care unit|Device|false|false||ICUnull|intensive care unit|Entity|false|false||ICUnull|Recovery - healing process|Finding|false|false|C0228479|recoverynull|null|Event|false|false|C0228479|recoverynull|recovery - adjustment|LabModifier|false|false||recoverynull|Postoperative Period|Time|false|false||post-operativenull|CAT scan of head|Procedure|false|false|C0018670;C0152336|head CTnull|Problems with head|Disorder|false|false|C0018670;C0152336|headnull|Procedure on head|Procedure|false|false|C0018670;C0152336|headnull|Structure of head of caudate nucleus|Anatomy|false|false|C0392747;C0362076;C0202691;C0876917;C0241311|head
null|Head|Anatomy|false|false|C0392747;C0362076;C0202691;C0876917;C0241311|headnull|Head Device|Device|false|false||headnull|post operative (finding)|Finding|false|false|C0018670;C0152336|post operativenull|Operative|Time|false|false||operativenull|Changing|Finding|false|false|C0018670;C0152336|changesnull|Changed status|LabModifier|false|false||changesnull|Query Status Code - new|Finding|true|false||new
null|Act Status - new|Finding|true|false||newnull|Newar Language|Entity|true|false||newnull|New|Modifier|false|false||newnull|Chairs|Device|false|false||chairnull|Chairperson|Subject|false|false||chairnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Floor (anatomic)|Anatomy|false|false||floornull|floor (object)|Device|false|false||floornull|Floor - story of building|Entity|false|false||floornull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Communicable Diseases|Disorder|false|false||Infectious Diseasenull|Infectious Disease Medicine|Title|false|false||Infectious Diseasenull|Communicable Diseases|Disorder|false|false||Infectiousnull|infectious - Entity Risk|Modifier|false|false||Infectiousnull|Disease|Disorder|false|false||Diseasenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|vancomycin|Drug|false|false||vancomycin
null|vancomycin|Drug|false|false||vancomycinnull|Vancomycin measurement|Procedure|false|false||vancomycinnull|INJECTION, MEROPENEM, 100 MG ADMINISTERED|Drug|false|false||meropenem
null|meropenem|Drug|false|false||meropenem
null|meropenem|Drug|false|false||meropenemnull|Culture Dose Form|Drug|false|false||culturenull|Culture (Anthropological)|Finding|false|false||culture
null|Cultural aspects|Finding|false|false||culturenull|Microbial culture (procedure)|Procedure|false|false||culture
null|Laboratory culture|Procedure|false|false||culturenull|Data|Finding|false|false||datanull|Data call receiving device|Device|false|false||datanull|Data <Amphipyrinae>|Entity|false|false||datanull|Problems with head|Disorder|false|false|C0018670;C0152336|headnull|Procedure on head|Procedure|false|false|C0018670;C0152336|headnull|Structure of head of caudate nucleus|Anatomy|false|false|C3263723;C0043251;C0043250;C0876917;C1549529;C1547965;C1550680;C0362076|head
null|Head|Anatomy|false|false|C3263723;C0043251;C0043250;C0876917;C1549529;C1547965;C1550680;C0362076|headnull|Head Device|Device|false|false||headnull|Traumatic Wound|Disorder|false|false|C0018670;C0152336|wound
null|Wounds and Injuries|Disorder|false|false|C0018670;C0152336|wound
null|Traumatic injury|Disorder|false|false|C0018670;C0152336|woundnull|Route of Administration - Wound|Finding|false|false|C0018670;C0152336|wound
null|null|Finding|false|false|C0018670;C0152336|wound
null|Specimen Type - Wound|Finding|false|false|C0018670;C0152336|woundnull|Culture (Anthropological)|Finding|false|false||culturesnull|Growth & development aspects|Finding|true|false||growth
null|Tissue Growth|Finding|true|false||growth
null|Growth|Finding|true|false||growth
null|growth aspects|Finding|true|false||growthnull|Growth action|Phenomenon|true|false||growthnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|vancomycin|Drug|false|false||Vancomycin
null|vancomycin|Drug|false|false||Vancomycinnull|Vancomycin measurement|Procedure|false|false||Vancomycinnull|INJECTION, MEROPENEM, 100 MG ADMINISTERED|Drug|false|false||meropenem
null|meropenem|Drug|false|false||meropenem
null|meropenem|Drug|false|false||meropenemnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Residual|Modifier|false|false||residualnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Weakness|Finding|false|false||weakness
null|Asthenia|Finding|false|false||weaknessnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Numbness|Finding|false|false||numbness
null|Hypesthesia|Finding|false|false||numbnessnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Problems with head|Disorder|false|false|C0018670;C0152336|headnull|Procedure on head|Procedure|false|false|C0018670;C0152336|headnull|Structure of head of caudate nucleus|Anatomy|false|false|C0876917;C0362076|head
null|Head|Anatomy|false|false|C0876917;C0362076|headnull|Head Device|Device|false|false||headnull|Contrast Media|Drug|false|false||contrastnull|Contrast|Modifier|false|false||contrastnull|Driving While Intoxicated|Finding|false|false||DWInull|Diffusion weighted imaging|Procedure|false|false||DWInull|Intensity and Distress 1|Finding|false|false||slightnull|Slight (qualifier value)|Modifier|false|false||slight
null|Mild (qualifier value)|Modifier|false|false||slightnull|Improvement|Finding|false|false||improvementnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Appropriate|Modifier|false|false||appropriatenull|Follow-up status|Finding|false|false||follow-upnull|follow-up|Procedure|false|false||follow-upnull|Follow - dosing instruction imperative|Finding|false|false||follow
null|Follow|Finding|false|false||follownull|Followed by|Time|false|false||follownull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|MEDICATION LIST|Finding|false|false||Medication listnull|Pharmaceutical Preparations|Drug|false|false||Medicationnull|medication - HL7 publishing domain|Finding|false|false||Medication
null|Medications|Finding|false|false||Medicationnull|List|Finding|false|false||list
null|Sequence Data Type|Finding|false|false||listnull|Accurate (qualifier value)|Modifier|false|false||accuratenull|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||completenull|Completion Status for valid values - Complete|Finding|false|false||complete
null|Data operation - complete|Finding|false|false||complete
null|Finish - dosing instruction imperative|Finding|false|false||completenull|Complete|Modifier|false|false||completenull|ceftriaxone|Drug|false|false||CeftriaXONE
null|ceftriaxone|Drug|false|false||CeftriaXONEnull|Every twelve hours|Time|false|false||Q12Hnull|metronidazole|Drug|false|false||MetRONIDAZOLE
null|metronidazole|Drug|false|false||MetRONIDAZOLEnull|Flagyl|Drug|false|false||FLagyl
null|Flagyl|Drug|false|false||FLagylnull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|oxycodone|Drug|false|false||OxycoDONE
null|oxycodone|Drug|false|false||OxycoDONEnull|Oxycodone measurement|Procedure|false|false||OxycoDONEnull|Immediate Release Dosage Form|Drug|false|false||Immediate Releasenull|Query Priority - Immediate|Finding|false|false||Immediate
null|immediate - ResponseCode|Finding|false|false||Immediatenull|Immediate|Time|false|false||Immediate
null|Stat (do immediately)|Time|false|false||Immediatenull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|levetiracetam|Drug|false|false||LeVETiracetam
null|levetiracetam|Drug|false|false||LeVETiracetamnull|Measurement of levetiracetam|Procedure|false|false||LeVETiracetamnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|ADMIN.FACILITY|Finding|false|false||Facilitynull|Facility (object)|Device|false|false||Facilitynull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Brain Abscess|Disorder|false|false|C4266577;C0006104|Brain Abscess
null|Cerebral abscess|Disorder|false|false|C4266577;C0006104|Brain Abscessnull|Brain Diseases|Disorder|false|false|C4266577;C0006104|Brainnull|Head>Brain|Anatomy|false|false|C0006111;C0000833;C0006105;C1510428;C1546533|Brain
null|Brain|Anatomy|false|false|C0006111;C0000833;C0006105;C1510428;C1546533|Brainnull|Abscess|Disorder|false|false|C4266577;C0006104|Abscessnull|null|Finding|false|false|C4266577;C0006104|Abscessnull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Coordination of Benefits - Independent|Finding|false|false||Independent
null|Religious Affiliation - Independent|Finding|false|false||Independent
null|Independence|Finding|false|false||Independent
null|Independently able|Finding|false|false||Independentnull|Staple, Surgical|Device|false|false||staplesnull|Cleaning (activity)|Event|false|false||cleannull|Relationship - Friend|Finding|false|false||friendnull|friend|Subject|false|false||friendnull|Family member|Subject|false|false||family membernull|Entity Name Part Type - family|Finding|false|false||family
null|Last Name|Finding|false|false||family
null|Living Arrangement - Family|Finding|false|false||family
null|Family (taxonomic)|Finding|false|false||family
null|Family Collection|Finding|false|false||familynull|Family|Subject|false|false||familynull|Member Organization|Subject|false|false||member
null|Role Class - member|Subject|false|false||member
null|member|Subject|false|false||membernull|Traumatic Wound|Disorder|false|false||wound
null|Wounds and Injuries|Disorder|false|false||wound
null|Traumatic injury|Disorder|false|false||woundnull|Route of Administration - Wound|Finding|false|false||wound
null|null|Finding|false|false||wound
null|Specimen Type - Wound|Finding|false|false||woundnull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|Erythema|Disorder|false|false||rednessnull|Redness|Finding|false|false||rednessnull|Red color|Modifier|false|false||rednessnull|Body Substance Discharge|Finding|false|false||drainage
null|Body Fluid Discharge|Finding|false|false||drainagenull|Drainage procedure|Procedure|false|false||drainagenull|Daily|Time|false|false||dailynull|Analgesics|Drug|false|false||pain medicine
null|Analgesics|Drug|false|false||pain medicine
null|Analgesics|Drug|false|false||pain medicinenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicinenull|Medicine|Title|false|false||medicinenull|Have Pain|Finding|false|false||have painnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Exercise|Finding|false|false||Exercisenull|Exercise Pain Management|Procedure|false|false||Exercisenull|history of recreational walking|Finding|false|false||walking
null|walking - neurological symptom|Finding|false|false||walking
null|Walking (function)|Finding|false|false||walkingnull|Lifting|Event|true|false||liftingnull|Straining (finding)|Finding|false|false||strainingnull|Excessive (qualifier value)|Modifier|false|false||excessivenull|Decompression Sickness|Disorder|false|false||bendingnull|Bending - Changing basic body position|Finding|false|false||bending
null|Does bend|Finding|false|false||bendingnull|Bent|Modifier|false|false||bendingnull|Intake|Finding|false|false|C1304649|intakenull|Measurement of fluid intake|Procedure|false|false|C1304649|intake
null|Intake (treatment)|Procedure|false|false|C1304649|intakenull|Liquid substance|Drug|false|false||fluidsnull|Mouse Body Fluid or Substance|Finding|false|false||fluidsnull|Fluid Therapy|Procedure|false|false||fluidsnull|Fiber brand of calcium polycarbophil|Drug|false|false|C1304649|fiber
null|fiber|Drug|false|false|C1304649|fiber
null|fiber|Drug|false|false|C1304649|fiber
null|Fiber brand of calcium polycarbophil|Drug|false|false|C1304649|fibernull|Tissue fiber|Anatomy|false|false|C4521161;C3251814;C1512806;C0225326;C1321801|fibernull|Fiber Device|Device|false|false||fibernull|Animal in fiber production|Entity|false|false||fiber
null|Plant fiber|Entity|false|false||fibernull|Narcotics|Drug|false|false||narcotic
null|Narcotics|Drug|false|false||narcoticnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicinenull|Medicine|Title|false|false||medicinenull|Constipation|Finding|false|false||constipationnull|Drugs, Non-Prescription|Drug|false|false||over the counternull|Counter brand of Terbufos|Drug|false|false||counter
null|Counter brand of Terbufos|Drug|false|false||counternull|Counter device|Device|false|false||counternull|Stool Softener brand of docusate sodium|Drug|false|false||stool softener
null|Stool Softener brand of docusate sodium|Drug|false|false||stool softener
null|Stool Softener|Drug|false|false||stool softenernull|Feces|Finding|false|false||stoolnull|Stool seat|Device|false|false||stoolnull|docusate|Drug|false|false||Docusate
null|docusate|Drug|false|false||Docusatenull|Colace|Drug|false|false||Colace
null|Colace|Drug|false|false||Colacenull|Narcotics|Drug|false|false||narcotic
null|Narcotics|Drug|false|false||narcoticnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Anti-Inflammatory Agents|Drug|false|false||anti-inflammatorynull|Anti-inflammatory effect|Modifier|false|false||anti-inflammatorynull|Pharmaceutical Preparations|Drug|false|false||medicinesnull|Motrin|Drug|false|false||Motrin
null|Motrin|Drug|false|false||Motrinnull|aspirin|Drug|false|false||Aspirin
null|aspirin|Drug|false|false||Aspirinnull|Advil|Drug|false|false||Advil
null|Advil|Drug|false|false||Advilnull|AVIL gene|Finding|false|false||Advilnull|ibuprofen|Drug|false|false||Ibuprofen
null|ibuprofen|Drug|false|false||Ibuprofennull|Follow-up status|Finding|false|false||follow upnull|follow-up|Procedure|false|false||follow upnull|Follow - dosing instruction imperative|Finding|false|false||follow
null|Follow|Finding|false|false||follownull|Followed by|Time|false|false||follownull|Keppra|Drug|false|false||Keppra
null|Keppra|Drug|false|false||Keppranull|levetiracetam|Drug|false|false||Levetiracetam
null|levetiracetam|Drug|false|false||Levetiracetamnull|Measurement of levetiracetam|Procedure|false|false||Levetiracetamnull|Pharmaceutical Preparations|Drug|false|false||medicinenull|Medicine|Title|false|false||medicinenull|Blood and lymphatic system disorders|Disorder|true|false||bloodnull|peripheral blood|Finding|true|false||blood
null|Blood|Finding|true|false||blood
null|In Blood|Finding|true|false||bloodnull|Work|Event|true|false||worknull|Preventive monitoring|Procedure|false|false||monitoringnull|null|Event|false|false||monitoringnull|Follow-up status|Finding|false|false||follow upnull|follow-up|Procedure|false|false||follow upnull|Follow - dosing instruction imperative|Finding|false|false||follow
null|Follow|Finding|false|false||follownull|Followed by|Time|false|false||follownull|Appointments|Event|false|false||appointmentnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions