 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
_|27,28
_|28,29
_|29,30
No|31,33
:|33,34
_|37,38
_|38,39
_|39,40
<EOL>|40,41
<EOL>|42,43
Admission|43,52
Date|53,57
:|57,58
_|60,61
_|61,62
_|62,63
Discharge|77,86
Date|87,91
:|91,92
_|95,96
_|96,97
_|97,98
<EOL>|98,99
<EOL>|100,101
Date|101,105
of|106,108
Birth|109,114
:|114,115
_|117,118
_|118,119
_|119,120
Sex|133,136
:|136,137
F|140,141
<EOL>|141,142
<EOL>|143,144
Service|144,151
:|151,152
NEUROLOGY|153,162
<EOL>|162,163
<EOL>|164,165
Sulfa|177,182
(|183,184
Sulfonamides|184,196
)|196,197
/|198,199
Penicillins|200,211
<EOL>|211,212
<EOL>|213,214
Attending|214,223
:|223,224
_|225,226
_|226,227
_|227,228
<EOL>|228,229
<EOL>|230,231
Facial|248,254
weakness|255,263
<EOL>|263,264
<EOL>|265,266
Major|266,271
Surgical|272,280
or|281,283
Invasive|284,292
Procedure|293,302
:|302,303
<EOL>|303,304
None|304,308
<EOL>|308,309
<EOL>|310,311
HPI|339,342
:|342,343
_|344,345
_|345,346
_|346,347
RHF|348,351
w|352,353
/|353,354
hx|355,357
GERD|358,362
,|362,363
mild|364,368
depression|369,379
,|379,380
and|381,384
prior|385,390
migraines|391,400
,|400,401
<EOL>|401,402
presents|402,410
now|411,414
with|415,419
episode|420,427
of|428,430
facial|431,437
numbness|438,446
.|446,447
She|448,451
had|452,455
been|456,460
lying|461,466
<EOL>|466,467
on|467,469
her|470,473
left|474,478
face|479,483
,|483,484
watching|485,493
TV|494,496
,|496,497
and|498,501
noticed|502,509
when|510,514
she|515,518
got|519,522
up|523,525
that|526,530
<EOL>|530,531
her|531,534
left|535,539
face|540,544
was|545,548
numb|549,553
as|554,556
if|557,559
she|560,563
were|564,568
injected|569,577
with|578,582
novacaine|583,592
,|592,593
<EOL>|594,595
in|595,597
<EOL>|597,598
a|598,599
distribution|600,612
that|613,617
she|618,621
traces|622,628
along|629,634
mid-V2|635,641
down|642,646
to|647,649
her|650,653
jaw|654,657
<EOL>|658,659
line|659,663
.|663,664
<EOL>|664,665
She|665,668
initially|669,678
thought|679,686
it|687,689
was|690,693
_|694,695
_|695,696
_|696,697
the|698,701
way|702,705
she|706,709
was|710,713
lying|714,719
,|719,720
but|721,724
<EOL>|724,725
became|725,731
concerned|732,741
when|742,746
it|747,749
persisted|750,759
.|759,760
She|761,764
endorsed|765,773
a|774,775
mild|776,780
diffuse|781,788
<EOL>|788,789
dull|789,793
HA|794,796
that|797,801
is|802,804
not|805,808
unusual|809,816
for|817,820
her|821,824
.|824,825
She|826,829
states|830,836
in|837,839
some|840,844
ways|845,849
,|849,850
it|851,853
<EOL>|853,854
felt|854,858
as|859,861
though|862,868
a|869,870
migraine|871,879
were|880,884
coming|885,891
on|892,894
,|894,895
though|896,902
the|903,906
HA|907,909
she|910,913
had|914,917
<EOL>|917,918
was|918,921
not|922,925
typical|926,933
of|934,936
her|937,940
past|941,945
migraines|946,955
.|955,956
The|957,960
numbness|961,969
lasted|970,976
90|977,979
<EOL>|979,980
minutes|980,987
,|987,988
and|989,992
has|993,996
now|997,1000
resolved|1001,1009
completely|1010,1020
.|1020,1021
There|1022,1027
was|1028,1031
no|1032,1034
<EOL>|1035,1036
associated|1036,1046
<EOL>|1046,1047
weakness|1047,1055
,|1055,1056
no|1057,1059
sensory|1060,1067
changes|1068,1075
outside|1076,1083
of|1084,1086
her|1087,1090
face|1091,1095
,|1095,1096
no|1097,1099
VC|1100,1102
,|1102,1103
<EOL>|1104,1105
vertigo|1105,1112
,|1112,1113
<EOL>|1113,1114
or|1114,1116
language|1117,1125
impairment|1126,1136
.|1136,1137
She|1138,1141
can|1142,1145
not|1145,1148
recall|1149,1155
something|1156,1165
like|1166,1170
this|1171,1175
<EOL>|1175,1176
happening|1176,1185
before|1186,1192
,|1192,1193
and|1194,1197
states|1198,1204
that|1205,1209
her|1210,1213
day|1214,1217
was|1218,1221
otherwise|1222,1231
routine|1232,1239
.|1239,1240
<EOL>|1240,1241
On|1241,1243
ROS|1244,1247
,|1247,1248
she|1249,1252
notes|1253,1258
that|1259,1263
about|1264,1269
2|1270,1271
weeks|1272,1277
ago|1278,1281
she|1282,1285
had|1286,1289
diarrhea|1290,1298
for|1299,1302
1|1303,1304
<EOL>|1304,1305
week|1305,1309
which|1310,1315
resolved|1316,1324
spontaneously|1325,1338
.|1338,1339
She|1340,1343
also|1344,1348
endorses|1349,1357
feeling|1358,1365
<EOL>|1365,1366
"|1366,1367
achey|1367,1372
"|1372,1373
4|1374,1375
days|1376,1380
ago|1381,1384
,|1384,1385
otherwise|1386,1395
,|1395,1396
her|1397,1400
health|1401,1407
has|1408,1411
been|1412,1416
normal|1417,1423
.|1423,1424
<EOL>|1425,1426
<EOL>|1426,1427
<EOL>|1428,1429
GERD|1451,1455
<EOL>|1456,1457
mild|1457,1461
depression|1462,1472
<EOL>|1472,1473
migraines|1473,1482
(|1483,1484
throbing|1484,1492
HA|1493,1495
's|1495,1497
assoc|1498,1503
with|1504,1508
visual|1509,1515
flashes|1516,1523
of|1524,1526
light|1527,1532
)|1532,1533
,|1533,1534
<EOL>|1534,1535
last|1535,1539
_|1540,1541
_|1541,1542
_|1542,1543
years|1544,1549
ago|1550,1553
<EOL>|1554,1555
bunions|1555,1562
<EOL>|1562,1563
<EOL>|1564,1565
:|1579,1580
<EOL>|1580,1581
_|1581,1582
_|1582,1583
_|1583,1584
<EOL>|1584,1585
:|1599,1600
<EOL>|1600,1601
Father|1601,1607
with|1608,1612
HD|1613,1615
,|1615,1616
sustained|1617,1626
a|1627,1628
stroke|1629,1635
after|1636,1641
a|1642,1643
cardiac|1644,1651
cath|1652,1656
.|1656,1657
Later|1658,1663
<EOL>|1664,1665
in|1665,1667
<EOL>|1667,1668
life|1668,1672
father|1673,1679
developed|1680,1689
a|1690,1691
meningioma|1692,1702
and|1703,1706
subsequent|1707,1717
seizures|1718,1726
.|1726,1727
<EOL>|1728,1729
<EOL>|1729,1730
<EOL>|1731,1732
98.4|1747,1751
F|1751,1752
69|1753,1755
134|1756,1759
/|1759,1760
79|1760,1762
15|1763,1765
100|1766,1769
%|1769,1770
RA|1770,1772
<EOL>|1773,1774
<EOL>|1774,1775
Gen|1775,1778
:|1778,1779
Lying|1780,1785
in|1786,1788
bed|1789,1792
,|1792,1793
NAD|1794,1797
<EOL>|1797,1798
HEENT|1798,1803
:|1803,1804
NC|1805,1807
/|1807,1808
AT|1808,1810
,|1810,1811
moist|1812,1817
oral|1818,1822
mucosa|1823,1829
<EOL>|1832,1833
Neck|1833,1837
:|1837,1838
No|1839,1841
tenderness|1842,1852
to|1853,1855
palpation|1856,1865
,|1865,1866
normal|1867,1873
ROM|1874,1877
,|1877,1878
supple|1879,1885
,|1885,1886
no|1887,1889
carotid|1890,1897
<EOL>|1897,1898
or|1898,1900
vertebral|1901,1910
bruit|1911,1916
<EOL>|1916,1917
CV|1917,1919
:|1919,1920
RRR|1921,1924
,|1924,1925
Nl|1926,1928
S1|1929,1931
and|1932,1935
S2|1936,1938
,|1938,1939
no|1940,1942
murmurs|1943,1950
/|1950,1951
gallops|1951,1958
/|1958,1959
rubs|1959,1963
<EOL>|1964,1965
Lung|1965,1969
:|1969,1970
Clear|1971,1976
to|1977,1979
auscultation|1980,1992
bilaterally|1993,2004
<EOL>|2005,2006
aBd|2006,2009
:|2009,2010
+|2011,2012
BS|2012,2014
soft|2015,2019
,|2019,2020
nontender|2021,2030
<EOL>|2031,2032
ext|2032,2035
:|2035,2036
no|2037,2039
c|2040,2041
/|2041,2042
c|2042,2043
/|2043,2044
e|2044,2045
;|2045,2046
equal|2047,2052
radial|2053,2059
and|2060,2063
pedal|2064,2069
pulses|2070,2076
B|2077,2078
/|2078,2079
L|2079,2080
.|2080,2081
<EOL>|2082,2083
<EOL>|2083,2084
<EOL>|2085,2086
Neurologic|2086,2096
examination|2097,2108
:|2108,2109
<EOL>|2110,2111
Mental|2111,2117
status|2118,2124
:|2124,2125
Awake|2126,2131
and|2132,2135
alert|2136,2141
,|2141,2142
cooperative|2143,2154
with|2155,2159
exam|2160,2164
,|2164,2165
normal|2166,2172
<EOL>|2173,2174
affect|2174,2180
.|2180,2181
Oriented|2183,2191
to|2192,2194
person|2195,2201
,|2201,2202
place|2203,2208
,|2208,2209
and|2210,2213
date|2214,2218
.|2218,2219
Attentive|2221,2230
,|2230,2231
says|2232,2236
<EOL>|2236,2237
_|2237,2238
_|2238,2239
_|2239,2240
backwards|2241,2250
.|2250,2251
Speech|2253,2259
is|2260,2262
fluent|2263,2269
with|2270,2274
normal|2275,2281
comprehension|2282,2295
and|2296,2299
<EOL>|2299,2300
repetition|2300,2310
;|2310,2311
naming|2312,2318
intact|2319,2325
.|2325,2326
No|2327,2329
dysarthria|2330,2340
.|2340,2341
Reading|2342,2349
intact|2350,2356
.|2356,2357
No|2358,2360
<EOL>|2360,2361
right|2361,2366
left|2367,2371
confusion|2372,2381
.|2381,2382
No|2383,2385
evidence|2386,2394
of|2395,2397
apraxia|2398,2405
or|2406,2408
neglect|2409,2416
.|2416,2417
<EOL>|2417,2418
<EOL>|2419,2420
Cranial|2420,2427
Nerves|2428,2434
:|2434,2435
<EOL>|2437,2438
Pupils|2438,2444
equally|2445,2452
round|2453,2458
and|2459,2462
reactive|2463,2471
to|2472,2474
light|2475,2480
,|2480,2481
4|2482,2483
to|2484,2486
2|2487,2488
mm|2489,2491
<EOL>|2491,2492
bilaterally|2492,2503
.|2503,2504
Visual|2505,2511
fields|2512,2518
are|2519,2522
full|2523,2527
to|2528,2530
confrontation|2531,2544
.|2544,2545
Retinas|2546,2553
<EOL>|2553,2554
with|2554,2558
sharp|2559,2564
disc|2565,2569
margins|2570,2577
B|2578,2579
/|2579,2580
L|2580,2581
.|2581,2582
Extraocular|2583,2594
movements|2595,2604
intact|2605,2611
<EOL>|2611,2612
bilaterally|2612,2623
,|2623,2624
no|2625,2627
nystagmus|2628,2637
.|2637,2638
Sensation|2639,2648
intact|2649,2655
V1|2656,2658
-|2658,2659
V3|2659,2661
to|2662,2664
both|2665,2669
LT|2670,2672
and|2673,2676
<EOL>|2676,2677
PP|2677,2679
.|2679,2680
Facial|2682,2688
movement|2689,2697
symmetric|2698,2707
.|2707,2708
Hearing|2710,2717
intact|2718,2724
to|2725,2727
finger|2728,2734
rub|2735,2738
<EOL>|2738,2739
bilaterally|2739,2750
.|2750,2751
Palate|2753,2759
elevation|2760,2769
symmetrical|2770,2781
.|2781,2782
Sternocleidomastoid|2784,2803
<EOL>|2803,2804
and|2804,2807
trapezius|2808,2817
normal|2818,2824
bilaterally|2825,2836
.|2836,2837
Tongue|2838,2844
midline|2845,2852
,|2852,2853
movements|2854,2863
<EOL>|2863,2864
intact|2864,2870
<EOL>|2870,2871
<EOL>|2872,2873
Motor|2873,2878
:|2878,2879
<EOL>|2880,2881
Normal|2881,2887
bulk|2888,2892
bilaterally|2893,2904
.|2904,2905
Tone|2906,2910
normal|2911,2917
.|2917,2918
No|2919,2921
observed|2922,2930
myoclonus|2931,2940
or|2941,2943
<EOL>|2943,2944
tremor|2944,2950
<EOL>|2950,2951
No|2951,2953
pronator|2954,2962
drift|2963,2968
<EOL>|2968,2969
Del|2971,2974
Tri|2975,2978
Bi|2979,2981
WF|2983,2985
WE|2986,2988
FE|2989,2991
FF|2992,2994
IP|2996,2998
H|3000,3001
Q|3003,3004
DF|3005,3007
PF|3008,3010
TE|3011,3013
TF|3014,3016
<EOL>|3016,3017
R|3017,3018
_|3020,3021
_|3021,3022
_|3022,3023
_|3025,3026
_|3026,3027
_|3027,3028
_|3030,3031
_|3031,3032
_|3032,3033
_|3035,3036
_|3036,3037
_|3037,3038
5|3040,3041
5|3043,3044
<EOL>|3044,3045
L|3045,3046
_|3048,3049
_|3049,3050
_|3050,3051
_|3053,3054
_|3054,3055
_|3055,3056
_|3058,3059
_|3059,3060
_|3060,3061
_|3063,3064
_|3064,3065
_|3065,3066
5|3068,3069
5|3071,3072
<EOL>|3074,3075
<EOL>|3075,3076
Sensation|3076,3085
:|3085,3086
Intact|3087,3093
to|3094,3096
light|3097,3102
touch|3103,3108
,|3108,3109
pinprick|3110,3118
,|3118,3119
and|3120,3123
proprioception|3124,3138
<EOL>|3138,3139
throughout|3139,3149
.|3149,3150
<EOL>|3151,3152
<EOL>|3152,3153
Reflexes|3153,3161
:|3161,3162
<EOL>|3163,3164
+|3164,3165
2|3165,3166
and|3167,3170
symmetric|3171,3180
throughout|3181,3191
.|3191,3192
<EOL>|3194,3195
Toes|3195,3199
downgoing|3200,3209
bilaterally|3210,3221
<EOL>|3222,3223
<EOL>|3224,3225
Coordination|3225,3237
:|3237,3238
finger|3239,3245
-|3245,3246
nose|3246,3250
-|3250,3251
finger|3251,3257
normal|3258,3264
,|3264,3265
heel|3266,3270
to|3271,3273
shin|3274,3278
normal|3279,3285
,|3285,3286
FT|3287,3289
<EOL>|3289,3290
and|3290,3293
RAMs|3294,3298
normal|3299,3305
.|3305,3306
<EOL>|3307,3308
<EOL>|3309,3310
Gait|3310,3314
:|3314,3315
Narrow|3316,3322
based|3323,3328
,|3328,3329
steady|3330,3336
.|3336,3337
Able|3338,3342
to|3343,3345
tandem|3346,3352
walk|3353,3357
without|3358,3365
<EOL>|3365,3366
difficulty|3366,3376
<EOL>|3376,3377
<EOL>|3377,3378
Romberg|3378,3385
:|3385,3386
Negative|3387,3395
<EOL>|3395,3396
<EOL>|3396,3397
<EOL>|3398,3399
Pertinent|3399,3408
Results|3409,3416
:|3416,3417
<EOL>|3417,3418
_|3418,3419
_|3419,3420
_|3420,3421
06|3422,3424
:|3424,3425
10AM|3425,3429
BLOOD|3430,3435
WBC|3436,3439
-|3439,3440
5.3|3440,3443
RBC|3444,3447
-|3447,3448
4|3448,3449
.|3449,3450
38|3450,3452
Hgb|3453,3456
-|3456,3457
11|3457,3459
.|3459,3460
5|3460,3461
*|3461,3462
Hct|3463,3466
-|3466,3467
36.1|3467,3471
<EOL>|3472,3473
MCV|3473,3476
-|3476,3477
82|3477,3479
MCH|3480,3483
-|3483,3484
26|3484,3486
.|3486,3487
2|3487,3488
*|3488,3489
MCHC|3490,3494
-|3494,3495
31.8|3495,3499
RDW|3500,3503
-|3503,3504
13.3|3504,3508
Plt|3509,3512
_|3513,3514
_|3514,3515
_|3515,3516
<EOL>|3516,3517
_|3517,3518
_|3518,3519
_|3519,3520
11|3521,3523
:|3523,3524
14PM|3524,3528
BLOOD|3529,3534
Neuts|3535,3540
-|3540,3541
52.1|3541,3545
_|3546,3547
_|3547,3548
_|3548,3549
Monos|3550,3555
-|3555,3556
4.7|3556,3559
Eos|3560,3563
-|3563,3564
2.0|3564,3567
<EOL>|3568,3569
Baso|3569,3573
-|3573,3574
0.5|3574,3577
<EOL>|3577,3578
_|3578,3579
_|3579,3580
_|3580,3581
11|3582,3584
:|3584,3585
14PM|3585,3589
BLOOD|3590,3595
_|3596,3597
_|3597,3598
_|3598,3599
PTT|3600,3603
-|3603,3604
33.7|3604,3608
_|3609,3610
_|3610,3611
_|3611,3612
<EOL>|3612,3613
_|3613,3614
_|3614,3615
_|3615,3616
06|3617,3619
:|3619,3620
10AM|3620,3624
BLOOD|3625,3630
Glucose|3631,3638
-|3638,3639
82|3639,3641
UreaN|3642,3647
-|3647,3648
16|3648,3650
Creat|3651,3656
-|3656,3657
0.8|3657,3660
Na|3661,3663
-|3663,3664
140|3664,3667
<EOL>|3668,3669
K|3669,3670
-|3670,3671
4.0|3671,3674
Cl|3675,3677
-|3677,3678
105|3678,3681
HCO3|3682,3686
-|3686,3687
26|3687,3689
AnGap|3690,3695
-|3695,3696
13|3696,3698
<EOL>|3698,3699
_|3699,3700
_|3700,3701
_|3701,3702
11|3703,3705
:|3705,3706
14PM|3706,3710
BLOOD|3711,3716
ALT|3717,3720
-|3720,3721
13|3721,3723
AST|3724,3727
-|3727,3728
19|3728,3730
CK|3731,3733
(|3733,3734
CPK|3734,3737
)|3737,3738
-|3738,3739
69|3739,3741
AlkPhos|3742,3749
-|3749,3750
70|3750,3752
<EOL>|3753,3754
TotBili|3754,3761
-|3761,3762
0.2|3762,3765
<EOL>|3765,3766
_|3766,3767
_|3767,3768
_|3768,3769
11|3770,3772
:|3772,3773
14PM|3773,3777
BLOOD|3778,3783
CK|3784,3786
-|3786,3787
MB|3787,3789
-|3789,3790
NotDone|3790,3797
cTropnT|3798,3805
-|3805,3806
<|3806,3807
0|3807,3808
.|3808,3809
01|3809,3811
<EOL>|3811,3812
_|3812,3813
_|3813,3814
_|3814,3815
11|3816,3818
:|3818,3819
14PM|3819,3823
BLOOD|3824,3829
TotProt|3830,3837
-|3837,3838
7.1|3838,3841
Albumin|3842,3849
-|3849,3850
4.5|3850,3853
Globuln|3854,3861
-|3861,3862
2.6|3862,3865
<EOL>|3866,3867
Calcium|3867,3874
-|3874,3875
9.5|3875,3878
Phos|3879,3883
-|3883,3884
3.7|3884,3887
Mg|3888,3890
-|3890,3891
2.1|3891,3894
<EOL>|3894,3895
_|3895,3896
_|3896,3897
_|3897,3898
02|3899,3901
:|3901,3902
26AM|3902,3906
BLOOD|3907,3912
%|3913,3914
HbA1c|3914,3919
-|3919,3920
5.7|3920,3923
<EOL>|3923,3924
_|3924,3925
_|3925,3926
_|3926,3927
11|3928,3930
:|3930,3931
14PM|3931,3935
BLOOD|3936,3941
ASA|3942,3945
-|3945,3946
NEG|3946,3949
Ethanol|3950,3957
-|3957,3958
NEG|3958,3961
Acetmnp|3962,3969
-|3969,3970
NEG|3970,3973
<EOL>|3974,3975
Bnzodzp|3975,3982
-|3982,3983
NEG|3983,3986
Barbitr|3987,3994
-|3994,3995
NEG|3995,3998
Tricycl|3999,4006
-|4006,4007
NEG|4007,4010
<EOL>|4010,4011
<EOL>|4011,4012
Radiology|4012,4021
Report|4022,4028
MRA|4029,4032
BRAIN|4033,4038
W|4039,4040
/|4040,4041
O|4041,4042
CONTRAST|4043,4051
Study|4052,4057
Date|4058,4062
of|4063,4065
_|4066,4067
_|4067,4068
_|4068,4069
<EOL>|4070,4071
9|4071,4072
:|4072,4073
44|4073,4075
AM|4076,4078
<EOL>|4079,4080
1|4080,4081
.|4081,4082
No|4083,4085
acute|4086,4091
intracranial|4092,4104
abnormality|4105,4116
;|4116,4117
specifically|4118,4130
,|4130,4131
there|4132,4137
is|4138,4140
no|4141,4143
<EOL>|4144,4145
evidence|4145,4153
of|4154,4156
<EOL>|4157,4158
either|4158,4164
acute|4165,4170
or|4171,4173
previous|4174,4182
ischemic|4183,4191
event|4192,4197
.|4197,4198
<EOL>|4199,4200
2.|4200,4202
Normal|4203,4209
cranial|4210,4217
and|4218,4221
cervical|4222,4230
MRA|4231,4234
,|4234,4235
with|4236,4240
no|4241,4243
significant|4244,4255
mural|4256,4261
<EOL>|4262,4263
irregularity|4263,4275
or|4276,4278
<EOL>|4279,4280
flow|4280,4284
-|4284,4285
limiting|4285,4293
stenosis|4294,4302
.|4302,4303
<EOL>|4304,4305
<EOL>|4305,4306
<EOL>|4307,4308
Ms.|4331,4334
_|4335,4336
_|4336,4337
_|4337,4338
is|4339,4341
a|4342,4343
_|4344,4345
_|4345,4346
_|4346,4347
yo|4348,4350
woman|4351,4356
with|4357,4361
a|4362,4363
hx|4364,4366
of|4367,4369
depression|4370,4380
,|4380,4381
GERD|4382,4386
and|4387,4390
<EOL>|4391,4392
migraines|4392,4401
,|4401,4402
presenting|4403,4413
with|4414,4418
an|4419,4421
episode|4422,4429
of|4430,4432
facial|4433,4439
numbness|4440,4448
.|4448,4449
<EOL>|4449,4450
<EOL>|4450,4451
1.|4451,4453
Facial|4454,4460
numbness|4461,4469
.|4469,4470
As|4472,4474
this|4475,4479
episode|4480,4487
preceeded|4488,4497
a|4498,4499
headache|4500,4508
,|4508,4509
<EOL>|4510,4511
suspect|4511,4518
likely|4519,4525
due|4526,4529
to|4530,4532
a|4533,4534
migraine|4535,4543
equivalent|4544,4554
,|4554,4555
however|4556,4563
episode|4564,4571
<EOL>|4572,4573
could|4573,4578
also|4579,4583
be|4584,4586
due|4587,4590
to|4591,4593
a|4594,4595
TIA|4596,4599
in|4600,4602
the|4603,4606
thalamus|4607,4615
.|4615,4616
The|4618,4621
patient|4622,4629
had|4630,4633
an|4634,4636
<EOL>|4637,4638
MRI|4638,4641
,|4641,4642
which|4643,4648
showed|4649,4655
no|4656,4658
signs|4659,4664
of|4665,4667
ischemia|4668,4676
,|4676,4677
and|4678,4681
normal|4682,4688
vasculature|4689,4700
,|4700,4701
<EOL>|4702,4703
making|4703,4709
migraine|4710,4718
equivalent|4719,4729
a|4730,4731
much|4732,4736
more|4737,4741
likely|4742,4748
diagnosis|4749,4758
.|4758,4759
<EOL>|4761,4762
However|4762,4769
,|4769,4770
given|4771,4776
the|4777,4780
possibility|4781,4792
of|4793,4795
TIA|4796,4799
,|4799,4800
she|4801,4804
has|4805,4808
been|4809,4813
started|4814,4821
on|4822,4824
a|4825,4826
<EOL>|4827,4828
daily|4828,4833
aspirin|4834,4841
for|4842,4845
future|4846,4852
stroke|4853,4859
prophylaxis|4860,4871
.|4871,4872
Exam|4874,4878
on|4879,4881
discharge|4882,4891
<EOL>|4892,4893
was|4893,4896
notable|4897,4904
for|4905,4908
mild|4909,4913
symmetric|4914,4923
hyperreflexia|4924,4937
in|4938,4940
the|4941,4944
lower|4945,4950
<EOL>|4951,4952
extremities|4952,4963
,|4963,4964
but|4965,4968
otherwise|4969,4978
normal|4979,4985
neurological|4986,4998
exam|4999,5003
,|5003,5004
with|5005,5009
no|5010,5012
<EOL>|5013,5014
residual|5014,5022
sensory|5023,5030
deficits|5031,5039
.|5039,5040
<EOL>|5040,5041
<EOL>|5042,5043
Medications|5043,5054
on|5055,5057
Admission|5058,5067
:|5067,5068
<EOL>|5068,5069
NEXIUM|5069,5075
40|5076,5078
mg|5079,5081
-|5081,5082
-|5082,5083
1|5083,5084
capsule|5085,5092
(|5092,5093
s|5093,5094
)|5094,5095
by|5096,5098
mouth|5099,5104
once|5105,5109
a|5110,5111
day|5112,5115
<EOL>|5115,5116
PROZAC|5116,5122
20|5123,5125
mg|5126,5128
-|5128,5129
-|5129,5130
1|5130,5131
capsule|5132,5139
(|5139,5140
s|5140,5141
)|5141,5142
by|5143,5145
mouth|5146,5151
once|5152,5156
a|5157,5158
day|5159,5162
<EOL>|5162,5163
<EOL>|5163,5164
<EOL>|5165,5166
Discharge|5166,5175
Medications|5176,5187
:|5187,5188
<EOL>|5188,5189
1.|5189,5191
Pantoprazole|5192,5204
40|5205,5207
mg|5208,5210
Tablet|5211,5217
,|5217,5218
Delayed|5219,5226
Release|5227,5234
(|5235,5236
E.C|5236,5239
.|5239,5240
)|5240,5241
Sig|5242,5245
:|5245,5246
One|5247,5250
<EOL>|5251,5252
(|5252,5253
1|5253,5254
)|5254,5255
Tablet|5256,5262
,|5262,5263
Delayed|5264,5271
Release|5272,5279
(|5280,5281
E.C|5281,5284
.|5284,5285
)|5285,5286
PO|5287,5289
Q24H|5290,5294
(|5295,5296
every|5296,5301
24|5302,5304
hours|5305,5310
)|5310,5311
.|5311,5312
<EOL>|5314,5315
2.|5315,5317
Fluoxetine|5318,5328
20|5329,5331
mg|5332,5334
Capsule|5335,5342
Sig|5343,5346
:|5346,5347
One|5348,5351
(|5352,5353
1|5353,5354
)|5354,5355
Capsule|5356,5363
PO|5364,5366
DAILY|5367,5372
<EOL>|5373,5374
(|5374,5375
Daily|5375,5380
)|5380,5381
.|5381,5382
<EOL>|5384,5385
3.|5385,5387
Aspirin|5388,5395
81|5396,5398
mg|5399,5401
Tablet|5402,5408
,|5408,5409
Delayed|5410,5417
Release|5418,5425
(|5426,5427
E.C|5427,5430
.|5430,5431
)|5431,5432
Sig|5433,5436
:|5436,5437
One|5438,5441
(|5442,5443
1|5443,5444
)|5444,5445
<EOL>|5446,5447
Tablet|5447,5453
,|5453,5454
Delayed|5455,5462
Release|5463,5470
(|5471,5472
E.C|5472,5475
.|5475,5476
)|5476,5477
PO|5478,5480
DAILY|5481,5486
(|5487,5488
Daily|5488,5493
)|5493,5494
.|5494,5495
<EOL>|5497,5498
<EOL>|5498,5499
<EOL>|5500,5501
Discharge|5501,5510
Disposition|5511,5522
:|5522,5523
<EOL>|5523,5524
Home|5524,5528
<EOL>|5528,5529
<EOL>|5530,5531
Discharge|5531,5540
Diagnosis|5541,5550
:|5550,5551
<EOL>|5551,5552
Migraine|5552,5560
<EOL>|5561,5562
<EOL>|5563,5564
Mild|5585,5589
symmetric|5590,5599
hyperreflexia|5600,5613
in|5614,5616
the|5617,5620
lower|5621,5626
extremities|5627,5638
,|5638,5639
otherwise|5640,5649
<EOL>|5650,5651
normal|5651,5657
neurological|5658,5670
exam|5671,5675
.|5675,5676
<EOL>|5676,5677
<EOL>|5677,5678
<EOL>|5679,5680
You|5704,5707
were|5708,5712
admitted|5713,5721
for|5722,5725
left|5726,5730
sided|5731,5736
facial|5737,5743
numbness|5744,5752
.|5752,5753
You|5755,5758
had|5759,5762
an|5763,5765
<EOL>|5766,5767
MRI|5767,5770
which|5771,5776
showed|5777,5783
no|5784,5786
signs|5787,5792
of|5793,5795
ischemia|5796,5804
.|5804,5805
It|5807,5809
is|5810,5812
suspected|5813,5822
that|5823,5827
<EOL>|5828,5829
this|5829,5833
was|5834,5837
related|5838,5845
to|5846,5848
migraine|5849,5857
headaches|5858,5867
,|5867,5868
but|5869,5872
we|5873,5875
recommend|5876,5885
that|5886,5890
<EOL>|5891,5892
you|5892,5895
start|5896,5901
taking|5902,5908
a|5909,5910
full|5911,5915
dose|5916,5920
of|5921,5923
aspirin|5924,5931
.|5931,5932
<EOL>|5932,5933
<EOL>|5933,5934
If|5934,5936
you|5937,5940
notice|5941,5947
new|5948,5951
numbness|5952,5960
,|5960,5961
weakness|5962,5970
,|5970,5971
worsening|5972,5981
headaches|5982,5991
,|5991,5992
or|5993,5995
<EOL>|5996,5997
other|5997,6002
new|6003,6006
concerning|6007,6017
symptoms|6018,6026
,|6026,6027
please|6028,6034
return|6035,6041
to|6042,6044
the|6045,6048
nearest|6049,6056
ED|6057,6059
<EOL>|6060,6061
for|6061,6064
further|6065,6072
evaluation|6073,6083
.|6083,6084
<EOL>|6084,6085
<EOL>|6086,6087
Followup|6087,6095
Instructions|6096,6108
:|6108,6109
<EOL>|6109,6110
_|6110,6111
_|6111,6112
_|6112,6113
<EOL>|6113,6114

