 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|30,34
No|35,37
:|37,38
_|41,42
_|42,43
_|43,44
<EOL>|44,45
<EOL>|46,47
Admission|47,56
Date|57,61
:|61,62
_|64,65
_|65,66
_|66,67
Discharge|81,90
Date|91,95
:|95,96
_|99,100
_|100,101
_|101,102
<EOL>|102,103
<EOL>|104,105
Date|105,109
of|110,112
Birth|113,118
:|118,119
_|121,122
_|122,123
_|123,124
Sex|137,140
:|140,141
M|144,145
<EOL>|145,146
<EOL>|147,148
Service|148,155
:|155,156
SURGERY|157,164
<EOL>|164,165
<EOL>|166,167
No|179,181
Known|182,187
Allergies|188,197
/|198,199
Adverse|200,207
Drug|208,212
Reactions|213,222
<EOL>|222,223
<EOL>|224,225
Attending|225,234
:|234,235
_|236,237
_|237,238
_|238,239
.|239,240
<EOL>|240,241
<EOL>|242,243
Locally|260,267
advanced|268,276
gastric|277,284
carcinoma|285,294
<EOL>|294,295
<EOL>|296,297
Major|297,302
Surgical|303,311
or|312,314
Invasive|315,323
Procedure|324,333
:|333,334
<EOL>|334,335
Cystoscopy|335,345
for|346,349
foley|350,355
catheter|356,364
placement|365,374
;|374,375
Laparoscopy|376,387
with|388,392
<EOL>|393,394
biopsy|394,400
;|400,401
Gastroscopy|402,413
<EOL>|413,414
<EOL>|414,415
<EOL>|416,417
Mr.|445,448
_|449,450
_|450,451
_|451,452
is|453,455
a|456,457
_|458,459
_|459,460
_|460,461
year|462,466
old|467,470
male|471,475
with|476,480
locally|481,488
advanced|489,497
gastric|498,505
<EOL>|506,507
cancer|507,513
(|514,515
stage|515,520
II|521,523
[|524,525
T3N2|525,529
]|529,530
)|530,531
who|532,535
arrives|536,543
to|544,546
_|547,548
_|548,549
_|549,550
for|551,554
<EOL>|555,556
curative|556,564
-|564,565
intent|565,571
surgical|572,580
resection|581,590
after|591,596
completion|597,607
of|608,610
induction|611,620
<EOL>|621,622
chemotherapy|622,634
.|634,635
<EOL>|636,637
<EOL>|637,638
He|638,640
was|641,644
started|645,652
on|653,655
neoadjuvant|656,667
chemotherapy|668,680
with|681,685
FLOT4|686,691
on|692,694
<EOL>|694,695
_|695,696
_|696,697
_|697,698
.|698,699
Overall|700,707
he|708,710
tolerated|711,720
the|721,724
chemotherapy|725,737
well|738,742
without|743,750
any|751,754
<EOL>|755,756
significant|756,767
side|768,772
effects|773,780
.|780,781
However|782,789
,|789,790
last|791,795
<EOL>|795,796
month|796,801
he|802,804
developed|805,814
right|815,820
upper|821,826
extremity|827,836
edema|837,842
and|843,846
was|847,850
noted|851,856
to|857,859
<EOL>|859,860
have|860,864
a|865,866
thrombosis|867,877
in|878,880
the|881,884
R|885,886
SVC.|887,891
He|892,894
was|895,898
started|899,906
on|907,909
Lovenox|910,917
1|918,919
<EOL>|920,921
mg|921,923
/|923,924
kg|924,926
<EOL>|926,927
BID|927,930
,|930,931
which|932,937
he|938,940
is|941,943
compliant|944,953
with|954,958
.|958,959
Denies|960,966
any|967,970
fever|971,976
,|976,977
nausea|978,984
,|984,985
<EOL>|985,986
emesis|986,992
,|992,993
chills|994,1000
,|1000,1001
weight|1002,1008
loss|1009,1013
,|1013,1014
melena|1015,1021
,|1021,1022
hematochezia|1023,1035
or|1036,1038
hematuria|1039,1048
.|1048,1049
<EOL>|1050,1051
<EOL>|1051,1052
He|1052,1054
comes|1055,1060
after|1061,1066
recent|1067,1073
repeat|1074,1080
staging|1081,1088
(|1089,1090
_|1090,1091
_|1091,1092
_|1092,1093
)|1093,1094
with|1095,1099
torso|1100,1105
CT|1106,1108
<EOL>|1108,1109
scan|1109,1113
demonstrating|1114,1127
no|1128,1130
evidence|1131,1139
of|1140,1142
disease|1143,1150
.|1150,1151
He|1152,1154
is|1155,1157
now|1158,1161
now|1162,1165
taken|1166,1171
<EOL>|1171,1172
to|1172,1174
the|1175,1178
operating|1179,1188
room|1189,1193
for|1194,1197
minimally|1198,1207
invasive|1208,1216
and|1217,1220
possibly|1221,1229
open|1230,1234
<EOL>|1234,1235
radical|1235,1242
distal|1243,1249
gastrectomy|1250,1261
with|1262,1266
lymphadenectomy|1267,1282
.|1282,1283
The|1285,1288
risks|1289,1294
<EOL>|1294,1295
and|1295,1298
benefits|1299,1307
of|1308,1310
surgery|1311,1318
have|1319,1323
been|1324,1328
described|1329,1338
with|1339,1343
the|1344,1347
patient|1348,1355
<EOL>|1355,1356
in|1356,1358
detail|1359,1365
and|1366,1369
are|1370,1373
documented|1374,1384
by|1385,1387
Dr.|1388,1391
_|1392,1393
_|1393,1394
_|1394,1395
in|1396,1398
a|1399,1400
separate|1401,1409
<EOL>|1409,1410
note|1410,1414
.|1414,1415
<EOL>|1415,1416
<EOL>|1417,1418
Past|1440,1444
Medical|1445,1452
History|1453,1460
:|1460,1461
Prostate|1462,1470
cancer|1471,1477
,|1477,1478
Thyroid|1479,1486
nodule|1487,1493
,|1493,1494
<EOL>|1494,1495
Hypothyroid|1495,1506
,|1506,1507
GERD|1508,1512
mild|1513,1517
,|1517,1518
Diverticulosis|1519,1533
on|1534,1536
colonoscopy|1537,1548
_|1549,1550
_|1550,1551
_|1551,1552
<EOL>|1552,1553
anemia|1553,1559
iron|1560,1564
def|1565,1568
.|1568,1569
anemia|1570,1576
which|1577,1582
resolved|1583,1591
and|1592,1595
no|1596,1598
workup|1599,1605
<EOL>|1605,1606
<EOL>|1606,1607
Past|1607,1611
Surgical|1612,1620
History|1621,1628
:|1628,1629
Prostate|1630,1638
cancer|1639,1645
external|1646,1654
beam|1655,1659
_|1660,1661
_|1661,1662
_|1662,1663
,|1663,1664
<EOL>|1664,1665
Achilles|1665,1673
tendon|1674,1680
repair|1681,1687
_|1688,1689
_|1689,1690
_|1690,1691
,|1691,1692
Shattered|1693,1702
right|1703,1708
tibia|1709,1714
and|1715,1718
fibula|1719,1725
,|1725,1726
<EOL>|1726,1727
Tonsillectomy|1727,1740
age|1741,1744
_|1745,1746
_|1746,1747
_|1747,1748
.|1748,1749
<EOL>|1749,1750
<EOL>|1751,1752
:|1766,1767
<EOL>|1767,1768
_|1768,1769
_|1769,1770
_|1770,1771
<EOL>|1771,1772
:|1786,1787
<EOL>|1787,1788
Father|1788,1794
died|1795,1799
at|1800,1802
_|1803,1804
_|1804,1805
_|1805,1806
from|1807,1811
Lymphoma|1812,1820
.|1820,1821
Mother|1822,1828
died|1829,1833
at|1834,1836
_|1837,1838
_|1838,1839
_|1839,1840
with|1841,1845
type|1846,1850
II|1851,1853
<EOL>|1854,1855
DM|1855,1857
,|1857,1858
Dementia|1859,1867
.|1867,1868
<EOL>|1870,1871
<EOL>|1872,1873
VS|1888,1890
:|1890,1891
24|1892,1894
HR|1895,1897
Data|1898,1902
(|1903,1904
last|1904,1908
updated|1909,1916
_|1917,1918
_|1918,1919
_|1919,1920
@|1921,1922
1118|1923,1927
)|1927,1928
<EOL>|1928,1929
Temp|1933,1937
:|1937,1938
98.1|1939,1943
(|1944,1945
Tm|1945,1947
98.9|1948,1952
)|1952,1953
,|1953,1954
BP|1955,1957
:|1957,1958
116|1959,1962
/|1962,1963
73|1963,1965
(|1966,1967
108|1967,1970
-|1970,1971
118|1971,1974
/|1974,1975
59|1975,1977
-|1977,1978
77|1978,1980
)|1980,1981
,|1981,1982
HR|1983,1985
:|1985,1986
79|1987,1989
<EOL>|1990,1991
(|1991,1992
77|1992,1994
-|1994,1995
86|1995,1997
)|1997,1998
,|1998,1999
RR|2000,2002
:|2002,2003
18|2004,2006
(|2007,2008
_|2008,2009
_|2009,2010
_|2010,2011
)|2011,2012
,|2012,2013
O2|2014,2016
sat|2017,2020
:|2020,2021
99|2022,2024
%|2024,2025
(|2026,2027
97|2027,2029
-|2029,2030
99|2030,2032
)|2032,2033
,|2033,2034
O2|2035,2037
delivery|2038,2046
:|2046,2047
Ra|2048,2050
<EOL>|2052,2053
GEN|2053,2056
:|2056,2057
A|2058,2059
&|2059,2060
Ox3|2060,2063
,|2063,2064
NAD|2065,2068
,|2068,2069
resting|2070,2077
comfortably|2078,2089
<EOL>|2090,2091
HEENT|2091,2096
:|2096,2097
NCAT|2098,2102
,|2102,2103
EOMI|2104,2108
,|2108,2109
sclera|2110,2116
anicteric|2117,2126
<EOL>|2126,2127
CV|2127,2129
:|2129,2130
RRR|2131,2134
<EOL>|2134,2135
PULM|2135,2139
:|2139,2140
no|2141,2143
respiratory|2144,2155
distress|2156,2164
<EOL>|2164,2165
ABD|2165,2168
:|2168,2169
soft|2170,2174
,|2174,2175
NT|2176,2178
,|2178,2179
ND|2180,2182
,|2182,2183
no|2184,2186
rebound|2187,2194
or|2195,2197
guarding|2198,2206
<EOL>|2207,2208
EXT|2208,2211
:|2211,2212
warm|2213,2217
,|2217,2218
well|2219,2223
-|2223,2224
perfused|2224,2232
,|2232,2233
no|2234,2236
edema|2237,2242
<EOL>|2243,2244
PSYCH|2244,2249
:|2249,2250
normal|2251,2257
insight|2258,2265
,|2265,2266
memory|2267,2273
,|2273,2274
and|2275,2278
mood|2279,2283
<EOL>|2283,2284
WOUND|2284,2289
(|2289,2290
S|2290,2291
)|2291,2292
:|2292,2293
Incision|2294,2302
c|2303,2304
/|2304,2305
d|2305,2306
/|2306,2307
i|2307,2308
<EOL>|2308,2309
<EOL>|2310,2311
Mr.|2334,2337
_|2338,2339
_|2339,2340
_|2340,2341
is|2342,2344
a|2345,2346
_|2347,2348
_|2348,2349
_|2349,2350
year|2351,2355
old|2356,2359
Male|2360,2364
who|2365,2368
presented|2369,2378
on|2379,2381
_|2382,2383
_|2383,2384
_|2384,2385
for|2386,2389
<EOL>|2390,2391
a|2391,2392
planned|2393,2400
minimally|2401,2410
invasive|2411,2419
and|2420,2423
possibly|2424,2432
open|2433,2437
radical|2438,2445
distal|2446,2452
<EOL>|2453,2454
gastrectomy|2454,2465
with|2466,2470
lymphadenectomy|2471,2486
for|2487,2490
locally|2491,2498
advanced|2499,2507
gastric|2508,2515
<EOL>|2516,2517
carcinoma|2517,2526
after|2527,2532
chemotherapy|2533,2545
.|2545,2546
After|2547,2552
placement|2553,2562
of|2563,2565
the|2566,2569
Right|2570,2575
upper|2576,2581
<EOL>|2582,2583
quadrant|2583,2591
port|2592,2596
,|2596,2597
insufflation|2598,2610
revealed|2611,2619
the|2620,2623
right|2624,2629
upper|2630,2635
quadrant|2636,2644
<EOL>|2645,2646
port|2646,2650
to|2651,2653
be|2654,2656
penetrating|2657,2668
the|2669,2672
omentum|2673,2680
.|2680,2681
It|2682,2684
appeared|2685,2693
to|2694,2696
miss|2697,2701
the|2702,2705
<EOL>|2706,2707
transverse|2707,2717
mesocolon|2718,2727
as|2728,2730
well|2731,2735
as|2736,2738
the|2739,2742
colon|2743,2748
itself|2749,2755
.|2755,2756
During|2757,2763
the|2764,2767
<EOL>|2768,2769
surgery|2769,2776
,|2776,2777
there|2778,2783
were|2784,2788
visually|2789,2797
obvious|2798,2805
peritoneal|2806,2816
deposits|2817,2825
on|2826,2828
all|2829,2832
<EOL>|2833,2834
peritoneal|2834,2844
surfaces|2845,2853
in|2854,2856
all|2857,2860
four|2861,2865
quadrants|2866,2875
,|2875,2876
which|2877,2882
demonstrated|2883,2895
<EOL>|2896,2897
undetected|2897,2907
carcinomatosis|2908,2922
,|2922,2923
poorly|2924,2930
-|2931,2932
differentiated|2932,2946
adenocarcinoma|2947,2961
<EOL>|2962,2963
involving|2963,2972
the|2973,2976
peritoneum|2977,2987
.|2987,2988
For|2989,2992
this|2993,2997
reason|2998,3004
,|3004,3005
the|3006,3009
procedure|3010,3019
was|3020,3023
<EOL>|3024,3025
then|3025,3029
aborted|3030,3037
.|3037,3038
Post-operatively|3039,3055
the|3056,3059
patient|3060,3067
was|3068,3071
taken|3072,3077
to|3078,3080
the|3081,3084
PACU|3085,3089
<EOL>|3090,3091
until|3091,3096
stable|3097,3103
and|3104,3107
then|3108,3112
transferred|3113,3124
to|3125,3127
the|3128,3131
wards|3132,3137
until|3138,3143
stable|3144,3150
to|3151,3153
<EOL>|3154,3155
go|3155,3157
home|3158,3162
.|3162,3163
<EOL>|3164,3165
<EOL>|3165,3166
#|3166,3167
NEURO|3167,3172
:|3172,3173
The|3174,3177
patient|3178,3185
was|3186,3189
alert|3190,3195
and|3196,3199
oriented|3200,3208
throughout|3209,3219
<EOL>|3220,3221
hospitalization|3221,3236
;|3236,3237
pain|3238,3242
was|3243,3246
initially|3247,3256
managed|3257,3264
with|3265,3269
dilaudid|3270,3278
PCA|3279,3282
<EOL>|3283,3284
which|3284,3289
he|3290,3292
was|3293,3296
not|3297,3300
using|3301,3306
and|3307,3310
then|3311,3315
transitioned|3316,3328
to|3329,3331
tramadol|3332,3340
which|3341,3346
<EOL>|3347,3348
he|3348,3350
got|3351,3354
only|3355,3359
one|3360,3363
dose|3364,3368
.|3368,3369
Pain|3370,3374
was|3375,3378
very|3379,3383
well|3384,3388
controlled|3389,3399
.|3399,3400
<EOL>|3400,3401
<EOL>|3401,3402
#|3402,3403
CV|3403,3405
:|3405,3406
The|3407,3410
patient|3411,3418
remained|3419,3427
stable|3428,3434
from|3435,3439
a|3440,3441
cardiovascular|3442,3456
<EOL>|3457,3458
standpoint|3458,3468
;|3468,3469
vital|3470,3475
signs|3476,3481
were|3482,3486
routinely|3487,3496
monitored|3497,3506
.|3506,3507
<EOL>|3509,3510
<EOL>|3510,3511
#|3511,3512
PULMONARY|3512,3521
:|3521,3522
The|3523,3526
patient|3527,3534
remained|3535,3543
stable|3544,3550
from|3551,3555
a|3556,3557
pulmonary|3558,3567
<EOL>|3568,3569
standpoint|3569,3579
;|3579,3580
vital|3581,3586
signs|3587,3592
were|3593,3597
routinely|3598,3607
monitored|3608,3617
.|3617,3618
Good|3619,3623
pulmonary|3624,3633
<EOL>|3634,3635
toilet|3635,3641
,|3641,3642
early|3643,3648
ambulation|3649,3659
and|3660,3663
incentive|3664,3673
spirometry|3674,3684
were|3685,3689
<EOL>|3690,3691
encouraged|3691,3701
throughout|3702,3712
hospitalization|3713,3728
.|3728,3729
<EOL>|3731,3732
<EOL>|3732,3733
#|3733,3734
GI|3734,3736
/|3736,3737
GU|3737,3739
/|3739,3740
FEN|3740,3743
:|3743,3744
Before|3745,3751
the|3752,3755
procedure|3756,3765
started|3766,3773
,|3773,3774
OR|3775,3777
nurse|3778,3783
was|3784,3787
unable|3788,3794
to|3795,3797
<EOL>|3798,3799
pass|3799,3803
Foley|3804,3809
after|3810,3815
attempt|3816,3823
with|3824,3828
standard|3829,3837
and|3838,3841
coude|3842,3847
type|3848,3852
.|3852,3853
PA|3854,3856
<EOL>|3857,3858
_|3858,3859
_|3859,3860
_|3860,3861
,|3861,3862
with|3863,3867
usual|3868,3873
sterile|3874,3881
technique|3882,3891
,|3891,3892
re-attempted|3893,3905
foley|3906,3911
<EOL>|3912,3913
placement|3913,3922
after|3923,3928
10cc|3929,3933
urojet|3934,3940
application|3941,3952
with|3953,3957
_|3958,3959
_|3959,3960
_|3960,3961
and|3962,3965
_|3966,3967
_|3967,3968
_|3968,3969
<EOL>|3970,3971
coude|3971,3976
-|3976,3977
type|3977,3981
catheters|3982,3991
but|3992,3995
was|3996,3999
also|4000,4004
unable|4005,4011
to|4012,4014
get|4015,4018
passed|4019,4025
the|4026,4029
<EOL>|4030,4031
prostate|4031,4039
.|4039,4040
Urology|4041,4048
was|4049,4052
consulted|4053,4062
and|4063,4066
they|4067,4071
performed|4072,4081
a|4082,4083
flexible|4084,4092
<EOL>|4093,4094
cystoscope|4094,4104
demonstrating|4105,4118
a|4119,4120
normal|4121,4127
urethra|4128,4135
.|4135,4136
Using|4137,4142
a|4143,4144
flexible|4145,4153
<EOL>|4154,4155
guidewire|4155,4164
,|4164,4165
cystoscope|4166,4176
was|4177,4180
advanced|4181,4189
into|4190,4194
the|4195,4198
bladder|4199,4206
.|4206,4207
The|4208,4211
scope|4212,4217
<EOL>|4218,4219
was|4219,4222
withdrawn|4223,4232
and|4233,4236
a|4237,4238
_|4239,4240
_|4240,4241
_|4241,4242
council|4243,4250
was|4251,4254
advanced|4255,4263
over|4264,4268
the|4269,4272
wire|4273,4277
,|4277,4278
<EOL>|4279,4280
passed|4280,4286
the|4287,4290
prostate|4291,4299
and|4300,4303
into|4304,4308
the|4309,4312
bladder|4313,4320
.|4320,4321
The|4322,4325
patient|4326,4333
was|4334,4337
<EOL>|4338,4339
discharged|4339,4349
with|4350,4354
the|4355,4358
Foley|4359,4364
in|4365,4367
place|4368,4373
with|4374,4378
instructions|4379,4391
to|4392,4394
<EOL>|4395,4396
follow|4396,4402
-|4402,4403
up|4403,4405
with|4406,4410
urology|4411,4418
as|4419,4421
outpatient|4422,4432
in|4433,4435
5|4436,4437
to|4438,4440
7|4441,4442
days|4443,4447
for|4448,4451
a|4452,4453
<EOL>|4454,4455
voiding|4455,4462
trial|4463,4468
.|4468,4469
No|4470,4472
antibiotics|4473,4484
were|4485,4489
administered|4490,4502
.|4502,4503
The|4504,4507
patient|4508,4515
was|4516,4519
<EOL>|4520,4521
tolerating|4521,4531
a|4532,4533
regular|4534,4541
diet|4542,4546
prior|4547,4552
to|4553,4555
discharge|4556,4565
.|4565,4566
<EOL>|4567,4568
<EOL>|4568,4569
#|4569,4570
ID|4570,4572
:|4572,4573
The|4574,4577
patient|4578,4585
's|4585,4587
fever|4588,4593
curves|4594,4600
were|4601,4605
closely|4606,4613
watched|4614,4621
for|4622,4625
signs|4626,4631
<EOL>|4632,4633
of|4633,4635
infection|4636,4645
,|4645,4646
of|4647,4649
which|4650,4655
there|4656,4661
were|4662,4666
none|4667,4671
.|4671,4672
<EOL>|4674,4675
<EOL>|4675,4676
#|4676,4677
HEME|4677,4681
:|4681,4682
Patient|4683,4690
received|4691,4699
BID|4700,4703
SQH|4704,4707
for|4708,4711
DVT|4712,4715
prophylaxis|4716,4727
,|4727,4728
in|4729,4731
addition|4732,4740
<EOL>|4741,4742
to|4742,4744
encouraging|4745,4756
early|4757,4762
ambulation|4763,4773
and|4774,4777
Venodyne|4778,4786
compression|4787,4798
<EOL>|4799,4800
devices|4800,4807
.|4807,4808
On|4809,4811
POD1|4812,4816
the|4817,4820
patient|4821,4828
was|4829,4832
restarted|4833,4842
on|4843,4845
his|4846,4849
home|4850,4854
<EOL>|4855,4856
enoxaparin|4856,4866
before|4867,4873
discharge|4874,4883
.|4883,4884
<EOL>|4884,4885
<EOL>|4885,4886
#|4886,4887
TRANSITIONAL|4887,4899
ISSUES|4900,4906
<EOL>|4906,4907
-|4907,4908
-|4908,4909
-|4909,4910
-|4910,4911
-|4911,4912
-|4912,4913
-|4913,4914
-|4914,4915
-|4915,4916
-|4916,4917
-|4917,4918
-|4918,4919
-|4919,4920
-|4920,4921
-|4921,4922
-|4922,4923
-|4923,4924
-|4924,4925
-|4925,4926
-|4926,4927
<EOL>|4927,4928
<EOL>|4928,4929
At|4929,4931
the|4932,4935
time|4936,4940
of|4941,4943
discharge|4944,4953
,|4953,4954
the|4955,4958
patient|4959,4966
was|4967,4970
doing|4971,4976
well|4977,4981
,|4981,4982
afebrile|4983,4991
<EOL>|4992,4993
with|4993,4997
stable|4998,5004
vital|5005,5010
signs|5011,5016
.|5016,5017
The|5018,5021
patient|5022,5029
was|5030,5033
tolerating|5034,5044
diet|5045,5049
as|5050,5052
<EOL>|5053,5054
above|5054,5059
per|5060,5063
oral|5064,5068
,|5068,5069
ambulating|5070,5080
,|5080,5081
and|5082,5085
pain|5086,5090
was|5091,5094
well|5095,5099
controlled|5100,5110
.|5110,5111
The|5112,5115
<EOL>|5116,5117
patient|5117,5124
was|5125,5128
discharged|5129,5139
home|5140,5144
with|5145,5149
the|5150,5153
Foley|5154,5159
catheter|5160,5168
with|5169,5173
<EOL>|5174,5175
appropriate|5175,5186
teaching|5187,5195
for|5196,5199
care|5200,5204
.|5204,5205
The|5206,5209
patient|5210,5217
received|5218,5226
discharge|5227,5236
<EOL>|5237,5238
teaching|5238,5246
and|5247,5250
follow|5251,5257
-|5257,5258
up|5258,5260
instructions|5261,5273
with|5274,5278
understanding|5279,5292
<EOL>|5293,5294
verbalized|5294,5304
and|5305,5308
agreement|5309,5318
with|5319,5323
the|5324,5327
discharge|5328,5337
plan|5338,5342
.|5342,5343
<EOL>|5343,5344
<EOL>|5345,5346
Medications|5346,5357
on|5358,5360
Admission|5361,5370
:|5370,5371
<EOL>|5371,5372
Medications|5372,5383
-|5384,5385
Prescription|5386,5398
<EOL>|5398,5399
BIO-THROID|5399,5409
-|5410,5411
Bio-Throid|5412,5422
.|5424,5425
65|5426,5428
mg|5429,5431
.|5431,5432
once|5433,5437
a|5438,5439
day|5440,5443
-|5444,5445
(|5447,5448
Prescribed|5448,5458
by|5459,5461
<EOL>|5462,5463
Other|5463,5468
Provider|5469,5477
)|5477,5478
<EOL>|5478,5479
ENOXAPARIN|5479,5489
-|5490,5491
enoxaparin|5492,5502
120|5503,5506
mg|5507,5509
/|5509,5510
0.8|5510,5513
mL|5514,5516
subcutaneous|5517,5529
syringe|5530,5537
.|5537,5538
120|5539,5542
<EOL>|5543,5544
mg|5544,5546
SC|5547,5549
daily|5550,5555
<EOL>|5555,5556
OMEPRAZOLE|5556,5566
-|5567,5568
omeprazole|5569,5579
20|5580,5582
mg|5583,5585
capsule|5586,5593
,|5593,5594
delayed|5594,5601
release.|5602,5610
1|5611,5612
<EOL>|5613,5614
capsule|5614,5621
(|5621,5622
s|5622,5623
)|5623,5624
by|5625,5627
mouth|5628,5633
twice|5634,5639
daily|5640,5645
<EOL>|5645,5646
UBIQUINOL|5646,5655
-|5656,5657
ubiquinol|5658,5667
.|5669,5670
(|5671,5672
100|5672,5675
mg|5676,5678
)|5678,5679
2|5680,5681
tabs|5682,5686
mouth|5687,5692
twice|5693,5698
a|5699,5700
day|5701,5704
-|5705,5706
<EOL>|5708,5709
(|5709,5710
Prescribed|5710,5720
by|5721,5723
Other|5724,5729
Provider|5730,5738
)|5738,5739
<EOL>|5739,5740
<EOL>|5741,5742
Medications|5742,5753
-|5754,5755
OTC|5756,5759
<EOL>|5759,5760
FERROUS|5760,5767
SULFATE|5768,5775
-|5776,5777
ferrous|5778,5785
sulfate|5786,5793
325|5794,5797
mg|5798,5800
(|5801,5802
65|5802,5804
mg|5805,5807
iron|5808,5812
)|5812,5813
tablet.|5814,5821
1|5822,5823
<EOL>|5824,5825
tablet|5825,5831
(|5831,5832
s|5832,5833
)|5833,5834
by|5835,5837
mouth|5838,5843
twice|5844,5849
a|5850,5851
day|5852,5855
-|5856,5857
(|5859,5860
Prescribed|5860,5870
by|5871,5873
Other|5874,5879
Provider|5880,5888
)|5888,5889
<EOL>|5889,5890
LACTOBACILLUS|5890,5903
COMBINATION|5904,5915
NO|5916,5918
.4|5918,5920
[|5921,5922
PROBIOTIC|5922,5931
]|5931,5932
-|5933,5934
Dosage|5935,5941
uncertain|5942,5951
-|5952,5953
<EOL>|5955,5956
(|5956,5957
Prescribed|5957,5967
by|5968,5970
Other|5971,5976
Provider|5977,5985
;|5985,5986
daily|5987,5992
)|5992,5993
<EOL>|5993,5994
<EOL>|5995,5996
Discharge|5996,6005
Medications|6006,6017
:|6017,6018
<EOL>|6018,6019
1.|6019,6021
Acetaminophen|6023,6036
1000|6037,6041
mg|6042,6044
PO|6045,6047
TID|6048,6051
<EOL>|6053,6054
2.|6054,6056
Docusate|6058,6066
Sodium|6067,6073
100|6074,6077
mg|6078,6080
PO|6081,6083
BID|6084,6087
<EOL>|6089,6090
3.|6090,6092
Senna|6094,6099
8.6|6100,6103
mg|6104,6106
PO|6107,6109
BID|6110,6113
:|6113,6114
PRN|6114,6117
Constipation|6118,6130
-|6131,6132
First|6133,6138
Line|6139,6143
<EOL>|6145,6146
4.|6146,6148
TraMADol|6150,6158
50|6159,6161
mg|6162,6164
PO|6165,6167
Q6H|6168,6171
:|6171,6172
PRN|6172,6175
Pain|6176,6180
-|6181,6182
Moderate|6183,6191
<EOL>|6192,6193
This|6193,6197
medication|6198,6208
is|6209,6211
a|6212,6213
low|6214,6217
dose|6218,6222
narcotic|6223,6231
and|6232,6235
may|6236,6239
cause|6240,6245
<EOL>|6246,6247
constipation|6247,6259
.|6259,6260
<EOL>|6261,6262
RX|6262,6264
*|6265,6266
tramadol|6266,6274
50|6275,6277
mg|6278,6280
1|6281,6282
(|6283,6284
One|6284,6287
)|6287,6288
tablet|6289,6295
(|6295,6296
s|6296,6297
)|6297,6298
by|6299,6301
mouth|6302,6307
every|6308,6313
six|6314,6317
(|6318,6319
6|6319,6320
)|6320,6321
<EOL>|6322,6323
hours|6323,6328
Disp|6329,6333
#|6334,6335
*|6335,6336
20|6336,6338
Tablet|6339,6345
Refills|6346,6353
:|6353,6354
*|6354,6355
0|6355,6356
<EOL>|6357,6358
5.|6358,6360
Enoxaparin|6362,6372
Sodium|6373,6379
120|6380,6383
mg|6384,6386
SC|6387,6389
DAILY|6390,6395
<EOL>|6397,6398
<EOL>|6398,6399
<EOL>|6400,6401
Discharge|6401,6410
Disposition|6411,6422
:|6422,6423
<EOL>|6423,6424
Home|6424,6428
<EOL>|6428,6429
<EOL>|6430,6431
Discharge|6431,6440
Diagnosis|6441,6450
:|6450,6451
<EOL>|6451,6452
Metastatic|6452,6462
gastric|6463,6470
cancer|6471,6477
(|6478,6479
stage|6479,6484
IV|6485,6487
[|6488,6489
T3N2M1|6489,6495
]|6495,6496
)|6496,6497
<EOL>|6497,6498
Urethral|6498,6506
stricture|6507,6516
<EOL>|6516,6517
<EOL>|6518,6519
Mental|6540,6546
Status|6547,6553
:|6553,6554
Clear|6555,6560
and|6561,6564
coherent|6565,6573
.|6573,6574
<EOL>|6574,6575
Level|6575,6580
of|6581,6583
Consciousness|6584,6597
:|6597,6598
Alert|6599,6604
and|6605,6608
interactive|6609,6620
.|6620,6621
<EOL>|6621,6622
Activity|6622,6630
Status|6631,6637
:|6637,6638
Ambulatory|6639,6649
-|6650,6651
Independent|6652,6663
.|6663,6664
<EOL>|6664,6665
<EOL>|6665,6666
<EOL>|6667,6668
Dear|6692,6696
Mr.|6697,6700
_|6701,6702
_|6702,6703
_|6703,6704
,|6704,6705
<EOL>|6705,6706
<EOL>|6706,6707
It|6707,6709
was|6710,6713
a|6714,6715
pleasure|6716,6724
taking|6725,6731
care|6732,6736
of|6737,6739
you|6740,6743
here|6744,6748
at|6749,6751
_|6752,6753
_|6753,6754
_|6754,6755
<EOL>|6756,6757
_|6757,6758
_|6758,6759
_|6759,6760
.|6760,6761
You|6762,6765
were|6766,6770
admitted|6771,6779
to|6780,6782
our|6783,6786
hospital|6787,6795
for|6796,6799
<EOL>|6800,6801
gastric|6801,6808
cancer|6809,6815
.|6815,6816
You|6817,6820
had|6821,6824
an|6825,6827
attempted|6828,6837
Robot|6838,6843
-|6843,6844
assisted|6844,6852
laparoscopic|6853,6865
<EOL>|6866,6867
partial|6867,6874
gastrectomy|6875,6886
and|6887,6890
gastroscopy|6891,6902
on|6903,6905
_|6906,6907
_|6907,6908
_|6908,6909
without|6910,6917
<EOL>|6918,6919
complications|6919,6932
.|6932,6933
You|6934,6937
tolerated|6938,6947
the|6948,6951
procedure|6952,6961
well|6962,6966
and|6967,6970
are|6971,6974
<EOL>|6975,6976
ambulating|6976,6986
,|6986,6987
stooling|6988,6996
,|6996,6997
tolerating|6998,7008
a|7009,7010
regular|7011,7018
diet|7019,7023
,|7023,7024
and|7025,7028
your|7029,7033
pain|7034,7038
<EOL>|7039,7040
is|7040,7042
controlled|7043,7053
by|7054,7056
pain|7057,7061
medications|7062,7073
by|7074,7076
mouth|7077,7082
.|7082,7083
You|7084,7087
are|7088,7091
now|7092,7095
ready|7096,7101
to|7102,7104
<EOL>|7105,7106
be|7106,7108
discharged|7109,7119
to|7120,7122
home|7123,7127
.|7127,7128
Please|7129,7135
follow|7136,7142
the|7143,7146
recommendations|7147,7162
below|7163,7168
<EOL>|7169,7170
to|7170,7172
ensure|7173,7179
a|7180,7181
speedy|7182,7188
and|7189,7192
uneventful|7193,7203
recovery|7204,7212
.|7212,7213
<EOL>|7214,7215
<EOL>|7215,7216
ACTIVITY|7216,7224
:|7224,7225
<EOL>|7225,7226
-|7226,7227
Do|7228,7230
not|7231,7234
drive|7235,7240
until|7241,7246
you|7247,7250
have|7251,7255
stopped|7256,7263
taking|7264,7270
pain|7271,7275
medicine|7276,7284
and|7285,7288
<EOL>|7289,7290
feel|7290,7294
you|7295,7298
could|7299,7304
respond|7305,7312
in|7313,7315
an|7316,7318
emergency|7319,7328
.|7328,7329
<EOL>|7329,7330
-|7330,7331
You|7332,7335
may|7336,7339
climb|7340,7345
stairs|7346,7352
.|7352,7353
You|7354,7357
should|7358,7364
continue|7365,7373
to|7374,7376
walk|7377,7381
several|7382,7389
<EOL>|7390,7391
times|7391,7396
a|7397,7398
day|7399,7402
.|7402,7403
<EOL>|7404,7405
-|7405,7406
You|7407,7410
may|7411,7414
go|7415,7417
outside|7418,7425
,|7425,7426
but|7427,7430
avoid|7431,7436
traveling|7437,7446
long|7447,7451
distances|7452,7461
until|7462,7467
<EOL>|7468,7469
you|7469,7472
see|7473,7476
your|7477,7481
surgeon|7482,7489
at|7490,7492
your|7493,7497
next|7498,7502
visit|7503,7508
.|7508,7509
<EOL>|7510,7511
-|7511,7512
You|7513,7516
may|7517,7520
start|7521,7526
some|7527,7531
light|7532,7537
exercise|7538,7546
when|7547,7551
you|7552,7555
feel|7556,7560
comfortable|7561,7572
.|7572,7573
<EOL>|7574,7575
Slowly|7575,7581
increase|7582,7590
your|7591,7595
activity|7596,7604
back|7605,7609
to|7610,7612
your|7613,7617
baseline|7618,7626
as|7627,7629
<EOL>|7630,7631
tolerated|7631,7640
.|7640,7641
<EOL>|7641,7642
-|7642,7643
Heavy|7644,7649
exercise|7650,7658
may|7659,7662
be|7663,7665
started|7666,7673
after|7674,7679
6|7680,7681
weeks|7682,7687
,|7687,7688
but|7689,7692
use|7693,7696
common|7697,7703
<EOL>|7704,7705
sense|7705,7710
and|7711,7714
go|7715,7717
slowly|7718,7724
at|7725,7727
first|7728,7733
.|7733,7734
<EOL>|7735,7736
-|7736,7737
No|7738,7740
heavy|7741,7746
lifting|7747,7754
(|7755,7756
10|7756,7758
pounds|7759,7765
or|7766,7768
more|7769,7773
)|7773,7774
until|7775,7780
cleared|7781,7788
by|7789,7791
your|7792,7796
<EOL>|7797,7798
surgeon|7798,7805
,|7805,7806
usually|7807,7814
about|7815,7820
6|7821,7822
weeks|7823,7828
.|7828,7829
<EOL>|7830,7831
-|7831,7832
You|7833,7836
may|7837,7840
resume|7841,7847
sexual|7848,7854
activity|7855,7863
unless|7864,7870
your|7871,7875
doctor|7876,7882
has|7883,7886
told|7887,7891
you|7892,7895
<EOL>|7896,7897
otherwise|7897,7906
.|7906,7907
<EOL>|7907,7908
<EOL>|7908,7909
HOW|7909,7912
YOU|7913,7916
MAY|7917,7920
FEEL|7921,7925
:|7925,7926
<EOL>|7927,7928
-|7928,7929
You|7930,7933
may|7934,7937
feel|7938,7942
weak|7943,7947
or|7948,7950
"|7951,7952
washed|7952,7958
out|7959,7962
"|7962,7963
for|7964,7967
6|7968,7969
weeks|7970,7975
.|7975,7976
You|7977,7980
might|7981,7986
want|7987,7991
<EOL>|7992,7993
to|7993,7995
nap|7996,7999
often|8000,8005
.|8005,8006
Simple|8007,8013
tasks|8014,8019
may|8020,8023
exhaust|8024,8031
you|8032,8035
.|8035,8036
<EOL>|8036,8037
-|8037,8038
You|8039,8042
may|8043,8046
have|8047,8051
a|8052,8053
sore|8054,8058
throat|8059,8065
because|8066,8073
of|8074,8076
a|8077,8078
tube|8079,8083
that|8084,8088
was|8089,8092
in|8093,8095
your|8096,8100
<EOL>|8101,8102
throat|8102,8108
during|8109,8115
the|8116,8119
surgery|8120,8127
.|8127,8128
<EOL>|8128,8129
<EOL>|8129,8130
YOUR|8130,8134
BOWELS|8135,8141
:|8141,8142
<EOL>|8142,8143
-|8143,8144
Constipation|8145,8157
is|8158,8160
a|8161,8162
common|8163,8169
side|8170,8174
effect|8175,8181
of|8182,8184
narcotic|8185,8193
pain|8194,8198
medicine|8199,8207
<EOL>|8208,8209
such|8209,8213
as|8214,8216
oxycodone|8217,8226
.|8226,8227
If|8228,8230
needed|8231,8237
,|8237,8238
you|8239,8242
may|8243,8246
take|8247,8251
a|8252,8253
stool|8254,8259
softener|8260,8268
<EOL>|8269,8270
(|8270,8271
such|8271,8275
as|8276,8278
Colace|8279,8285
,|8285,8286
one|8287,8290
capsule|8291,8298
)|8298,8299
or|8300,8302
gentle|8303,8309
laxative|8310,8318
(|8319,8320
such|8320,8324
as|8325,8327
milk|8328,8332
<EOL>|8333,8334
of|8334,8336
magnesia|8337,8345
,|8345,8346
1|8347,8348
tbs|8349,8352
)|8352,8353
twice|8354,8359
a|8360,8361
day|8362,8365
.|8365,8366
You|8367,8370
can|8371,8374
get|8375,8378
both|8379,8383
of|8384,8386
these|8387,8392
<EOL>|8393,8394
medicines|8394,8403
without|8404,8411
a|8412,8413
prescription|8414,8426
.|8426,8427
<EOL>|8427,8428
-|8428,8429
If|8430,8432
you|8433,8436
go|8437,8439
48|8440,8442
hours|8443,8448
without|8449,8456
a|8457,8458
bowel|8459,8464
movement|8465,8473
,|8473,8474
or|8475,8477
have|8478,8482
pain|8483,8487
<EOL>|8488,8489
moving|8489,8495
the|8496,8499
bowels|8500,8506
,|8506,8507
call|8508,8512
your|8513,8517
surgeon|8518,8525
.|8525,8526
<EOL>|8526,8527
-|8527,8528
After|8529,8534
some|8535,8539
operations|8540,8550
,|8550,8551
diarrhea|8552,8560
can|8561,8564
occur|8565,8570
.|8570,8571
If|8572,8574
you|8575,8578
get|8579,8582
<EOL>|8583,8584
diarrhea|8584,8592
,|8592,8593
do|8594,8596
n't|8596,8599
take|8600,8604
anti-diarrhea|8605,8618
medicines|8619,8628
.|8628,8629
Drink|8630,8635
plenty|8636,8642
of|8643,8645
<EOL>|8646,8647
fluids|8647,8653
and|8654,8657
see|8658,8661
if|8662,8664
it|8665,8667
goes|8668,8672
away|8673,8677
.|8677,8678
If|8679,8681
it|8682,8684
does|8685,8689
not|8690,8693
go|8694,8696
away|8697,8701
,|8701,8702
or|8703,8705
is|8706,8708
<EOL>|8709,8710
severe|8710,8716
and|8717,8720
you|8721,8724
feel|8725,8729
ill|8730,8733
,|8733,8734
please|8735,8741
call|8742,8746
your|8747,8751
surgeon|8752,8759
.|8759,8760
<EOL>|8760,8761
<EOL>|8761,8762
PAIN|8762,8766
MANAGEMENT|8767,8777
:|8777,8778
<EOL>|8778,8779
-|8779,8780
You|8781,8784
are|8785,8788
being|8789,8794
discharged|8795,8805
with|8806,8810
a|8811,8812
prescription|8813,8825
for|8826,8829
*|8830,8831
*|8831,8832
oxycodone|8832,8841
<EOL>|8842,8843
for|8843,8846
pain|8847,8851
control|8852,8859
.|8859,8860
You|8861,8864
may|8865,8868
take|8869,8873
Tylenol|8874,8881
as|8882,8884
directed|8885,8893
,|8893,8894
not|8895,8898
to|8899,8901
<EOL>|8902,8903
exceed|8903,8909
3500mg|8910,8916
in|8917,8919
24|8920,8922
hours|8923,8928
.|8928,8929
Take|8930,8934
regularly|8935,8944
for|8945,8948
a|8949,8950
few|8951,8954
days|8955,8959
after|8960,8965
<EOL>|8966,8967
surgery|8967,8974
but|8975,8978
you|8979,8982
may|8983,8986
skip|8987,8991
a|8992,8993
dose|8994,8998
or|8999,9001
increase|9002,9010
time|9011,9015
between|9016,9023
doses|9024,9029
<EOL>|9030,9031
if|9031,9033
you|9034,9037
are|9038,9041
not|9042,9045
having|9046,9052
pain|9053,9057
until|9058,9063
you|9064,9067
no|9068,9070
longer|9071,9077
need|9078,9082
it|9083,9085
.|9085,9086
You|9087,9090
may|9091,9094
<EOL>|9095,9096
take|9096,9100
the|9101,9104
oxycodone|9105,9114
for|9115,9118
moderate|9119,9127
and|9128,9131
severe|9132,9138
pain|9139,9143
not|9144,9147
controlled|9148,9158
<EOL>|9159,9160
by|9160,9162
the|9163,9166
Tylenol|9167,9174
.|9174,9175
You|9176,9179
may|9180,9183
take|9184,9188
a|9189,9190
stool|9191,9196
softener|9197,9205
while|9206,9211
on|9212,9214
narcotics|9215,9224
<EOL>|9225,9226
to|9226,9228
help|9229,9233
prevent|9234,9241
the|9242,9245
constipation|9246,9258
that|9259,9263
they|9264,9268
may|9269,9272
cause|9273,9278
.|9278,9279
Slowly|9280,9286
<EOL>|9287,9288
wean|9288,9292
off|9293,9296
these|9297,9302
medications|9303,9314
as|9315,9317
tolerated|9318,9327
.|9327,9328
<EOL>|9329,9330
-|9330,9331
Your|9332,9336
pain|9337,9341
should|9342,9348
get|9349,9352
better|9353,9359
day|9360,9363
by|9364,9366
day|9367,9370
.|9370,9371
If|9372,9374
you|9375,9378
find|9379,9383
the|9384,9387
pain|9388,9392
<EOL>|9393,9394
is|9394,9396
getting|9397,9404
worse|9405,9410
instead|9411,9418
of|9419,9421
better|9422,9428
,|9428,9429
please|9430,9436
contact|9437,9444
your|9445,9449
surgeon|9450,9457
.|9457,9458
<EOL>|9458,9459
<EOL>|9459,9460
If|9460,9462
you|9463,9466
experience|9467,9477
any|9478,9481
of|9482,9484
the|9485,9488
following|9489,9498
,|9498,9499
please|9500,9506
contact|9507,9514
your|9515,9519
<EOL>|9520,9521
surgeon|9521,9528
:|9528,9529
<EOL>|9530,9531
-|9531,9532
sharp|9533,9538
pain|9539,9543
or|9544,9546
any|9547,9550
severe|9551,9557
pain|9558,9562
that|9563,9567
lasts|9568,9573
several|9574,9581
hours|9582,9587
<EOL>|9587,9588
-|9588,9589
chest|9590,9595
pain|9596,9600
,|9600,9601
pressure|9602,9610
,|9610,9611
squeezing|9612,9621
,|9621,9622
or|9623,9625
tightness|9626,9635
<EOL>|9635,9636
-|9636,9637
cough|9638,9643
,|9643,9644
shortness|9645,9654
of|9655,9657
breath|9658,9664
,|9664,9665
wheezing|9666,9674
<EOL>|9674,9675
-|9675,9676
pain|9677,9681
that|9682,9686
is|9687,9689
getting|9690,9697
worse|9698,9703
over|9704,9708
time|9709,9713
or|9714,9716
pain|9717,9721
with|9722,9726
fever|9727,9732
<EOL>|9732,9733
-|9733,9734
shaking|9735,9742
chills|9743,9749
,|9749,9750
fever|9751,9756
of|9757,9759
more|9760,9764
than|9765,9769
101|9770,9773
<EOL>|9773,9774
-|9774,9775
a|9776,9777
drastic|9778,9785
change|9786,9792
in|9793,9795
nature|9796,9802
or|9803,9805
quality|9806,9813
of|9814,9816
your|9817,9821
pain|9822,9826
<EOL>|9826,9827
-|9827,9828
nausea|9829,9835
and|9836,9839
vomiting|9840,9848
,|9848,9849
inability|9850,9859
to|9860,9862
tolerate|9863,9871
fluids|9872,9878
,|9878,9879
food|9880,9884
,|9884,9885
or|9886,9888
<EOL>|9889,9890
your|9890,9894
medications|9895,9906
<EOL>|9906,9907
-|9907,9908
if|9909,9911
you|9912,9915
are|9916,9919
getting|9920,9927
dehydrated|9928,9938
(|9939,9940
dry|9940,9943
mouth|9944,9949
,|9949,9950
rapid|9951,9956
heart|9957,9962
beat|9963,9967
,|9967,9968
<EOL>|9969,9970
feeling|9970,9977
dizzy|9978,9983
or|9984,9986
faint|9987,9992
especially|9993,10003
while|10004,10009
standing|10010,10018
)|10018,10019
<EOL>|10019,10020
-|10020,10021
any|10021,10024
change|10025,10031
in|10032,10034
your|10035,10039
symptoms|10040,10048
or|10049,10051
any|10052,10055
symptoms|10056,10064
that|10065,10069
concern|10070,10077
you|10078,10081
<EOL>|10081,10082
<EOL>|10082,10083
Additional|10083,10093
:|10093,10094
<EOL>|10095,10096
*|10096,10097
-|10097,10098
pain|10099,10103
that|10104,10108
is|10109,10111
getting|10112,10119
worse|10120,10125
over|10126,10130
time|10131,10135
,|10135,10136
or|10137,10139
going|10140,10145
to|10146,10148
your|10149,10153
chest|10154,10159
<EOL>|10160,10161
or|10161,10163
back|10164,10168
<EOL>|10168,10169
*|10169,10170
-|10170,10171
urinary|10172,10179
:|10179,10180
burning|10182,10189
or|10190,10192
blood|10193,10198
in|10199,10201
your|10202,10206
urine|10207,10212
or|10213,10215
the|10216,10219
inability|10220,10229
to|10230,10232
<EOL>|10233,10234
urinate|10234,10241
<EOL>|10241,10242
<EOL>|10242,10243
-|10256,10257
Take|10258,10262
all|10263,10266
the|10267,10270
medicines|10271,10280
you|10281,10284
were|10285,10289
on|10290,10292
before|10293,10299
the|10300,10303
operation|10304,10313
just|10314,10318
<EOL>|10319,10320
as|10320,10322
you|10323,10326
did|10327,10330
before|10331,10337
,|10337,10338
unless|10339,10345
you|10346,10349
have|10350,10354
been|10355,10359
told|10360,10364
differently|10365,10376
.|10376,10377
<EOL>|10377,10378
-|10378,10379
If|10380,10382
you|10383,10386
have|10387,10391
any|10392,10395
questions|10396,10405
about|10406,10411
what|10412,10416
medicine|10417,10425
to|10426,10428
take|10429,10433
or|10434,10436
not|10437,10440
<EOL>|10441,10442
to|10442,10444
take|10445,10449
,|10449,10450
please|10451,10457
call|10458,10462
your|10463,10467
surgeon|10468,10475
.|10475,10476
<EOL>|10477,10478
<EOL>|10478,10479
WOUND|10479,10484
CARE|10485,10489
:|10489,10490
<EOL>|10491,10492
-|10492,10493
dressing|10494,10502
removal|10503,10510
:|10510,10511
<EOL>|10511,10512
-|10512,10513
You|10514,10517
may|10518,10521
remove|10522,10528
your|10529,10533
dressings|10534,10543
tomorrow|10544,10552
_|10553,10554
_|10554,10555
_|10555,10556
and|10557,10560
shower|10561,10567
that|10568,10572
<EOL>|10573,10574
same|10574,10578
day|10579,10582
with|10583,10587
any|10588,10591
bandage|10592,10599
strips|10600,10606
that|10607,10611
may|10612,10615
be|10616,10618
covering|10619,10627
your|10628,10632
<EOL>|10633,10634
wound.|10634,10640
Do|10641,10643
not|10644,10647
scrub|10648,10653
and|10654,10657
do|10658,10660
not|10661,10664
soak|10665,10669
or|10670,10672
swim|10673,10677
,|10677,10678
and|10679,10682
pat|10683,10686
the|10687,10690
<EOL>|10691,10692
incision|10692,10700
dry|10701,10704
.|10704,10705
If|10706,10708
you|10709,10712
have|10713,10717
steri|10718,10723
strips|10724,10730
,|10730,10731
they|10732,10736
will|10737,10741
fall|10742,10746
off|10747,10750
by|10751,10753
<EOL>|10754,10755
themselves|10755,10765
in|10766,10768
_|10769,10770
_|10770,10771
_|10771,10772
weeks|10773,10778
.|10778,10779
If|10780,10782
any|10783,10786
are|10787,10790
still|10791,10796
on|10797,10799
in|10800,10802
two|10803,10806
weeks|10807,10812
and|10813,10816
<EOL>|10817,10818
the|10818,10821
edges|10822,10827
are|10828,10831
curling|10832,10839
up|10840,10842
,|10842,10843
you|10844,10847
may|10848,10851
carefully|10852,10861
peel|10862,10866
them|10867,10871
off|10872,10875
.|10875,10876
<EOL>|10876,10877
Do|10878,10880
not|10881,10884
take|10885,10889
baths|10890,10895
,|10895,10896
soak|10897,10901
,|10901,10902
or|10903,10905
swim|10906,10910
for|10911,10914
6|10915,10916
weeks|10917,10922
after|10923,10928
surgery|10929,10936
<EOL>|10937,10938
unless|10938,10944
told|10945,10949
otherwise|10950,10959
by|10960,10962
your|10963,10967
surgical|10968,10976
team|10977,10981
.|10981,10982
<EOL>|10983,10984
-|10984,10985
Notify|10985,10991
your|10992,10996
surgeon|10997,11004
is|11005,11007
you|11008,11011
notice|11012,11018
abnormal|11019,11027
(|11028,11029
foul|11029,11033
smelling|11034,11042
,|11042,11043
<EOL>|11044,11045
bloody|11045,11051
,|11051,11052
pus|11053,11056
,|11056,11057
etc|11058,11061
)|11061,11062
or|11063,11065
increased|11066,11075
drainage|11076,11084
from|11085,11089
your|11090,11094
incision|11095,11103
site|11104,11108
,|11108,11109
<EOL>|11110,11111
opening|11111,11118
of|11119,11121
your|11122,11126
incision|11127,11135
,|11135,11136
or|11137,11139
increased|11140,11149
pain|11150,11154
or|11155,11157
bruising|11158,11166
.|11166,11167
Watch|11168,11173
<EOL>|11174,11175
for|11175,11178
signs|11179,11184
of|11185,11187
infection|11188,11197
such|11198,11202
as|11203,11205
redness|11206,11213
,|11213,11214
streaking|11215,11224
of|11225,11227
your|11228,11232
skin|11233,11237
,|11237,11238
<EOL>|11239,11240
swelling|11240,11248
,|11248,11249
increased|11250,11259
pain|11260,11264
,|11264,11265
or|11266,11268
increased|11269,11278
drainage|11279,11287
.|11287,11288
<EOL>|11289,11290
<EOL>|11290,11291
Please|11291,11297
call|11298,11302
with|11303,11307
any|11308,11311
questions|11312,11321
or|11322,11324
concerns|11325,11333
.|11333,11334
Thank|11335,11340
you|11341,11344
for|11345,11348
<EOL>|11349,11350
allowing|11350,11358
us|11359,11361
to|11362,11364
participate|11365,11376
in|11377,11379
your|11380,11384
care|11385,11389
.|11389,11390
We|11391,11393
hope|11394,11398
you|11399,11402
have|11403,11407
a|11408,11409
<EOL>|11410,11411
quick|11411,11416
return|11417,11423
to|11424,11426
your|11427,11431
usual|11432,11437
life|11438,11442
and|11443,11446
activities|11447,11457
.|11457,11458
<EOL>|11458,11459
<EOL>|11459,11460
Home|11460,11464
with|11465,11469
_|11470,11471
_|11471,11472
_|11472,11473
:|11473,11474
<EOL>|11474,11475
You|11475,11478
had|11479,11482
a|11483,11484
Foley|11485,11490
catheter|11491,11499
in|11500,11502
your|11503,11507
bladder|11508,11515
placed|11516,11522
by|11523,11525
urology|11526,11533
on|11534,11536
<EOL>|11537,11538
the|11538,11541
day|11542,11545
of|11546,11548
your|11549,11553
surgery|11554,11561
after|11562,11567
difficulty|11568,11578
trying|11579,11585
to|11586,11588
place|11589,11594
it|11595,11597
.|11597,11598
<EOL>|11598,11599
You|11599,11602
will|11603,11607
keep|11608,11612
the|11613,11616
catheter|11617,11625
until|11626,11631
your|11632,11636
appointment|11637,11648
with|11649,11653
Urology|11654,11661
<EOL>|11662,11663
in|11663,11665
5|11666,11667
days|11668,11672
(|11673,11674
please|11674,11680
call|11681,11685
the|11686,11689
number|11690,11696
below|11697,11702
to|11703,11705
schedule|11706,11714
your|11715,11719
<EOL>|11720,11721
appointment|11721,11732
)|11732,11733
,|11733,11734
who|11735,11738
will|11739,11743
decide|11744,11750
if|11751,11753
you|11754,11757
need|11758,11762
it|11763,11765
longer|11766,11772
or|11773,11775
attempt|11776,11783
<EOL>|11784,11785
to|11785,11787
remove|11788,11794
it|11795,11797
and|11798,11801
see|11802,11805
if|11806,11808
you|11809,11812
are|11813,11816
able|11817,11821
to|11822,11824
void|11825,11829
.|11829,11830
<EOL>|11830,11831
Empty|11832,11837
the|11838,11841
bag|11842,11845
as|11846,11848
needed|11849,11855
and|11856,11859
as|11860,11862
shown|11863,11868
to|11869,11871
you|11872,11875
by|11876,11878
nursing|11879,11886
staff|11887,11892
.|11892,11893
<EOL>|11894,11895
You|11895,11898
will|11899,11903
be|11904,11906
given|11907,11912
a|11913,11914
leg|11915,11918
bag|11919,11922
before|11923,11929
your|11930,11934
discharge|11935,11944
,|11944,11945
that|11946,11950
you|11951,11954
may|11955,11958
<EOL>|11959,11960
use|11960,11963
for|11964,11967
short|11968,11973
trips|11974,11979
.|11979,11980
This|11981,11985
is|11986,11988
a|11989,11990
smaller|11991,11998
bag|11999,12002
that|12003,12007
straps|12008,12014
to|12015,12017
your|12018,12022
<EOL>|12023,12024
leg|12024,12027
,|12027,12028
to|12029,12031
take|12032,12036
home|12037,12041
and|12042,12045
wear|12046,12050
if|12051,12053
you|12054,12057
are|12058,12061
traveling|12062,12071
outside|12072,12079
your|12080,12084
<EOL>|12085,12086
home|12086,12090
.|12090,12091
This|12092,12096
holds|12097,12102
a|12103,12104
smaller|12105,12112
amount|12113,12119
than|12120,12124
the|12125,12128
bag|12129,12132
you|12133,12136
have|12137,12141
now|12142,12145
,|12145,12146
so|12147,12149
<EOL>|12150,12151
it|12151,12153
needs|12154,12159
to|12160,12162
be|12163,12165
emptied|12166,12173
more|12174,12178
often|12179,12184
.|12184,12185
Some|12186,12190
people|12191,12197
find|12198,12202
it|12203,12205
easier|12206,12212
to|12213,12215
<EOL>|12216,12217
use|12217,12220
the|12221,12224
larger|12225,12231
bad|12232,12235
when|12236,12240
they|12241,12245
are|12246,12249
at|12250,12252
home|12253,12257
or|12258,12260
carry|12261,12266
it|12267,12269
with|12270,12274
them|12275,12279
.|12279,12280
<EOL>|12281,12282
<EOL>|12282,12283
-|12283,12284
-|12284,12285
Your|12286,12290
_|12291,12292
_|12292,12293
_|12293,12294
Care|12295,12299
Team|12300,12304
<EOL>|12304,12305
<EOL>|12306,12307
Followup|12307,12315
Instructions|12316,12328
:|12328,12329
<EOL>|12329,12330
_|12330,12331
_|12331,12332
_|12332,12333
<EOL>|12333,12334

