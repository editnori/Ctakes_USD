 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|45,54|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|45,54|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|45,59|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|79,88|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|79,88|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|79,88|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|79,88|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|79,88|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|79,93|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|111,116|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|111,116|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|111,116|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|135,138|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|135,138|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|135,138|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|135,138|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|135,138|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|146,153|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|146,153|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Event|Event|SIMPLE_SEGMENT|155,162|false|false|false|||SURGERY
Finding|Finding|SIMPLE_SEGMENT|155,162|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|SURGERY
Finding|Functional Concept|SIMPLE_SEGMENT|155,162|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|SURGERY
Finding|Idea or Concept|SIMPLE_SEGMENT|155,162|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|SURGERY
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|155,162|false|false|false|C0543467|Operative Surgical Procedures|SURGERY
Drug|Organic Chemical|Allergies|177,184|false|false|false|C0009214|codeine|Codeine
Drug|Pharmacologic Substance|Allergies|177,184|false|false|false|C0009214|codeine|Codeine
Drug|Antibiotic|Allergies|187,196|false|false|false|C0591132|Augmentin|Augmentin
Drug|Organic Chemical|Allergies|187,196|false|false|false|C0591132|Augmentin|Augmentin
Drug|Organic Chemical|Allergies|199,206|false|false|false|C0723778|Topamax|Topamax
Drug|Pharmacologic Substance|Allergies|199,206|false|false|false|C0723778|Topamax|Topamax
Event|Event|Allergies|209,218|false|false|false|||Attending
Finding|Functional Concept|Allergies|209,218|false|false|false|C1999232|Attending (action)|Attending
Attribute|Clinical Attribute|Allergies|230,239|false|false|false|C3864418||Complaint
Event|Event|Allergies|230,239|false|false|false|||Complaint
Finding|Finding|Allergies|230,239|false|false|false|C5441521|Complaint (finding)|Complaint
Finding|Functional Concept|Allergies|241,245|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Allergies|241,252|false|false|false|C0222601|Left breast|left breast
Finding|Sign or Symptom|Allergies|241,261|false|false|false|C2127345|localized swelling in left breast|left breast swelling
Anatomy|Body Part, Organ, or Organ Component|Allergies|246,252|false|false|false|C0006141|Breast|breast
Disorder|Neoplastic Process|Allergies|246,252|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|breast
Event|Event|Allergies|246,252|false|false|false|||breast
Finding|Finding|Allergies|246,252|false|false|false|C0567499|Breast problem|breast
Procedure|Therapeutic or Preventive Procedure|Allergies|246,252|false|false|false|C0191838|Procedures on breast|breast
Finding|Finding|Allergies|246,261|false|false|false|C0006152|Swelling of breast|breast swelling
Event|Event|Allergies|253,261|false|false|false|||swelling
Finding|Finding|Allergies|253,261|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|Allergies|253,261|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Attribute|Clinical Attribute|Allergies|266,270|false|false|false|C2598155||pain
Event|Event|Allergies|266,270|false|false|false|||pain
Finding|Functional Concept|Allergies|266,270|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Allergies|266,270|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Classification|Allergies|273,278|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Allergies|279,287|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Allergies|279,287|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Allergies|291,309|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Allergies|300,309|false|false|false|C0945766||Procedure
Event|Event|Allergies|300,309|false|false|false|||Procedure
Event|Occupational Activity|Allergies|300,309|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Allergies|300,309|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Allergies|300,309|false|false|false|C0184661|Interventional procedure|Procedure
Event|Event|Allergies|311,321|false|false|false|||Evacuation
Procedure|Therapeutic or Preventive Procedure|Allergies|311,321|false|false|false|C1282573|Evacuation procedure|Evacuation
Procedure|Therapeutic or Preventive Procedure|Allergies|311,333|false|false|false|C1261965|Evacuation of hematoma|Evacuation of hematoma
Event|Event|Allergies|325,333|false|false|false|||hematoma
Finding|Pathologic Function|Allergies|325,333|false|false|false|C0018944|Hematoma|hematoma
Event|Event|History of Present Illness|379,394|false|false|false|||anticoagulation
Finding|Finding|History of Present Illness|379,394|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Finding|Physiologic Function|History of Present Illness|379,394|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|379,394|false|false|false|C0003281|Anticoagulation Therapy|anticoagulation
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|402,408|false|false|false|C0006141|Breast|breast
Disorder|Neoplastic Process|History of Present Illness|402,408|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|breast
Event|Event|History of Present Illness|402,408|false|false|false|||breast
Finding|Finding|History of Present Illness|402,408|false|false|false|C0567499|Breast problem|breast
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|402,408|false|false|false|C0191838|Procedures on breast|breast
Disorder|Disease or Syndrome|History of Present Illness|409,412|false|false|false|C1449563|Cardiomyopathy, Familial Idiopathic|IDC
Event|Event|History of Present Illness|409,412|false|false|false|||IDC
Finding|Gene or Genome|History of Present Illness|409,412|false|false|false|C1881349|LMNA wt Allele|IDC
Finding|Classification|History of Present Illness|413,418|false|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|Grade
Finding|Finding|History of Present Illness|413,418|false|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|Grade
Finding|Classification|History of Present Illness|413,420|false|false|false|C0450094;C0475271;C0687697;C4283820|Grade three rank;Simpson Grade 3;Tumor grade G3;grade 3 education level|Grade 3
Finding|Finding|History of Present Illness|413,420|false|false|false|C0450094;C0475271;C0687697;C4283820|Grade three rank;Simpson Grade 3;Tumor grade G3;grade 3 education level|Grade 3
Finding|Intellectual Product|History of Present Illness|413,420|false|false|false|C0450094;C0475271;C0687697;C4283820|Grade three rank;Simpson Grade 3;Tumor grade G3;grade 3 education level|Grade 3
Event|Event|History of Present Illness|419,420|false|false|false|||3
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|432,438|false|false|false|C0006141|Breast|breast
Disorder|Neoplastic Process|History of Present Illness|432,438|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|breast
Event|Event|History of Present Illness|432,438|false|false|false|||breast
Finding|Finding|History of Present Illness|432,438|false|false|false|C0567499|Breast problem|breast
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|432,438|false|false|false|C0191838|Procedures on breast|breast
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|432,449|false|false|false|C0851238|Lumpectomy of breast|breast lumpectomy
Event|Event|History of Present Illness|439,449|false|false|false|||lumpectomy
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|439,449|false|false|false|C0851238;C1262070|Excision of mass (procedure);Lumpectomy of breast|lumpectomy
Event|Event|History of Present Illness|454,458|false|false|false|||SLNB
Procedure|Diagnostic Procedure|History of Present Illness|454,458|false|false|false|C0796693|Sentinel Lymph Node Biopsy|SLNB
Finding|Functional Concept|History of Present Illness|464,468|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|464,475|false|false|false|C0222601|Left breast|left breast
Finding|Sign or Symptom|History of Present Illness|464,484|false|false|false|C2127345|localized swelling in left breast|left breast swelling
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|469,475|false|false|false|C0006141|Breast|breast
Disorder|Neoplastic Process|History of Present Illness|469,475|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|breast
Finding|Finding|History of Present Illness|469,475|false|false|false|C0567499|Breast problem|breast
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|469,475|false|false|false|C0191838|Procedures on breast|breast
Finding|Finding|History of Present Illness|469,484|false|false|false|C0006152|Swelling of breast|breast swelling
Event|Event|History of Present Illness|476,484|false|false|false|||swelling
Finding|Finding|History of Present Illness|476,484|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|History of Present Illness|476,484|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Attribute|Clinical Attribute|History of Present Illness|490,494|false|false|false|C2598155||pain
Event|Event|History of Present Illness|490,494|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|490,494|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|490,494|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|History of Present Illness|512,520|false|false|false|||hematoma
Finding|Pathologic Function|History of Present Illness|512,520|false|false|false|C0018944|Hematoma|hematoma
Disorder|Disease or Syndrome|Past Medical History|547,559|false|false|false|C0242339|Dyslipidemias|Dyslipidemia
Event|Event|Past Medical History|547,559|false|false|false|||Dyslipidemia
Disorder|Disease or Syndrome|Past Medical History|561,575|false|false|false|C0042345|Varicosity|varicose veins
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|570,575|false|false|false|C0042449|Veins|veins
Event|Event|Past Medical History|570,575|false|false|false|||veins
Procedure|Therapeutic or Preventive Procedure|Past Medical History|570,575|false|false|false|C0398102|Procedure on vein|veins
Event|Event|Past Medical History|586,594|false|false|false|||ligation
Procedure|Therapeutic or Preventive Procedure|Past Medical History|586,594|false|false|false|C0023690|Ligation|ligation
Disorder|Disease or Syndrome|Past Medical History|596,600|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Past Medical History|596,600|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Past Medical History|596,600|false|false|false|||COPD
Finding|Gene or Genome|Past Medical History|596,600|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|Past Medical History|602,605|false|false|false|C0520679|Sleep Apnea, Obstructive|OSA
Drug|Amino Acid, Peptide, or Protein|Past Medical History|602,605|false|false|false|C0764906|OSA protein, Drosophila|OSA
Drug|Biologically Active Substance|Past Medical History|602,605|false|false|false|C0764906|OSA protein, Drosophila|OSA
Event|Event|Past Medical History|602,605|false|false|false|||OSA
Event|Event|Past Medical History|609,613|false|false|false|||CPap
Finding|Gene or Genome|Past Medical History|609,613|false|false|false|C1424863|CENPJ gene|CPap
Procedure|Therapeutic or Preventive Procedure|Past Medical History|609,613|false|false|false|C0199451|Continuous Positive Airway Pressure|CPap
Finding|Finding|Past Medical History|616,626|false|false|false|C2169609|recent upper respiratory infection|recent URI
Disorder|Disease or Syndrome|Past Medical History|623,626|false|false|false|C0041912|Upper Respiratory Infections|URI
Event|Event|Past Medical History|623,626|false|false|false|||URI
Finding|Gene or Genome|Past Medical History|623,626|false|false|false|C1421895;C1548524;C3272713|URI1 gene;URI1 wt Allele;Uniform Resource Identifier|URI
Finding|Intellectual Product|Past Medical History|623,626|false|false|false|C1421895;C1548524;C3272713|URI1 gene;URI1 wt Allele;Uniform Resource Identifier|URI
Event|Event|Past Medical History|637,643|false|false|false|||course
Drug|Antibiotic|Past Medical History|647,656|false|false|false|C0678143|Zithromax|Zithromax
Drug|Organic Chemical|Past Medical History|647,656|false|false|false|C0678143|Zithromax|Zithromax
Event|Event|Past Medical History|647,656|false|false|false|||Zithromax
Event|Event|Past Medical History|659,668|false|false|false|||bilateral
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|670,673|false|false|false|C0016504;C0687080;C1690938;C3853547|Foot;Hindfoot of quadruped;Paw;Structure of ankle and/or foot (body structure)|PEs
Finding|Gene or Genome|Past Medical History|670,673|false|false|false|C0687136;C1418467|PES1 gene;Personal Experience Scales|PEs
Finding|Intellectual Product|Past Medical History|670,673|false|false|false|C0687136;C1418467|PES1 gene;Personal Experience Scales|PEs
Drug|Amino Acid, Peptide, or Protein|Past Medical History|681,706|false|false|false|C0162595|Antiphospholipid Antibodies|antiphospholipid antibody
Drug|Immunologic Factor|Past Medical History|681,706|false|false|false|C0162595|Antiphospholipid Antibodies|antiphospholipid antibody
Finding|Finding|Past Medical History|681,706|false|false|false|C4019436|Antiphospholipid antibody positivity|antiphospholipid antibody
Disorder|Disease or Syndrome|Past Medical History|681,715|false|false|false|C0085278|Antiphospholipid Syndrome|antiphospholipid antibody syndrome
Anatomy|Cell Component|Past Medical History|698,706|false|false|false|C1167408;C3665580|Immunoglobulin complex location, circulating;immunoglobulin complex location|antibody
Drug|Amino Acid, Peptide, or Protein|Past Medical History|698,706|false|false|false|C0003241;C0021027|Antibodies;Immunoglobulins|antibody
Drug|Immunologic Factor|Past Medical History|698,706|false|false|false|C0003241;C0021027|Antibodies;Immunoglobulins|antibody
Drug|Pharmacologic Substance|Past Medical History|698,706|false|false|false|C0003241;C0021027|Antibodies;Immunoglobulins|antibody
Procedure|Laboratory Procedure|Past Medical History|698,706|false|false|false|C4551530|Antibody (immunoassay)|antibody
Disorder|Disease or Syndrome|Past Medical History|707,715|false|false|false|C0039082|Syndrome|syndrome
Event|Event|Past Medical History|707,715|false|false|false|||syndrome
Event|Event|Past Medical History|730,745|false|false|false|||anticoagulation
Finding|Finding|Past Medical History|730,745|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Finding|Physiologic Function|Past Medical History|730,745|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Procedure|Therapeutic or Preventive Procedure|Past Medical History|730,745|false|false|false|C0003281|Anticoagulation Therapy|anticoagulation
Event|Event|Past Medical History|759,762|false|false|false|||A1C
Finding|Classification|Past Medical History|759,762|false|false|false|C4521595|United States Military enlisted E3 (qualifier value)|A1C
Procedure|Laboratory Procedure|Past Medical History|759,762|false|false|false|C0474680|Hemoglobin A1c measurement|A1C
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|775,783|false|false|false|C0006104;C0228174|Brain;Cerebral hemisphere structure (body structure)|cerebral
Event|Event|Past Medical History|785,793|false|false|false|||aneurysm
Finding|Pathologic Function|Past Medical History|785,793|false|false|false|C0002940|Aneurysm|aneurysm
Finding|Finding|Past Medical History|816,825|false|false|false|C0442739||unchanged
Disorder|Disease or Syndrome|Past Medical History|828,832|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Event|Event|Past Medical History|828,832|false|false|false|||GERD
Disorder|Disease or Syndrome|Past Medical History|835,849|false|false|false|C1510475|Diverticulosis|diverticulosis
Event|Event|Past Medical History|835,849|false|false|false|||diverticulosis
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|855,860|false|false|false|C0009368;C4071907|Abdomen+Pelvis>Colon;Colon structure (body structure)|colon
Disorder|Disease or Syndrome|Past Medical History|855,860|true|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Disorder|Neoplastic Process|Past Medical History|855,860|true|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Finding|Finding|Past Medical History|855,860|true|false|false|C0750873|COLON PROBLEM|colon
Disorder|Anatomical Abnormality|Past Medical History|855,867|true|false|false|C0009376|Colonic Polyps|colon polyps
Disorder|Anatomical Abnormality|Past Medical History|861,867|false|false|false|C0032584|polyps|polyps
Event|Event|Past Medical History|861,867|false|false|false|||polyps
Finding|Intellectual Product|Past Medical History|861,867|false|false|false|C1546747||polyps
Disorder|Mental or Behavioral Dysfunction|Past Medical History|869,879|false|false|false|C0011570;C0011581;C0344315;C0812393|Cancer patients and suicide and depression;Depressed mood;Depressive disorder;Mental Depression|depression
Event|Event|Past Medical History|869,879|false|false|false|||depression
Finding|Functional Concept|Past Medical History|869,879|false|false|false|C0460137;C1579931|Depression - motion|depression
Finding|Sign or Symptom|Past Medical History|869,879|false|false|false|C0460137;C1579931|Depression - motion|depression
Finding|Functional Concept|Past Medical History|885,890|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Cell|Past Medical History|891,894|false|false|false|C3890599|Circulating Melanoma Cell|CMC
Disorder|Congenital Abnormality|Past Medical History|891,894|false|false|false|C0006845;C0340803|Candidiasis, Chronic Mucocutaneous;Capillary malformation (disorder)|CMC
Disorder|Disease or Syndrome|Past Medical History|891,894|false|false|false|C0006845;C0340803|Candidiasis, Chronic Mucocutaneous;Capillary malformation (disorder)|CMC
Event|Event|Past Medical History|891,894|false|false|false|||CMC
Procedure|Therapeutic or Preventive Procedure|Past Medical History|891,894|false|false|false|C0065772|MCC protocol|CMC
Anatomy|Body Space or Junction|Past Medical History|896,901|false|false|false|C0022417;C0392905;C1269611|Articular system;Joints|joint
Anatomy|Body System|Past Medical History|896,901|false|false|false|C0022417;C0392905;C1269611|Articular system;Joints|joint
Finding|Finding|Past Medical History|896,901|false|false|false|C0575044|Joint problem|joint
Procedure|Therapeutic or Preventive Procedure|Past Medical History|896,914|false|false|false|C0003893|Arthroplasty|joint arthroplasty
Event|Event|Past Medical History|902,914|false|false|false|||arthroplasty
Procedure|Therapeutic or Preventive Procedure|Past Medical History|902,914|false|false|false|C0003893;C0700235;C5887062|Arthroplasty;Reconstruction of joint;Temporomandibular joint arthroplasty by dentist|arthroplasty
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|920,932|false|false|false|C0085515|Rotator Cuff|rotator cuff
Procedure|Therapeutic or Preventive Procedure|Past Medical History|920,939|false|false|false|C0186666|Repair of musculotendinous cuff of shoulder|rotator cuff repair
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|928,932|false|false|false|C1550244|Cuff - body part|cuff
Finding|Pathologic Function|Past Medical History|928,932|false|false|false|C3668885|Cuffing (morphologic abnormality)|cuff
Event|Event|Past Medical History|933,939|false|false|false|||repair
Finding|Functional Concept|Past Medical History|933,939|false|false|false|C0043240;C4319951|Repair;Wound Healing|repair
Finding|Organism Function|Past Medical History|933,939|false|false|false|C0043240;C4319951|Repair;Wound Healing|repair
Procedure|Health Care Activity|Past Medical History|933,939|false|false|false|C0374711;C1705181|Repair - Remedial Action;Surgical repair|repair
Procedure|Therapeutic or Preventive Procedure|Past Medical History|933,939|false|false|false|C0374711;C1705181|Repair - Remedial Action;Surgical repair|repair
Procedure|Therapeutic or Preventive Procedure|Past Medical History|941,949|false|false|false|C0015252;C0728940|Excision;removal technique|excision
Finding|Functional Concept|Past Medical History|950,955|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|961,966|false|false|false|C0582802|Digit structure|digit
Finding|Gene or Genome|Past Medical History|961,966|false|false|false|C4761764|GSC-DT gene|digit
Event|Event|Past Medical History|967,971|false|false|false|||mass
Finding|Finding|Past Medical History|967,971|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|Past Medical History|967,971|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|Past Medical History|967,971|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Event|Event|Past Medical History|973,976|false|false|false|||CCY
Event|Event|Past Medical History|979,984|false|false|false|||stone
Finding|Body Substance|Past Medical History|979,984|false|false|false|C0006736|Calculi|stone
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|987,997|false|false|false|C0030274|Pancreas|pancreatic
Drug|Amino Acid, Peptide, or Protein|Past Medical History|987,997|false|false|false|C0030292|Pancreatic Hormones|pancreatic
Drug|Hormone|Past Medical History|987,997|false|false|false|C0030292|Pancreatic Hormones|pancreatic
Drug|Pharmacologic Substance|Past Medical History|987,997|false|false|false|C0030292|Pancreatic Hormones|pancreatic
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|987,1002|false|false|false|C0030288;C4482304|Abdomen>Pancreatic duct;Pancreatic duct|pancreatic duct
Disorder|Neoplastic Process|Past Medical History|987,1002|false|false|false|C0153461|Malignant neoplasm of pancreatic duct|pancreatic duct
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|998,1002|false|false|false|C0687028;C1550227|Duct (organ) structure;canal [body parts]|duct
Event|Event|Past Medical History|1003,1014|false|false|false|||exploration
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1003,1014|false|false|false|C1280903|Exploration procedure|exploration
Event|Event|Past Medical History|1023,1035|false|false|false|||hysterectomy
Finding|Finding|Past Medical History|1023,1035|false|false|false|C1548863|Consent Type - Hysterectomy|hysterectomy
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1023,1035|false|false|false|C0020699|Hysterectomy|hysterectomy
Event|Event|Past Medical History|1037,1050|false|false|false|||tonsillectomy
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1037,1050|false|false|false|C0040423|Tonsillectomy|tonsillectomy
Finding|Classification|Family Medical History|1093,1099|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|Family Medical History|1093,1099|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|Family Medical History|1093,1099|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|Family Medical History|1093,1099|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Anatomy|Body Location or Region|Family Medical History|1106,1109|true|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|Family Medical History|1106,1109|true|false|false|C2926618||DVT
Disorder|Disease or Syndrome|Family Medical History|1106,1109|true|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Event|Event|Family Medical History|1106,1109|true|false|false|||DVT
Event|Event|Family Medical History|1113,1115|true|false|false|||PE
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1134,1140|false|false|false|C0018792|Heart Atrium|atrial
Attribute|Clinical Attribute|Family Medical History|1134,1153|false|false|false|C2926591||atrial fibrillation
Disorder|Disease or Syndrome|Family Medical History|1134,1153|false|false|false|C0004238|Atrial Fibrillation|atrial fibrillation
Lab|Laboratory or Test Result|Family Medical History|1134,1153|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|atrial fibrillation
Disorder|Disease or Syndrome|Family Medical History|1141,1153|false|false|false|C0232197|Fibrillation|fibrillation
Event|Event|Family Medical History|1141,1153|false|false|false|||fibrillation
Event|Event|General Exam|1204,1208|false|false|false|||Temp
Finding|Gene or Genome|General Exam|1204,1208|false|false|false|C1823816|C1orf210 gene|Temp
Procedure|Therapeutic or Preventive Procedure|General Exam|1204,1208|false|false|false|C0279848|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Temp
Event|Event|General Exam|1257,1265|false|false|false|||delivery
Finding|Finding|General Exam|1257,1265|false|false|false|C1314680;C1705822;C2053584|Transfer Technique;delivery (history)|delivery
Finding|Functional Concept|General Exam|1257,1265|false|false|false|C1314680;C1705822;C2053584|Transfer Technique;delivery (history)|delivery
Finding|Organism Function|General Exam|1257,1265|false|false|false|C1314680;C1705822;C2053584|Transfer Technique;delivery (history)|delivery
Procedure|Therapeutic or Preventive Procedure|General Exam|1257,1265|false|false|false|C0011209|Obstetric Delivery|delivery
Event|Event|General Exam|1271,1274|false|false|false|||GEN
Finding|Classification|General Exam|1271,1274|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|GEN
Finding|Gene or Genome|General Exam|1271,1274|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|GEN
Disorder|Disease or Syndrome|General Exam|1276,1279|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|General Exam|1276,1279|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|General Exam|1276,1279|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|1276,1279|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|General Exam|1276,1279|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|General Exam|1276,1279|false|false|false|||NAD
Finding|Finding|General Exam|1276,1279|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Event|Event|General Exam|1281,1289|false|false|false|||pleasant
Finding|Mental Process|General Exam|1281,1289|false|false|false|C2987187|Pleasant|pleasant
Anatomy|Body Location or Region|General Exam|1303,1308|false|false|false|C1512338|HEENT|HEENT
Event|Event|General Exam|1310,1314|false|false|false|||NCAT
Event|Event|General Exam|1316,1320|false|false|false|||EOMI
Anatomy|Body Part, Organ, or Organ Component|General Exam|1322,1328|false|false|false|C0036410|Sclera|sclera
Disorder|Disease or Syndrome|General Exam|1322,1328|false|false|false|C0036412|Scleral Diseases|sclera
Event|Event|General Exam|1322,1328|false|false|false|||sclera
Procedure|Health Care Activity|General Exam|1322,1328|false|false|false|C2228481|examination of sclera|sclera
Event|Event|General Exam|1329,1338|false|false|false|||anicteric
Finding|Finding|General Exam|1329,1338|false|false|false|C0205180|Anicteric|anicteric
Event|Event|General Exam|1343,1346|false|false|false|||RRR
Event|Event|General Exam|1347,1351|false|false|false|||PULM
Procedure|Health Care Activity|General Exam|1347,1351|false|false|false|C1315068|Pulmonary ventilator management|PULM
Event|Event|General Exam|1356,1365|true|false|false|||increased
Finding|Finding|General Exam|1356,1365|true|false|false|C0442805;C5236002|Increase;Increased (finding)|increased
Finding|Functional Concept|General Exam|1356,1365|true|false|false|C0442805;C5236002|Increase;Increased (finding)|increased
Finding|Sign or Symptom|General Exam|1356,1383|true|false|false|C0859927|Increased work of breathing|increased work of breathing
Event|Event|General Exam|1366,1370|true|false|false|||work
Event|Occupational Activity|General Exam|1366,1370|true|false|false|C0043227|Work|work
Finding|Organ or Tissue Function|General Exam|1366,1383|true|false|false|C0043229|Work of Breathing|work of breathing
Attribute|Clinical Attribute|General Exam|1374,1383|true|false|false|C5885990||breathing
Event|Event|General Exam|1374,1383|true|false|false|||breathing
Finding|Finding|General Exam|1374,1383|true|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|General Exam|1374,1383|true|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|General Exam|1374,1383|true|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|General Exam|1374,1383|true|false|false|C1160636|respiratory system process|breathing
Event|Event|General Exam|1385,1396|true|false|false|||comfortable
Finding|Finding|General Exam|1385,1396|true|false|false|C5546696|Feeling comfortable|comfortable
Event|Event|General Exam|1400,1402|false|false|false|||RA
Anatomy|Body Part, Organ, or Organ Component|General Exam|1403,1409|false|false|false|C0006141|Breast|BREAST
Disorder|Neoplastic Process|General Exam|1403,1409|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|BREAST
Event|Event|General Exam|1403,1409|false|false|false|||BREAST
Finding|Finding|General Exam|1403,1409|false|false|false|C0567499|Breast problem|BREAST
Procedure|Therapeutic or Preventive Procedure|General Exam|1403,1409|false|false|false|C0191838|Procedures on breast|BREAST
Anatomy|Body Part, Organ, or Organ Component|General Exam|1413,1419|false|false|false|C0006141|Breast|breast
Disorder|Neoplastic Process|General Exam|1413,1419|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|breast
Event|Event|General Exam|1413,1419|false|false|false|||breast
Finding|Finding|General Exam|1413,1419|false|false|false|C0567499|Breast problem|breast
Procedure|Therapeutic or Preventive Procedure|General Exam|1413,1419|false|false|false|C0191838|Procedures on breast|breast
Finding|Functional Concept|General Exam|1425,1434|false|false|false|C3244310|dependent|dependent
Event|Event|General Exam|1435,1445|false|false|false|||ecchymosis
Finding|Finding|General Exam|1435,1445|false|false|false|C0013491;C3812660|Ecchymosis;Skin Bruise|ecchymosis
Finding|Pathologic Function|General Exam|1435,1445|false|false|false|C0013491;C3812660|Ecchymosis;Skin Bruise|ecchymosis
Event|Event|General Exam|1458,1466|false|false|false|||inferior
Finding|Social Behavior|General Exam|1458,1466|false|false|false|C0678975|inferiority|inferior
Anatomy|Body Part, Organ, or Organ Component|General Exam|1467,1473|false|false|false|C0006141|Breast|breast
Disorder|Neoplastic Process|General Exam|1467,1473|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|breast
Event|Event|General Exam|1467,1473|false|false|false|||breast
Finding|Finding|General Exam|1467,1473|false|false|false|C0567499|Breast problem|breast
Procedure|Therapeutic or Preventive Procedure|General Exam|1467,1473|false|false|false|C0191838|Procedures on breast|breast
Anatomy|Body Location or Region|General Exam|1475,1483|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|General Exam|1475,1483|false|false|false|C0332803|Surgical wound|incision
Event|Event|General Exam|1475,1483|false|false|false|||incision
Procedure|Therapeutic or Preventive Procedure|General Exam|1475,1483|false|false|false|C0184898|Surgical incisions|incision
Drug|Substance|General Exam|1494,1499|false|false|false|C1550628|Drain - SpecimenType|drain
Event|Event|General Exam|1494,1499|false|false|false|||drain
Finding|Intellectual Product|General Exam|1494,1499|false|false|false|C1546604|Drain Specimen Code|drain
Event|Event|General Exam|1521,1527|false|false|false|||output
Finding|Conceptual Entity|General Exam|1521,1527|false|false|false|C1709366|system output|output
Procedure|Health Care Activity|General Exam|1521,1527|false|false|false|C3251815|Measurement of fluid output|output
Anatomy|Body Location or Region|General Exam|1530,1533|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|ABD
Disorder|Cell or Molecular Dysfunction|General Exam|1530,1533|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|ABD
Event|Event|General Exam|1530,1533|false|false|false|||ABD
Disorder|Disease or Syndrome|General Exam|1535,1539|true|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|General Exam|1535,1539|true|false|false|||soft
Event|Event|General Exam|1571,1577|true|false|false|||masses
Disorder|Anatomical Abnormality|General Exam|1581,1587|true|false|false|C0019270|Hernia|hernia
Event|Event|General Exam|1581,1587|true|false|false|||hernia
Disorder|Congenital Abnormality|General Exam|1588,1591|true|false|false|C0015306|Hereditary Multiple Exostoses|EXT
Event|Event|General Exam|1588,1591|true|false|false|||EXT
Finding|Gene or Genome|General Exam|1588,1591|true|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|EXT
Event|Event|General Exam|1593,1597|true|false|false|||Warm
Finding|Finding|General Exam|1593,1597|true|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|General Exam|1593,1597|true|false|false|C0687712|warming process|Warm
Finding|Finding|General Exam|1599,1603|true|false|false|C5575035|Well (answer to question)|well
Event|Event|General Exam|1604,1612|true|false|false|||perfused
Attribute|Clinical Attribute|General Exam|1617,1622|true|false|false|C1717255||edema
Event|Event|General Exam|1617,1622|true|false|false|||edema
Finding|Pathologic Function|General Exam|1617,1622|true|false|false|C0013604|Edema|edema
Event|Event|General Exam|1627,1637|true|false|false|||tenderness
Finding|Mental Process|General Exam|1627,1637|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|General Exam|1627,1637|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Finding|General Exam|1656,1681|true|false|false|C0746857|Focal Neurologic Deficits|focal neurologic deficits
Finding|Finding|General Exam|1662,1681|true|false|false|C0521654|Neurologic Deficits|neurologic deficits
Event|Event|General Exam|1673,1681|true|false|false|||deficits
Disorder|Mental or Behavioral Dysfunction|General Exam|1682,1687|true|false|false|C0004936;C1306597|Mental disorders;Psychiatric problem|PSYCH
Event|Event|General Exam|1682,1687|true|false|false|||PSYCH
Event|Event|General Exam|1696,1704|false|false|false|||judgment
Finding|Mental Process|General Exam|1696,1704|false|false|false|C0022423|Judgment|judgment
Finding|Mental Process|General Exam|1705,1712|false|false|false|C0233820|Insight|insight
Event|Event|General Exam|1721,1727|false|false|false|||memory
Finding|Finding|General Exam|1721,1727|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Finding|Intellectual Product|General Exam|1721,1727|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Finding|Mental Process|General Exam|1721,1727|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Event|Event|General Exam|1729,1735|false|false|false|||normal
Attribute|Clinical Attribute|General Exam|1737,1741|false|false|false|C2713234||mood
Event|Event|General Exam|1737,1741|false|false|false|||mood
Finding|Conceptual Entity|General Exam|1737,1741|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|mood
Finding|Finding|General Exam|1737,1741|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|mood
Finding|Mental Process|General Exam|1737,1741|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|mood
Event|Event|General Exam|1742,1748|false|false|false|||affect
Finding|Mental Process|General Exam|1742,1748|false|false|false|C0001721|Affect (mental function)|affect
Procedure|Health Care Activity|General Exam|1742,1748|false|false|false|C2237113|assessment of affect|affect
Disorder|Disease or Syndrome|General Exam|1782,1787|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|1782,1787|false|false|false|||BLOOD
Finding|Body Substance|General Exam|1782,1787|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|1788,1791|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|1796,1799|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|1796,1799|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|1796,1799|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|1806,1809|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|1806,1809|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|1806,1809|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|1806,1809|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|1815,1818|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|1815,1818|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|1826,1829|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|1826,1829|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|1826,1829|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|1826,1829|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|1826,1829|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|1833,1836|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|1833,1836|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|1833,1836|false|false|false|||MCH
Finding|Gene or Genome|General Exam|1833,1836|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|1833,1836|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|1833,1836|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|General Exam|1842,1846|false|false|false|||MCHC
Procedure|Laboratory Procedure|General Exam|1842,1846|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|1874,1877|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|1894,1899|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|1894,1899|false|false|false|||BLOOD
Finding|Body Substance|General Exam|1894,1899|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|1904,1907|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|General Exam|1904,1907|false|false|false|||PTT
Procedure|Laboratory Procedure|General Exam|1904,1907|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|General Exam|1929,1934|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|1929,1934|false|false|false|||BLOOD
Finding|Body Substance|General Exam|1929,1934|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|1929,1942|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|1929,1942|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|1929,1942|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|1935,1942|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|1935,1942|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|1935,1942|false|false|false|C0017725|glucose|Glucose
Event|Event|General Exam|1935,1942|false|false|false|||Glucose
Lab|Laboratory or Test Result|General Exam|1935,1942|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|1935,1942|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|General Exam|1987,1991|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|1987,1991|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|General Exam|1987,1991|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|General Exam|2016,2021|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|2016,2021|false|false|false|||BLOOD
Finding|Body Substance|General Exam|2016,2021|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|2016,2029|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|General Exam|2022,2029|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|General Exam|2022,2029|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|General Exam|2022,2029|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|General Exam|2022,2029|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|General Exam|2022,2029|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|General Exam|2022,2029|false|false|false|||Calcium
Finding|Physiologic Function|General Exam|2022,2029|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|General Exam|2022,2029|false|false|false|C0201925|Calcium measurement|Calcium
Event|Activity|General Exam|2052,2063|false|false|false|C4321457|Examination|EXAMINATION
Event|Event|General Exam|2052,2063|false|false|false|||EXAMINATION
Procedure|Health Care Activity|General Exam|2052,2063|false|false|false|C0031809;C0582103|Medical Examination;Physical Examination|EXAMINATION
Drug|Amino Acid, Peptide, or Protein|General Exam|2066,2069|false|false|false|C3813556|Cancer/Testis Antigen|CTA
Event|Event|General Exam|2066,2069|false|false|false|||CTA
Finding|Gene or Genome|General Exam|2066,2069|false|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|General Exam|2066,2069|false|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Anatomy|Body Location or Region|General Exam|2070,2075|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|CHEST
Event|Event|General Exam|2070,2075|false|false|false|||CHEST
Finding|Finding|General Exam|2070,2075|false|false|false|C0741025|Chest problem|CHEST
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|2081,2089|false|false|false|C0009924|Contrast Media|CONTRAST
Event|Event|General Exam|2081,2089|false|false|false|||CONTRAST
Event|Activity|General Exam|2092,2102|false|false|false|C1707455|Comparison|COMPARISON
Event|Event|General Exam|2092,2102|false|false|false|||COMPARISON
Anatomy|Body Location or Region|General Exam|2105,2110|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|General Exam|2105,2110|false|false|false|C0741025|Chest problem|Chest
Procedure|Diagnostic Procedure|General Exam|2105,2113|false|false|false|C0202823|Chest CT|Chest CT
Event|Event|General Exam|2111,2113|false|false|false|||CT
Anatomy|Body Part, Organ, or Organ Component|Findings|2144,2149|false|false|false|C0018787;C4037974|Chest>Heart;Heart|HEART
Disorder|Neoplastic Process|Findings|2144,2149|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|HEART
Event|Event|Findings|2144,2149|false|false|false|||HEART
Finding|Sign or Symptom|Findings|2144,2149|false|false|false|C0795691|HEART PROBLEM|HEART
Anatomy|Anatomical Structure|Findings|2154,2165|false|false|false|C3714653|Vasculature|VASCULATURE
Drug|Pharmacologic Substance|Findings|2179,2186|true|false|false|C0719205|Central brand of multivitamin with minerals|central
Drug|Vitamin|Findings|2179,2186|true|false|false|C0719205|Central brand of multivitamin with minerals|central
Event|Event|Findings|2179,2186|true|false|false|||central
Procedure|Laboratory Procedure|Findings|2179,2186|true|false|false|C1879652|Central Minus|central
Anatomy|Body Part, Organ, or Organ Component|Findings|2187,2196|true|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Findings|2187,2196|true|false|false|C2707265||pulmonary
Finding|Finding|Findings|2187,2196|true|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|Findings|2187,2205|true|false|false|C0034065|Pulmonary Embolism|pulmonary embolism
Event|Event|Findings|2197,2205|true|false|false|||embolism
Finding|Finding|Findings|2197,2205|true|false|false|C0013922;C1704212|Embolism;Embolus|embolism
Finding|Pathologic Function|Findings|2197,2205|true|false|false|C0013922;C1704212|Embolism;Embolus|embolism
Anatomy|Body Location or Region|Findings|2213,2221|true|false|false|C0817096|Chest|thoracic
Disorder|Disease or Syndrome|Findings|2213,2221|true|false|false|C5779551|Dissecting Thoracic Aortic Aneurysm|thoracic
Anatomy|Body Part, Organ, or Organ Component|Findings|2223,2228|true|false|false|C0003483;C4037978|Aorta;Chest+Abdomen>Aorta|aorta
Event|Event|Findings|2223,2228|true|false|false|||aorta
Procedure|Health Care Activity|Findings|2223,2228|true|false|false|C0869784|Procedure on aorta|aorta
Event|Event|Findings|2232,2238|true|false|false|||normal
Event|Event|Findings|2242,2249|true|false|false|||caliber
Event|Event|Findings|2258,2266|true|false|false|||evidence
Finding|Idea or Concept|Findings|2258,2266|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Findings|2258,2269|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Event|Event|Findings|2270,2280|true|false|false|||dissection
Finding|Pathologic Function|Findings|2270,2280|true|false|false|C0333288|Dissecting hemorrhage|dissection
Procedure|Therapeutic or Preventive Procedure|Findings|2270,2280|true|false|false|C0012737|Tissue Dissection|dissection
Event|Event|Findings|2297,2305|false|false|false|||hematoma
Finding|Pathologic Function|Findings|2297,2305|false|false|false|C0018944|Hematoma|hematoma
Anatomy|Body Part, Organ, or Organ Component|Findings|2312,2317|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Findings|2312,2317|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Event|Event|Findings|2312,2317|false|false|false|||heart
Finding|Sign or Symptom|Findings|2312,2317|false|false|false|C0795691|HEART PROBLEM|heart
Anatomy|Body Part, Organ, or Organ Component|Findings|2319,2330|false|false|false|C0031050|Pericardial sac structure|pericardium
Finding|Gene or Genome|Findings|2336,2341|false|false|false|C1424898|RXFP2 gene|great
Anatomy|Body Part, Organ, or Organ Component|Findings|2336,2349|false|false|false|C0225991|Structure of great blood vessel (organ)|great vessels
Anatomy|Body Part, Organ, or Organ Component|Findings|2342,2349|false|false|false|C0005847|Blood Vessel|vessels
Event|Event|Findings|2369,2375|false|false|false|||limits
Finding|Functional Concept|Findings|2369,2375|false|false|false|C0439801|Limited (extensiveness)|limits
Anatomy|Body Location or Region|Findings|2381,2392|true|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Anatomy|Body Part, Organ, or Organ Component|Findings|2381,2392|true|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Disorder|Disease or Syndrome|Findings|2381,2401|true|false|false|C0031039|Pericardial effusion|pericardial effusion
Finding|Body Substance|Findings|2381,2401|true|false|false|C1253937|Pericardial effusion body substance|pericardial effusion
Event|Event|Findings|2393,2401|true|false|false|||effusion
Finding|Body Substance|Findings|2393,2401|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|Findings|2393,2401|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|Findings|2393,2401|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Event|Event|Findings|2405,2409|true|false|false|||seen
Anatomy|Body Location or Region|Findings|2415,2421|false|false|false|C0004454|Axilla|AXILLA
Event|Event|Findings|2423,2427|false|false|false|||HILA
Anatomy|Body Location or Region|Findings|2433,2444|false|false|false|C0025066;C4037971|Chest>Mediastinum;Mediastinum|MEDIASTINUM
Anatomy|Body Part, Organ, or Organ Component|Findings|2433,2444|false|false|false|C0025066;C4037971|Chest>Mediastinum;Mediastinum|MEDIASTINUM
Disorder|Neoplastic Process|Findings|2433,2444|false|false|false|C0153956;C0496915|Benign tumor of mediastinum;Neoplasm of uncertain or unknown behavior of mediastinum|MEDIASTINUM
Event|Event|Findings|2477,2487|false|false|false|||collection
Finding|Conceptual Entity|Findings|2477,2487|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|Findings|2477,2487|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|Findings|2477,2487|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|Findings|2477,2487|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|Findings|2496,2500|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Findings|2496,2507|false|false|false|C0222601|Left breast|left breast
Anatomy|Body Part, Organ, or Organ Component|Findings|2501,2507|false|false|false|C0006141|Breast|breast
Disorder|Neoplastic Process|Findings|2501,2507|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|breast
Event|Event|Findings|2501,2507|false|false|false|||breast
Finding|Finding|Findings|2501,2507|false|false|false|C0567499|Breast problem|breast
Procedure|Therapeutic or Preventive Procedure|Findings|2501,2507|false|false|false|C0191838|Procedures on breast|breast
Event|Event|Findings|2514,2521|false|false|false|||density
Event|Event|Findings|2522,2531|false|false|false|||measuring
Event|Event|Findings|2554,2564|false|false|false|||consistent
Finding|Idea or Concept|Findings|2554,2564|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|Findings|2554,2569|false|false|false|C0332290|Consistent with|consistent with
Event|Event|Findings|2571,2579|false|false|false|||hematoma
Finding|Pathologic Function|Findings|2571,2579|false|false|false|C0018944|Hematoma|hematoma
Event|Event|Findings|2596,2600|false|false|false|||foci
Finding|Finding|Findings|2596,2600|false|false|false|C4321394|Foci|foci
Drug|Inorganic Chemical|Findings|2604,2607|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|Findings|2604,2607|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|Findings|2604,2607|false|false|false|C0001861;C3536832|Air (substance);air|air
Event|Event|Findings|2604,2607|false|false|false|||air
Finding|Finding|Findings|2604,2607|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|Findings|2604,2607|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|Findings|2604,2607|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Event|Event|Findings|2619,2629|false|false|false|||collection
Finding|Conceptual Entity|Findings|2619,2629|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|Findings|2619,2629|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|Findings|2619,2629|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|Findings|2619,2629|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Finding|Findings|2632,2638|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Findings|2632,2638|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Disorder|Injury or Poisoning|Findings|2651,2661|false|false|false|C1720922|Respiratory Aspiration|aspiration
Event|Event|Findings|2651,2661|false|false|false|||aspiration
Finding|Finding|Findings|2651,2661|false|false|false|C0220787;C0700198;C2712334|Aspiration into respiratory tract;Endotracheal aspiration;Pulmonary aspiration|aspiration
Finding|Organ or Tissue Function|Findings|2651,2661|false|false|false|C0220787;C0700198;C2712334|Aspiration into respiratory tract;Endotracheal aspiration;Pulmonary aspiration|aspiration
Finding|Pathologic Function|Findings|2651,2661|false|false|false|C0220787;C0700198;C2712334|Aspiration into respiratory tract;Endotracheal aspiration;Pulmonary aspiration|aspiration
Procedure|Therapeutic or Preventive Procedure|Findings|2651,2661|false|false|false|C0349707||aspiration
Finding|Finding|Findings|2666,2670|false|false|false|C5575035|Well (answer to question)|well
Event|Event|Findings|2687,2701|false|false|false|||hyperdensities
Event|Event|Findings|2710,2719|false|false|false|||periphery
Anatomy|Body Location or Region|Findings|2726,2734|true|false|false|C0004454|Axilla|axillary
Anatomy|Body Location or Region|Findings|2736,2747|true|false|false|C0025066|Mediastinum|mediastinal
Disorder|Disease or Syndrome|Findings|2752,2773|true|false|false|C0456973|Hilar lymphadenopathy|hilar lymphadenopathy
Disorder|Disease or Syndrome|Findings|2758,2773|false|false|false|C0497156|Lymphadenopathy|lymphadenopathy
Event|Event|Findings|2758,2773|false|false|false|||lymphadenopathy
Finding|Sign or Symptom|Findings|2758,2773|false|false|false|C4282165|Swollen Lymph Node|lymphadenopathy
Event|Event|Findings|2777,2784|false|false|false|||present
Finding|Finding|Findings|2777,2784|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|Findings|2777,2784|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Functional Concept|Findings|2792,2797|true|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|Findings|2792,2804|true|false|false|C0230337|Structure of right axillary region|right axilla
Anatomy|Body Location or Region|Findings|2798,2804|true|false|false|C0004454|Axilla|axilla
Event|Event|Findings|2813,2821|true|false|false|||included
Event|Event|Findings|2829,2834|true|false|false|||study
Finding|Intellectual Product|Findings|2829,2834|true|false|false|C1705923|Study Object|study
Procedure|Research Activity|Findings|2829,2834|true|false|false|C0008972;C0947630;C2603343|Clinical Research;Scientific Study;Study|study
Anatomy|Body Location or Region|Findings|2840,2851|true|false|false|C0025066|Mediastinum|mediastinal
Finding|Finding|Findings|2840,2856|true|false|false|C0240318|Mediastinal mass|mediastinal mass
Event|Event|Findings|2852,2856|true|false|false|||mass
Finding|Finding|Findings|2852,2856|true|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|Findings|2852,2856|true|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|Findings|2852,2856|true|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Anatomy|Tissue|Findings|2862,2869|false|false|false|C0032225|Pleura|PLEURAL
Disorder|Disease or Syndrome|Findings|2862,2869|false|false|false|C0032226|Pleural Diseases|PLEURAL
Anatomy|Body Space or Junction|Findings|2862,2876|false|false|false|C0178802|Pleural cavity|PLEURAL SPACES
Anatomy|Tissue|Findings|2881,2888|true|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|Findings|2881,2888|true|false|false|C0032226|Pleural Diseases|pleural
Finding|Body Substance|Findings|2881,2897|true|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Finding|Finding|Findings|2881,2897|true|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Finding|Pathologic Function|Findings|2881,2897|true|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Event|Event|Findings|2889,2897|true|false|false|||effusion
Finding|Body Substance|Findings|2889,2897|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|Findings|2889,2897|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|Findings|2889,2897|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Disorder|Disease or Syndrome|Findings|2901,2913|true|false|false|C0032326|Pneumothorax|pneumothorax
Event|Event|Findings|2901,2913|true|false|false|||pneumothorax
Anatomy|Body Part, Organ, or Organ Component|Findings|2919,2924|false|false|false|C0024109|Lung|LUNGS
Anatomy|Body Part, Organ, or Organ Component|Findings|2925,2932|false|false|false|C0458827|Airway structure|AIRWAYS
Anatomy|Body Part, Organ, or Organ Component|Findings|2955,2960|true|false|false|C0024109|Lung|lungs
Event|Event|Findings|2965,2970|true|false|false|||clear
Finding|Idea or Concept|Findings|2965,2970|true|false|false|C1550016|Remote control command - Clear|clear
Event|Event|Findings|2980,2986|true|false|false|||masses
Event|Event|Findings|2990,2995|true|false|false|||areas
Event|Event|Findings|3012,3025|false|false|false|||opacification
Anatomy|Body Part, Organ, or Organ Component|Findings|3032,3039|false|false|false|C0458827|Airway structure|airways
Event|Event|Findings|3044,3050|false|false|false|||patent
Finding|Intellectual Product|Findings|3044,3050|false|false|false|C0030650|Legal patent|patent
Anatomy|Body Part, Organ, or Organ Component|Findings|3083,3090|false|false|false|C0006255|Bronchi|bronchi
Anatomy|Body Location or Region|Findings|3108,3112|false|false|false|C2987514|Anatomical base|BASE
Drug|Biomedical or Dental Material|Findings|3108,3112|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|BASE
Drug|Chemical Viewed Functionally|Findings|3108,3112|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|BASE
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Findings|3108,3112|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|BASE
Event|Event|Findings|3108,3112|false|false|false|||BASE
Finding|Gene or Genome|Findings|3108,3112|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|BASE
Finding|Idea or Concept|Findings|3108,3112|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|BASE
Anatomy|Body Location or Region|Findings|3108,3120|false|false|false|C3686666|Base of neck|BASE OF NECK
Anatomy|Body Location or Region|Findings|3116,3120|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|Findings|3116,3120|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|Findings|3116,3120|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Finding|Functional Concept|Findings|3122,3132|false|false|false|C0234621|Visual|Visualized
Event|Event|Findings|3133,3141|false|false|false|||portions
Anatomy|Body Location or Region|Findings|3149,3153|true|false|false|C2987514|Anatomical base|base
Drug|Biomedical or Dental Material|Findings|3149,3153|true|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Chemical Viewed Functionally|Findings|3149,3153|true|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Findings|3149,3153|true|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Finding|Gene or Genome|Findings|3149,3153|true|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Finding|Idea or Concept|Findings|3149,3153|true|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Anatomy|Body Location or Region|Findings|3161,3165|true|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|Findings|3161,3165|true|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|Findings|3161,3165|true|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Disorder|Congenital Abnormality|Findings|3175,3186|true|false|false|C0000768|Congenital Abnormality|abnormality
Event|Event|Findings|3175,3186|true|false|false|||abnormality
Finding|Finding|Findings|3175,3186|true|false|false|C1704258|Abnormality|abnormality
Anatomy|Body Part, Organ, or Organ Component|Findings|3192,3197|false|false|false|C0262950;C1442209|Skeletal bone;XXX bone|BONES
Anatomy|Body Part, Organ, or Organ Component|Findings|3213,3220|true|false|false|C0262950;C4520924|Bone Tissue, Human;Skeletal bone|osseous
Anatomy|Tissue|Findings|3213,3220|true|false|false|C0262950;C4520924|Bone Tissue, Human;Skeletal bone|osseous
Disorder|Congenital Abnormality|Findings|3221,3232|true|false|false|C0000768|Congenital Abnormality|abnormality
Event|Event|Findings|3221,3232|true|false|false|||abnormality
Finding|Finding|Findings|3221,3232|true|false|false|C1704258|Abnormality|abnormality
Event|Event|Findings|3236,3240|true|false|false|||seen
Finding|Intellectual Product|Findings|3256,3261|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Disorder|Injury or Poisoning|Findings|3262,3270|true|false|false|C0016658|Fracture|fracture
Event|Event|Findings|3262,3270|true|false|false|||fracture
Finding|Functional Concept|Impression|3312,3316|true|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Impression|3312,3323|true|false|false|C0222601|Left breast|left breast
Anatomy|Body Part, Organ, or Organ Component|Impression|3317,3323|true|false|false|C0006141|Breast|breast
Disorder|Neoplastic Process|Impression|3317,3323|true|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|breast
Finding|Finding|Impression|3317,3323|true|false|false|C0567499|Breast problem|breast
Procedure|Therapeutic or Preventive Procedure|Impression|3317,3323|true|false|false|C0191838|Procedures on breast|breast
Finding|Pathologic Function|Impression|3317,3332|true|false|false|C0342095|Breast hematoma|breast hematoma
Event|Event|Impression|3324,3332|true|false|false|||hematoma
Finding|Pathologic Function|Impression|3324,3332|true|false|false|C0018944|Hematoma|hematoma
Event|Event|Impression|3342,3350|true|false|false|||evidence
Finding|Idea or Concept|Impression|3342,3350|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Impression|3342,3353|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Event|Event|Impression|3362,3367|true|false|false|||bleed
Finding|Pathologic Function|Impression|3362,3367|true|false|false|C0019080|Hemorrhage|bleed
Event|Event|Impression|3378,3382|false|false|false|||note
Event|Event|Impression|3384,3390|false|false|false|||timing
Finding|Intellectual Product|Impression|3384,3390|false|false|false|C1704250|Timing, LOINC Axis 3|timing
Event|Event|Impression|3395,3405|false|false|false|||suboptimal
Finding|Body Substance|Impression|3413,3420|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Impression|3413,3420|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Impression|3413,3420|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Impression|3421,3427|false|false|false|||needed
Event|Event|Impression|3446,3449|false|false|false|||due
Finding|Functional Concept|Impression|3446,3449|false|false|false|C0678226;C3146286|Due;Due to|due
Finding|Idea or Concept|Impression|3446,3449|false|false|false|C0678226;C3146286|Due;Due to|due
Finding|Idea or Concept|Impression|3454,3464|false|false|false|C1548386|Document Completion - incomplete|incomplete
Event|Event|Impression|3465,3470|false|false|false|||field
Finding|Conceptual Entity|Impression|3465,3470|false|false|false|C1521738;C2346620;C2349184|Field;Force Field;Knowledge Field|field
Procedure|Health Care Activity|Impression|3465,3470|false|false|false|C1553496|field - patient encounter|field
Finding|Idea or Concept|Impression|3482,3489|false|false|false|C1555582|Initial (abbreviation)|initial
Event|Event|Impression|3490,3496|false|false|false|||images
Event|Event|Impression|3512,3519|false|false|false|||density
Event|Event|Impression|3528,3538|false|false|false|||collection
Finding|Conceptual Entity|Impression|3528,3538|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|Impression|3528,3538|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|Impression|3528,3538|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|Impression|3528,3538|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Event|Event|Impression|3543,3552|false|false|false|||unchanged
Finding|Finding|Impression|3543,3552|false|false|false|C0442739||unchanged
Event|Event|Hospital Course|3626,3634|false|false|false|||admitted
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|3643,3649|false|false|false|C0006141|Breast|breast
Disorder|Neoplastic Process|Hospital Course|3643,3649|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|breast
Event|Event|Hospital Course|3643,3649|false|false|false|||breast
Finding|Finding|Hospital Course|3643,3649|false|false|false|C0567499|Breast problem|breast
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3643,3649|false|false|false|C0191838|Procedures on breast|breast
Event|Occupational Activity|Hospital Course|3650,3657|false|false|false|C0557854|Services|service
Finding|Idea or Concept|Hospital Course|3650,3657|false|false|false|C3245478|ActInformationPrivacyReason - service|service
Finding|Functional Concept|Hospital Course|3670,3674|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|3670,3681|false|false|false|C0222601|Left breast|left breast
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3670,3692|false|false|true|C2140215|Lumpectomy of left breast|left breast lumpectomy
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|3675,3681|false|false|false|C0006141|Breast|breast
Disorder|Neoplastic Process|Hospital Course|3675,3681|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|breast
Finding|Finding|Hospital Course|3675,3681|false|false|false|C0567499|Breast problem|breast
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3675,3681|false|false|false|C0191838|Procedures on breast|breast
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3675,3692|false|false|true|C0851238|Lumpectomy of breast|breast lumpectomy
Event|Event|Hospital Course|3682,3692|false|false|false|||lumpectomy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3682,3692|false|false|false|C0851238;C1262070|Excision of mass (procedure);Lumpectomy of breast|lumpectomy
Disorder|Neoplastic Process|Hospital Course|3707,3716|false|false|false|C0007097|Carcinoma|carcinoma
Event|Event|Hospital Course|3707,3716|false|false|false|||carcinoma
Event|Event|Hospital Course|3739,3748|false|false|false|||presented
Event|Event|Hospital Course|3756,3765|false|false|false|||recurrent
Finding|Functional Concept|Hospital Course|3767,3771|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|3767,3778|false|false|false|C0222601|Left breast|left breast
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|3772,3778|false|false|false|C0006141|Breast|breast
Disorder|Neoplastic Process|Hospital Course|3772,3778|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|breast
Event|Event|Hospital Course|3772,3778|false|false|false|||breast
Finding|Finding|Hospital Course|3772,3778|false|false|false|C0567499|Breast problem|breast
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3772,3778|false|false|false|C0191838|Procedures on breast|breast
Finding|Pathologic Function|Hospital Course|3772,3787|false|false|false|C0342095|Breast hematoma|breast hematoma
Event|Event|Hospital Course|3779,3787|false|false|false|||hematoma
Finding|Pathologic Function|Hospital Course|3779,3787|false|false|false|C0018944|Hematoma|hematoma
Event|Event|Hospital Course|3801,3810|false|false|false|||evacuated
Finding|Intellectual Product|Hospital Course|3814,3820|false|false|false|C1546717||needle
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3814,3831|false|false|false|C2243017||needle aspiration
Disorder|Injury or Poisoning|Hospital Course|3821,3831|false|false|false|C1720922|Respiratory Aspiration|aspiration
Event|Event|Hospital Course|3821,3831|false|false|false|||aspiration
Finding|Finding|Hospital Course|3821,3831|false|false|false|C0220787;C0700198;C2712334|Aspiration into respiratory tract;Endotracheal aspiration;Pulmonary aspiration|aspiration
Finding|Organ or Tissue Function|Hospital Course|3821,3831|false|false|false|C0220787;C0700198;C2712334|Aspiration into respiratory tract;Endotracheal aspiration;Pulmonary aspiration|aspiration
Finding|Pathologic Function|Hospital Course|3821,3831|false|false|false|C0220787;C0700198;C2712334|Aspiration into respiratory tract;Endotracheal aspiration;Pulmonary aspiration|aspiration
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3821,3831|false|false|false|C0349707||aspiration
Event|Event|Hospital Course|3859,3867|false|false|false|||admitted
Event|Event|Hospital Course|3872,3883|false|false|false|||observation
Finding|Finding|Hospital Course|3872,3883|false|false|false|C0478530;C1548358;C1554188;C5890437|Examination and observation for unspecified reason;Observation (finding)|observation
Finding|Idea or Concept|Hospital Course|3872,3883|false|false|false|C0478530;C1548358;C1554188;C5890437|Examination and observation for unspecified reason;Observation (finding)|observation
Procedure|Diagnostic Procedure|Hospital Course|3872,3883|false|false|false|C0302523;C0700325;C1964257|Observation - diagnostic procedure;Observation in research;Patient observation|observation
Procedure|Health Care Activity|Hospital Course|3872,3883|false|false|false|C0302523;C0700325;C1964257|Observation - diagnostic procedure;Observation in research;Patient observation|observation
Procedure|Research Activity|Hospital Course|3872,3883|false|false|false|C0302523;C0700325;C1964257|Observation - diagnostic procedure;Observation in research;Patient observation|observation
Procedure|Health Care Activity|Hospital Course|3889,3897|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3889,3897|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Event|Event|Hospital Course|3898,3908|false|false|false|||evacuation
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3898,3908|false|false|false|C1282573|Evacuation procedure|evacuation
Event|Event|Hospital Course|3916,3924|false|false|false|||hematoma
Finding|Pathologic Function|Hospital Course|3916,3924|false|false|false|C0018944|Hematoma|hematoma
Event|Event|Hospital Course|3943,3950|false|false|false|||brought
Finding|Finding|Hospital Course|3958,3967|false|false|false|C4738506|Operating|operating
Event|Event|Hospital Course|3977,3987|false|false|false|||evacuation
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3977,3987|false|false|false|C1282573|Evacuation procedure|evacuation
Finding|Functional Concept|Hospital Course|3996,4000|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Event|Event|Hospital Course|4005,4013|false|false|false|||hematoma
Finding|Pathologic Function|Hospital Course|4005,4013|false|false|false|C0018944|Hematoma|hematoma
Event|Event|Hospital Course|4018,4027|false|false|false|||placement
Procedure|Health Care Activity|Hospital Course|4018,4027|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4018,4027|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Health Care Activity|Hospital Course|4033,4041|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4033,4041|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Drug|Substance|Hospital Course|4042,4047|false|false|false|C1550628|Drain - SpecimenType|drain
Event|Event|Hospital Course|4042,4047|false|false|false|||drain
Finding|Intellectual Product|Hospital Course|4042,4047|false|false|false|C1546604|Drain Specimen Code|drain
Finding|Idea or Concept|Hospital Course|4050,4058|false|false|false|C1547192|Organization unit type - Hospital|Hospital
Attribute|Clinical Attribute|Hospital Course|4050,4065|false|false|false|C0488549||Hospital course
Finding|Finding|Hospital Course|4050,4065|false|false|false|C0489547|Hospital course|Hospital course
Event|Event|Hospital Course|4059,4065|false|false|false|||course
Event|Event|Hospital Course|4069,4077|false|false|false|||detailed
Attribute|Clinical Attribute|Hospital Course|4093,4097|false|false|false|C2598155||pain
Event|Event|Hospital Course|4093,4097|false|false|false|||pain
Finding|Functional Concept|Hospital Course|4093,4097|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|4093,4097|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|4102,4112|false|false|false|||controlled
Anatomy|Body Space or Junction|Hospital Course|4118,4122|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|4118,4122|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|4118,4122|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|4118,4122|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Sign or Symptom|Hospital Course|4118,4127|false|false|false|C0221776|Oral pain|oral pain
Attribute|Clinical Attribute|Hospital Course|4123,4127|false|false|false|C2598155||pain
Event|Event|Hospital Course|4123,4127|false|false|false|||pain
Finding|Functional Concept|Hospital Course|4123,4127|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|4123,4127|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Pharmacologic Substance|Hospital Course|4128,4138|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Hospital Course|4128,4138|false|false|false|||medication
Finding|Intellectual Product|Hospital Course|4128,4138|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Drug|Organic Chemical|Hospital Course|4150,4163|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Drug|Pharmacologic Substance|Hospital Course|4150,4163|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Event|Event|Hospital Course|4150,4163|false|false|false|||acetaminophen
Procedure|Laboratory Procedure|Hospital Course|4150,4163|false|false|false|C0373527|Acetaminophen measurement|acetaminophen
Drug|Organic Chemical|Hospital Course|4168,4176|false|false|false|C0040610|tramadol|tramadol
Drug|Pharmacologic Substance|Hospital Course|4168,4176|false|false|false|C0040610|tramadol|tramadol
Event|Event|Hospital Course|4168,4176|false|false|false|||tramadol
Procedure|Laboratory Procedure|Hospital Course|4168,4176|false|false|false|C1266765|Tramadol measurement (procedure)|tramadol
Drug|Food|Hospital Course|4185,4190|false|false|false|C1875856|Vital High Nitrogen Enteral Nutrition|Vital
Attribute|Clinical Attribute|Hospital Course|4185,4196|false|false|false|C0488614;C0518766|Vital signs|Vital signs
Procedure|Health Care Activity|Hospital Course|4185,4196|false|false|false|C0150404|Taking vital signs|Vital signs
Event|Event|Hospital Course|4191,4196|false|false|false|||signs
Finding|Finding|Hospital Course|4191,4196|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|Hospital Course|4191,4196|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Event|Event|Hospital Course|4202,4211|false|false|false|||monitored
Finding|Finding|Hospital Course|4212,4224|false|false|false|C1698058;C5551028|On Protocol Therapy;per protocol|per protocol
Finding|Functional Concept|Hospital Course|4212,4224|false|false|false|C1698058;C5551028|On Protocol Therapy;per protocol|per protocol
Event|Event|Hospital Course|4216,4224|false|false|false|||protocol
Finding|Finding|Hospital Course|4216,4224|false|false|false|C0442711;C1507394;C1522729;C2348563;C3715209|Clinical trial protocol document;Library Protocol;Protocol - answer to question;Protocols documentation;Study Protocol|protocol
Finding|Intellectual Product|Hospital Course|4216,4224|false|false|false|C0442711;C1507394;C1522729;C2348563;C3715209|Clinical trial protocol document;Library Protocol;Protocol - answer to question;Protocols documentation;Study Protocol|protocol
Event|Event|Hospital Course|4234,4243|false|false|false|||continued
Finding|Idea or Concept|Hospital Course|4252,4256|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|4252,4256|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|4252,4256|false|false|false|C1553498|home health encounter|home
Attribute|Clinical Attribute|Hospital Course|4257,4268|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Hospital Course|4257,4268|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Hospital Course|4257,4268|false|false|false|||medications
Finding|Intellectual Product|Hospital Course|4257,4268|false|false|false|C4284232|Medications|medications
Attribute|Clinical Attribute|Hospital Course|4272,4276|false|false|false|C0231832|Respiratory rate|Resp
Disorder|Disease or Syndrome|Hospital Course|4272,4276|false|false|false|C0851355|Respiratory, thoracic and mediastinal disorders|Resp
Event|Event|Hospital Course|4272,4276|false|false|false|||Resp
Event|Event|Hospital Course|4286,4295|false|false|false|||continued
Finding|Idea or Concept|Hospital Course|4303,4307|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|4303,4307|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|4303,4307|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Hospital Course|4308,4317|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|Hospital Course|4308,4317|false|false|false|C0001927|albuterol|albuterol
Attribute|Clinical Attribute|Hospital Course|4318,4329|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Hospital Course|4318,4329|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Hospital Course|4318,4329|false|false|false|||medications
Finding|Intellectual Product|Hospital Course|4318,4329|false|false|false|C4284232|Medications|medications
Event|Event|Hospital Course|4331,4334|false|false|false|||FEN
Event|Event|Hospital Course|4347,4356|false|false|false|||continued
Finding|Daily or Recreational Activity|Hospital Course|4362,4374|false|false|false|C0184625||regular diet
Drug|Food|Hospital Course|4370,4374|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|Hospital Course|4370,4374|false|false|false|||diet
Finding|Functional Concept|Hospital Course|4370,4374|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|Hospital Course|4370,4374|false|false|false|C0012159|Diet therapy|diet
Event|Event|Hospital Course|4391,4400|false|false|false|||admission
Procedure|Health Care Activity|Hospital Course|4391,4400|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|Hospital Course|4423,4426|false|false|false|||NPO
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4423,4426|false|false|false|C0419179|NPO - Nothing by mouth|NPO
Finding|Finding|Hospital Course|4435,4444|false|false|false|C4738506|Operating|operating
Event|Event|Hospital Course|4455,4463|false|false|false|||hydrated
Drug|Substance|Hospital Course|4472,4478|false|false|false|C0302908|Liquid substance|fluids
Event|Event|Hospital Course|4472,4478|false|false|false|||fluids
Finding|Body Substance|Hospital Course|4472,4478|false|false|false|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4472,4478|false|false|false|C0016286|Fluid Therapy|fluids
Event|Event|Hospital Course|4500,4506|false|false|false|||period
Finding|Organism Function|Hospital Course|4500,4506|false|false|false|C0025344|Menstruation|period
Procedure|Research Activity|Hospital Course|4500,4506|false|false|false|C2347804|Clinical Trial Period|period
Event|Event|Hospital Course|4518,4524|true|false|false|||voided
Event|Activity|Hospital Course|4533,4538|true|false|false|C5966184|Issue (action)|issue
Event|Event|Hospital Course|4533,4538|true|false|false|||issue
Finding|Finding|Hospital Course|4533,4538|true|false|false|C0033213;C1706387|Issue (document);Problem|issue
Finding|Intellectual Product|Hospital Course|4533,4538|true|false|false|C0033213;C1706387|Issue (document);Problem|issue
Finding|Idea or Concept|Hospital Course|4554,4562|true|false|false|C1547192|Organization unit type - Hospital|hospital
Attribute|Clinical Attribute|Hospital Course|4554,4569|true|false|false|C0488549||hospital course
Finding|Finding|Hospital Course|4554,4569|true|false|false|C0489547|Hospital course|hospital course
Event|Event|Hospital Course|4563,4569|true|false|false|||course
Drug|Biologically Active Substance|Hospital Course|4571,4575|false|false|false|C0018966|Heme|Heme
Drug|Organic Chemical|Hospital Course|4571,4575|false|false|false|C0018966|Heme|Heme
Event|Event|Hospital Course|4571,4575|false|false|false|||Heme
Event|Event|Hospital Course|4593,4602|false|false|false|||monitored
Lab|Laboratory or Test Result|Hospital Course|4614,4618|false|false|false|C0587081|Laboratory test finding|labs
Event|Event|Hospital Course|4623,4628|false|false|false|||found
Event|Event|Hospital Course|4636,4642|false|false|false|||stable
Finding|Intellectual Product|Hospital Course|4636,4642|false|false|false|C1547311|Patient Condition Code - Stable|stable
Finding|Idea or Concept|Hospital Course|4648,4652|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|4648,4652|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|4648,4652|false|false|false|C1553498|home health encounter|home
Event|Event|Hospital Course|4653,4668|false|false|false|||anticoagulation
Finding|Finding|Hospital Course|4653,4668|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Finding|Physiologic Function|Hospital Course|4653,4668|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4653,4668|false|false|false|C0003281|Anticoagulation Therapy|anticoagulation
Event|Event|Hospital Course|4673,4677|false|false|false|||held
Event|Event|Hospital Course|4689,4697|false|false|false|||hospital
Finding|Idea or Concept|Hospital Course|4689,4697|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|Hospital Course|4699,4705|false|false|false|||course
Event|Event|Hospital Course|4715,4722|false|false|false|||resumed
Finding|Idea or Concept|Hospital Course|4730,4734|true|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|4730,4734|true|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|4730,4734|true|false|false|C1553498|home health encounter|home
Event|Event|Hospital Course|4735,4739|true|false|false|||dose
Drug|Hazardous or Poisonous Substance|Hospital Course|4743,4751|true|false|false|C0043031|warfarin|warfarin
Drug|Organic Chemical|Hospital Course|4743,4751|true|false|false|C0043031|warfarin|warfarin
Drug|Pharmacologic Substance|Hospital Course|4743,4751|true|false|false|C0043031|warfarin|warfarin
Event|Event|Hospital Course|4743,4751|true|false|false|||warfarin
Event|Event|Hospital Course|4756,4765|true|false|false|||discharge
Finding|Body Substance|Hospital Course|4756,4765|true|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|4756,4765|true|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|4756,4765|true|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|4756,4765|true|false|false|C0030685|Patient Discharge|discharge
Drug|Organic Chemical|Hospital Course|4776,4783|true|false|false|C0728963|Lovenox|lovenox
Drug|Pharmacologic Substance|Hospital Course|4776,4783|true|false|false|C0728963|Lovenox|lovenox
Event|Event|Hospital Course|4784,4790|true|false|false|||bridge
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4784,4790|true|false|false|C0399080|Fixation of dental bridge|bridge
Event|Event|Hospital Course|4796,4804|false|false|false|||remained
Event|Event|Hospital Course|4808,4819|false|false|false|||compression
Finding|Functional Concept|Hospital Course|4808,4819|false|false|false|C0332459;C4551657|Compressed structure|compression
Phenomenon|Natural Phenomenon or Process|Hospital Course|4808,4819|false|false|false|C0728907|Compression|compression
Procedure|Machine Activity|Hospital Course|4808,4819|false|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4808,4819|false|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Event|Event|Hospital Course|4821,4826|false|false|false|||boots
Finding|Idea or Concept|Hospital Course|4838,4846|false|false|false|C1547192|Organization unit type - Hospital|hospital
Attribute|Clinical Attribute|Hospital Course|4838,4853|false|false|false|C0488549||hospital course
Finding|Finding|Hospital Course|4838,4853|false|false|false|C0489547|Hospital course|hospital course
Event|Event|Hospital Course|4847,4853|false|false|false|||course
Event|Event|Hospital Course|4857,4864|false|false|false|||prevent
Disorder|Disease or Syndrome|Hospital Course|4865,4869|false|false|false|C0151950|Deep thrombophlebitis|DVTs
Event|Event|Hospital Course|4865,4869|false|false|false|||DVTs
Drug|Antibiotic|Hospital Course|4890,4895|false|false|false|C0700926|Ancef|ancef
Drug|Organic Chemical|Hospital Course|4890,4895|false|false|false|C0700926|Ancef|ancef
Event|Event|Hospital Course|4903,4908|false|false|false|||Q8hrs
Event|Event|Hospital Course|4913,4924|false|false|false|||prophylaxis
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4913,4924|false|false|false|C0199176|Prophylactic treatment|prophylaxis
Event|Event|Hospital Course|4931,4939|true|false|false|||remained
Event|Event|Hospital Course|4940,4948|true|false|false|||afebrile
Finding|Finding|Hospital Course|4940,4948|true|false|false|C0277797|Apyrexial|afebrile
Event|Event|Hospital Course|4961,4968|true|false|false|||develop
Disorder|Disease or Syndrome|Hospital Course|4971,4983|true|true|false|C0023518|Leukocytosis|leukocytosis
Event|Event|Hospital Course|4971,4983|true|false|false|||leukocytosis
Finding|Finding|Hospital Course|4971,4983|true|true|false|C0750426|Blood leukocyte number above reference range|leukocytosis
Finding|Idea or Concept|Hospital Course|4996,5004|true|false|false|C1547192|Organization unit type - Hospital|hospital
Attribute|Clinical Attribute|Hospital Course|4996,5011|true|false|false|C0488549||hospital course
Finding|Finding|Hospital Course|4996,5011|true|false|false|C0489547|Hospital course|hospital course
Event|Event|Hospital Course|5005,5011|false|false|false|||course
Disorder|Disease or Syndrome|Hospital Course|5015,5019|false|false|false|C0014130;C0014175|Endocrine System Diseases;Endometriosis|Endo
Event|Event|Hospital Course|5015,5019|false|false|false|||Endo
Finding|Gene or Genome|Hospital Course|5015,5019|false|false|false|C1427293|MANEA gene|Endo
Event|Event|Hospital Course|5030,5037|false|false|false|||history
Finding|Conceptual Entity|Hospital Course|5030,5037|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|5030,5037|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Hospital Course|5030,5037|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|5030,5040|false|false|false|C0262926|Medical History|history of
Event|Event|Hospital Course|5041,5050|false|false|false|||metabolic
Finding|Cell Function|Hospital Course|5041,5050|false|false|false|C0311400;C1524026|Metabolic;Metabolic Process, Cellular|metabolic
Finding|Functional Concept|Hospital Course|5041,5050|false|false|false|C0311400;C1524026|Metabolic;Metabolic Process, Cellular|metabolic
Procedure|Diagnostic Procedure|Hospital Course|5041,5050|false|false|false|C4263342|Multisection metabolic|metabolic
Disorder|Disease or Syndrome|Hospital Course|5041,5059|false|false|false|C0524620|Metabolic Syndrome X|metabolic syndrome
Disorder|Disease or Syndrome|Hospital Course|5051,5059|false|false|false|C0039082|Syndrome|syndrome
Event|Event|Hospital Course|5051,5059|false|false|false|||syndrome
Disorder|Disease or Syndrome|Hospital Course|5064,5076|false|false|false|C0362046|Prediabetes syndrome|pre-diabetes
Event|Event|Hospital Course|5086,5090|false|false|false|||kept
Finding|Intellectual Product|Hospital Course|5096,5104|false|false|false|C1720529|Constant - dosing instruction fragment|constant
Drug|Organic Chemical|Hospital Course|5105,5117|false|false|false|C0007004|Carbohydrates|carbohydrate
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5105,5122|false|false|false|C0301577|Carbohydrate diet|carbohydrate diet
Drug|Food|Hospital Course|5118,5122|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|Hospital Course|5118,5122|false|false|false|||diet
Finding|Functional Concept|Hospital Course|5118,5122|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|Hospital Course|5118,5122|false|false|false|C0012159|Diet therapy|diet
Finding|Idea or Concept|Hospital Course|5133,5136|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|5133,5136|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Hospital Course|5140,5149|false|false|false|||discharge
Finding|Body Substance|Hospital Course|5140,5149|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|5140,5149|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|5140,5149|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|5140,5149|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|Hospital Course|5158,5168|false|false|false|||tolerating
Finding|Daily or Recreational Activity|Hospital Course|5171,5183|false|false|false|C0184625||regular diet
Drug|Food|Hospital Course|5179,5183|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|Hospital Course|5179,5183|false|false|false|||diet
Finding|Functional Concept|Hospital Course|5179,5183|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|Hospital Course|5179,5183|false|false|false|C0012159|Diet therapy|diet
Attribute|Clinical Attribute|Hospital Course|5189,5195|false|false|false|C4255480||nausea
Event|Event|Hospital Course|5189,5195|false|false|false|||nausea
Finding|Sign or Symptom|Hospital Course|5189,5195|false|false|false|C0027497|Nausea|nausea
Event|Event|Hospital Course|5199,5205|false|false|false|||emesis
Finding|Body Substance|Hospital Course|5199,5205|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Finding|Physiologic Function|Hospital Course|5199,5205|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Finding|Sign or Symptom|Hospital Course|5199,5205|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Event|Event|Hospital Course|5215,5225|false|false|false|||ambulating
Attribute|Clinical Attribute|Hospital Course|5245,5249|false|false|false|C2598155||pain
Event|Event|Hospital Course|5245,5249|false|false|false|||pain
Finding|Functional Concept|Hospital Course|5245,5249|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|5245,5249|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|5255,5265|false|false|false|||controlled
Anatomy|Body Space or Junction|Hospital Course|5271,5275|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|5271,5275|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|5271,5275|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|5271,5275|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Sign or Symptom|Hospital Course|5271,5280|false|false|false|C0221776|Oral pain|oral pain
Attribute|Clinical Attribute|Hospital Course|5276,5280|false|false|false|C2598155||pain
Event|Event|Hospital Course|5276,5280|false|false|false|||pain
Finding|Functional Concept|Hospital Course|5276,5280|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|5276,5280|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|Hospital Course|5281,5292|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Hospital Course|5281,5292|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Hospital Course|5281,5292|false|false|false|||medications
Finding|Intellectual Product|Hospital Course|5281,5292|false|false|false|C4284232|Medications|medications
Event|Event|Hospital Course|5302,5310|true|false|false|||afebrile
Finding|Finding|Hospital Course|5302,5310|true|false|false|C0277797|Apyrexial|afebrile
Disorder|Disease or Syndrome|Hospital Course|5331,5343|true|true|false|C0023518|Leukocytosis|leukocytosis
Event|Event|Hospital Course|5331,5343|true|false|false|||leukocytosis
Finding|Finding|Hospital Course|5331,5343|true|true|false|C0750426|Blood leukocyte number above reference range|leukocytosis
Drug|Antibiotic|Hospital Course|5349,5360|true|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|Hospital Course|5349,5360|true|false|false|||antibiotics
Event|Event|Hospital Course|5366,5378|false|false|false|||discontinued
Event|Event|Hospital Course|5389,5399|false|false|false|||discharged
Event|Event|Hospital Course|5400,5404|false|false|false|||home
Finding|Idea or Concept|Hospital Course|5400,5404|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|5400,5404|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|5400,5404|false|false|false|C1553498|home health encounter|home
Drug|Substance|Hospital Course|5418,5423|false|false|false|C1550628|Drain - SpecimenType|drain
Finding|Intellectual Product|Hospital Course|5418,5423|false|false|false|C1546604|Drain Specimen Code|drain
Event|Event|Hospital Course|5424,5434|false|false|false|||management
Event|Occupational Activity|Hospital Course|5424,5434|false|false|false|C0001554;C1273870|Administration occupational activities;Management procedure|management
Procedure|Health Care Activity|Hospital Course|5424,5434|false|false|false|C0376636|Disease Management|management
Event|Event|Hospital Course|5439,5444|false|false|false|||close
Finding|Finding|Hospital Course|5439,5444|false|false|false|C0587267;C3810854|Close;Closed|close
Finding|Functional Concept|Hospital Course|5439,5444|false|false|false|C0587267;C3810854|Close;Closed|close
Event|Event|Hospital Course|5446,5452|false|false|false|||follow
Drug|Substance|Hospital Course|5483,5488|false|false|false|C1550628|Drain - SpecimenType|drain
Finding|Intellectual Product|Hospital Course|5483,5488|false|false|false|C1546604|Drain Specimen Code|drain
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5483,5496|false|false|false|C0411815|Removal of drain|drain removal
Event|Activity|Hospital Course|5489,5496|false|false|false|C1883720|Removing (action)|removal
Event|Event|Hospital Course|5489,5496|false|false|false|||removal
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5489,5496|false|false|false|C0015252;C0185115;C0728940|Excision;Extraction;removal technique|removal
Event|Event|Hospital Course|5513,5519|false|false|false|||follow
Event|Event|Hospital Course|5564,5571|false|false|false|||routine
Finding|Idea or Concept|Hospital Course|5564,5571|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|routine
Finding|Intellectual Product|Hospital Course|5564,5571|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|routine
Procedure|Laboratory Procedure|Hospital Course|5564,5571|false|false|false|C1979801|Routine coag|routine
Event|Event|Hospital Course|5572,5578|false|false|false|||follow
Attribute|Clinical Attribute|Hospital Course|5587,5598|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|5587,5598|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|5587,5598|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|5587,5598|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|5587,5611|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|Hospital Course|5602,5611|false|false|false|||Admission
Procedure|Health Care Activity|Hospital Course|5602,5611|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Finding|Intellectual Product|Hospital Course|5613,5635|false|false|false|C5885264|Active medication list|Active Medication list
Drug|Pharmacologic Substance|Hospital Course|5620,5630|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Event|Event|Hospital Course|5620,5630|false|false|false|||Medication
Finding|Intellectual Product|Hospital Course|5620,5630|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|Hospital Course|5620,5635|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|Hospital Course|5631,5635|false|false|false|||list
Finding|Intellectual Product|Hospital Course|5631,5635|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Attribute|Clinical Attribute|Hospital Course|5649,5660|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|5649,5660|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|5649,5660|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|5649,5660|false|false|false|C4284232|Medications|Medications
Attribute|Clinical Attribute|Hospital Course|5663,5675|false|false|false|C5886759|Prescription (attribute)|Prescription
Event|Event|Hospital Course|5663,5675|false|false|false|||Prescription
Finding|Intellectual Product|Hospital Course|5663,5675|false|false|false|C1521941|prescription document|Prescription
Procedure|Health Care Activity|Hospital Course|5663,5675|false|false|false|C0033080|Prescription (procedure)|Prescription
Drug|Organic Chemical|Hospital Course|5676,5685|false|false|false|C0001927|albuterol|ALBUTEROL
Drug|Pharmacologic Substance|Hospital Course|5676,5685|false|false|false|C0001927|albuterol|ALBUTEROL
Drug|Organic Chemical|Hospital Course|5676,5693|false|false|false|C0543495|albuterol sulfate|ALBUTEROL SULFATE
Drug|Pharmacologic Substance|Hospital Course|5676,5693|false|false|false|C0543495|albuterol sulfate|ALBUTEROL SULFATE
Drug|Element, Ion, or Isotope|Hospital Course|5686,5693|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|SULFATE
Drug|Inorganic Chemical|Hospital Course|5686,5693|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|SULFATE
Drug|Pharmacologic Substance|Hospital Course|5686,5693|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|SULFATE
Event|Event|Hospital Course|5686,5693|false|false|false|||SULFATE
Drug|Organic Chemical|Hospital Course|5696,5705|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|Hospital Course|5696,5705|false|false|false|C0001927|albuterol|albuterol
Event|Event|Hospital Course|5696,5705|false|false|false|||albuterol
Drug|Organic Chemical|Hospital Course|5696,5713|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Pharmacologic Substance|Hospital Course|5696,5713|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Element, Ion, or Isotope|Hospital Course|5706,5713|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Inorganic Chemical|Hospital Course|5706,5713|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Pharmacologic Substance|Hospital Course|5706,5713|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Event|Event|Hospital Course|5706,5713|false|false|false|||sulfate
Drug|Biomedical or Dental Material|Hospital Course|5736,5744|false|false|false|C0037633;C0525069;C1382100|Pharmaceutical Solutions;Solution Dosage Form;Solutions|solution
Drug|Substance|Hospital Course|5736,5744|false|false|false|C0037633;C0525069;C1382100|Pharmaceutical Solutions;Solution Dosage Form;Solutions|solution
Event|Event|Hospital Course|5736,5744|false|false|false|||solution
Finding|Conceptual Entity|Hospital Course|5736,5744|false|false|false|C2699488|Resolution|solution
Event|Event|Hospital Course|5749,5761|false|false|false|||nebulization
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5749,5761|false|false|false|C1659427|nebulization-mediated drug administration|nebulization
Disorder|Disease or Syndrome|Hospital Course|5784,5789|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|Hospital Course|5792,5795|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|5792,5795|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Hospital Course|5799,5805|false|false|false|||needed
Drug|Organic Chemical|Hospital Course|5810,5815|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|Hospital Course|5810,5815|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|Hospital Course|5810,5815|false|false|false|||cough
Finding|Sign or Symptom|Hospital Course|5810,5815|false|false|false|C0010200|Coughing|cough
Event|Event|Hospital Course|5817,5823|false|false|false|||wheeze
Finding|Sign or Symptom|Hospital Course|5817,5823|false|false|false|C0043144|Wheezing|wheeze
Drug|Organic Chemical|Hospital Course|5824,5833|false|false|false|C0001927|albuterol|ALBUTEROL
Drug|Pharmacologic Substance|Hospital Course|5824,5833|false|false|false|C0001927|albuterol|ALBUTEROL
Drug|Organic Chemical|Hospital Course|5824,5841|false|false|false|C0543495|albuterol sulfate|ALBUTEROL SULFATE
Drug|Pharmacologic Substance|Hospital Course|5824,5841|false|false|false|C0543495|albuterol sulfate|ALBUTEROL SULFATE
Drug|Element, Ion, or Isotope|Hospital Course|5834,5841|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|SULFATE
Drug|Inorganic Chemical|Hospital Course|5834,5841|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|SULFATE
Drug|Pharmacologic Substance|Hospital Course|5834,5841|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|SULFATE
Drug|Organic Chemical|Hospital Course|5843,5849|false|false|false|C0162684;C1739179|Pro-Air Procaterol;ProAir|PROAIR
Drug|Pharmacologic Substance|Hospital Course|5843,5849|false|false|false|C0162684;C1739179|Pro-Air Procaterol;ProAir|PROAIR
Drug|Organic Chemical|Hospital Course|5843,5853|false|false|false|C1739179|ProAir|PROAIR HFA
Drug|Pharmacologic Substance|Hospital Course|5843,5853|false|false|false|C1739179|ProAir|PROAIR HFA
Disorder|Disease or Syndrome|Hospital Course|5850,5853|false|false|false|C0015458|Facial Hemiatrophy|HFA
Event|Event|Hospital Course|5850,5853|false|false|false|||HFA
Procedure|Diagnostic Procedure|Hospital Course|5850,5853|false|false|false|C0430649|High frequency audiometry|HFA
Drug|Organic Chemical|Hospital Course|5857,5863|false|false|false|C0162684;C1739179|Pro-Air Procaterol;ProAir|ProAir
Drug|Pharmacologic Substance|Hospital Course|5857,5863|false|false|false|C0162684;C1739179|Pro-Air Procaterol;ProAir|ProAir
Drug|Organic Chemical|Hospital Course|5857,5867|false|false|false|C1739179|ProAir|ProAir HFA
Drug|Pharmacologic Substance|Hospital Course|5857,5867|false|false|false|C1739179|ProAir|ProAir HFA
Disorder|Disease or Syndrome|Hospital Course|5864,5867|false|false|false|C0015458|Facial Hemiatrophy|HFA
Event|Event|Hospital Course|5864,5867|false|false|false|||HFA
Procedure|Diagnostic Procedure|Hospital Course|5864,5867|false|false|false|C0430649|High frequency audiometry|HFA
Drug|Biomedical or Dental Material|Hospital Course|5885,5892|false|false|false|C1112870|Aerosol Dose Form|aerosol
Event|Event|Hospital Course|5910,5920|false|false|false|||inhalation
Finding|Functional Concept|Hospital Course|5910,5920|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Finding|Organism Function|Hospital Course|5910,5920|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Event|Event|Hospital Course|5935,5941|false|false|false|||needed
Drug|Organic Chemical|Hospital Course|5946,5951|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|Hospital Course|5946,5951|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|Hospital Course|5946,5951|false|false|false|||cough
Finding|Sign or Symptom|Hospital Course|5946,5951|false|false|false|C0010200|Coughing|cough
Event|Event|Hospital Course|5952,5958|false|false|false|||wheeze
Finding|Sign or Symptom|Hospital Course|5952,5958|false|false|false|C0043144|Wheezing|wheeze
Drug|Organic Chemical|Hospital Course|5959,5971|false|false|false|C0286651|atorvastatin|ATORVASTATIN
Drug|Pharmacologic Substance|Hospital Course|5959,5971|false|false|false|C0286651|atorvastatin|ATORVASTATIN
Drug|Organic Chemical|Hospital Course|5974,5986|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|Hospital Course|5974,5986|false|false|false|C0286651|atorvastatin|atorvastatin
Event|Event|Hospital Course|5974,5986|false|false|false|||atorvastatin
Drug|Biomedical or Dental Material|Hospital Course|6009,6015|false|false|false|C0039225|Tablet Dosage Form|tablet
Event|Event|Hospital Course|6009,6015|false|false|false|||tablet
Anatomy|Body Location or Region|Hospital Course|6022,6027|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|6022,6027|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Event|Event|Hospital Course|6043,6053|false|false|false|||Prescribed
Finding|Functional Concept|Hospital Course|6063,6071|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|Provider
Finding|Intellectual Product|Hospital Course|6063,6071|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|Provider
Event|Event|Hospital Course|6078,6088|true|false|false|||adjustment
Finding|Classification|Hospital Course|6078,6088|true|false|false|C0376209;C0456081;C0678219;C0683269;C1546424|Adjustment - classification term;Personal Adjustment;Psychological adjustment;Transaction Type - Adjustment|adjustment
Finding|Functional Concept|Hospital Course|6078,6088|true|false|false|C0376209;C0456081;C0678219;C0683269;C1546424|Adjustment - classification term;Personal Adjustment;Psychological adjustment;Transaction Type - Adjustment|adjustment
Finding|Idea or Concept|Hospital Course|6078,6088|true|false|false|C0376209;C0456081;C0678219;C0683269;C1546424|Adjustment - classification term;Personal Adjustment;Psychological adjustment;Transaction Type - Adjustment|adjustment
Finding|Individual Behavior|Hospital Course|6078,6088|true|false|false|C0376209;C0456081;C0678219;C0683269;C1546424|Adjustment - classification term;Personal Adjustment;Psychological adjustment;Transaction Type - Adjustment|adjustment
Finding|Finding|Hospital Course|6094,6097|true|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Hospital Course|6094,6097|true|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Drug|Organic Chemical|Hospital Course|6102,6112|false|false|false|C0206460|enoxaparin|ENOXAPARIN
Drug|Pharmacologic Substance|Hospital Course|6102,6112|false|false|false|C0206460|enoxaparin|ENOXAPARIN
Event|Event|Hospital Course|6102,6112|false|false|false|||ENOXAPARIN
Drug|Organic Chemical|Hospital Course|6115,6125|false|false|false|C0206460|enoxaparin|enoxaparin
Drug|Pharmacologic Substance|Hospital Course|6115,6125|false|false|false|C0206460|enoxaparin|enoxaparin
Event|Event|Hospital Course|6115,6125|false|false|false|||enoxaparin
Finding|Functional Concept|Hospital Course|6136,6148|false|false|false|C1522438|Subcutaneous Route of Administration|subcutaneous
Event|Event|Hospital Course|6149,6156|false|false|false|||syringe
Event|Event|Hospital Course|6216,6221|false|false|false|||start
Event|Event|Hospital Course|6250,6260|false|false|false|||Prescribed
Finding|Functional Concept|Hospital Course|6270,6278|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|Provider
Finding|Intellectual Product|Hospital Course|6270,6278|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|Provider
Event|Event|Hospital Course|6285,6295|true|false|false|||adjustment
Finding|Classification|Hospital Course|6285,6295|true|false|false|C0376209;C0456081;C0678219;C0683269;C1546424|Adjustment - classification term;Personal Adjustment;Psychological adjustment;Transaction Type - Adjustment|adjustment
Finding|Functional Concept|Hospital Course|6285,6295|true|false|false|C0376209;C0456081;C0678219;C0683269;C1546424|Adjustment - classification term;Personal Adjustment;Psychological adjustment;Transaction Type - Adjustment|adjustment
Finding|Idea or Concept|Hospital Course|6285,6295|true|false|false|C0376209;C0456081;C0678219;C0683269;C1546424|Adjustment - classification term;Personal Adjustment;Psychological adjustment;Transaction Type - Adjustment|adjustment
Finding|Individual Behavior|Hospital Course|6285,6295|true|false|false|C0376209;C0456081;C0678219;C0683269;C1546424|Adjustment - classification term;Personal Adjustment;Psychological adjustment;Transaction Type - Adjustment|adjustment
Finding|Finding|Hospital Course|6301,6304|true|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Hospital Course|6301,6304|true|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Drug|Antibiotic|Hospital Course|6309,6321|false|false|false|C0014806|erythromycin|ERYTHROMYCIN
Drug|Organic Chemical|Hospital Course|6309,6321|false|false|false|C0014806|erythromycin|ERYTHROMYCIN
Event|Event|Hospital Course|6309,6321|false|false|false|||ERYTHROMYCIN
Drug|Antibiotic|Hospital Course|6324,6336|false|false|false|C0014806|erythromycin|erythromycin
Drug|Organic Chemical|Hospital Course|6324,6336|false|false|false|C0014806|erythromycin|erythromycin
Event|Event|Hospital Course|6324,6336|false|false|false|||erythromycin
Anatomy|Body Location or Region|Hospital Course|6355,6358|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|eye
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6355,6358|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|eye
Disorder|Disease or Syndrome|Hospital Course|6355,6358|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|eye
Disorder|Neoplastic Process|Hospital Course|6355,6358|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|eye
Finding|Body Substance|Hospital Course|6355,6358|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Finding|Hospital Course|6355,6358|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Intellectual Product|Hospital Course|6355,6358|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Drug|Biomedical or Dental Material|Hospital Course|6355,6367|false|false|false|C0304651|Ophthalmic Ointment|eye ointment
Drug|Biomedical or Dental Material|Hospital Course|6359,6367|false|false|false|C0028912|Ointments|ointment
Event|Event|Hospital Course|6359,6367|false|false|false|||ointment
Finding|Functional Concept|Hospital Course|6370,6375|false|false|false|C1632850;C1879355;C4048755;C4521676|Apply;Apply (administration method);Apply (instruction)|Apply
Anatomy|Body Location or Region|Hospital Course|6394,6397|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|eye
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6394,6397|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|eye
Disorder|Disease or Syndrome|Hospital Course|6394,6397|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|eye
Disorder|Neoplastic Process|Hospital Course|6394,6397|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|eye
Finding|Body Substance|Hospital Course|6394,6397|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Finding|Hospital Course|6394,6397|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Intellectual Product|Hospital Course|6394,6397|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Disorder|Disease or Syndrome|Hospital Course|6403,6408|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|Hospital Course|6411,6414|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|6411,6414|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|Hospital Course|6415,6425|false|false|false|C0016860|furosemide|FUROSEMIDE
Drug|Pharmacologic Substance|Hospital Course|6415,6425|false|false|false|C0016860|furosemide|FUROSEMIDE
Event|Event|Hospital Course|6415,6425|false|false|false|||FUROSEMIDE
Drug|Organic Chemical|Hospital Course|6428,6438|false|false|false|C0016860|furosemide|furosemide
Drug|Pharmacologic Substance|Hospital Course|6428,6438|false|false|false|C0016860|furosemide|furosemide
Event|Event|Hospital Course|6428,6438|false|false|false|||furosemide
Drug|Biomedical or Dental Material|Hospital Course|6445,6451|false|false|false|C0039225|Tablet Dosage Form|tablet
Drug|Biomedical or Dental Material|Hospital Course|6457,6463|false|false|false|C0039225|Tablet Dosage Form|tablet
Event|Event|Hospital Course|6457,6463|false|false|false|||tablet
Finding|Functional Concept|Hospital Course|6467,6475|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|6470,6475|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|6470,6475|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Intellectual Product|Hospital Course|6476,6480|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|Hospital Course|6476,6486|false|false|false|C3537736|Once A Day|once a day
Event|Event|Hospital Course|6483,6486|false|false|false|||day
Finding|Idea or Concept|Hospital Course|6483,6486|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|6483,6486|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Hospital Course|6490,6496|false|false|false|||needed
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6501,6504|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Finding|Pathologic Function|Hospital Course|6501,6513|false|false|false|C0581394|Swelling of lower limb|leg swelling
Event|Event|Hospital Course|6505,6513|false|false|false|||swelling
Finding|Finding|Hospital Course|6505,6513|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|Hospital Course|6505,6513|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Drug|Organic Chemical|Hospital Course|6514,6527|false|false|false|C0012306|hydromorphone|HYDROMORPHONE
Drug|Pharmacologic Substance|Hospital Course|6514,6527|false|false|false|C0012306|hydromorphone|HYDROMORPHONE
Event|Event|Hospital Course|6514,6527|false|false|false|||HYDROMORPHONE
Drug|Organic Chemical|Hospital Course|6530,6543|false|false|false|C0012306|hydromorphone|hydromorphone
Drug|Pharmacologic Substance|Hospital Course|6530,6543|false|false|false|C0012306|hydromorphone|hydromorphone
Event|Event|Hospital Course|6530,6543|false|false|false|||hydromorphone
Drug|Biomedical or Dental Material|Hospital Course|6549,6555|false|false|false|C0039225|Tablet Dosage Form|tablet
Drug|Biomedical or Dental Material|Hospital Course|6561,6567|false|false|false|C0039225|Tablet Dosage Form|tablet
Event|Event|Hospital Course|6561,6567|false|false|false|||tablet
Anatomy|Body Location or Region|Hospital Course|6574,6579|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|6574,6579|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Event|Event|Hospital Course|6604,6610|true|false|false|||needed
Finding|Finding|Hospital Course|6615,6621|true|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|Hospital Course|6615,6621|true|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Finding|Hospital Course|6615,6626|true|false|false|C0278140;C4050465;C4521229|Neck Pain Score 6;Severe Extremity Pain;Severe pain|severe pain
Attribute|Clinical Attribute|Hospital Course|6622,6626|true|false|false|C2598155||pain
Event|Event|Hospital Course|6622,6626|true|false|false|||pain
Finding|Functional Concept|Hospital Course|6622,6626|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|6622,6626|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Food|Hospital Course|6635,6640|true|false|false|C0452428|Drink (dietary substance)|drink
Event|Event|Hospital Course|6635,6640|true|false|false|||drink
Drug|Organic Chemical|Hospital Course|6641,6648|true|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Drug|Pharmacologic Substance|Hospital Course|6641,6648|true|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Event|Event|Hospital Course|6641,6648|true|false|false|||alcohol
Finding|Intellectual Product|Hospital Course|6641,6648|true|false|false|C1547288|Alcohol - Recreational Drug Use Code|alcohol
Event|Event|Hospital Course|6652,6657|true|false|false|||drive
Event|Event|Hospital Course|6664,6670|false|false|false|||taking
Drug|Pharmacologic Substance|Hospital Course|6676,6686|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Hospital Course|6676,6686|false|false|false|||medication
Finding|Intellectual Product|Hospital Course|6676,6686|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|Hospital Course|6701,6711|false|false|false|||COMPRESSOR
Drug|Biomedical or Dental Material|Hospital Course|6732,6738|false|false|false|C5671121|System (basic dose form)|SYSTEM
Event|Event|Hospital Course|6732,6738|false|false|false|||SYSTEM
Finding|Functional Concept|Hospital Course|6732,6738|false|false|false|C0449913;C5441654|System;System, LOINC Axis 4|SYSTEM
Drug|Biomedical or Dental Material|Hospital Course|6761,6767|false|false|false|C5671121|System (basic dose form)|System
Event|Event|Hospital Course|6761,6767|false|false|false|||System
Finding|Functional Concept|Hospital Course|6761,6767|false|false|false|C0449913;C5441654|System;System, LOINC Axis 4|System
Event|Event|Hospital Course|6769,6772|false|false|false|||Use
Finding|Functional Concept|Hospital Course|6769,6772|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|Use
Finding|Intellectual Product|Hospital Course|6769,6772|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|Use
Drug|Organic Chemical|Hospital Course|6778,6787|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|Hospital Course|6778,6787|false|false|false|C0001927|albuterol|albuterol
Event|Event|Hospital Course|6788,6797|false|false|false|||nebulizer
Disorder|Disease or Syndrome|Hospital Course|6808,6813|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|Hospital Course|6816,6819|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|6816,6819|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Hospital Course|6823,6829|false|false|false|||needed
Drug|Organic Chemical|Hospital Course|6834,6839|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|Hospital Course|6834,6839|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|Hospital Course|6834,6839|false|false|false|||cough
Finding|Sign or Symptom|Hospital Course|6834,6839|false|false|false|C0010200|Coughing|cough
Event|Event|Hospital Course|6840,6846|false|false|false|||wheeze
Finding|Sign or Symptom|Hospital Course|6840,6846|false|false|false|C0043144|Wheezing|wheeze
Drug|Organic Chemical|Hospital Course|6847,6857|false|false|false|C0028978|omeprazole|OMEPRAZOLE
Drug|Pharmacologic Substance|Hospital Course|6847,6857|false|false|false|C0028978|omeprazole|OMEPRAZOLE
Drug|Organic Chemical|Hospital Course|6860,6870|false|false|false|C0028978|omeprazole|omeprazole
Drug|Pharmacologic Substance|Hospital Course|6860,6870|false|false|false|C0028978|omeprazole|omeprazole
Event|Event|Hospital Course|6860,6870|false|false|false|||omeprazole
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6877,6884|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Anatomy|Cell Component|Hospital Course|6877,6884|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Drug|Biomedical or Dental Material|Hospital Course|6877,6884|false|false|false|C0006935|capsule (pharmacologic)|capsule
Event|Event|Hospital Course|6893,6900|false|false|false|||release
Finding|Functional Concept|Hospital Course|6893,6900|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|release
Procedure|Health Care Activity|Hospital Course|6893,6900|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6893,6900|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|release
Event|Event|Hospital Course|6902,6906|false|false|false|||TAKE
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6909,6916|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|CAPSULE
Anatomy|Cell Component|Hospital Course|6909,6916|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|CAPSULE
Drug|Biomedical or Dental Material|Hospital Course|6909,6916|false|false|false|C0006935|capsule (pharmacologic)|CAPSULE
Anatomy|Body Location or Region|Hospital Course|6933,6949|false|false|false|C0744316|gastroesophageal|GASTROESOPHAGEAL
Drug|Organic Chemical|Hospital Course|6964,6974|false|false|false|C0074393|sertraline|SERTRALINE
Drug|Pharmacologic Substance|Hospital Course|6964,6974|false|false|false|C0074393|sertraline|SERTRALINE
Event|Event|Hospital Course|6964,6974|false|false|false|||SERTRALINE
Drug|Organic Chemical|Hospital Course|6977,6987|false|false|false|C0074393|sertraline|sertraline
Drug|Pharmacologic Substance|Hospital Course|6977,6987|false|false|false|C0074393|sertraline|sertraline
Event|Event|Hospital Course|6977,6987|false|false|false|||sertraline
Drug|Biomedical or Dental Material|Hospital Course|6995,7001|false|false|false|C0039225|Tablet Dosage Form|tablet
Event|Event|Hospital Course|6995,7001|false|false|false|||tablet
Drug|Biomedical or Dental Material|Hospital Course|7007,7013|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|Hospital Course|7017,7025|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|7020,7025|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|7020,7025|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Intellectual Product|Hospital Course|7026,7030|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|Hospital Course|7026,7036|false|false|false|C3537736|Once A Day|once a day
Event|Event|Hospital Course|7033,7036|false|false|false|||day
Finding|Idea or Concept|Hospital Course|7033,7036|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|7033,7036|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|Hospital Course|7037,7045|false|false|false|C0040610|tramadol|TRAMADOL
Drug|Pharmacologic Substance|Hospital Course|7037,7045|false|false|false|C0040610|tramadol|TRAMADOL
Event|Event|Hospital Course|7037,7045|false|false|false|||TRAMADOL
Procedure|Laboratory Procedure|Hospital Course|7037,7045|false|false|false|C1266765|Tramadol measurement (procedure)|TRAMADOL
Drug|Organic Chemical|Hospital Course|7048,7056|false|false|false|C0040610|tramadol|tramadol
Drug|Pharmacologic Substance|Hospital Course|7048,7056|false|false|false|C0040610|tramadol|tramadol
Event|Event|Hospital Course|7048,7056|false|false|false|||tramadol
Procedure|Laboratory Procedure|Hospital Course|7048,7056|false|false|false|C1266765|Tramadol measurement (procedure)|tramadol
Drug|Biomedical or Dental Material|Hospital Course|7075,7081|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|Hospital Course|7085,7093|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|7088,7093|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|7088,7093|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Disorder|Disease or Syndrome|Hospital Course|7100,7105|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Event|Event|Hospital Course|7100,7105|false|false|false|||times
Finding|Idea or Concept|Hospital Course|7108,7111|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|7108,7111|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|Hospital Course|7112,7121|false|false|false|C0040805|trazodone|TRAZODONE
Drug|Pharmacologic Substance|Hospital Course|7112,7121|false|false|false|C0040805|trazodone|TRAZODONE
Drug|Organic Chemical|Hospital Course|7124,7133|false|false|false|C0040805|trazodone|trazodone
Drug|Pharmacologic Substance|Hospital Course|7124,7133|false|false|false|C0040805|trazodone|trazodone
Event|Event|Hospital Course|7124,7133|false|false|false|||trazodone
Drug|Biomedical or Dental Material|Hospital Course|7150,7156|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|Hospital Course|7160,7168|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|7163,7168|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|7163,7168|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Event|Event|Hospital Course|7172,7179|false|false|false|||bedtime
Event|Event|Hospital Course|7183,7189|false|false|false|||needed
Event|Event|Hospital Course|7194,7201|false|false|false|||insomia
Drug|Hazardous or Poisonous Substance|Hospital Course|7202,7210|false|false|false|C0043031|warfarin|WARFARIN
Drug|Organic Chemical|Hospital Course|7202,7210|false|false|false|C0043031|warfarin|WARFARIN
Drug|Pharmacologic Substance|Hospital Course|7202,7210|false|false|false|C0043031|warfarin|WARFARIN
Event|Event|Hospital Course|7202,7210|false|false|false|||WARFARIN
Drug|Hazardous or Poisonous Substance|Hospital Course|7213,7221|false|false|false|C0043031|warfarin|warfarin
Drug|Organic Chemical|Hospital Course|7213,7221|false|false|false|C0043031|warfarin|warfarin
Drug|Pharmacologic Substance|Hospital Course|7213,7221|false|false|false|C0043031|warfarin|warfarin
Event|Event|Hospital Course|7213,7221|false|false|false|||warfarin
Drug|Biomedical or Dental Material|Hospital Course|7243,7249|false|false|false|C0039225|Tablet Dosage Form|tablet
Event|Event|Hospital Course|7243,7249|false|false|false|||tablet
Finding|Functional Concept|Hospital Course|7253,7261|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|7256,7261|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|7256,7261|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Disorder|Disease or Syndrome|Hospital Course|7264,7269|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Disorder|Disease or Syndrome|Hospital Course|7291,7296|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Event|Event|Hospital Course|7291,7296|false|false|false|||times
Finding|Intellectual Product|Hospital Course|7299,7303|false|false|false|C1561540|Transaction counts and value totals - week|week
Anatomy|Body Location or Region|Hospital Course|7315,7318|false|false|false|C0449201|PER (body structure)|per
Disorder|Disease or Syndrome|Hospital Course|7315,7318|false|false|false|C1861457|PROGRESSIVE ENCEPHALOMYELITIS WITH RIGIDITY|per
Finding|Functional Concept|Hospital Course|7315,7318|false|false|false|C1418464;C1704764;C3273590;C4281991|Follow;PER1 gene;PER1 wt Allele;Per - dosing instruction fragment|per
Finding|Gene or Genome|Hospital Course|7315,7318|false|false|false|C1418464;C1704764;C3273590;C4281991|Follow;PER1 gene;PER1 wt Allele;Per - dosing instruction fragment|per
Finding|Intellectual Product|Hospital Course|7315,7318|false|false|false|C1418464;C1704764;C3273590;C4281991|Follow;PER1 gene;PER1 wt Allele;Per - dosing instruction fragment|per
Event|Event|Hospital Course|7338,7348|false|false|false|||Prescribed
Finding|Functional Concept|Hospital Course|7358,7366|false|true|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|Provider
Finding|Intellectual Product|Hospital Course|7358,7366|false|true|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|Provider
Event|Event|Hospital Course|7373,7383|true|false|false|||adjustment
Finding|Classification|Hospital Course|7373,7383|true|false|false|C0376209;C0456081;C0678219;C0683269;C1546424|Adjustment - classification term;Personal Adjustment;Psychological adjustment;Transaction Type - Adjustment|adjustment
Finding|Functional Concept|Hospital Course|7373,7383|true|false|false|C0376209;C0456081;C0678219;C0683269;C1546424|Adjustment - classification term;Personal Adjustment;Psychological adjustment;Transaction Type - Adjustment|adjustment
Finding|Idea or Concept|Hospital Course|7373,7383|true|false|false|C0376209;C0456081;C0678219;C0683269;C1546424|Adjustment - classification term;Personal Adjustment;Psychological adjustment;Transaction Type - Adjustment|adjustment
Finding|Individual Behavior|Hospital Course|7373,7383|true|false|false|C0376209;C0456081;C0678219;C0683269;C1546424|Adjustment - classification term;Personal Adjustment;Psychological adjustment;Transaction Type - Adjustment|adjustment
Finding|Finding|Hospital Course|7389,7392|true|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Hospital Course|7389,7392|true|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Attribute|Clinical Attribute|Hospital Course|7399,7410|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|7399,7410|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|7399,7410|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|7399,7410|false|false|false|C4284232|Medications|Medications
Drug|Pharmacologic Substance|Hospital Course|7413,7416|false|false|false|C0013231|Drugs, Non-Prescription|OTC
Event|Event|Hospital Course|7413,7416|false|false|false|||OTC
Finding|Gene or Genome|Hospital Course|7413,7416|false|false|false|C1418193|OTC gene|OTC
Drug|Organic Chemical|Hospital Course|7417,7430|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|ACETAMINOPHEN
Drug|Pharmacologic Substance|Hospital Course|7417,7430|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|ACETAMINOPHEN
Event|Event|Hospital Course|7417,7430|false|false|false|||ACETAMINOPHEN
Procedure|Laboratory Procedure|Hospital Course|7417,7430|false|false|false|C0373527|Acetaminophen measurement|ACETAMINOPHEN
Drug|Organic Chemical|Hospital Course|7433,7446|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Drug|Pharmacologic Substance|Hospital Course|7433,7446|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Event|Event|Hospital Course|7433,7446|false|false|false|||acetaminophen
Procedure|Laboratory Procedure|Hospital Course|7433,7446|false|false|false|C0373527|Acetaminophen measurement|acetaminophen
Drug|Biomedical or Dental Material|Hospital Course|7464,7470|false|false|false|C0039225|Tablet Dosage Form|tablet
Anatomy|Body Location or Region|Hospital Course|7478,7483|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|7478,7483|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Finding|Hospital Course|7484,7491|false|false|false|C4035626|3 times|3 times
Disorder|Disease or Syndrome|Hospital Course|7486,7491|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Event|Event|Hospital Course|7486,7491|false|false|false|||times
Event|Event|Hospital Course|7501,7507|false|false|false|||needed
Attribute|Clinical Attribute|Hospital Course|7512,7516|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|7512,7516|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|7512,7516|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Disorder|Congenital Abnormality|Hospital Course|7527,7530|false|false|false|C0026760|Multiple Epiphyseal Dysplasia|med
Finding|Gene or Genome|Hospital Course|7527,7530|false|false|false|C1413596;C1413597;C1419866;C1456376;C1549978;C4321267;C5781216|COL9A2 gene;COL9A3 gene;COMP gene;COMP wt Allele;Master of Education;SCN8A gene;SCN8A wt Allele|med
Finding|Intellectual Product|Hospital Course|7527,7530|false|false|false|C1413596;C1413597;C1419866;C1456376;C1549978;C4321267;C5781216|COL9A2 gene;COL9A3 gene;COMP gene;COMP wt Allele;Master of Education;SCN8A gene;SCN8A wt Allele|med
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7531,7534|false|false|false|C2606415|ZDHHC2 protein, human|rec
Drug|Enzyme|Hospital Course|7531,7534|false|false|false|C2606415|ZDHHC2 protein, human|rec
Finding|Gene or Genome|Hospital Course|7531,7534|false|false|false|C1422148;C1424025|MCM8 gene;RBPJP4 gene|rec
Drug|Organic Chemical|Hospital Course|7536,7551|false|false|false|C0008318|cholecalciferol|CHOLECALCIFEROL
Drug|Pharmacologic Substance|Hospital Course|7536,7551|false|false|false|C0008318|cholecalciferol|CHOLECALCIFEROL
Drug|Vitamin|Hospital Course|7536,7551|false|false|false|C0008318|cholecalciferol|CHOLECALCIFEROL
Event|Event|Hospital Course|7536,7551|false|false|false|||CHOLECALCIFEROL
Drug|Organic Chemical|Hospital Course|7536,7564|false|false|false|C0008318|cholecalciferol|CHOLECALCIFEROL (VITAMIN D3)
Drug|Pharmacologic Substance|Hospital Course|7536,7564|false|false|false|C0008318|cholecalciferol|CHOLECALCIFEROL (VITAMIN D3)
Drug|Vitamin|Hospital Course|7536,7564|false|false|false|C0008318|cholecalciferol|CHOLECALCIFEROL (VITAMIN D3)
Drug|Organic Chemical|Hospital Course|7553,7560|false|false|false|C0042890|Vitamins|VITAMIN
Drug|Pharmacologic Substance|Hospital Course|7553,7560|false|false|false|C0042890|Vitamins|VITAMIN
Drug|Vitamin|Hospital Course|7553,7560|false|false|false|C0042890|Vitamins|VITAMIN
Event|Event|Hospital Course|7553,7560|false|false|false|||VITAMIN
Drug|Organic Chemical|Hospital Course|7553,7563|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|VITAMIN D3
Drug|Pharmacologic Substance|Hospital Course|7553,7563|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|VITAMIN D3
Drug|Vitamin|Hospital Course|7553,7563|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|VITAMIN D3
Drug|Organic Chemical|Hospital Course|7567,7582|false|false|false|C0008318|cholecalciferol|cholecalciferol
Drug|Pharmacologic Substance|Hospital Course|7567,7582|false|false|false|C0008318|cholecalciferol|cholecalciferol
Drug|Vitamin|Hospital Course|7567,7582|false|false|false|C0008318|cholecalciferol|cholecalciferol
Event|Event|Hospital Course|7567,7582|false|false|false|||cholecalciferol
Drug|Organic Chemical|Hospital Course|7567,7595|false|false|false|C0008318|cholecalciferol|cholecalciferol (vitamin D3)
Drug|Pharmacologic Substance|Hospital Course|7567,7595|false|false|false|C0008318|cholecalciferol|cholecalciferol (vitamin D3)
Drug|Vitamin|Hospital Course|7567,7595|false|false|false|C0008318|cholecalciferol|cholecalciferol (vitamin D3)
Drug|Organic Chemical|Hospital Course|7584,7591|false|false|false|C0042890|Vitamins|vitamin
Drug|Pharmacologic Substance|Hospital Course|7584,7591|false|false|false|C0042890|Vitamins|vitamin
Drug|Vitamin|Hospital Course|7584,7591|false|false|false|C0042890|Vitamins|vitamin
Event|Event|Hospital Course|7584,7591|false|false|false|||vitamin
Drug|Organic Chemical|Hospital Course|7584,7594|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Drug|Pharmacologic Substance|Hospital Course|7584,7594|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Drug|Vitamin|Hospital Course|7584,7594|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Drug|Biomedical or Dental Material|Hospital Course|7618,7624|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|Hospital Course|7628,7636|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|7631,7636|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|7631,7636|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Intellectual Product|Hospital Course|7637,7641|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|Hospital Course|7637,7647|false|false|false|C3537736|Once A Day|once a day
Finding|Idea or Concept|Hospital Course|7644,7647|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|7644,7647|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Pharmacologic Substance|Hospital Course|7652,7655|false|false|false|C0013231|Drugs, Non-Prescription|OTC
Event|Event|Hospital Course|7652,7655|false|false|false|||OTC
Finding|Gene or Genome|Hospital Course|7652,7655|false|false|false|C1418193|OTC gene|OTC
Drug|Biomedical or Dental Material|Hospital Course|7657,7669|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|POLYETHYLENE
Drug|Organic Chemical|Hospital Course|7657,7669|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|POLYETHYLENE
Drug|Organic Chemical|Hospital Course|7657,7676|false|false|false|C0032483|polyethylene glycols|POLYETHYLENE GLYCOL
Drug|Pharmacologic Substance|Hospital Course|7657,7676|false|false|false|C0032483|polyethylene glycols|POLYETHYLENE GLYCOL
Drug|Organic Chemical|Hospital Course|7657,7681|false|false|false|C0724672|polyethylene glycol 3350|POLYETHYLENE GLYCOL 3350
Drug|Pharmacologic Substance|Hospital Course|7657,7681|false|false|false|C0724672|polyethylene glycol 3350|POLYETHYLENE GLYCOL 3350
Drug|Hazardous or Poisonous Substance|Hospital Course|7670,7676|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|GLYCOL
Drug|Organic Chemical|Hospital Course|7670,7676|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|GLYCOL
Drug|Organic Chemical|Hospital Course|7683,7690|false|false|false|C0876088|Miralax|MIRALAX
Drug|Pharmacologic Substance|Hospital Course|7683,7690|false|false|false|C0876088|Miralax|MIRALAX
Event|Event|Hospital Course|7683,7690|false|false|false|||MIRALAX
Drug|Organic Chemical|Hospital Course|7694,7701|false|false|false|C0876088|Miralax|Miralax
Drug|Pharmacologic Substance|Hospital Course|7694,7701|false|false|false|C0876088|Miralax|Miralax
Anatomy|Body Space or Junction|Hospital Course|7715,7719|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|7715,7719|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|7715,7719|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|7715,7719|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Drug|Biomedical or Dental Material|Hospital Course|7730,7736|false|false|false|C0032861;C1382110|Powder dose form;powder physical state|powder
Drug|Substance|Hospital Course|7730,7736|false|false|false|C0032861;C1382110|Powder dose form;powder physical state|powder
Finding|Functional Concept|Hospital Course|7740,7748|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|7743,7748|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|7743,7748|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Intellectual Product|Hospital Course|7749,7753|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|Hospital Course|7749,7759|false|false|false|C3537736|Once A Day|once a day
Event|Event|Hospital Course|7756,7759|false|false|false|||day
Finding|Idea or Concept|Hospital Course|7756,7759|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|7756,7759|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Hospital Course|7763,7769|false|false|false|||needed
Event|Event|Hospital Course|7774,7786|false|false|false|||constipation
Finding|Sign or Symptom|Hospital Course|7774,7786|false|false|false|C0009806|Constipation|constipation
Event|Event|Hospital Course|7791,7801|false|false|false|||Prescribed
Finding|Functional Concept|Hospital Course|7811,7819|false|true|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|Provider
Finding|Intellectual Product|Hospital Course|7811,7819|false|true|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|Provider
Procedure|Health Care Activity|Hospital Course|7821,7836|true|false|false|C2826232|Dose Adjustment|Dose adjustment
Event|Event|Hospital Course|7826,7836|true|false|false|||adjustment
Finding|Classification|Hospital Course|7826,7836|true|false|false|C0376209;C0456081;C0678219;C0683269;C1546424|Adjustment - classification term;Personal Adjustment;Psychological adjustment;Transaction Type - Adjustment|adjustment
Finding|Functional Concept|Hospital Course|7826,7836|true|false|false|C0376209;C0456081;C0678219;C0683269;C1546424|Adjustment - classification term;Personal Adjustment;Psychological adjustment;Transaction Type - Adjustment|adjustment
Finding|Idea or Concept|Hospital Course|7826,7836|true|false|false|C0376209;C0456081;C0678219;C0683269;C1546424|Adjustment - classification term;Personal Adjustment;Psychological adjustment;Transaction Type - Adjustment|adjustment
Finding|Individual Behavior|Hospital Course|7826,7836|true|false|false|C0376209;C0456081;C0678219;C0683269;C1546424|Adjustment - classification term;Personal Adjustment;Psychological adjustment;Transaction Type - Adjustment|adjustment
Finding|Finding|Hospital Course|7842,7845|true|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Hospital Course|7842,7845|true|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Drug|Organic Chemical|Hospital Course|7850,7860|false|false|false|C3489575|sennosides, USP|SENNOSIDES
Drug|Pharmacologic Substance|Hospital Course|7850,7860|false|false|false|C3489575|sennosides, USP|SENNOSIDES
Event|Event|Hospital Course|7850,7860|false|false|false|||SENNOSIDES
Drug|Organic Chemical|Hospital Course|7862,7867|false|false|false|C3489575|sennosides, USP|SENNA
Drug|Pharmacologic Substance|Hospital Course|7862,7867|false|false|false|C3489575|sennosides, USP|SENNA
Event|Event|Hospital Course|7862,7867|false|false|false|||SENNA
Drug|Organic Chemical|Hospital Course|7871,7876|false|false|false|C3489575|sennosides, USP|senna
Drug|Pharmacologic Substance|Hospital Course|7871,7876|false|false|false|C3489575|sennosides, USP|senna
Drug|Biomedical or Dental Material|Hospital Course|7894,7900|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|Hospital Course|7904,7912|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|7907,7912|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|7907,7912|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Intellectual Product|Hospital Course|7913,7917|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|Hospital Course|7913,7923|false|false|false|C3537736|Once A Day|once a day
Event|Event|Hospital Course|7920,7923|false|false|false|||day
Finding|Idea or Concept|Hospital Course|7920,7923|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|7920,7923|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Hospital Course|7927,7933|false|false|false|||needed
Event|Event|Hospital Course|7938,7950|false|false|false|||constipation
Finding|Sign or Symptom|Hospital Course|7938,7950|false|false|false|C0009806|Constipation|constipation
Drug|Pharmacologic Substance|Hospital Course|7955,7958|false|false|false|C0013231|Drugs, Non-Prescription|OTC
Event|Event|Hospital Course|7955,7958|false|false|false|||OTC
Finding|Gene or Genome|Hospital Course|7955,7958|false|false|false|C1418193|OTC gene|OTC
Event|Event|Hospital Course|7963,7972|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|7963,7972|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|7963,7972|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|7963,7972|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|7963,7972|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|7963,7984|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|7973,7984|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|7973,7984|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|7973,7984|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|7973,7984|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Hospital Course|7990,7998|false|false|false|C0040610|tramadol|TraMADol
Drug|Pharmacologic Substance|Hospital Course|7990,7998|false|false|false|C0040610|tramadol|TraMADol
Event|Event|Hospital Course|7990,7998|false|false|false|||TraMADol
Procedure|Laboratory Procedure|Hospital Course|7990,7998|false|false|false|C1266765|Tramadol measurement (procedure)|TraMADol
Finding|Gene or Genome|Hospital Course|8012,8015|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|8016,8020|false|false|false|C2598155||Pain
Event|Event|Hospital Course|8016,8020|false|false|false|||Pain
Finding|Functional Concept|Hospital Course|8016,8020|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|Hospital Course|8016,8020|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Finding|Hospital Course|8023,8031|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Intellectual Product|Hospital Course|8023,8031|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Event|Event|Hospital Course|8035,8041|false|false|false|||Reason
Finding|Idea or Concept|Hospital Course|8035,8041|false|false|false|C0392360|Indication of (contextual qualifier)|Reason
Finding|Idea or Concept|Hospital Course|8035,8045|false|false|false|C0392360|Indication of (contextual qualifier)|Reason for
Finding|Gene or Genome|Hospital Course|8046,8049|false|false|false|C1422467|CIAO3 gene|PRN
Event|Activity|Hospital Course|8050,8059|false|false|false|C1883725|Replicate|duplicate
Finding|Functional Concept|Hospital Course|8050,8059|false|false|false|C0205173;C3539942|Double (qualifier value);Duplicate component (foundation metadata concept)|duplicate
Finding|Intellectual Product|Hospital Course|8050,8059|false|false|false|C0205173;C3539942|Double (qualifier value);Duplicate component (foundation metadata concept)|duplicate
Event|Event|Hospital Course|8060,8068|false|false|false|||override
Finding|Functional Concept|Hospital Course|8060,8068|false|false|false|C1547671|Override|override
Event|Event|Hospital Course|8082,8088|false|false|false|||agents
Drug|Organic Chemical|Hospital Course|8115,8123|false|false|false|C0040610|tramadol|tramadol
Drug|Pharmacologic Substance|Hospital Course|8115,8123|false|false|false|C0040610|tramadol|tramadol
Event|Event|Hospital Course|8115,8123|false|false|false|||tramadol
Procedure|Laboratory Procedure|Hospital Course|8115,8123|false|false|false|C1266765|Tramadol measurement (procedure)|tramadol
Drug|Biomedical or Dental Material|Hospital Course|8132,8138|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|Hospital Course|8142,8150|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|8145,8150|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|8145,8150|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Gene or Genome|Hospital Course|8156,8159|false|false|false|C1422467|CIAO3 gene|prn
Drug|Biomedical or Dental Material|Hospital Course|8169,8175|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|8169,8175|false|false|false|||Tablet
Event|Event|Hospital Course|8177,8184|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|8177,8184|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|8193,8205|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|Hospital Course|8193,8205|false|false|false|C0286651|atorvastatin|Atorvastatin
Event|Event|Hospital Course|8215,8218|false|false|false|||QPM
Drug|Organic Chemical|Hospital Course|8225,8233|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|Hospital Course|8225,8233|false|false|false|C1692318|docusate|Docusate
Event|Event|Hospital Course|8225,8233|false|false|false|||Docusate
Drug|Organic Chemical|Hospital Course|8225,8240|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|Hospital Course|8225,8240|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|Hospital Course|8234,8240|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|8234,8240|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|8234,8240|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|Hospital Course|8234,8240|false|false|false|||Sodium
Finding|Physiologic Function|Hospital Course|8234,8240|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|8234,8240|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8251,8254|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8251,8254|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|8251,8254|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|8251,8254|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|8251,8254|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|8261,8271|false|false|false|C0028978|omeprazole|Omeprazole
Drug|Pharmacologic Substance|Hospital Course|8261,8271|false|false|false|C0028978|omeprazole|Omeprazole
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8281,8284|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8281,8284|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|8281,8284|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|8281,8284|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|8281,8284|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|8291,8296|false|false|false|C3489575|sennosides, USP|Senna
Drug|Pharmacologic Substance|Hospital Course|8291,8296|false|false|false|C3489575|sennosides, USP|Senna
Drug|Organic Chemical|Hospital Course|8317,8327|false|false|false|C0074393|sertraline|Sertraline
Drug|Pharmacologic Substance|Hospital Course|8317,8327|false|false|false|C0074393|sertraline|Sertraline
Drug|Organic Chemical|Hospital Course|8350,8359|false|false|false|C0040805|trazodone|TraZODone
Drug|Pharmacologic Substance|Hospital Course|8350,8359|false|false|false|C0040805|trazodone|TraZODone
Finding|Gene or Genome|Hospital Course|8373,8376|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Organic Chemical|Hospital Course|8377,8382|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Drug|Pharmacologic Substance|Hospital Course|8377,8382|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Event|Event|Hospital Course|8377,8382|false|false|false|||sleep
Finding|Organism Function|Hospital Course|8377,8382|false|false|false|C0037313|Sleep|sleep
Event|Event|Hospital Course|8388,8397|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|8388,8397|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|8388,8397|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|8388,8397|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|8388,8397|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|8388,8409|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|8388,8409|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|8398,8409|false|false|false|C2926604||Disposition
Event|Event|Hospital Course|8398,8409|false|false|false|||Disposition
Procedure|Health Care Activity|Hospital Course|8398,8409|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|Hospital Course|8411,8415|false|false|false|||Home
Finding|Idea or Concept|Hospital Course|8411,8415|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|8411,8415|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|8411,8415|false|false|false|C1553498|home health encounter|Home
Event|Occupational Activity|Hospital Course|8421,8428|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|Hospital Course|8421,8428|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Event|Event|Hospital Course|8431,8439|false|false|false|||Facility
Finding|Intellectual Product|Hospital Course|8431,8439|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|Hospital Course|8447,8456|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|8447,8456|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|8447,8456|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|8447,8456|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|8447,8456|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|8447,8466|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|8457,8466|false|false|false|C0945731||Diagnosis
Event|Event|Hospital Course|8457,8466|false|false|false|||Diagnosis
Finding|Classification|Hospital Course|8457,8466|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|8457,8466|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|8457,8466|false|false|false|C0011900|Diagnosis|Diagnosis
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8468,8474|false|false|false|C0006141|Breast|breast
Disorder|Neoplastic Process|Hospital Course|8468,8474|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|breast
Event|Event|Hospital Course|8468,8474|false|false|false|||breast
Finding|Finding|Hospital Course|8468,8474|false|false|false|C0567499|Breast problem|breast
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8468,8474|false|false|false|C0191838|Procedures on breast|breast
Finding|Pathologic Function|Hospital Course|8468,8483|false|false|false|C0342095|Breast hematoma|breast hematoma
Event|Event|Hospital Course|8475,8483|false|false|false|||hematoma
Finding|Pathologic Function|Hospital Course|8475,8483|false|false|false|C0018944|Hematoma|hematoma
Finding|Mental Process|Discharge Condition|8509,8515|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|8509,8522|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|8509,8522|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|8516,8522|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|8516,8522|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|8524,8529|false|false|false|||Clear
Finding|Idea or Concept|Discharge Condition|8524,8529|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|Discharge Condition|8534,8542|false|false|false|||coherent
Finding|Finding|Discharge Condition|8534,8542|false|false|false|C4068804|Coherent|coherent
Event|Event|Discharge Condition|8544,8549|false|false|false|||Level
Attribute|Clinical Attribute|Discharge Condition|8544,8566|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|8544,8566|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|Discharge Condition|8553,8566|false|false|false|||Consciousness
Finding|Finding|Discharge Condition|8553,8566|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|8553,8566|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|8568,8573|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|8568,8573|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|8568,8573|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|Discharge Condition|8568,8573|false|false|false|||Alert
Finding|Finding|Discharge Condition|8568,8573|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|8568,8573|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|8568,8573|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|Discharge Condition|8578,8589|false|false|false|||interactive
Finding|Functional Concept|Discharge Condition|8578,8589|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|8591,8599|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|8591,8599|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|8591,8599|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|8600,8606|false|false|false|C5889824||Status
Event|Event|Discharge Condition|8600,8606|false|false|false|||Status
Finding|Idea or Concept|Discharge Condition|8600,8606|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|8608,8618|false|false|false|||Ambulatory
Finding|Functional Concept|Discharge Condition|8608,8618|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|Discharge Condition|8608,8618|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|Discharge Condition|8608,8618|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|Discharge Condition|8608,8618|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|Discharge Condition|8621,8632|false|false|false|||Independent
Finding|Finding|Discharge Condition|8621,8632|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|Discharge Condition|8621,8632|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Daily or Recreational Activity|Discharge Instructions|8661,8674|false|false|false|C0036592|Self-care interventions|Personal Care
Event|Activity|Discharge Instructions|8670,8674|false|false|false|C1947933|care activity|Care
Finding|Finding|Discharge Instructions|8670,8674|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|Discharge Instructions|8670,8674|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Event|Event|Discharge Instructions|8689,8693|false|false|false|||keep
Event|Event|Discharge Instructions|8699,8708|false|false|false|||incisions
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|8699,8708|false|false|false|C0184898|Surgical incisions|incisions
Drug|Inorganic Chemical|Discharge Instructions|8717,8720|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|Discharge Instructions|8717,8720|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|Discharge Instructions|8717,8720|false|false|false|C0001861;C3536832|Air (substance);air|air
Event|Event|Discharge Instructions|8717,8720|false|false|false|||air
Finding|Finding|Discharge Instructions|8717,8720|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|Discharge Instructions|8717,8720|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|Discharge Instructions|8717,8720|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Event|Event|Discharge Instructions|8724,8731|false|false|false|||covered
Event|Activity|Discharge Instructions|8740,8745|false|false|false|C1947930|Cleaning (activity)|clean
Finding|Finding|Discharge Instructions|8747,8754|false|false|false|C0021359;C4074771|Infertility;Sterility, Reproductive|sterile
Finding|Pathologic Function|Discharge Instructions|8747,8754|false|false|false|C0021359;C4074771|Infertility;Sterility, Reproductive|sterile
Event|Event|Discharge Instructions|8770,8776|false|false|false|||change
Event|Activity|Discharge Instructions|8787,8792|false|false|false|C1947930|Cleaning (activity)|Clean
Drug|Substance|Discharge Instructions|8804,8809|false|false|false|C1550628|Drain - SpecimenType|drain
Event|Event|Discharge Instructions|8804,8809|false|false|false|||drain
Finding|Intellectual Product|Discharge Instructions|8804,8809|false|false|false|C1546604|Drain Specimen Code|drain
Anatomy|Body Location or Region|Discharge Instructions|8810,8814|false|false|false|C1515974|Anatomic Site|site
Finding|Intellectual Product|Discharge Instructions|8810,8814|false|false|false|C1546778||site
Event|Event|Discharge Instructions|8836,8841|false|false|false|||exits
Anatomy|Body System|Discharge Instructions|8847,8851|false|false|false|C1123023;C4520765|Skin;Skin, Human|skin
Disorder|Disease or Syndrome|Discharge Instructions|8847,8851|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Disorder|Neoplastic Process|Discharge Instructions|8847,8851|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Event|Event|Discharge Instructions|8847,8851|false|false|false|||skin
Finding|Body Substance|Discharge Instructions|8847,8851|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Finding|Intellectual Product|Discharge Instructions|8847,8851|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Drug|Biomedical or Dental Material|Discharge Instructions|8858,8862|false|false|false|C1705308|Soap Dosage Form|soap
Event|Event|Discharge Instructions|8858,8862|false|false|false|||soap
Drug|Inorganic Chemical|Discharge Instructions|8867,8872|false|false|false|C0043047;C1550678|Water Specimen;water|water
Drug|Pharmacologic Substance|Discharge Instructions|8867,8872|false|false|false|C0043047;C1550678|Water Specimen;water|water
Event|Event|Discharge Instructions|8867,8872|false|false|false|||water
Finding|Intellectual Product|Discharge Instructions|8867,8872|false|false|false|C1547961|Water - Specimen Source Codes|water
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|8867,8872|false|false|false|C0020311|Hydrotherapy|water
Drug|Biomedical or Dental Material|Discharge Instructions|8879,8884|false|false|false|C1555557;C3241918|Compliance Package - Strip;Strip Dosage Form|Strip
Drug|Substance|Discharge Instructions|8885,8890|false|false|false|C1550628|Drain - SpecimenType|drain
Event|Event|Discharge Instructions|8885,8890|false|false|false|||drain
Finding|Intellectual Product|Discharge Instructions|8885,8890|false|false|false|C1546604|Drain Specimen Code|drain
Event|Event|Discharge Instructions|8891,8897|false|false|false|||tubing
Finding|Functional Concept|Discharge Instructions|8899,8904|false|false|false|C5848602|Exhausted|empty
Anatomy|Anatomical Structure|Discharge Instructions|8905,8909|false|false|false|C0025148;C1947952|Medulla Oblongata;anatomical bulb|bulb
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|8905,8909|false|false|false|C0025148;C1947952|Medulla Oblongata;anatomical bulb|bulb
Finding|Intellectual Product|Discharge Instructions|8918,8924|false|false|false|C0034869|Records|record
Event|Event|Discharge Instructions|8925,8931|false|false|false|||output
Finding|Conceptual Entity|Discharge Instructions|8925,8931|false|false|false|C1709366|system output|output
Procedure|Health Care Activity|Discharge Instructions|8925,8931|false|false|false|C3251815|Measurement of fluid output|output
Disorder|Disease or Syndrome|Discharge Instructions|8940,8945|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Event|Event|Discharge Instructions|8940,8945|false|false|false|||times
Finding|Idea or Concept|Discharge Instructions|8950,8953|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Discharge Instructions|8950,8953|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Functional Concept|Discharge Instructions|8962,8969|false|false|false|C1547186;C1576874|Written - Consent Mode;written - ParticipationMode|written
Finding|Idea or Concept|Discharge Instructions|8962,8969|false|false|false|C1547186;C1576874|Written - Consent Mode;written - ParticipationMode|written
Event|Event|Discharge Instructions|8970,8976|false|false|false|||record
Finding|Intellectual Product|Discharge Instructions|8970,8976|false|false|false|C0034869|Records|record
Event|Event|Discharge Instructions|8990,8996|false|false|false|||output
Finding|Conceptual Entity|Discharge Instructions|8990,8996|false|false|false|C1709366|system output|output
Procedure|Health Care Activity|Discharge Instructions|8990,8996|false|false|false|C3251815|Measurement of fluid output|output
Drug|Substance|Discharge Instructions|9007,9012|false|false|false|C1550628|Drain - SpecimenType|drain
Finding|Intellectual Product|Discharge Instructions|9007,9012|false|false|false|C1546604|Drain Specimen Code|drain
Event|Event|Discharge Instructions|9013,9019|false|false|false|||should
Event|Event|Discharge Instructions|9024,9031|false|false|false|||brought
Event|Event|Discharge Instructions|9041,9047|false|false|false|||follow
Finding|Functional Concept|Discharge Instructions|9041,9047|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|Discharge Instructions|9041,9047|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|Discharge Instructions|9041,9050|false|false|false|C0589120|Follow-up status|follow-up
Procedure|Health Care Activity|Discharge Instructions|9041,9050|false|false|false|C1522577|follow-up|follow-up
Event|Activity|Discharge Instructions|9051,9062|false|false|false|C0003629|Appointments|appointment
Event|Event|Discharge Instructions|9051,9062|false|false|false|||appointment
Event|Event|Discharge Instructions|9069,9075|false|false|false|||drains
Event|Event|Discharge Instructions|9085,9092|false|false|false|||removed
Finding|Finding|Discharge Instructions|9104,9112|false|false|false|C0332149|Possible|possible
Event|Event|Discharge Instructions|9128,9134|false|false|false|||output
Finding|Conceptual Entity|Discharge Instructions|9128,9134|false|false|false|C1709366|system output|output
Procedure|Health Care Activity|Discharge Instructions|9128,9134|false|false|false|C3251815|Measurement of fluid output|output
Event|Event|Discharge Instructions|9135,9141|false|false|false|||tapers
Event|Event|Discharge Instructions|9164,9170|false|false|false|||amount
Finding|Intellectual Product|Discharge Instructions|9164,9170|false|false|false|C1561574|Amount class - Amount|amount
Event|Event|Discharge Instructions|9185,9189|false|false|false|||wear
Procedure|Health Care Activity|Discharge Instructions|9192,9200|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|9192,9200|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|9201,9204|false|false|false|C0006104|Brain|bra
Disorder|Disease or Syndrome|Discharge Instructions|9208,9212|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|Discharge Instructions|9208,9212|false|false|false|||soft
Drug|Organic Chemical|Discharge Instructions|9234,9241|false|false|false|C1310585|Comfort brand of hydroxyethyl cellulose|comfort
Drug|Pharmacologic Substance|Discharge Instructions|9234,9241|false|false|false|C1310585|Comfort brand of hydroxyethyl cellulose|comfort
Event|Event|Discharge Instructions|9234,9241|false|false|false|||comfort
Finding|Mental Process|Discharge Instructions|9234,9241|false|false|false|C1331418|Comfort|comfort
Event|Event|Discharge Instructions|9255,9261|true|false|false|||shower
Drug|Substance|Discharge Instructions|9273,9278|false|false|false|C1550628|Drain - SpecimenType|drain
Event|Event|Discharge Instructions|9273,9278|false|false|false|||drain
Finding|Intellectual Product|Discharge Instructions|9273,9278|false|false|false|C1546604|Drain Specimen Code|drain
Event|Activity|Discharge Instructions|9285,9290|false|false|false|C1882509|put - instruction imperative|place
Event|Event|Discharge Instructions|9285,9290|false|false|false|||place
Finding|Functional Concept|Discharge Instructions|9285,9290|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|Discharge Instructions|9285,9290|false|false|false|C1533810||place
Drug|Biomedical or Dental Material|Discharge Instructions|9300,9309|false|false|false|C1530215|DERMABOND|Dermabond
Drug|Organic Chemical|Discharge Instructions|9300,9309|false|false|false|C1530215|DERMABOND|Dermabond
Anatomy|Body System|Discharge Instructions|9310,9314|false|false|false|C1123023;C4520765|Skin;Skin, Human|skin
Disorder|Disease or Syndrome|Discharge Instructions|9310,9314|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Disorder|Neoplastic Process|Discharge Instructions|9310,9314|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Finding|Body Substance|Discharge Instructions|9310,9314|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Finding|Intellectual Product|Discharge Instructions|9310,9314|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Drug|Substance|Discharge Instructions|9315,9319|false|false|false|C0017780|Glues|glue
Event|Event|Discharge Instructions|9315,9319|false|false|false|||glue
Event|Event|Discharge Instructions|9325,9330|false|false|false|||begin
Event|Event|Discharge Instructions|9334,9339|false|false|false|||flake
Event|Activity|Discharge Instructions|9367,9375|false|false|false|C0441655|Activities|Activity
Event|Event|Discharge Instructions|9367,9375|false|false|false|||Activity
Finding|Daily or Recreational Activity|Discharge Instructions|9367,9375|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Instructions|9367,9375|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Event|Event|Discharge Instructions|9390,9396|false|false|false|||resume
Finding|Daily or Recreational Activity|Discharge Instructions|9402,9414|false|false|false|C0184625||regular diet
Drug|Food|Discharge Instructions|9410,9414|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|Discharge Instructions|9410,9414|false|false|false|||diet
Finding|Functional Concept|Discharge Instructions|9410,9414|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|Discharge Instructions|9410,9414|false|false|false|C0012159|Diet therapy|diet
Finding|Daily or Recreational Activity|Discharge Instructions|9421,9425|false|false|false|C0080331|Walking (function)|Walk
Disorder|Disease or Syndrome|Discharge Instructions|9434,9439|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|Discharge Instructions|9442,9445|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Discharge Instructions|9442,9445|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Discharge Instructions|9459,9463|true|false|false|||lift
Finding|Daily or Recreational Activity|Discharge Instructions|9509,9527|false|false|false|C1514989|Strenuous Exercise|strenuous activity
Event|Activity|Discharge Instructions|9519,9527|false|false|false|C0441655|Activities|activity
Event|Event|Discharge Instructions|9519,9527|false|false|false|||activity
Finding|Daily or Recreational Activity|Discharge Instructions|9519,9527|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|activity
Finding|Finding|Discharge Instructions|9519,9527|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|activity
Event|Event|Discharge Instructions|9550,9557|false|false|false|||surgery
Finding|Finding|Discharge Instructions|9550,9557|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|Discharge Instructions|9550,9557|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|Discharge Instructions|9550,9557|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|9550,9557|false|false|false|C0543467|Operative Surgical Procedures|surgery
Event|Event|Medications|9579,9585|false|false|false|||Resume
Finding|Functional Concept|Medications|9579,9585|false|false|false|C1550028;C1880201;C3242342|Curriculum Vitae;Resume - Remote control command;resume - DataOperation|Resume
Finding|Idea or Concept|Medications|9579,9585|false|false|false|C1550028;C1880201;C3242342|Curriculum Vitae;Resume - Remote control command;resume - DataOperation|Resume
Finding|Intellectual Product|Medications|9579,9585|false|false|false|C1550028;C1880201;C3242342|Curriculum Vitae;Resume - Remote control command;resume - DataOperation|Resume
Attribute|Clinical Attribute|Medications|9599,9610|true|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Medications|9599,9610|true|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Medications|9599,9610|true|false|false|||medications
Finding|Intellectual Product|Medications|9599,9610|true|false|false|C4284232|Medications|medications
Event|Event|Medications|9618,9628|true|false|false|||instructed
Event|Event|Medications|9644,9648|true|false|false|||take
Finding|Finding|Medications|9653,9656|true|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Medications|9653,9656|true|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Disorder|Disease or Syndrome|Medications|9657,9661|true|false|false|C3280240|MICROCEPHALY, EPILEPSY, AND DIABETES SYNDROME 1|meds
Event|Event|Medications|9657,9661|true|false|false|||meds
Finding|Intellectual Product|Medications|9657,9661|true|false|false|C4284232|Medications|meds
Event|Event|Medications|9665,9672|true|false|false|||ordered
Event|Event|Medications|9688,9692|false|false|false|||take
Event|Event|Medications|9698,9708|false|false|false|||prescribed
Attribute|Clinical Attribute|Medications|9709,9713|false|false|false|C2598155||pain
Finding|Functional Concept|Medications|9709,9713|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Medications|9709,9713|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Pharmacologic Substance|Medications|9714,9724|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Medications|9714,9724|false|false|false|||medication
Finding|Intellectual Product|Medications|9714,9724|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|Medications|9729,9737|false|false|false|||moderate
Finding|Finding|Medications|9729,9737|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|Medications|9729,9737|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Finding|Medications|9742,9748|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|Medications|9742,9748|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Finding|Medications|9742,9753|false|false|false|C0278140;C4050465;C4521229|Neck Pain Score 6;Severe Extremity Pain;Severe pain|severe pain
Attribute|Clinical Attribute|Medications|9749,9753|false|false|false|C2598155||pain
Event|Event|Medications|9749,9753|false|false|false|||pain
Finding|Functional Concept|Medications|9749,9753|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Medications|9749,9753|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Medications|9763,9769|false|false|false|||switch
Drug|Organic Chemical|Medications|9773,9780|false|false|false|C0699142|Tylenol|Tylenol
Drug|Pharmacologic Substance|Medications|9773,9780|false|false|false|C0699142|Tylenol|Tylenol
Event|Event|Medications|9773,9780|false|false|false|||Tylenol
Drug|Organic Chemical|Medications|9784,9806|false|false|false|C0724019|Tylenol Extra Strength|Extra Strength Tylenol
Drug|Pharmacologic Substance|Medications|9784,9806|false|false|false|C0724019|Tylenol Extra Strength|Extra Strength Tylenol
Finding|Idea or Concept|Medications|9790,9798|false|false|false|C0808080|Strength (attribute)|Strength
Drug|Organic Chemical|Medications|9799,9806|false|false|false|C0699142|Tylenol|Tylenol
Drug|Pharmacologic Substance|Medications|9799,9806|false|false|false|C0699142|Tylenol|Tylenol
Event|Event|Medications|9799,9806|false|false|false|||Tylenol
Finding|Intellectual Product|Medications|9812,9816|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Finding|Medications|9812,9821|false|false|false|C0278138;C4522280|Mild pain;Neck Pain Score 2|mild pain
Attribute|Clinical Attribute|Medications|9817,9821|false|false|false|C2598155||pain
Event|Event|Medications|9817,9821|false|false|false|||pain
Finding|Functional Concept|Medications|9817,9821|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Medications|9817,9821|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Medications|9825,9833|false|false|false|||directed
Event|Activity|Medications|9841,9850|false|false|false|C2828395|Packing (action)|packaging
Phenomenon|Human-caused Phenomenon or Process|Medications|9841,9850|false|false|false|C0030176|Packaging|packaging
Event|Event|Medications|9859,9863|false|false|false|||note
Drug|Organic Chemical|Medications|9870,9878|false|false|false|C0086787|Percocet|Percocet
Drug|Pharmacologic Substance|Medications|9870,9878|false|false|false|C0086787|Percocet|Percocet
Drug|Organic Chemical|Medications|9883,9890|false|false|false|C0483514|Vicodin|Vicodin
Drug|Pharmacologic Substance|Medications|9883,9890|false|false|false|C0483514|Vicodin|Vicodin
Drug|Organic Chemical|Medications|9896,9903|false|false|false|C0699142|Tylenol|Tylenol
Drug|Pharmacologic Substance|Medications|9896,9903|false|false|false|C0699142|Tylenol|Tylenol
Event|Event|Medications|9896,9903|false|false|false|||Tylenol
Drug|Chemical Viewed Functionally|Medications|9910,9927|true|false|false|C1372955|Active ingredient|active ingredient
Drug|Chemical Viewed Functionally|Medications|9917,9927|true|false|false|C1550600|Ingredient|ingredient
Event|Event|Medications|9917,9927|true|false|false|||ingredient
Event|Event|Medications|9939,9943|true|false|false|||take
Disorder|Disease or Syndrome|Medications|9950,9954|true|false|false|C3280240|MICROCEPHALY, EPILEPSY, AND DIABETES SYNDROME 1|meds
Event|Event|Medications|9950,9954|true|false|false|||meds
Finding|Intellectual Product|Medications|9950,9954|true|false|false|C4284232|Medications|meds
Finding|Functional Concept|Medications|9960,9970|true|false|false|C1524062|Additional|additional
Drug|Organic Chemical|Medications|9971,9978|true|false|false|C0699142|Tylenol|Tylenol
Drug|Pharmacologic Substance|Medications|9971,9978|true|false|false|C0699142|Tylenol|Tylenol
Event|Event|Medications|9985,9989|true|false|false|||Take
Attribute|Clinical Attribute|Medications|9990,10002|true|false|false|C5886759|Prescription (attribute)|prescription
Event|Event|Medications|9990,10002|true|false|false|||prescription
Finding|Intellectual Product|Medications|9990,10002|true|false|false|C1521941|prescription document|prescription
Procedure|Health Care Activity|Medications|9990,10002|true|false|false|C0033080|Prescription (procedure)|prescription
Attribute|Clinical Attribute|Medications|10003,10007|true|false|false|C2598155||pain
Finding|Functional Concept|Medications|10003,10007|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Medications|10003,10007|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|Medications|10008,10019|true|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Medications|10008,10019|true|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Medications|10008,10019|true|false|false|||medications
Finding|Intellectual Product|Medications|10008,10019|true|false|false|C4284232|Medications|medications
Attribute|Clinical Attribute|Medications|10024,10028|true|false|false|C2598155||pain
Event|Event|Medications|10024,10028|true|false|false|||pain
Finding|Functional Concept|Medications|10024,10028|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Medications|10024,10028|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Medications|10033,10041|true|false|false|||relieved
Drug|Organic Chemical|Medications|10046,10053|true|false|false|C0699142|Tylenol|Tylenol
Drug|Pharmacologic Substance|Medications|10046,10053|true|false|false|C0699142|Tylenol|Tylenol
Event|Event|Medications|10060,10064|false|false|false|||Take
Drug|Organic Chemical|Medications|10065,10071|false|false|false|C0282139|Colace|Colace
Drug|Pharmacologic Substance|Medications|10065,10071|false|false|false|C0282139|Colace|Colace
Event|Event|Medications|10065,10071|false|false|false|||Colace
Finding|Functional Concept|Medications|10080,10088|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Medications|10083,10088|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Medications|10083,10088|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Finding|Medications|10089,10096|false|false|false|C4035627|2 times|2 times
Finding|Finding|Medications|10089,10104|false|false|false|C3844164|2 times per day|2 times per day
Disorder|Disease or Syndrome|Medications|10091,10096|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Event|Event|Medications|10091,10096|false|false|false|||times
Finding|Idea or Concept|Medications|10101,10104|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Medications|10101,10104|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Medications|10112,10118|false|false|false|||taking
Attribute|Clinical Attribute|Medications|10124,10136|false|false|false|C5886759|Prescription (attribute)|prescription
Event|Event|Medications|10124,10136|false|false|false|||prescription
Finding|Intellectual Product|Medications|10124,10136|false|false|false|C1521941|prescription document|prescription
Procedure|Health Care Activity|Medications|10124,10136|false|false|false|C0033080|Prescription (procedure)|prescription
Attribute|Clinical Attribute|Medications|10137,10141|false|false|false|C2598155||pain
Finding|Functional Concept|Medications|10137,10141|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Medications|10137,10141|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Pharmacologic Substance|Medications|10142,10152|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Medications|10142,10152|false|false|false|||medication
Finding|Intellectual Product|Medications|10142,10152|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|Medications|10162,10165|false|false|false|||use
Event|Event|Medications|10168,10177|false|false|false|||different
Drug|Hazardous or Poisonous Substance|Medications|10188,10195|false|false|false|C0702263|Counter brand of Terbufos|counter
Drug|Organic Chemical|Medications|10188,10195|false|false|false|C0702263|Counter brand of Terbufos|counter
Finding|Body Substance|Medications|10196,10201|false|false|false|C0015733|Feces|stool
Drug|Organic Chemical|Medications|10196,10210|false|false|false|C0301470;C1154263|Stool Softener;Stool Softener brand of docusate sodium|stool softener
Drug|Pharmacologic Substance|Medications|10196,10210|false|false|false|C0301470;C1154263|Stool Softener;Stool Softener brand of docusate sodium|stool softener
Event|Event|Medications|10202,10210|false|false|false|||softener
Event|Event|Medications|10218,10222|false|false|false|||wish
Event|Event|Medications|10236,10241|true|false|false|||drive
Event|Event|Medications|10245,10252|true|false|false|||operate
Disorder|Injury or Poisoning|Medications|10259,10268|true|false|false|C0337246|Contact with machinery|machinery
Event|Event|Medications|10259,10268|true|false|false|||machinery
Drug|Hazardous or Poisonous Substance|Medications|10287,10295|true|false|false|C0027415|Narcotics|narcotic
Drug|Pharmacologic Substance|Medications|10287,10295|true|false|false|C0027415|Narcotics|narcotic
Event|Event|Medications|10287,10295|true|false|false|||narcotic
Attribute|Clinical Attribute|Medications|10296,10300|true|false|false|C2598155||pain
Event|Event|Medications|10296,10300|true|false|false|||pain
Finding|Functional Concept|Medications|10296,10300|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Medications|10296,10300|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Pharmacologic Substance|Medications|10301,10311|true|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Medications|10301,10311|true|false|false|||medication
Finding|Intellectual Product|Medications|10301,10311|true|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Finding|Intellectual Product|Medications|10321,10338|false|false|false|C3641755|Have Constipation|have constipation
Event|Event|Medications|10326,10338|false|false|false|||constipation
Finding|Sign or Symptom|Medications|10326,10338|false|false|false|C0009806|Constipation|constipation
Drug|Hazardous or Poisonous Substance|Medications|10352,10360|false|false|false|C0027415|Narcotics|narcotic
Drug|Pharmacologic Substance|Medications|10352,10360|false|false|false|C0027415|Narcotics|narcotic
Attribute|Clinical Attribute|Medications|10361,10365|false|false|false|C2598155||pain
Event|Event|Medications|10361,10365|false|false|false|||pain
Finding|Functional Concept|Medications|10361,10365|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Medications|10361,10365|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|Medications|10366,10377|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Medications|10366,10377|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Medications|10366,10377|false|false|false|||medications
Finding|Intellectual Product|Medications|10366,10377|false|false|false|C4284232|Medications|medications
Drug|Organic Chemical|Medications|10379,10388|false|false|false|C0030049|oxycodone|oxycodone
Drug|Pharmacologic Substance|Medications|10379,10388|false|false|false|C0030049|oxycodone|oxycodone
Event|Event|Medications|10379,10388|false|false|false|||oxycodone
Procedure|Laboratory Procedure|Medications|10379,10388|false|false|false|C0524222|Oxycodone measurement|oxycodone
Drug|Organic Chemical|Medications|10390,10398|false|false|false|C0086787|Percocet|percocet
Drug|Pharmacologic Substance|Medications|10390,10398|false|false|false|C0086787|Percocet|percocet
Event|Event|Medications|10390,10398|false|false|false|||percocet
Drug|Organic Chemical|Medications|10400,10407|false|false|false|C0483514|Vicodin|vicodin
Drug|Pharmacologic Substance|Medications|10400,10407|false|false|false|C0483514|Vicodin|vicodin
Event|Event|Medications|10400,10407|false|false|false|||vicodin
Drug|Organic Chemical|Medications|10410,10421|false|false|false|C0020264|hydrocodone|hydrocodone
Drug|Pharmacologic Substance|Medications|10410,10421|false|false|false|C0020264|hydrocodone|hydrocodone
Event|Event|Medications|10410,10421|false|false|false|||hydrocodone
Drug|Organic Chemical|Medications|10423,10431|false|false|false|C0728755|Dilaudid|dilaudid
Drug|Pharmacologic Substance|Medications|10423,10431|false|false|false|C0728755|Dilaudid|dilaudid
Event|Event|Medications|10423,10431|false|false|false|||dilaudid
Event|Event|Medications|10433,10436|false|false|false|||etc
Finding|Idea or Concept|Medications|10433,10436|false|false|false|C1548556|Etc.|etc
Event|Event|Medications|10451,10459|false|false|false|||continue
Event|Event|Medications|10460,10468|false|false|false|||drinking
Finding|Individual Behavior|Medications|10460,10468|false|false|false|C0001948;C0684271|Alcohol consumption;Drinking (function)|drinking
Finding|Organism Function|Medications|10460,10468|false|false|false|C0001948;C0684271|Alcohol consumption;Drinking (function)|drinking
Drug|Substance|Medications|10470,10476|false|false|false|C0302908|Liquid substance|fluids
Event|Event|Medications|10470,10476|false|false|false|||fluids
Finding|Body Substance|Medications|10470,10476|false|false|false|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|Medications|10470,10476|false|false|false|C0016286|Fluid Therapy|fluids
Finding|Body Substance|Medications|10491,10496|false|false|false|C0015733|Feces|stool
Drug|Pharmacologic Substance|Medications|10491,10506|false|false|false|C0301470|Stool Softener|stool softeners
Event|Event|Medications|10497,10506|false|false|false|||softeners
Event|Event|Medications|10519,10522|false|false|false|||eat
Drug|Food|Medications|10523,10528|false|false|false|C0016452|Food|foods
Event|Event|Medications|10523,10528|false|false|false|||foods
Event|Event|Medications|10539,10543|false|false|false|||high
Finding|Finding|Medications|10539,10543|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|Medications|10539,10543|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|Medications|10539,10543|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Anatomy|Tissue|Medications|10547,10552|false|false|false|C1304649|Tissue fiber|fiber
Drug|Organic Chemical|Medications|10547,10552|false|false|false|C0225326;C1321801|Fiber brand of calcium polycarbophil;fiber|fiber
Drug|Pharmacologic Substance|Medications|10547,10552|false|false|false|C0225326;C1321801|Fiber brand of calcium polycarbophil;fiber|fiber
Event|Event|Medications|10557,10561|false|false|false|||Call
Event|Event|Medications|10566,10572|false|false|false|||office
Finding|Idea or Concept|Medications|10566,10572|false|false|false|C1549636|Address type - Office|office
Event|Event|Medications|10624,10629|false|false|false|||Signs
Finding|Finding|Medications|10624,10629|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|Signs
Finding|Functional Concept|Medications|10624,10629|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|Signs
Disorder|Disease or Syndrome|Medications|10633,10642|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|Medications|10633,10642|false|false|false|||infection
Finding|Pathologic Function|Medications|10633,10642|false|false|false|C3714514|Infection|infection
Event|Event|Medications|10644,10649|false|false|false|||fever
Finding|Finding|Medications|10644,10649|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|Medications|10644,10649|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|Medications|10644,10661|false|false|false|C0085594|Fever with chills|fever with chills
Event|Event|Medications|10655,10661|false|false|false|||chills
Finding|Sign or Symptom|Medications|10655,10661|false|false|false|C0085593|Chills|chills
Event|Event|Medications|10663,10672|false|false|false|||increased
Disorder|Disease or Syndrome|Medications|10673,10680|false|false|false|C0041834|Erythema|redness
Event|Event|Medications|10673,10680|false|false|false|||redness
Finding|Finding|Medications|10673,10680|false|false|false|C0332575|Redness|redness
Event|Event|Medications|10683,10691|false|false|false|||swelling
Finding|Finding|Medications|10683,10691|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|Medications|10683,10691|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Event|Event|Medications|10693,10699|false|false|false|||warmth
Finding|Finding|Medications|10693,10699|false|false|false|C0392197;C0518610|Physiologic warmth;Social warmth|warmth
Finding|Physiologic Function|Medications|10693,10699|false|false|false|C0392197;C0518610|Physiologic warmth;Social warmth|warmth
Event|Event|Medications|10703,10713|false|false|false|||tenderness
Finding|Mental Process|Medications|10703,10713|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|Medications|10703,10713|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Procedure|Health Care Activity|Medications|10721,10729|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Procedure|Therapeutic or Preventive Procedure|Medications|10721,10729|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Anatomy|Body Location or Region|Medications|10730,10734|false|false|false|C1515974|Anatomic Site|site
Finding|Intellectual Product|Medications|10730,10734|false|false|false|C1546778||site
Event|Event|Medications|10739,10746|false|false|false|||unusual
Event|Event|Medications|10748,10756|false|false|false|||drainage
Finding|Body Substance|Medications|10748,10756|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Finding|Sign or Symptom|Medications|10748,10756|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Procedure|Therapeutic or Preventive Procedure|Medications|10748,10756|false|false|false|C0013103|Drainage procedure|drainage
Anatomy|Body Location or Region|Medications|10766,10774|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|Medications|10766,10774|false|false|false|C0332803|Surgical wound|incision
Procedure|Therapeutic or Preventive Procedure|Medications|10766,10774|false|false|false|C0184898|Surgical incisions|incision
Finding|Gene or Genome|Medications|10786,10791|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Finding|Intellectual Product|Medications|10792,10798|false|false|false|C1561574|Amount class - Amount|amount
Event|Event|Medications|10802,10810|false|false|false|||bleeding
Finding|Pathologic Function|Medications|10802,10810|false|false|false|C0019080|Hemorrhage|bleeding
Anatomy|Body Location or Region|Medications|10820,10828|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|Medications|10820,10828|false|false|false|C0332803|Surgical wound|incision
Procedure|Therapeutic or Preventive Procedure|Medications|10820,10828|false|false|false|C0184898|Surgical incisions|incision
Drug|Substance|Medications|10835,10840|false|false|false|C1550628|Drain - SpecimenType|drain
Event|Event|Medications|10835,10840|false|false|false|||drain
Finding|Intellectual Product|Medications|10835,10840|false|false|false|C1546604|Drain Specimen Code|drain
Event|Event|Medications|10851,10856|false|false|false|||Fever
Finding|Finding|Medications|10851,10856|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|Fever
Finding|Sign or Symptom|Medications|10851,10856|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|Fever
Finding|Finding|Medications|10884,10890|true|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|Severe
Finding|Intellectual Product|Medications|10884,10890|true|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|Severe
Finding|Finding|Medications|10884,10895|true|false|false|C0278140;C4050465;C4521229|Neck Pain Score 6;Severe Extremity Pain;Severe pain|Severe pain
Attribute|Clinical Attribute|Medications|10891,10895|true|false|false|C2598155||pain
Event|Event|Medications|10891,10895|true|false|false|||pain
Finding|Functional Concept|Medications|10891,10895|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Medications|10891,10895|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Medications|10900,10908|true|false|false|||relieved
Drug|Pharmacologic Substance|Medications|10917,10927|true|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Medications|10917,10927|true|false|false|||medication
Finding|Intellectual Product|Medications|10917,10927|true|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|Medications|10934,10940|false|false|false|||Return
Event|Event|Medications|10970,10978|true|false|false|||vomiting
Finding|Sign or Symptom|Medications|10970,10978|true|false|false|C0042963|Vomiting|vomiting
Event|Event|Medications|10990,10994|true|false|false|||keep
Drug|Substance|Medications|10998,11004|true|false|true|C0302908|Liquid substance|fluids
Event|Event|Medications|10998,11004|true|false|false|||fluids
Finding|Body Substance|Medications|10998,11004|true|false|true|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|Medications|10998,11004|true|false|true|C0016286|Fluid Therapy|fluids
Attribute|Clinical Attribute|Medications|11014,11025|true|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Medications|11014,11025|true|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Medications|11014,11025|true|false|false|||medications
Finding|Intellectual Product|Medications|11014,11025|true|false|false|C4284232|Medications|medications
Event|Event|Medications|11051,11057|false|false|false|||chills
Finding|Sign or Symptom|Medications|11051,11057|false|false|false|C0085593|Chills|chills
Event|Event|Medications|11059,11064|false|false|false|||fever
Finding|Finding|Medications|11059,11064|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|Medications|11059,11064|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Event|Event|Medications|11089,11096|false|false|false|||degrees
Finding|Intellectual Product|Medications|11089,11096|false|false|false|C0542560|Academic degree|degrees
Event|Event|Medications|11107,11114|false|false|false|||degrees
Finding|Intellectual Product|Medications|11107,11114|false|false|false|C0542560|Academic degree|degrees
Finding|Finding|Medications|11116,11125|false|false|false|C0442805;C5236002|Increase;Increased (finding)|increased
Finding|Functional Concept|Medications|11116,11125|false|false|false|C0442805;C5236002|Increase;Increased (finding)|increased
Disorder|Disease or Syndrome|Medications|11126,11133|false|false|false|C0041834|Erythema|redness
Event|Event|Medications|11126,11133|false|false|false|||redness
Finding|Finding|Medications|11126,11133|false|false|false|C0332575|Redness|redness
Event|Event|Medications|11135,11143|false|false|false|||swelling
Finding|Finding|Medications|11135,11143|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|Medications|11135,11143|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Event|Event|Medications|11148,11157|false|false|false|||discharge
Finding|Body Substance|Medications|11148,11157|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Medications|11148,11157|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Medications|11148,11157|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Medications|11148,11157|false|false|false|C0030685|Patient Discharge|discharge
Anatomy|Body Location or Region|Medications|11163,11171|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|Medications|11163,11171|false|false|false|C0332803|Surgical wound|incision
Event|Event|Medications|11163,11171|false|false|false|||incision
Procedure|Therapeutic or Preventive Procedure|Medications|11163,11171|false|false|false|C0184898|Surgical incisions|incision
Anatomy|Body Location or Region|Medications|11173,11178|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Medications|11173,11178|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Medications|11173,11183|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|Medications|11173,11183|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Medications|11179,11183|false|false|false|C2598155||pain
Event|Event|Medications|11179,11183|false|false|false|||pain
Finding|Functional Concept|Medications|11179,11183|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Medications|11179,11183|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Medications|11185,11194|false|false|false|||shortness
Attribute|Clinical Attribute|Medications|11185,11204|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|Medications|11185,11204|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|Medications|11198,11204|false|false|false|C0225386|Breath|breath
Event|Event|Medications|11219,11223|false|false|false|||else
Finding|Finding|Medications|11219,11223|false|false|false|C3842296|Else|else
Event|Event|Medications|11232,11241|false|false|false|||troubling
Finding|Finding|Medications|11255,11262|true|false|false|C1551395;C1552745;C1561576|Alert level - Serious;Device Alert Level - Serious;Equipment Alert Level - Serious|serious
Finding|Idea or Concept|Medications|11255,11262|true|false|false|C1551395;C1552745;C1561576|Alert level - Serious;Device Alert Level - Serious;Equipment Alert Level - Serious|serious
Event|Event|Medications|11263,11269|true|false|false|||change
Finding|Functional Concept|Medications|11263,11269|true|false|false|C0392747|Changing|change
Procedure|Therapeutic or Preventive Procedure|Medications|11263,11269|true|false|false|C4319952|Change - procedure|change
Finding|Functional Concept|Medications|11263,11272|true|false|false|C0392747|Changing|change in
Event|Event|Medications|11278,11286|true|false|false|||symptoms
Finding|Functional Concept|Medications|11278,11286|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Medications|11278,11286|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Finding|Medications|11295,11298|true|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Medications|11295,11298|true|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Event|Event|Medications|11299,11307|true|false|false|||symptoms
Finding|Functional Concept|Medications|11299,11307|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Medications|11299,11307|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|Medications|11314,11321|true|false|false|||concern
Finding|Idea or Concept|Medications|11314,11321|true|false|false|C2699424|Concern|concern
Event|Event|Medications|11330,11345|false|false|false|||ANTICOAGULATION
Finding|Finding|Medications|11330,11345|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|ANTICOAGULATION
Finding|Physiologic Function|Medications|11330,11345|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|ANTICOAGULATION
Procedure|Therapeutic or Preventive Procedure|Medications|11330,11345|false|false|false|C0003281|Anticoagulation Therapy|ANTICOAGULATION
Event|Event|Medications|11358,11363|false|false|false|||begin
Event|Event|Medications|11364,11370|false|false|false|||taking
Finding|Idea or Concept|Medications|11376,11380|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Medications|11376,11380|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Medications|11376,11380|false|false|false|C1553498|home health encounter|home
Drug|Hazardous or Poisonous Substance|Medications|11381,11389|false|false|false|C0043031|warfarin|warfarin
Drug|Organic Chemical|Medications|11381,11389|false|false|false|C0043031|warfarin|warfarin
Drug|Pharmacologic Substance|Medications|11381,11389|false|false|false|C0043031|warfarin|warfarin
Attribute|Clinical Attribute|Medications|11381,11394|false|false|false|C4082242||warfarin dose
Procedure|Laboratory Procedure|Medications|11381,11394|false|false|false|C0366686|warfarin dose|warfarin dose
Event|Event|Medications|11390,11394|false|false|false|||dose
Event|Event|Medications|11419,11425|false|false|false|||resume
Finding|Functional Concept|Medications|11419,11425|false|false|false|C1550028;C1880201;C3242342|Curriculum Vitae;Resume - Remote control command;resume - DataOperation|resume
Finding|Idea or Concept|Medications|11419,11425|false|false|false|C1550028;C1880201;C3242342|Curriculum Vitae;Resume - Remote control command;resume - DataOperation|resume
Finding|Intellectual Product|Medications|11419,11425|false|false|false|C1550028;C1880201;C3242342|Curriculum Vitae;Resume - Remote control command;resume - DataOperation|resume
Drug|Hazardous or Poisonous Substance|Medications|11433,11441|false|false|false|C0043031|warfarin|warfarin
Drug|Organic Chemical|Medications|11433,11441|false|false|false|C0043031|warfarin|warfarin
Drug|Pharmacologic Substance|Medications|11433,11441|false|false|false|C0043031|warfarin|warfarin
Event|Event|Medications|11433,11441|false|false|false|||warfarin
Event|Event|Medications|11458,11467|false|false|false|||scheduled
Event|Event|Medications|11469,11474|false|false|false|||doses
Event|Event|Medications|11489,11493|true|false|false|||need
Procedure|Therapeutic or Preventive Procedure|Medications|11496,11502|true|false|false|C0399080|Fixation of dental bridge|bridge
Procedure|Therapeutic or Preventive Procedure|Medications|11496,11510|true|false|false|C5420848|Bridge Therapy|bridge therapy
Event|Event|Medications|11503,11510|true|false|false|||therapy
Finding|Finding|Medications|11503,11510|true|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|Medications|11503,11510|true|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|Medications|11503,11510|true|false|false|C0087111|Therapeutic procedure|therapy
Event|Event|Medications|11514,11519|true|false|false|||begin
Drug|Hazardous or Poisonous Substance|Medications|11520,11528|true|false|false|C0043031|warfarin|warfarin
Drug|Organic Chemical|Medications|11520,11528|true|false|false|C0043031|warfarin|warfarin
Drug|Pharmacologic Substance|Medications|11520,11528|true|false|false|C0043031|warfarin|warfarin
Event|Event|Medications|11520,11528|true|false|false|||warfarin
Drug|Substance|Medications|11532,11537|false|false|false|C1550628|Drain - SpecimenType|DRAIN
Event|Event|Medications|11532,11537|false|false|false|||DRAIN
Finding|Intellectual Product|Medications|11532,11537|false|false|false|C1546604|Drain Specimen Code|DRAIN
Finding|Body Substance|Medications|11538,11547|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|Medications|11538,11547|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|Medications|11538,11547|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|Medications|11538,11547|false|false|false|C0030685|Patient Discharge|DISCHARGE
Attribute|Clinical Attribute|Medications|11538,11560|false|false|false|C3669312||DISCHARGE INSTRUCTIONS
Finding|Intellectual Product|Medications|11538,11560|false|false|false|C4282220|Discharge instructions|DISCHARGE INSTRUCTIONS
Procedure|Health Care Activity|Medications|11538,11560|false|false|false|C2266673|hospital discharge instructions (treatment)|DISCHARGE INSTRUCTIONS
Attribute|Clinical Attribute|Medications|11548,11560|false|false|false|C3263700||INSTRUCTIONS
Event|Event|Medications|11548,11560|false|false|false|||INSTRUCTIONS
Finding|Intellectual Product|Medications|11548,11560|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|INSTRUCTIONS
Event|Event|Medications|11577,11587|false|false|false|||discharged
Event|Event|Medications|11593,11599|false|false|false|||drains
Event|Activity|Medications|11603,11608|false|false|false|C1882509|put - instruction imperative|place
Event|Event|Medications|11603,11608|false|false|false|||place
Finding|Functional Concept|Medications|11603,11608|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|Medications|11603,11608|false|false|false|C1533810||place
Drug|Substance|Medications|11610,11615|false|false|false|C1550628|Drain - SpecimenType|Drain
Finding|Intellectual Product|Medications|11610,11615|false|false|false|C1546604|Drain Specimen Code|Drain
Event|Activity|Medications|11616,11620|false|false|false|C1947933|care activity|care
Event|Event|Medications|11616,11620|false|false|false|||care
Finding|Finding|Medications|11616,11620|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Medications|11616,11620|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Event|Activity|Medications|11627,11632|false|false|false|C1947930|Cleaning (activity)|clean
Attribute|Clinical Attribute|Medications|11633,11642|false|false|false|C0945766||procedure
Event|Event|Medications|11633,11642|false|false|false|||procedure
Event|Occupational Activity|Medications|11633,11642|false|false|false|C1546467|Act Class - procedure|procedure
Finding|Functional Concept|Medications|11633,11642|false|false|false|C2700391|Procedure (set of actions)|procedure
Procedure|Therapeutic or Preventive Procedure|Medications|11633,11642|false|false|false|C0184661|Interventional procedure|procedure
Event|Event|Medications|11644,11648|false|false|false|||Wash
Anatomy|Body Part, Organ, or Organ Component|Medications|11654,11659|false|false|false|C0018563|Hand|hands
Finding|Intellectual Product|Medications|11660,11670|false|false|false|C4708903|Thoroughly|thoroughly
Drug|Biomedical or Dental Material|Medications|11676,11680|false|false|false|C1705308|Soap Dosage Form|soap
Event|Event|Medications|11676,11680|false|false|false|||soap
Event|Event|Medications|11685,11689|false|false|false|||warm
Finding|Finding|Medications|11685,11689|false|false|false|C0582051|Feels warm|warm
Phenomenon|Natural Phenomenon or Process|Medications|11685,11689|false|false|false|C0687712|warming process|warm
Drug|Inorganic Chemical|Medications|11691,11696|false|false|false|C0043047;C1550678|Water Specimen;water|water
Drug|Pharmacologic Substance|Medications|11691,11696|false|false|false|C0043047;C1550678|Water Specimen;water|water
Event|Event|Medications|11691,11696|false|false|false|||water
Finding|Intellectual Product|Medications|11691,11696|false|false|false|C1547961|Water - Specimen Source Codes|water
Procedure|Therapeutic or Preventive Procedure|Medications|11691,11696|false|false|false|C0020311|Hydrotherapy|water
Event|Event|Medications|11704,11714|false|false|false|||performing
Drug|Substance|Medications|11715,11720|false|false|false|C1550628|Drain - SpecimenType|drain
Finding|Intellectual Product|Medications|11715,11720|false|false|false|C1546604|Drain Specimen Code|drain
Event|Activity|Medications|11721,11725|false|false|false|C1947933|care activity|care
Event|Event|Medications|11721,11725|false|false|false|||care
Finding|Finding|Medications|11721,11725|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Medications|11721,11725|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Event|Event|Medications|11735,11743|false|false|false|||drainage
Finding|Body Substance|Medications|11735,11743|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Finding|Sign or Symptom|Medications|11735,11743|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Procedure|Therapeutic or Preventive Procedure|Medications|11735,11743|false|false|false|C0013103|Drainage procedure|drainage
Event|Activity|Medications|11744,11748|false|false|false|C1947933|care activity|care
Event|Event|Medications|11744,11748|false|false|false|||care
Finding|Finding|Medications|11744,11748|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Medications|11744,11748|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Idea or Concept|Medications|11758,11761|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Medications|11758,11761|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Functional Concept|Medications|11770,11775|false|false|false|C5848602|Exhausted|empty
Drug|Substance|Medications|11780,11785|false|false|false|C1550628|Drain - SpecimenType|drain
Event|Event|Medications|11780,11785|false|false|false|||drain
Finding|Intellectual Product|Medications|11780,11785|false|false|false|C1546604|Drain Specimen Code|drain
Finding|Finding|Medications|11798,11802|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Medications|11798,11802|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Medications|11798,11802|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Medications|11808,11811|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Medications|11808,11811|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Finding|Medications|11813,11817|false|false|false|C0580846|Does pull|Pull
Event|Event|Medications|11842,11850|false|false|false|||drainage
Finding|Body Substance|Medications|11842,11850|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Finding|Sign or Symptom|Medications|11842,11850|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Procedure|Therapeutic or Preventive Procedure|Medications|11842,11850|false|false|false|C0013103|Drainage procedure|drainage
Finding|Functional Concept|Medications|11862,11867|false|false|false|C5848602|Exhausted|empty
Event|Event|Medications|11872,11880|false|false|false|||drainage
Finding|Body Substance|Medications|11872,11880|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Finding|Sign or Symptom|Medications|11872,11880|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Procedure|Therapeutic or Preventive Procedure|Medications|11872,11880|false|false|false|C0013103|Drainage procedure|drainage
Drug|Substance|Medications|11882,11887|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|Medications|11882,11887|false|false|false|||fluid
Finding|Intellectual Product|Medications|11882,11887|false|false|false|C1546638|Fluid Specimen Code|fluid
Disorder|Neoplastic Process|Medications|11907,11910|false|false|false|C0220647|Carcinoma of unknown primary|cup
Event|Event|Medications|11912,11918|false|false|false|||Record
Event|Event|Medications|11923,11929|false|false|false|||amount
Finding|Intellectual Product|Medications|11923,11929|false|false|false|C1561574|Amount class - Amount|amount
Event|Event|Medications|11933,11941|false|false|false|||drainage
Finding|Body Substance|Medications|11933,11941|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Finding|Sign or Symptom|Medications|11933,11941|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Procedure|Therapeutic or Preventive Procedure|Medications|11933,11941|false|false|false|C0013103|Drainage procedure|drainage
Drug|Substance|Medications|11943,11948|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|Medications|11943,11948|false|false|false|||fluid
Finding|Intellectual Product|Medications|11943,11948|false|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Intellectual Product|Medications|11956,11962|false|false|false|C0034869|Records|record
Event|Event|Medications|11970,11981|false|false|false|||Reestablish
Drug|Substance|Medications|11982,11987|false|false|false|C1550628|Drain - SpecimenType|drain
Finding|Intellectual Product|Medications|11982,11987|false|false|false|C1546604|Drain Specimen Code|drain
Event|Event|Medications|11988,11995|false|false|false|||suction
Procedure|Therapeutic or Preventive Procedure|Medications|11988,11995|false|false|false|C0038638|Suction drainage|suction
Event|Event|Medications|12006,12012|false|false|false|||assist
Finding|Body Substance|Medications|12013,12020|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Medications|12013,12020|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Medications|12013,12020|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Substance|Medications|12026,12031|false|false|false|C1550628|Drain - SpecimenType|drain
Event|Event|Medications|12026,12031|false|false|false|||drain
Finding|Intellectual Product|Medications|12026,12031|false|false|false|C1546604|Drain Specimen Code|drain
Event|Activity|Medications|12032,12036|false|false|false|C1947933|care activity|care
Event|Event|Medications|12032,12036|false|false|false|||care
Finding|Finding|Medications|12032,12036|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Medications|12032,12036|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Anatomy|Body Part, Organ, or Organ Component|Medications|12046,12049|false|false|false|C0228228|lateral occipital gyrus (human only)|log
Finding|Intellectual Product|Medications|12046,12049|false|false|false|C1708728|Event Log|log
Event|Event|Medications|12053,12063|false|false|false|||individual
Finding|Idea or Concept|Medications|12053,12063|false|false|false|C3245468|Individual - insurance coverage level|individual
Drug|Substance|Medications|12065,12070|false|false|false|C1550628|Drain - SpecimenType|drain
Finding|Intellectual Product|Medications|12065,12070|false|false|false|C1546604|Drain Specimen Code|drain
Event|Event|Medications|12071,12078|false|false|false|||outputs
Event|Event|Medications|12089,12099|false|false|false|||maintained
Event|Event|Medications|12104,12111|false|false|false|||brought
Finding|Body Substance|Medications|12117,12124|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Medications|12117,12124|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Medications|12117,12124|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Medications|12129,12135|false|false|false|||follow
Event|Activity|Medications|12139,12150|false|false|false|C0003629|Appointments|appointment
Event|Event|Medications|12139,12150|false|false|false|||appointment
Attribute|Clinical Attribute|Medications|12161,12168|false|false|false|C5444295||surgeon
Procedure|Health Care Activity|Medications|12173,12181|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Medications|12182,12194|false|false|false|C3263700||Instructions
Event|Event|Medications|12182,12194|false|false|false|||Instructions
Finding|Intellectual Product|Medications|12182,12194|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

