 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|46,55|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|46,55|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|46,60|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|80,89|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|80,89|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|80,94|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|136,139|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|147,154|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|147,154|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|156,164|true|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Finding|Body Substance|Allergies|179,186|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Allergies|179,186|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Allergies|179,186|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Allergies|187,195|true|false|false|||recorded
Attribute|Clinical Attribute|Allergies|215,224|true|false|false|C1717415||Allergies
Event|Event|Allergies|215,224|true|false|false|||Allergies
Finding|Pathologic Function|Allergies|215,224|true|false|false|C0020517|Hypersensitivity|Allergies
Drug|Pharmacologic Substance|Allergies|228,233|true|false|false|C0013227|Pharmaceutical Preparations|Drugs
Event|Event|Allergies|228,233|true|false|false|||Drugs
Procedure|Therapeutic or Preventive Procedure|Allergies|228,233|true|false|false|C3687832|Drugs - dental services|Drugs
Event|Event|Allergies|236,245|true|false|false|||Attending
Finding|Functional Concept|Allergies|236,245|true|false|false|C1999232|Attending (action)|Attending
Finding|Classification|Chief Complaint|275,280|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|281,289|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|281,289|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|293,311|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|302,311|false|false|false|C0945766||Procedure
Event|Event|Chief Complaint|302,311|false|false|false|||Procedure
Event|Occupational Activity|Chief Complaint|302,311|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|302,311|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|302,311|false|false|false|C0184661|Interventional procedure|Procedure
Disorder|Disease or Syndrome|History of Present Illness|366,369|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|366,369|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|History of Present Illness|366,369|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|History of Present Illness|366,369|false|false|false|||CAD
Finding|Gene or Genome|History of Present Illness|366,369|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|History of Present Illness|366,369|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|History of Present Illness|366,369|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|366,369|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Disorder|Disease or Syndrome|History of Present Illness|371,374|false|false|false|C0006430|Burning Mouth Syndrome|BMS
Event|Event|History of Present Illness|371,374|false|false|false|||BMS
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|408,411|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|History of Present Illness|408,411|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Finding|Gene or Genome|History of Present Illness|408,411|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Finding|Functional Concept|History of Present Illness|415,432|false|false|false|C3853134|Poorly controlled|poorly controlled
Event|Event|History of Present Illness|422,432|false|false|false|||controlled
Finding|Gene or Genome|History of Present Illness|433,437|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Finding|Intellectual Product|History of Present Illness|433,437|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Finding|Classification|History of Present Illness|433,439|false|false|false|C0441730|Type 2|type 2
Disorder|Disease or Syndrome|History of Present Illness|440,444|false|false|false|C0011854|Diabetes Mellitus, Insulin-Dependent|IDDM
Event|Event|History of Present Illness|440,444|false|false|false|||IDDM
Disorder|Disease or Syndrome|History of Present Illness|446,449|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|History of Present Illness|446,449|false|false|false|||HTN
Event|Event|History of Present Illness|450,459|false|false|false|||presented
Disorder|Disease or Syndrome|History of Present Illness|463,466|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|463,466|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|History of Present Illness|463,466|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|463,466|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|History of Present Illness|463,466|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|History of Present Illness|463,466|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|History of Present Illness|463,466|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|History of Present Illness|463,466|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|History of Present Illness|463,466|false|false|false|||PCP
Finding|Gene or Genome|History of Present Illness|463,466|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|History of Present Illness|463,466|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Event|History of Present Illness|469,475|false|false|false|||office
Finding|Idea or Concept|History of Present Illness|469,475|false|false|false|C1549636|Address type - Office|office
Event|Event|History of Present Illness|485,494|false|false|false|||reporting
Event|Event|History of Present Illness|495,502|false|false|false|||episode
Finding|Intellectual Product|History of Present Illness|535,539|false|false|false|C1561540|Transaction counts and value totals - week|week
Finding|Body Substance|History of Present Illness|541,548|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|541,548|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|541,548|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|570,579|false|false|false|||increased
Event|Event|History of Present Illness|588,592|false|false|false|||felt
Event|Event|History of Present Illness|593,597|false|false|false|||weak
Finding|Intellectual Product|History of Present Illness|593,597|false|false|false|C3538976;C3714552|Feel Weak (question);Weakness|weak
Finding|Sign or Symptom|History of Present Illness|593,597|false|false|false|C3538976;C3714552|Feel Weak (question);Weakness|weak
Event|Event|History of Present Illness|603,611|false|false|false|||fatigued
Finding|Sign or Symptom|History of Present Illness|603,611|false|false|false|C0015672|Fatigue|fatigued
Event|Event|History of Present Illness|613,619|false|false|false|||Admits
Procedure|Health Care Activity|History of Present Illness|613,619|false|false|false|C0184666|Hospital admission|Admits
Event|Event|History of Present Illness|623,632|false|false|false|||radiation
Phenomenon|Natural Phenomenon or Process|History of Present Illness|623,632|false|false|false|C0034519;C0851346|Electromagnetic Radiation;Radiation|radiation
Procedure|Research Activity|History of Present Illness|623,632|false|false|false|C1522449;C1524020;C1524021|Radiation Ionizing Radiotherapy;Radiation therapy (procedure);Radiotherapy Research|radiation
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|623,632|false|false|false|C1522449;C1524020;C1524021|Radiation Ionizing Radiotherapy;Radiation therapy (procedure);Radiotherapy Research|radiation
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|636,641|false|false|false|C4048756|Right arm|R arm
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|638,641|false|false|false|C0446516;C1140618;C1269078|Upper Extremity;Upper arm|arm
Disorder|Anatomical Abnormality|History of Present Illness|638,641|false|false|false|C3495676|Anorectal Malformations|arm
Event|Event|History of Present Illness|638,641|false|false|false|||arm
Finding|Gene or Genome|History of Present Illness|638,641|false|false|false|C1824218;C3715044|AKR1A1 wt Allele;ARMC9 gene|arm
Procedure|Diagnostic Procedure|History of Present Illness|638,641|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Research Activity|History of Present Illness|638,641|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|638,641|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Finding|Body Substance|History of Present Illness|671,678|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|671,678|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|671,678|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|679,683|false|false|false|||felt
Finding|Sign or Symptom|History of Present Illness|679,689|false|false|false|C0581879|Felt faint|felt faint
Event|Event|History of Present Illness|684,689|false|false|false|||faint
Finding|Finding|History of Present Illness|684,689|false|false|false|C0039070;C4554554|Faint - appearance;Syncope|faint
Finding|Sign or Symptom|History of Present Illness|684,689|false|false|false|C0039070;C4554554|Faint - appearance;Syncope|faint
Anatomy|Body Location or Region|History of Present Illness|702,707|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|702,707|false|false|false|C0741025|Chest problem|chest
Finding|Sign or Symptom|History of Present Illness|702,717|false|false|false|C0232292|Chest tightness|chest tightness
Event|Event|History of Present Illness|708,717|false|false|false|||tightness
Event|Event|History of Present Illness|720,728|false|false|false|||relieved
Event|Event|History of Present Illness|739,742|false|false|false|||NTG
Finding|Finding|History of Present Illness|739,742|false|false|false|C1417953;C1847730;C5575300|GLAUCOMA, NORMAL TENSION, SUSCEPTIBILITY TO;OPA1 gene;OPA1 wt Allele|NTG
Finding|Gene or Genome|History of Present Illness|739,742|false|false|false|C1417953;C1847730;C5575300|GLAUCOMA, NORMAL TENSION, SUSCEPTIBILITY TO;OPA1 gene;OPA1 wt Allele|NTG
Event|Event|History of Present Illness|744,750|true|false|false|||Denies
Event|Event|History of Present Illness|766,769|true|false|false|||SOB
Finding|Sign or Symptom|History of Present Illness|766,769|true|false|false|C0013404|Dyspnea|SOB
Event|Event|History of Present Illness|771,782|true|false|false|||Diaphoresis
Finding|Finding|History of Present Illness|771,782|true|false|false|C0700590|Increased sweating|Diaphoresis
Finding|Body Substance|History of Present Illness|785,792|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|785,792|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|785,792|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|History of Present Illness|794,795|false|false|false|||/
Event|Event|History of Present Illness|826,831|false|false|false|||feels
Event|Event|History of Present Illness|839,842|false|false|false|||SOB
Finding|Sign or Symptom|History of Present Illness|839,842|false|false|false|C0013404|Dyspnea|SOB
Finding|Body Substance|History of Present Illness|857,864|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|857,864|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|857,864|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|867,869|false|false|false|||VS
Finding|Body Substance|History of Present Illness|910,917|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|910,917|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|910,917|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Organic Chemical|History of Present Illness|925,931|false|false|false|C0723011|Relief brand of phenylephrine|relief
Drug|Pharmacologic Substance|History of Present Illness|925,931|false|false|false|C0723011|Relief brand of phenylephrine|relief
Event|Event|History of Present Illness|925,931|false|false|false|||relief
Finding|Finding|History of Present Illness|925,931|false|false|false|C0564405|Feeling relief|relief
Event|Event|History of Present Illness|940,943|false|false|false|||NTG
Finding|Finding|History of Present Illness|940,943|false|false|false|C1417953;C1847730;C5575300|GLAUCOMA, NORMAL TENSION, SUSCEPTIBILITY TO;OPA1 gene;OPA1 wt Allele|NTG
Finding|Gene or Genome|History of Present Illness|940,943|false|false|false|C1417953;C1847730;C5575300|GLAUCOMA, NORMAL TENSION, SUSCEPTIBILITY TO;OPA1 gene;OPA1 wt Allele|NTG
Event|Event|History of Present Illness|948,956|true|false|false|||transfer
Finding|Functional Concept|History of Present Illness|948,956|true|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|History of Present Illness|948,956|true|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|History of Present Illness|948,956|true|false|false|C4706767|Transfer (immobility management)|transfer
Anatomy|Anatomical Structure|History of Present Illness|960,965|true|false|false|C3714591|Floor (anatomic)|floor
Finding|Body Substance|History of Present Illness|967,974|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|967,974|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|967,974|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Anatomy|Body Location or Region|History of Present Illness|983,988|true|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|983,988|true|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|History of Present Illness|983,993|true|false|false|C2926613||chest pain
Finding|Sign or Symptom|History of Present Illness|983,993|true|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|History of Present Illness|989,993|true|false|false|C2598155||pain
Event|Event|History of Present Illness|989,993|true|false|false|||pain
Finding|Functional Concept|History of Present Illness|989,993|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|989,993|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Body Substance|History of Present Illness|1001,1008|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|1001,1008|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|1001,1008|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|History of Present Illness|1009,1015|true|false|false|||denies
Event|Event|History of Present Illness|1020,1021|true|false|false|||N
Event|Event|History of Present Illness|1029,1031|true|false|false|||CP
Event|Event|History of Present Illness|1033,1036|false|false|false|||SOB
Finding|Sign or Symptom|History of Present Illness|1033,1036|true|false|false|C0013404|Dyspnea|SOB
Finding|Finding|History of Present Illness|1048,1057|false|false|false|C5425799|All other|All other
Anatomy|Body Space or Junction|History of Present Illness|1058,1061|false|false|false|C0262327|rostral sulcus|ROS
Drug|Biologically Active Substance|History of Present Illness|1058,1061|false|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Drug|Element, Ion, or Isotope|History of Present Illness|1058,1061|false|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Drug|Organic Chemical|History of Present Illness|1058,1061|false|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Drug|Pharmacologic Substance|History of Present Illness|1058,1061|false|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Event|Event|History of Present Illness|1058,1061|false|false|false|||ROS
Finding|Gene or Genome|History of Present Illness|1058,1061|false|false|false|C0812281;C1709820|ROS1 gene;ROS1 wt Allele|ROS
Procedure|Health Care Activity|History of Present Illness|1058,1061|false|false|false|C0489633|Review of systems (procedure)|ROS
Event|Event|History of Present Illness|1063,1071|false|false|false|||negative
Finding|Classification|History of Present Illness|1063,1071|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|History of Present Illness|1063,1071|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|History of Present Illness|1063,1071|false|false|false|C5237010|Expression Negative|negative
Event|Event|History of Present Illness|1089,1098|false|false|false|||specified
Disorder|Disease or Syndrome|Past Medical History|1125,1131|false|false|false|C0004096|Asthma|asthma
Event|Event|Past Medical History|1125,1131|false|false|false|||asthma
Disorder|Disease or Syndrome|Past Medical History|1133,1142|false|false|false|C0034067|Pulmonary Emphysema|emphysema
Event|Event|Past Medical History|1133,1142|false|false|false|||emphysema
Finding|Pathologic Function|Past Medical History|1133,1142|false|false|false|C0013990|Pathological accumulation of air in tissues|emphysema
Event|Event|Past Medical History|1144,1151|false|false|false|||chronic
Finding|Intellectual Product|Past Medical History|1144,1151|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|Past Medical History|1144,1151|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Disorder|Disease or Syndrome|Past Medical History|1144,1162|false|false|false|C0008677|Bronchitis, Chronic|chronic bronchitis
Disorder|Disease or Syndrome|Past Medical History|1152,1162|false|false|false|C0006277;C0149514|Acute bronchitis;Bronchitis|bronchitis
Event|Event|Past Medical History|1152,1162|false|false|false|||bronchitis
Disorder|Disease or Syndrome|Past Medical History|1164,1167|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|Past Medical History|1164,1167|false|false|false|||HTN
Disorder|Disease or Syndrome|Past Medical History|1169,1172|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Past Medical History|1169,1172|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Past Medical History|1169,1172|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|Past Medical History|1169,1172|false|false|false|||CAD
Finding|Gene or Genome|Past Medical History|1169,1172|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Past Medical History|1169,1172|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Past Medical History|1169,1172|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1169,1172|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Event|Event|Past Medical History|1174,1178|false|false|false|||MIx2
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1182,1189|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|Past Medical History|1182,1189|false|false|false|C1314974|Cardiac attachment|cardiac
Event|Event|Past Medical History|1190,1196|false|false|false|||stents
Disorder|Disease or Syndrome|Past Medical History|1202,1211|false|false|false|C0149931|Migraine Disorders|migraines
Event|Event|Past Medical History|1202,1211|false|false|false|||migraines
Disorder|Disease or Syndrome|Past Medical History|1213,1217|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Event|Event|Past Medical History|1213,1217|false|false|false|||GERD
Drug|Biomedical or Dental Material|Past Medical History|1229,1234|false|false|false|C0994475|Pills|pills
Event|Event|Past Medical History|1229,1234|false|false|false|||pills
Drug|Amino Acid, Peptide, or Protein|Past Medical History|1239,1246|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|Past Medical History|1239,1246|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|Past Medical History|1239,1246|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|Past Medical History|1239,1246|false|false|false|||insulin
Finding|Gene or Genome|Past Medical History|1239,1246|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|Past Medical History|1239,1246|false|false|false|C0202098|Insulin measurement|insulin
Disorder|Disease or Syndrome|Past Medical History|1249,1255|false|false|false|C0002871|Anemia|Anemia
Event|Event|Past Medical History|1249,1255|false|false|false|||Anemia
Disorder|Disease or Syndrome|Past Medical History|1257,1267|false|false|false|C0442874|Neuropathy|neuropathy
Event|Event|Past Medical History|1257,1267|false|false|false|||neuropathy
Disorder|Mental or Behavioral Dysfunction|Past Medical History|1269,1276|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Event|Event|Past Medical History|1269,1276|false|false|false|||anxiety
Finding|Sign or Symptom|Past Medical History|1269,1276|false|false|false|C0860603|Anxiety symptoms|anxiety
Event|Event|Family Medical History|1328,1333|true|false|false|||known
Disorder|Disease or Syndrome|Family Medical History|1344,1347|false|false|false|C0020538|Hypertensive disease|htn
Event|Event|Family Medical History|1344,1347|false|false|false|||htn
Event|Event|Family Medical History|1353,1361|false|false|false|||Physical
Finding|Finding|Family Medical History|1353,1361|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|Family Medical History|1353,1361|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|Family Medical History|1353,1361|false|false|false|C0031809|Physical Examination|Physical
Finding|Classification|Family Medical History|1402,1405|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Finding|Gene or Genome|Family Medical History|1402,1405|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Event|Event|Family Medical History|1412,1418|false|false|false|||middle
Finding|Intellectual Product|Family Medical History|1412,1418|false|false|false|C1552826|Table Cell Vertical Align - middle|middle
Event|Event|Family Medical History|1424,1428|false|false|false|||male
Finding|Finding|Family Medical History|1424,1428|false|false|false|C1706180|Male Gender|male
Disorder|Disease or Syndrome|Family Medical History|1432,1435|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|Family Medical History|1432,1435|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|Family Medical History|1432,1435|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Family Medical History|1432,1435|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|Family Medical History|1432,1435|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|Family Medical History|1432,1435|false|false|false|||NAD
Finding|Finding|Family Medical History|1432,1435|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Finding|Finding|Family Medical History|1437,1445|false|false|false|C1961028|Oriented to place|Oriented
Attribute|Clinical Attribute|Family Medical History|1450,1454|false|false|false|C2713234||Mood
Event|Event|Family Medical History|1450,1454|false|false|false|||Mood
Finding|Conceptual Entity|Family Medical History|1450,1454|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|Mood
Finding|Finding|Family Medical History|1450,1454|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|Mood
Finding|Mental Process|Family Medical History|1450,1454|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|Mood
Event|Event|Family Medical History|1456,1462|false|false|false|||affect
Finding|Mental Process|Family Medical History|1456,1462|false|false|false|C0001721|Affect (mental function)|affect
Procedure|Health Care Activity|Family Medical History|1456,1462|false|false|false|C2237113|assessment of affect|affect
Event|Event|Family Medical History|1464,1475|false|false|false|||appropriate
Anatomy|Body Location or Region|Family Medical History|1479,1484|false|false|false|C1512338|HEENT|HEENT
Event|Event|Family Medical History|1486,1490|false|false|false|||NCAT
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1492,1498|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|Family Medical History|1492,1498|false|false|false|C0036412|Scleral Diseases|Sclera
Event|Event|Family Medical History|1492,1498|false|false|false|||Sclera
Procedure|Health Care Activity|Family Medical History|1492,1498|false|false|false|C2228481|examination of sclera|Sclera
Event|Event|Family Medical History|1499,1508|false|false|false|||anicteric
Finding|Finding|Family Medical History|1499,1508|false|false|false|C0205180|Anicteric|anicteric
Event|Event|Family Medical History|1510,1515|false|false|false|||PERRL
Finding|Finding|Family Medical History|1510,1515|false|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Event|Event|Family Medical History|1517,1521|false|false|false|||EOMI
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1523,1534|true|false|false|C0009758;C0229274|Structure of palpebral conjunctiva;conjunctiva|Conjunctiva
Disorder|Disease or Syndrome|Family Medical History|1523,1534|true|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|Conjunctiva
Disorder|Neoplastic Process|Family Medical History|1523,1534|true|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|Conjunctiva
Event|Event|Family Medical History|1523,1534|true|false|false|||Conjunctiva
Finding|Body Substance|Family Medical History|1523,1534|true|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|Conjunctiva
Finding|Intellectual Product|Family Medical History|1523,1534|true|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|Conjunctiva
Procedure|Health Care Activity|Family Medical History|1523,1534|true|false|false|C0872390;C2228431|Procedure on conjunctiva;examination of conjunctiva|Conjunctiva
Event|Event|Family Medical History|1550,1556|true|false|false|||pallor
Finding|Finding|Family Medical History|1550,1556|true|false|false|C0241137|Pallor of skin|pallor
Event|Event|Family Medical History|1560,1568|true|false|false|||cyanosis
Finding|Sign or Symptom|Family Medical History|1560,1568|true|false|false|C0010520|Cyanosis|cyanosis
Anatomy|Body Space or Junction|Family Medical History|1576,1580|true|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Family Medical History|1576,1580|true|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Family Medical History|1576,1580|true|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Family Medical History|1576,1580|true|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1576,1587|true|false|false|C0026639|Oral mucous membrane structure|oral mucosa
Anatomy|Tissue|Family Medical History|1581,1587|true|false|false|C0026724|Mucous Membrane|mucosa
Finding|Intellectual Product|Family Medical History|1581,1587|true|false|false|C1561514||mucosa
Event|Event|Family Medical History|1592,1603|true|false|false|||xanthalesma
Anatomy|Body Location or Region|Family Medical History|1608,1612|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Anatomy|Cell Component|Family Medical History|1608,1612|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Finding|Finding|Family Medical History|1608,1612|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|Neck
Event|Event|Family Medical History|1617,1620|true|false|false|||JVD
Finding|Finding|Family Medical History|1617,1620|true|false|false|C0425687|Jugular venous engorgement|JVD
Event|Event|Family Medical History|1653,1654|true|false|false|||g
Event|Event|Family Medical History|1659,1666|true|false|false|||thrills
Finding|Finding|Family Medical History|1659,1666|true|false|false|C0232269|Cardiac thrill (finding)|thrills
Event|Event|Family Medical History|1668,1673|true|false|false|||lifts
Anatomy|Body Location or Region|Family Medical History|1691,1696|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|Family Medical History|1691,1696|false|false|false|C0741025|Chest problem|Chest
Drug|Organic Chemical|Family Medical History|1698,1702|true|false|false|C0951233|cetrimonium bromide|CTAB
Event|Event|Family Medical History|1698,1702|true|false|false|||CTAB
Event|Event|Family Medical History|1707,1715|true|false|false|||crackles
Finding|Finding|Family Medical History|1707,1715|true|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Event|Event|Family Medical History|1717,1724|true|false|false|||wheezes
Finding|Sign or Symptom|Family Medical History|1717,1724|true|false|false|C0043144|Wheezing|wheezes
Event|Event|Family Medical History|1728,1735|true|false|false|||rhonchi
Finding|Finding|Family Medical History|1728,1735|true|false|false|C0035508|Rhonchi|rhonchi
Anatomy|Body Location or Region|Family Medical History|1739,1742|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|Abd
Disorder|Cell or Molecular Dysfunction|Family Medical History|1739,1742|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|Abd
Disorder|Disease or Syndrome|Family Medical History|1744,1748|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Event|Event|Family Medical History|1744,1748|false|false|false|||Soft
Event|Event|Family Medical History|1750,1754|false|false|false|||NTND
Event|Event|Family Medical History|1759,1762|true|false|false|||HSM
Finding|Gene or Genome|Family Medical History|1759,1762|true|false|false|C1537594|LRRC4B gene|HSM
Event|Event|Family Medical History|1766,1776|true|false|false|||tenderness
Finding|Mental Process|Family Medical History|1766,1776|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|Family Medical History|1766,1776|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Anatomy|Body Location or Region|Family Medical History|1778,1781|true|false|false|C0000726;C0449202|ABD (body structure);Abdomen|Abd
Disorder|Cell or Molecular Dysfunction|Family Medical History|1778,1781|true|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|Abd
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1782,1787|true|false|false|C0003483;C4037978|Aorta;Chest+Abdomen>Aorta|aorta
Procedure|Health Care Activity|Family Medical History|1782,1787|true|false|false|C0869784|Procedure on aorta|aorta
Event|Event|Family Medical History|1792,1800|true|false|false|||enlarged
Event|Event|Family Medical History|1805,1814|true|false|false|||palpation
Procedure|Diagnostic Procedure|Family Medical History|1805,1814|true|false|false|C0030247|Palpation|palpation
Event|Event|Family Medical History|1830,1836|true|false|false|||bruits
Finding|Finding|Family Medical History|1830,1836|true|false|false|C0006318|Bruit|bruits
Disorder|Congenital Abnormality|Family Medical History|1840,1843|false|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Event|Event|Family Medical History|1840,1843|false|false|false|||Ext
Finding|Gene or Genome|Family Medical History|1840,1843|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1858,1865|true|false|false|C0015811|Femur|femoral
Event|Event|Family Medical History|1866,1872|true|false|false|||bruits
Finding|Finding|Family Medical History|1866,1872|true|false|false|C0006318|Bruit|bruits
Anatomy|Body System|Family Medical History|1876,1880|false|false|false|C1123023;C4520765|Skin;Skin, Human|Skin
Disorder|Disease or Syndrome|Family Medical History|1876,1880|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|Skin
Disorder|Neoplastic Process|Family Medical History|1876,1880|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|Skin
Finding|Body Substance|Family Medical History|1876,1880|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|Skin
Finding|Intellectual Product|Family Medical History|1876,1880|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|Skin
Finding|Pathologic Function|Family Medical History|1885,1891|true|false|false|C0333138|Stasis|stasis
Disorder|Disease or Syndrome|Family Medical History|1885,1902|true|false|false|C0011620|Stasis dermatitis|stasis dermatitis
Disorder|Disease or Syndrome|Family Medical History|1892,1902|true|false|false|C0011603|Dermatitis|dermatitis
Event|Event|Family Medical History|1892,1902|true|false|false|||dermatitis
Event|Event|Family Medical History|1904,1910|true|false|false|||ulcers
Finding|Pathologic Function|Family Medical History|1904,1910|true|false|false|C0041582|Ulcer|ulcers
Event|Event|Family Medical History|1912,1917|true|false|false|||scars
Finding|Finding|Family Medical History|1912,1917|true|false|false|C0241158;C2004491|Cicatrix;Scar Tissue|scars
Finding|Pathologic Function|Family Medical History|1912,1917|true|false|false|C0241158;C2004491|Cicatrix;Scar Tissue|scars
Disorder|Disease or Syndrome|Family Medical History|1922,1931|true|false|false|C0302314|Xanthoma|xanthomas
Event|Event|Family Medical History|1922,1931|false|false|false|||xanthomas
Drug|Food|Family Medical History|1939,1945|false|false|false|C5890763||Pulses
Event|Event|Family Medical History|1939,1945|false|false|false|||Pulses
Finding|Physiologic Function|Family Medical History|1939,1945|false|false|false|C0391850|Physiologic pulse|Pulses
Procedure|Health Care Activity|Family Medical History|1939,1945|false|false|false|C0034107|Pulse taking|Pulses
Finding|Functional Concept|Family Medical History|1949,1954|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1956,1963|false|false|false|C0007272|Carotid Arteries|Carotid
Finding|Functional Concept|Family Medical History|1982,1986|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1988,1995|false|false|false|C0007272|Carotid Arteries|Carotid
Attribute|Clinical Attribute|Family Medical History|2040,2046|false|false|false|C1718621|W stress|Stress
Drug|Organic Chemical|Family Medical History|2040,2046|false|false|false|C0723460|Stress bismuth subsalicylate|Stress
Drug|Pharmacologic Substance|Family Medical History|2040,2046|false|false|false|C0723460|Stress bismuth subsalicylate|Stress
Event|Event|Family Medical History|2040,2046|false|false|false|||Stress
Finding|Finding|Family Medical History|2040,2046|false|false|false|C0038435|Stress|Stress
Attribute|Clinical Attribute|Family Medical History|2047,2061|false|false|false|C3173575||INTERPRETATION
Event|Event|Family Medical History|2047,2061|false|false|false|||INTERPRETATION
Finding|Intellectual Product|Family Medical History|2047,2061|false|false|false|C0459471|Interpretation Process|INTERPRETATION
Finding|Gene or Genome|Family Medical History|2075,2079|false|true|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|Type
Finding|Intellectual Product|Family Medical History|2075,2079|false|true|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|Type
Disorder|Disease or Syndrome|Family Medical History|2083,2087|false|false|false|C0011854|Diabetes Mellitus, Insulin-Dependent|IDDM
Event|Event|Family Medical History|2083,2087|false|false|false|||IDDM
Event|Event|Family Medical History|2113,2118|false|false|false|||stent
Event|Event|Family Medical History|2130,2138|false|false|false|||referred
Event|Event|Family Medical History|2143,2153|false|false|false|||evaluation
Finding|Idea or Concept|Family Medical History|2143,2153|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|Family Medical History|2143,2153|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Anatomy|Body Location or Region|Family Medical History|2157,2162|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Family Medical History|2157,2162|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Family Medical History|2157,2167|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|Family Medical History|2157,2167|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Family Medical History|2163,2167|false|false|false|C2598155||pain
Event|Event|Family Medical History|2163,2167|false|false|false|||pain
Finding|Functional Concept|Family Medical History|2163,2167|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Family Medical History|2163,2167|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Body Substance|Family Medical History|2174,2181|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Family Medical History|2174,2181|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Family Medical History|2174,2181|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Family Medical History|2187,2194|false|false|false|||infused
Finding|Conceptual Entity|Family Medical History|2208,2214|false|false|false|C1532757|kg/min|kg/min
Drug|Organic Chemical|Family Medical History|2218,2228|false|false|false|C0700020|Persantine|persantine
Drug|Pharmacologic Substance|Family Medical History|2218,2228|false|false|false|C0700020|Persantine|persantine
Event|Event|Family Medical History|2218,2228|false|false|false|||persantine
Event|Event|Family Medical History|2254,2262|false|false|false|||infusion
Finding|Functional Concept|Family Medical History|2254,2262|false|false|false|C1827465|Infusion route|infusion
Procedure|Therapeutic or Preventive Procedure|Family Medical History|2254,2262|false|false|false|C0574032|Infusion procedures|infusion
Finding|Body Substance|Family Medical History|2268,2275|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Family Medical History|2268,2275|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Family Medical History|2268,2275|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Family Medical History|2276,2284|false|false|false|||reported
Anatomy|Body Location or Region|Family Medical History|2301,2306|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Family Medical History|2301,2306|false|false|false|C0741025|Chest problem|chest
Event|Event|Family Medical History|2308,2316|false|false|false|||pressure
Finding|Finding|Family Medical History|2308,2316|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|Family Medical History|2308,2316|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|Family Medical History|2308,2316|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|Family Medical History|2308,2316|false|false|false|C0033095||pressure
Event|Event|Family Medical History|2330,2339|false|false|false|||increased
Event|Event|Family Medical History|2354,2365|false|false|false|||inspiration
Finding|Organism Function|Family Medical History|2354,2365|false|false|false|C0004048|Inspiration (function)|inspiration
Attribute|Clinical Attribute|Family Medical History|2372,2379|false|false|false|C3854129||symptom
Event|Event|Family Medical History|2372,2379|false|false|false|||symptom
Finding|Sign or Symptom|Family Medical History|2372,2379|false|false|false|C1457887|Symptoms|symptom
Event|Event|Family Medical History|2385,2393|false|false|false|||relieved
Event|Event|Family Medical History|2401,2406|false|false|false|||125mg
Drug|Organic Chemical|Family Medical History|2413,2426|false|false|false|C0002575|aminophylline|aminophylline
Drug|Pharmacologic Substance|Family Medical History|2413,2426|false|false|false|C0002575|aminophylline|aminophylline
Event|Event|Family Medical History|2413,2426|false|false|false|||aminophylline
Finding|Finding|Family Medical History|2413,2436|false|false|false|C2024835||aminophylline was given
Event|Event|Family Medical History|2431,2436|false|false|false|||given
Drug|Biomedical or Dental Material|Family Medical History|2450,2459|false|false|false|C1272883|Injection|injection
Event|Event|Family Medical History|2450,2459|false|false|false|||injection
Finding|Functional Concept|Family Medical History|2450,2459|false|false|false|C1828121|Injection Route of Administration|injection
Procedure|Therapeutic or Preventive Procedure|Family Medical History|2450,2459|false|false|false|C0021485;C1533685|Injection of therapeutic agent;Injection procedure|injection
Finding|Idea or Concept|Family Medical History|2465,2476|true|false|false|C0750502|Significant|significant
Finding|Finding|Family Medical History|2477,2487|true|false|false|C0429029|ST segment|ST segment
Event|Event|Family Medical History|2488,2495|true|false|false|||changes
Finding|Functional Concept|Family Medical History|2488,2495|true|false|false|C0392747|Changing|changes
Event|Event|Family Medical History|2501,2506|true|false|false|||noted
Event|Event|Family Medical History|2512,2518|true|false|false|||rhythm
Finding|Finding|Family Medical History|2512,2518|true|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|Family Medical History|2512,2518|true|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Anatomy|Body Space or Junction|Family Medical History|2523,2528|true|false|false|C0030471;C1305231|Nasal sinus;Sinus - general anatomical term|sinus
Disorder|Anatomical Abnormality|Family Medical History|2523,2528|true|false|false|C0016169|pathologic fistula|sinus
Drug|Organic Chemical|Family Medical History|2523,2528|true|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Drug|Pharmacologic Substance|Family Medical History|2523,2528|true|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Event|Event|Family Medical History|2523,2528|true|false|false|||sinus
Event|Event|Family Medical History|2539,2545|true|false|false|||ectopy
Finding|Organ or Tissue Function|Family Medical History|2547,2558|false|false|false|C0019010|Hemodynamics|Hemodynamic
Procedure|Laboratory Procedure|Family Medical History|2547,2558|false|false|false|C4281788|hemodynamics (procedure)|Hemodynamic
Event|Event|Family Medical History|2559,2567|false|false|false|||response
Finding|Finding|Family Medical History|2559,2567|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Intellectual Product|Family Medical History|2559,2567|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Mental Process|Family Medical History|2559,2567|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Event|Event|Family Medical History|2571,2579|false|false|false|||infusion
Finding|Functional Concept|Family Medical History|2571,2579|false|false|false|C1827465|Infusion route|infusion
Procedure|Therapeutic or Preventive Procedure|Family Medical History|2571,2579|false|false|false|C0574032|Infusion procedures|infusion
Event|Event|Family Medical History|2584,2595|false|false|false|||appropriate
Event|Event|Family Medical History|2601,2611|false|false|false|||IMPRESSION
Finding|Intellectual Product|Family Medical History|2601,2611|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|Family Medical History|2601,2611|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Finding|Family Medical History|2613,2621|false|false|false|C0332149|Possible|Possible
Finding|Gene or Genome|Family Medical History|2630,2634|false|true|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Finding|Intellectual Product|Family Medical History|2630,2634|false|true|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Event|Event|Family Medical History|2635,2643|false|false|false|||symptoms
Finding|Functional Concept|Family Medical History|2635,2643|false|true|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Family Medical History|2635,2643|false|true|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Disorder|Anatomical Abnormality|Family Medical History|2651,2658|false|false|false|C1689985|Absence (morphologic abnormality)|absence
Event|Event|Family Medical History|2651,2658|false|false|false|||absence
Finding|Functional Concept|Family Medical History|2651,2658|false|false|false|C0332197|Absent|absence
Finding|Functional Concept|Family Medical History|2651,2661|false|false|false|C0332197|Absent|absence of
Finding|Functional Concept|Family Medical History|2663,2671|false|false|false|C0475224|Ischemic|ischemic
Event|Event|Family Medical History|2673,2676|false|false|false|||EKG
Finding|Intellectual Product|Family Medical History|2673,2676|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|Family Medical History|2673,2676|false|false|false|C1623258|Electrocardiography|EKG
Event|Event|Family Medical History|2677,2684|false|false|false|||changes
Finding|Functional Concept|Family Medical History|2677,2684|false|false|false|C0392747|Changing|changes
Attribute|Clinical Attribute|Family Medical History|2694,2700|false|false|false|C4255046||report
Event|Event|Family Medical History|2694,2700|false|false|false|||report
Finding|Intellectual Product|Family Medical History|2694,2700|false|false|false|C0684224|Report (document)|report
Procedure|Health Care Activity|Family Medical History|2694,2700|false|false|false|C0700287|Reporting|report
Event|Event|Family Medical History|2701,2705|false|false|false|||sent
Event|Event|Family Medical History|2722,2732|false|false|false|||IMPRESSION
Finding|Intellectual Product|Family Medical History|2722,2732|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|Family Medical History|2722,2732|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Anatomy|Tissue|Family Medical History|2741,2751|false|false|false|C0027061|Myocardium|myocardial
Event|Event|Family Medical History|2752,2761|false|false|false|||perfusion
Finding|Functional Concept|Family Medical History|2752,2761|false|false|false|C4281794;C4723760|Perfusion (biological);Perfusion route|perfusion
Finding|Organism Function|Family Medical History|2752,2761|false|false|false|C4281794;C4723760|Perfusion (biological);Perfusion route|perfusion
Procedure|Therapeutic or Preventive Procedure|Family Medical History|2752,2761|false|false|false|C0031001;C4721534|Chemotherapeutic Perfusion;Perfusion (procedure)|perfusion
Event|Event|Family Medical History|2766,2774|false|false|false|||function
Finding|Finding|Family Medical History|2766,2774|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|Family Medical History|2766,2774|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|Family Medical History|2766,2774|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|Family Medical History|2766,2774|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Disorder|Disease or Syndrome|Family Medical History|2798,2803|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|2798,2803|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|2798,2803|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|Family Medical History|2804,2807|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|Family Medical History|2812,2815|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|Family Medical History|2812,2815|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|Family Medical History|2812,2815|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|Family Medical History|2822,2825|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|Family Medical History|2822,2825|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|Family Medical History|2822,2825|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|Family Medical History|2822,2825|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|Family Medical History|2831,2834|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|Family Medical History|2831,2834|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|Family Medical History|2841,2844|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|Family Medical History|2841,2844|false|false|false|||MCV
Lab|Laboratory or Test Result|Family Medical History|2841,2844|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|Family Medical History|2841,2844|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|Family Medical History|2841,2844|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|Family Medical History|2848,2851|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|Family Medical History|2848,2851|false|false|false|C0600370|methacholine|MCH
Event|Event|Family Medical History|2848,2851|false|false|false|||MCH
Finding|Gene or Genome|Family Medical History|2848,2851|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|Family Medical History|2848,2851|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|Family Medical History|2848,2851|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|Family Medical History|2858,2862|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|Family Medical History|2878,2881|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|Family Medical History|2898,2903|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|2898,2903|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|2898,2903|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|Family Medical History|2904,2907|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|Family Medical History|2912,2915|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|Family Medical History|2912,2915|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|Family Medical History|2912,2915|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|Family Medical History|2922,2925|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|Family Medical History|2922,2925|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|Family Medical History|2922,2925|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|Family Medical History|2922,2925|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|Family Medical History|2931,2934|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|Family Medical History|2931,2934|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|Family Medical History|2942,2945|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|Family Medical History|2942,2945|false|false|false|||MCV
Lab|Laboratory or Test Result|Family Medical History|2942,2945|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|Family Medical History|2942,2945|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|Family Medical History|2942,2945|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|Family Medical History|2949,2952|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|Family Medical History|2949,2952|false|false|false|C0600370|methacholine|MCH
Event|Event|Family Medical History|2949,2952|false|false|false|||MCH
Finding|Gene or Genome|Family Medical History|2949,2952|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|Family Medical History|2949,2952|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|Family Medical History|2949,2952|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|Family Medical History|2959,2963|false|true|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|Family Medical History|2979,2982|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|Family Medical History|2999,3004|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|2999,3004|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|2999,3004|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|Family Medical History|3005,3008|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|Family Medical History|3013,3016|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|Family Medical History|3013,3016|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|Family Medical History|3013,3016|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|Family Medical History|3023,3026|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|Family Medical History|3023,3026|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|Family Medical History|3023,3026|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|Family Medical History|3023,3026|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|Family Medical History|3032,3035|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|Family Medical History|3032,3035|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|Family Medical History|3043,3046|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|Family Medical History|3043,3046|false|false|false|||MCV
Lab|Laboratory or Test Result|Family Medical History|3043,3046|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|Family Medical History|3043,3046|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|Family Medical History|3043,3046|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|Family Medical History|3050,3053|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|Family Medical History|3050,3053|false|false|false|C0600370|methacholine|MCH
Event|Event|Family Medical History|3050,3053|false|false|false|||MCH
Finding|Gene or Genome|Family Medical History|3050,3053|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|Family Medical History|3050,3053|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|Family Medical History|3050,3053|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|Family Medical History|3060,3064|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|Family Medical History|3080,3083|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|Family Medical History|3100,3105|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|3100,3105|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|3100,3105|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|Family Medical History|3106,3109|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|Family Medical History|3126,3131|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|Family Medical History|3126,3131|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|Family Medical History|3132,3135|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|Family Medical History|3152,3157|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|3152,3157|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|3152,3157|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|Family Medical History|3158,3161|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|Family Medical History|3178,3183|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|3178,3183|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|3178,3183|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|Family Medical History|3178,3191|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|Family Medical History|3178,3191|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|Family Medical History|3178,3191|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|Family Medical History|3184,3191|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|Family Medical History|3184,3191|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|Family Medical History|3184,3191|false|false|false|C0017725|glucose|Glucose
Event|Event|Family Medical History|3184,3191|false|false|false|||Glucose
Lab|Laboratory or Test Result|Family Medical History|3184,3191|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|Family Medical History|3184,3191|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|Family Medical History|3236,3240|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|Family Medical History|3236,3240|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|Family Medical History|3236,3240|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|Family Medical History|3265,3270|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|3265,3270|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|3265,3270|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|Family Medical History|3265,3278|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|Family Medical History|3265,3278|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|Family Medical History|3265,3278|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|Family Medical History|3271,3278|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|Family Medical History|3271,3278|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|Family Medical History|3271,3278|false|false|false|C0017725|glucose|Glucose
Event|Event|Family Medical History|3271,3278|false|false|false|||Glucose
Lab|Laboratory or Test Result|Family Medical History|3271,3278|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|Family Medical History|3271,3278|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|Family Medical History|3322,3326|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|Family Medical History|3322,3326|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|Family Medical History|3322,3326|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|Family Medical History|3351,3356|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|3351,3356|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|3351,3356|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|Family Medical History|3351,3364|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|Family Medical History|3351,3364|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|Family Medical History|3351,3364|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|Family Medical History|3357,3364|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|Family Medical History|3357,3364|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|Family Medical History|3357,3364|false|false|false|C0017725|glucose|Glucose
Event|Event|Family Medical History|3357,3364|false|false|false|||Glucose
Lab|Laboratory or Test Result|Family Medical History|3357,3364|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|Family Medical History|3357,3364|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|Family Medical History|3411,3415|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|Family Medical History|3411,3415|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|Family Medical History|3411,3415|false|false|false|C0202059|Bicarbonate measurement|HCO3
Finding|Body Substance|Hospital Course|3453,3460|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|3453,3460|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|3453,3460|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Hospital Course|3483,3490|false|false|false|||history
Finding|Conceptual Entity|Hospital Course|3483,3490|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|3483,3490|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Hospital Course|3483,3490|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|3483,3493|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|Hospital Course|3494,3497|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Hospital Course|3494,3497|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Hospital Course|3494,3497|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|Hospital Course|3494,3497|false|false|false|||CAD
Finding|Gene or Genome|Hospital Course|3494,3497|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Hospital Course|3494,3497|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Hospital Course|3494,3497|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3494,3497|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Disorder|Disease or Syndrome|Hospital Course|3503,3506|false|false|false|C0006430|Burning Mouth Syndrome|BMS
Event|Event|Hospital Course|3503,3506|false|false|false|||BMS
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|3541,3544|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|Hospital Course|3541,3544|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Finding|Gene or Genome|Hospital Course|3541,3544|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Disorder|Disease or Syndrome|Hospital Course|3550,3553|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|Hospital Course|3550,3553|false|false|false|||HTN
Disorder|Disease or Syndrome|Hospital Course|3555,3575|false|false|false|C0020443|Hypercholesterolemia|Hypercholesterolemia
Event|Event|Hospital Course|3555,3575|false|false|false|||Hypercholesterolemia
Finding|Finding|Hospital Course|3555,3575|false|false|false|C1522133|Hypercholesterolemia result|Hypercholesterolemia
Event|Event|Hospital Course|3581,3589|false|false|false|||presents
Finding|Finding|Hospital Course|3595,3603|false|false|false|C0741302|atypia morphology|atypical
Finding|Sign or Symptom|Hospital Course|3595,3614|false|false|false|C0262384|Atypical chest pain|atypical chest pain
Anatomy|Body Location or Region|Hospital Course|3604,3609|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Hospital Course|3604,3609|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Hospital Course|3604,3614|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|Hospital Course|3604,3614|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Hospital Course|3610,3614|false|false|false|C2598155||pain
Event|Event|Hospital Course|3610,3614|false|false|false|||pain
Finding|Functional Concept|Hospital Course|3610,3614|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|3610,3614|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Disorder|Disease or Syndrome|Hospital Course|3625,3628|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Hospital Course|3625,3628|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Hospital Course|3625,3628|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|Hospital Course|3625,3628|false|false|false|||CAD
Finding|Gene or Genome|Hospital Course|3625,3628|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Hospital Course|3625,3628|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Hospital Course|3625,3628|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3625,3628|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Disorder|Disease or Syndrome|Hospital Course|3641,3644|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Hospital Course|3641,3644|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Hospital Course|3641,3644|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|Hospital Course|3641,3644|false|false|false|||CAD
Finding|Gene or Genome|Hospital Course|3641,3644|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Hospital Course|3641,3644|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Hospital Course|3641,3644|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3641,3644|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Finding|Functional Concept|Hospital Course|3646,3663|false|false|false|C3853134|Poorly controlled|poorly controlled
Event|Event|Hospital Course|3653,3663|false|false|false|||controlled
Event|Event|Hospital Course|3668,3675|false|false|false|||episode
Event|Event|Hospital Course|3692,3701|false|false|false|||admission
Procedure|Health Care Activity|Hospital Course|3692,3701|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Attribute|Clinical Attribute|Hospital Course|3717,3723|false|false|false|C2926611||angina
Event|Event|Hospital Course|3717,3723|false|false|false|||angina
Finding|Finding|Hospital Course|3717,3723|false|false|false|C0002962;C2024883|Angina Pectoris|angina
Finding|Sign or Symptom|Hospital Course|3717,3723|false|false|false|C0002962;C2024883|Angina Pectoris|angina
Finding|Body Substance|Hospital Course|3726,3733|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|3726,3733|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|3726,3733|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Hospital Course|3736,3739|false|false|false|||EKG
Finding|Intellectual Product|Hospital Course|3736,3739|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|Hospital Course|3736,3739|false|false|false|C1623258|Electrocardiography|EKG
Event|Event|Hospital Course|3740,3746|false|false|false|||showed
Event|Event|Hospital Course|3755,3758|false|false|false|||AVL
Finding|Pathologic Function|Hospital Course|3755,3758|false|false|false|C5237386|Atypical Vascular Proliferation|AVL
Event|Event|Hospital Course|3767,3778|false|false|false|||nonspecific
Finding|Body Substance|Hospital Course|3780,3787|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|3780,3787|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|3780,3787|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Hospital Course|3788,3793|false|false|false|||ruled
Finding|Body Substance|Hospital Course|3808,3815|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|3808,3815|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|3808,3815|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Finding|Hospital Course|3830,3836|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Hospital Course|3830,3836|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|Hospital Course|3851,3857|false|false|false|||origin
Finding|Classification|Hospital Course|3851,3857|false|false|false|C0079946;C1550512|National origin;Participation Type - origin|origin
Finding|Intellectual Product|Hospital Course|3851,3857|false|false|false|C0079946;C1550512|National origin;Participation Type - origin|origin
Event|Event|Hospital Course|3879,3887|false|false|false|||episodes
Drug|Amino Acid, Peptide, or Protein|Hospital Course|3917,3921|false|false|false|C1742913|REST protein, human|rest
Drug|Biologically Active Substance|Hospital Course|3917,3921|false|false|false|C1742913|REST protein, human|rest
Event|Event|Hospital Course|3917,3921|false|false|false|||rest
Finding|Daily or Recreational Activity|Hospital Course|3917,3921|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Gene or Genome|Hospital Course|3917,3921|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Molecular Function|Hospital Course|3917,3921|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Event|Event|Hospital Course|3930,3938|false|false|false|||exertion
Finding|Organism Function|Hospital Course|3930,3938|false|false|false|C0015264|Exertion|exertion
Finding|Intellectual Product|Hospital Course|3952,3955|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|Hospital Course|3952,3955|false|false|false|C1623258|Electrocardiography|EKG
Event|Event|Hospital Course|3956,3963|false|false|false|||changes
Finding|Functional Concept|Hospital Course|3956,3963|false|false|false|C0392747|Changing|changes
Event|Event|Hospital Course|3968,3976|false|false|false|||negative
Finding|Classification|Hospital Course|3968,3976|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|3968,3976|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|3968,3976|false|false|false|C5237010|Expression Negative|negative
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|3977,3984|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|Hospital Course|3977,3984|false|false|false|C1314974|Cardiac attachment|cardiac
Attribute|Clinical Attribute|Hospital Course|3977,3992|false|false|false|C2926589||cardiac enzymes
Drug|Amino Acid, Peptide, or Protein|Hospital Course|3977,3992|false|false|false|C0443763|Cardiac enzymes|cardiac enzymes
Drug|Enzyme|Hospital Course|3977,3992|false|false|false|C0443763|Cardiac enzymes|cardiac enzymes
Procedure|Laboratory Procedure|Hospital Course|3977,3992|false|false|false|C0201934|Cardiac enzymes/isoenzymes measurement|cardiac enzymes
Drug|Amino Acid, Peptide, or Protein|Hospital Course|3985,3992|false|false|false|C0014442;C3540017;C3540048;C3540772;C3540790;C3541394;C3542456|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS;Enzymes;Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM;Enzymes for ALIMENTARY TRACT AND METABOLISM;Enzymes, antithrombotic;Enzymes, hematological;Enzymes, peripheral vasodilators|enzymes
Drug|Enzyme|Hospital Course|3985,3992|false|false|false|C0014442;C3540017;C3540048;C3540772;C3540790;C3541394;C3542456|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS;Enzymes;Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM;Enzymes for ALIMENTARY TRACT AND METABOLISM;Enzymes, antithrombotic;Enzymes, hematological;Enzymes, peripheral vasodilators|enzymes
Drug|Pharmacologic Substance|Hospital Course|3985,3992|false|false|false|C0014442;C3540017;C3540048;C3540772;C3540790;C3541394;C3542456|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS;Enzymes;Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM;Enzymes for ALIMENTARY TRACT AND METABOLISM;Enzymes, antithrombotic;Enzymes, hematological;Enzymes, peripheral vasodilators|enzymes
Event|Event|Hospital Course|3985,3992|false|false|false|||enzymes
Finding|Functional Concept|Hospital Course|3985,3992|false|false|false|C0014445|enzymology|enzymes
Finding|Body Substance|Hospital Course|3996,4003|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|3996,4003|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|3996,4003|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Attribute|Clinical Attribute|Hospital Course|4018,4024|false|false|false|C1718621|W stress|stress
Drug|Organic Chemical|Hospital Course|4018,4024|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|Hospital Course|4018,4024|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Event|Event|Hospital Course|4018,4024|false|false|false|||stress
Finding|Finding|Hospital Course|4018,4024|false|false|false|C0038435|Stress|stress
Event|Event|Hospital Course|4031,4040|true|false|false|||inpatient
Finding|Idea or Concept|Hospital Course|4031,4040|true|false|false|C1548438;C1549404|Patient Class - Inpatient;Referral category - Inpatient|inpatient
Procedure|Health Care Activity|Hospital Course|4031,4040|true|false|false|C1555324|inpatient encounter|inpatient
Event|Event|Hospital Course|4049,4057|true|false|false|||negative
Finding|Classification|Hospital Course|4049,4057|true|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|4049,4057|true|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|4049,4057|true|false|false|C5237010|Expression Negative|negative
Event|Event|Hospital Course|4067,4076|true|false|false|||perfusion
Finding|Functional Concept|Hospital Course|4067,4076|true|false|false|C4281794;C4723760|Perfusion (biological);Perfusion route|perfusion
Finding|Organism Function|Hospital Course|4067,4076|true|false|false|C4281794;C4723760|Perfusion (biological);Perfusion route|perfusion
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4067,4076|true|false|false|C0031001;C4721534|Chemotherapeutic Perfusion;Perfusion (procedure)|perfusion
Event|Event|Hospital Course|4077,4084|true|false|false|||defects
Finding|Functional Concept|Hospital Course|4077,4084|true|false|false|C0243067|defects aspect|defects
Event|Event|Hospital Course|4090,4098|false|false|false|||Continue
Finding|Idea or Concept|Hospital Course|4090,4098|false|false|false|C0549178|Continuous|Continue
Drug|Amino Acid, Peptide, or Protein|Hospital Course|4099,4102|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Enzyme|Hospital Course|4099,4102|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Organic Chemical|Hospital Course|4099,4102|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Pharmacologic Substance|Hospital Course|4099,4102|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Event|Event|Hospital Course|4099,4102|false|false|false|||ASA
Finding|Gene or Genome|Hospital Course|4099,4102|false|false|false|C1412553|ARSA gene|ASA
Drug|Organic Chemical|Hospital Course|4104,4110|false|false|false|C0633084|Plavix|Plavix
Drug|Pharmacologic Substance|Hospital Course|4104,4110|false|false|false|C0633084|Plavix|Plavix
Event|Event|Hospital Course|4104,4110|false|false|false|||Plavix
Drug|Amino Acid, Peptide, or Protein|Hospital Course|4123,4126|false|false|false|C1452534|ACE protein, human|ACE
Drug|Biologically Active Substance|Hospital Course|4123,4126|false|false|false|C1452534|ACE protein, human|ACE
Event|Event|Hospital Course|4123,4126|false|false|false|||ACE
Finding|Gene or Genome|Hospital Course|4123,4126|false|false|false|C1413931;C4284014|ACE gene;Adverse Childhood Experience questionnaire|ACE
Finding|Intellectual Product|Hospital Course|4123,4126|false|false|false|C1413931;C4284014|ACE gene;Adverse Childhood Experience questionnaire|ACE
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4123,4126|false|false|false|C0050385;C0108844;C0279078;C1879921|CDE Regimen;CDE protocol;cisplatin, cytarabine, and etoposide chemotherapy protocol;cyclophosphamide/doxorubicin protocol|ACE
Finding|Idea or Concept|Hospital Course|4135,4143|false|false|false|C0549178|Continuous|Continue
Drug|Organic Chemical|Hospital Course|4144,4150|false|false|false|C0360714|Hydroxymethylglutaryl-CoA Reductase Inhibitors|Statin
Drug|Pharmacologic Substance|Hospital Course|4144,4150|false|false|false|C0360714|Hydroxymethylglutaryl-CoA Reductase Inhibitors|Statin
Event|Event|Hospital Course|4144,4150|false|false|false|||Statin
Finding|Gene or Genome|Hospital Course|4144,4150|false|false|false|C1414273|EEF1A2 gene|Statin
Finding|Molecular Function|Hospital Course|4160,4164|false|false|false|C1150186|matrix metalloproteinase 7 activity|Pump
Event|Event|Hospital Course|4166,4175|false|false|false|||Euvolemic
Event|Event|Hospital Course|4179,4183|false|false|false|||exam
Finding|Functional Concept|Hospital Course|4179,4183|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|Hospital Course|4179,4183|false|false|false|C0582103|Medical Examination|exam
Finding|Finding|Hospital Course|4194,4200|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|Rhythm
Finding|Physiologic Function|Hospital Course|4194,4200|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|Rhythm
Event|Event|Hospital Course|4202,4205|false|false|false|||NSR
Finding|Molecular Function|Hospital Course|4202,4205|false|false|false|C1704493;C2700623|Neutral Sidebent Rotated|NSR
Finding|Pathologic Function|Hospital Course|4202,4205|false|false|false|C1704493;C2700623|Neutral Sidebent Rotated|NSR
Disorder|Disease or Syndrome|Hospital Course|4215,4218|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|Hospital Course|4215,4218|false|false|false|||HTN
Attribute|Clinical Attribute|Hospital Course|4220,4223|false|false|false|C0871470|Systolic Pressure|SBP
Drug|Amino Acid, Peptide, or Protein|Hospital Course|4220,4223|false|false|false|C0085805|Androgen Binding Protein|SBP
Drug|Biologically Active Substance|Hospital Course|4220,4223|false|false|false|C0085805|Androgen Binding Protein|SBP
Event|Event|Hospital Course|4220,4223|false|false|false|||SBP
Finding|Gene or Genome|Hospital Course|4220,4223|false|false|false|C1705296;C3274833|CCHCR1 wt Allele;SHBG wt Allele|SBP
Procedure|Diagnostic Procedure|Hospital Course|4220,4223|false|false|false|C1306620|Systolic blood pressure measurement|SBP
Event|Event|Hospital Course|4236,4245|false|false|false|||discharge
Finding|Body Substance|Hospital Course|4236,4245|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|4236,4245|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|4236,4245|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|4236,4245|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|Hospital Course|4248,4255|false|false|false|||Concern
Finding|Idea or Concept|Hospital Course|4248,4255|false|false|false|C2699424|Concern|Concern
Finding|Body Substance|Hospital Course|4261,4268|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|4261,4268|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|4261,4268|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|4281,4290|false|false|false|||compliant
Finding|Individual Behavior|Hospital Course|4281,4290|false|false|false|C1321605|Compliance behavior|compliant
Drug|Pharmacologic Substance|Hospital Course|4296,4306|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Hospital Course|4296,4306|false|false|false|||medication
Finding|Intellectual Product|Hospital Course|4296,4306|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4296,4314|false|false|false|C0237125|Medication Regimen|medication regimen
Event|Event|Hospital Course|4307,4314|false|false|false|||regimen
Finding|Intellectual Product|Hospital Course|4307,4314|false|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4307,4314|false|false|false|C0040808|Treatment Protocols|regimen
Finding|Body Substance|Hospital Course|4317,4324|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|4317,4324|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|4317,4324|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Hospital Course|4329,4336|false|false|false|||dropped
Attribute|Clinical Attribute|Hospital Course|4337,4340|false|false|false|C0871470|Systolic Pressure|SBP
Drug|Amino Acid, Peptide, or Protein|Hospital Course|4337,4340|false|false|false|C0085805|Androgen Binding Protein|SBP
Drug|Biologically Active Substance|Hospital Course|4337,4340|false|false|false|C0085805|Androgen Binding Protein|SBP
Event|Event|Hospital Course|4337,4340|false|false|false|||SBP
Finding|Gene or Genome|Hospital Course|4337,4340|false|false|false|C1705296;C3274833|CCHCR1 wt Allele;SHBG wt Allele|SBP
Procedure|Diagnostic Procedure|Hospital Course|4337,4340|false|false|false|C1306620|Systolic blood pressure measurement|SBP
Event|Event|Hospital Course|4354,4363|false|false|false|||admission
Procedure|Health Care Activity|Hospital Course|4354,4363|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Idea or Concept|Hospital Course|4369,4373|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|4369,4373|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|4369,4373|false|false|false|C1553498|home health encounter|home
Attribute|Clinical Attribute|Hospital Course|4374,4385|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Hospital Course|4374,4385|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Hospital Course|4374,4385|false|false|false|||medications
Finding|Intellectual Product|Hospital Course|4374,4385|false|false|false|C4284232|Medications|medications
Event|Event|Hospital Course|4391,4403|false|false|false|||administered
Drug|Organic Chemical|Hospital Course|4426,4431|false|false|false|C0590690|Imdur|Imdur
Drug|Pharmacologic Substance|Hospital Course|4426,4431|false|false|false|C0590690|Imdur|Imdur
Event|Event|Hospital Course|4442,4451|false|false|false|||decreased
Anatomy|Body Space or Junction|Hospital Course|4453,4457|false|false|false|C0228216|Structure of subparietal sulcus|SBPs
Event|Event|Hospital Course|4469,4479|false|false|false|||controlled
Event|Event|Hospital Course|4489,4493|false|false|false|||need
Finding|Classification|Hospital Course|4494,4504|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|4494,4504|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|Hospital Course|4505,4514|false|false|false|||titration
Procedure|Laboratory Procedure|Hospital Course|4505,4514|false|false|false|C0162621|Titration Method|titration
Event|Event|Hospital Course|4520,4528|false|false|false|||Continue
Disorder|Disease or Syndrome|Hospital Course|4532,4536|false|false|false|C3280240|MICROCEPHALY, EPILEPSY, AND DIABETES SYNDROME 1|meds
Event|Event|Hospital Course|4532,4536|false|false|false|||meds
Finding|Intellectual Product|Hospital Course|4532,4536|false|false|false|C4284232|Medications|meds
Event|Event|Hospital Course|4543,4544|false|false|false|||#
Drug|Amino Acid, Peptide, or Protein|Hospital Course|4551,4556|false|false|false|C0019018|Glycosylated hemoglobin A|HbA1c
Drug|Biologically Active Substance|Hospital Course|4551,4556|false|false|false|C0019018|Glycosylated hemoglobin A|HbA1c
Event|Event|Hospital Course|4551,4556|false|false|false|||HbA1c
Procedure|Laboratory Procedure|Hospital Course|4551,4556|false|false|false|C0202054|Glucohemoglobin measurement|HbA1c
Finding|Functional Concept|Hospital Course|4570,4587|false|false|false|C3853134|Poorly controlled|Poorly controlled
Event|Event|Hospital Course|4577,4587|false|false|false|||controlled
Drug|Amino Acid, Peptide, or Protein|Hospital Course|4603,4610|false|false|false|C1314782|Levemir|Levemir
Drug|Hormone|Hospital Course|4603,4610|false|false|false|C1314782|Levemir|Levemir
Drug|Pharmacologic Substance|Hospital Course|4603,4610|false|false|false|C1314782|Levemir|Levemir
Drug|Organic Chemical|Hospital Course|4641,4650|false|false|false|C0025598|metformin|Metformin
Drug|Pharmacologic Substance|Hospital Course|4641,4650|false|false|false|C0025598|metformin|Metformin
Event|Event|Hospital Course|4677,4686|true|false|false|||compliant
Finding|Individual Behavior|Hospital Course|4677,4686|true|false|false|C1321605|Compliance behavior|compliant
Finding|Idea or Concept|Hospital Course|4702,4710|false|false|false|C0549178|Continuous|Continue
Drug|Organic Chemical|Hospital Course|4711,4720|false|false|false|C0025598|metformin|metformin
Drug|Pharmacologic Substance|Hospital Course|4711,4720|false|false|false|C0025598|metformin|metformin
Event|Event|Hospital Course|4711,4720|false|false|false|||metformin
Event|Event|Hospital Course|4725,4733|false|false|false|||Continue
Finding|Idea or Concept|Hospital Course|4725,4733|false|false|false|C0549178|Continuous|Continue
Drug|Amino Acid, Peptide, or Protein|Hospital Course|4734,4740|false|false|false|C0876064|Lantus|Lantus
Drug|Pharmacologic Substance|Hospital Course|4734,4740|false|false|false|C0876064|Lantus|Lantus
Event|Event|Hospital Course|4734,4740|false|false|false|||Lantus
Disorder|Disease or Syndrome|Hospital Course|4766,4780|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|hyperlipidemia
Event|Event|Hospital Course|4766,4780|false|false|false|||hyperlipidemia
Finding|Finding|Hospital Course|4766,4780|false|false|false|C0428465|Serum lipids high (finding)|hyperlipidemia
Event|Event|Hospital Course|4783,4791|false|false|false|||Continue
Finding|Idea or Concept|Hospital Course|4783,4791|false|false|false|C0549178|Continuous|Continue
Drug|Organic Chemical|Hospital Course|4792,4799|false|false|false|C0593906|Lipitor|Lipitor
Drug|Pharmacologic Substance|Hospital Course|4792,4799|false|false|false|C0593906|Lipitor|Lipitor
Attribute|Clinical Attribute|Hospital Course|4817,4828|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|4817,4828|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|4817,4828|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|4817,4828|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|4817,4841|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|Hospital Course|4832,4841|false|false|false|||Admission
Procedure|Health Care Activity|Hospital Course|4832,4841|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Organic Chemical|Hospital Course|4843,4849|false|false|false|C0965130|Advair|Advair
Drug|Pharmacologic Substance|Hospital Course|4843,4849|false|false|false|C0965130|Advair|Advair
Drug|Organic Chemical|Hospital Course|4865,4874|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|Hospital Course|4865,4874|false|false|false|C0001927|albuterol|Albuterol
Drug|Biomedical or Dental Material|Hospital Course|4875,4882|false|false|false|C1112870|Aerosol Dose Form|Aerosol
Finding|Gene or Genome|Hospital Course|4883,4886|false|false|false|C1422467|CIAO3 gene|prn
Drug|Amino Acid, Peptide, or Protein|Hospital Course|4889,4892|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Enzyme|Hospital Course|4889,4892|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Organic Chemical|Hospital Course|4889,4892|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Pharmacologic Substance|Hospital Course|4889,4892|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Event|Event|Hospital Course|4889,4892|false|false|false|||ASA
Finding|Gene or Genome|Hospital Course|4889,4892|false|false|false|C1412553|ARSA gene|ASA
Drug|Organic Chemical|Hospital Course|4907,4915|false|false|false|C0004147|atenolol|Atenolol
Drug|Pharmacologic Substance|Hospital Course|4907,4915|false|false|false|C0004147|atenolol|Atenolol
Drug|Amino Acid, Peptide, or Protein|Hospital Course|4929,4936|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Hormone|Hospital Course|4929,4936|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Pharmacologic Substance|Hospital Course|4929,4936|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Event|Event|Hospital Course|4929,4936|false|false|false|||Insulin
Finding|Gene or Genome|Hospital Course|4929,4936|false|false|false|C1337112|INS gene|Insulin
Procedure|Laboratory Procedure|Hospital Course|4929,4936|false|false|false|C0202098|Insulin measurement|Insulin
Drug|Organic Chemical|Hospital Course|4974,4984|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Pharmacologic Substance|Hospital Course|4974,4984|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Organic Chemical|Hospital Course|4974,4996|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Drug|Pharmacologic Substance|Hospital Course|4974,4996|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Event|Event|Hospital Course|4997,5002|false|false|false|||120mg
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5011,5021|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Pharmacologic Substance|Hospital Course|5011,5021|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Organic Chemical|Hospital Course|5035,5044|false|false|false|C0025598|metformin|Metformin
Drug|Pharmacologic Substance|Hospital Course|5035,5044|false|false|false|C0025598|metformin|Metformin
Drug|Organic Chemical|Hospital Course|5059,5072|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Drug|Pharmacologic Substance|Hospital Course|5059,5072|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Drug|Organic Chemical|Hospital Course|5078,5088|false|false|false|C0028978|omeprazole|Omeprazole
Drug|Pharmacologic Substance|Hospital Course|5078,5088|false|false|false|C0028978|omeprazole|Omeprazole
Drug|Organic Chemical|Hospital Course|5103,5109|false|false|false|C0633084|Plavix|Plavix
Drug|Pharmacologic Substance|Hospital Course|5103,5109|false|false|false|C0633084|Plavix|Plavix
Drug|Biologically Active Substance|Hospital Course|5125,5134|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Element, Ion, or Isotope|Hospital Course|5125,5134|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Food|Hospital Course|5125,5134|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Inorganic Chemical|Hospital Course|5125,5134|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Pharmacologic Substance|Hospital Course|5125,5134|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Event|Event|Hospital Course|5125,5134|false|false|false|||Potassium
Finding|Physiologic Function|Hospital Course|5125,5134|false|false|false|C4553027|Potassium metabolic function|Potassium
Procedure|Laboratory Procedure|Hospital Course|5125,5134|false|false|false|C0202194|Potassium measurement|Potassium
Drug|Inorganic Chemical|Hospital Course|5125,5143|false|false|false|C0032825|potassium chloride|Potassium chloride
Drug|Pharmacologic Substance|Hospital Course|5125,5143|false|false|false|C0032825|potassium chloride|Potassium chloride
Drug|Element, Ion, or Isotope|Hospital Course|5135,5143|false|false|false|C0008203;C0596019|Chlorides;chloride ion|chloride
Event|Event|Hospital Course|5135,5143|false|false|false|||chloride
Finding|Physiologic Function|Hospital Course|5135,5143|false|false|false|C4553021|Chloride metabolic function|chloride
Procedure|Laboratory Procedure|Hospital Course|5135,5143|false|false|false|C0201952|Chloride measurement|chloride
Event|Event|Hospital Course|5147,5150|false|false|false|||mEq
Drug|Organic Chemical|Hospital Course|5153,5164|false|false|false|C0074554|simvastatin|Simvastatin
Drug|Pharmacologic Substance|Hospital Course|5153,5164|false|false|false|C0074554|simvastatin|Simvastatin
Event|Event|Hospital Course|5176,5185|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|5176,5185|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|5176,5185|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|5176,5185|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|5176,5185|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|5176,5197|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|5186,5197|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|5186,5197|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|5186,5197|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|5186,5197|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Hospital Course|5202,5213|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Hospital Course|5202,5213|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Hospital Course|5202,5224|false|false|false|C0939232|fluticasone / salmeterol|Fluticasone-Salmeterol
Drug|Organic Chemical|Hospital Course|5214,5224|false|false|false|C0073992|salmeterol|Salmeterol
Drug|Pharmacologic Substance|Hospital Course|5214,5224|false|false|false|C0073992|salmeterol|Salmeterol
Event|Event|Hospital Course|5214,5224|false|false|false|||Salmeterol
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5241,5245|false|false|false|C1556138|Disc - Body Part|Disk
Drug|Biomedical or Dental Material|Hospital Course|5241,5245|false|false|false|C0993608|Disk Drug Form|Disk
Finding|Functional Concept|Hospital Course|5251,5257|false|false|false|C1550509|Participation Type - device|Device
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5258,5261|false|false|false|C0262329|Short insular gyrus|Sig
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5258,5261|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Drug|Immunologic Factor|Hospital Course|5258,5261|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Finding|Receptor|Hospital Course|5258,5261|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5272,5276|false|false|false|C1556138|Disc - Body Part|Disk
Drug|Biomedical or Dental Material|Hospital Course|5272,5276|false|false|false|C0993608|Disk Drug Form|Disk
Finding|Functional Concept|Hospital Course|5282,5288|false|false|false|C1550509|Participation Type - device|Device
Event|Event|Hospital Course|5289,5299|false|false|false|||Inhalation
Finding|Functional Concept|Hospital Course|5289,5299|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Finding|Organism Function|Hospital Course|5289,5299|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Disorder|Mental or Behavioral Dysfunction|Hospital Course|5300,5303|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5300,5303|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|5300,5303|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|5300,5303|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|5300,5303|false|false|false|C1332410|BID gene|BID
Finding|Finding|Hospital Course|5305,5312|false|false|false|C4035627|2 times|2 times
Disorder|Disease or Syndrome|Hospital Course|5307,5312|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|Hospital Course|5315,5318|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|5315,5318|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|Hospital Course|5326,5333|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|Hospital Course|5326,5333|false|false|false|C0004057|aspirin|Aspirin
Drug|Biomedical or Dental Material|Hospital Course|5341,5347|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|5361,5367|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|5361,5367|false|false|false|||Tablet
Drug|Organic Chemical|Hospital Course|5391,5400|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|Hospital Course|5391,5400|false|false|false|C0001927|albuterol|Albuterol
Event|Event|Hospital Course|5391,5400|false|false|false|||Albuterol
Drug|Biomedical or Dental Material|Hospital Course|5418,5425|false|false|false|C1112870|Aerosol Dose Form|Aerosol
Event|Event|Hospital Course|5426,5429|false|false|false|||Sig
Event|Event|Hospital Course|5441,5451|false|false|false|||Inhalation
Finding|Functional Concept|Hospital Course|5441,5451|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Finding|Organism Function|Hospital Course|5441,5451|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Event|Event|Hospital Course|5476,5482|false|false|false|||needed
Drug|Organic Chemical|Hospital Course|5489,5500|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Pharmacologic Substance|Hospital Course|5489,5500|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Biomedical or Dental Material|Hospital Course|5507,5513|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|5527,5533|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|5527,5533|false|false|false|||Tablet
Drug|Organic Chemical|Hospital Course|5558,5569|false|false|false|C0074554|simvastatin|Simvastatin
Drug|Pharmacologic Substance|Hospital Course|5558,5569|false|false|false|C0074554|simvastatin|Simvastatin
Drug|Biomedical or Dental Material|Hospital Course|5576,5582|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|5596,5602|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|5603,5605|false|false|false|||PO
Drug|Organic Chemical|Hospital Course|5627,5637|false|false|false|C0028978|omeprazole|Omeprazole
Drug|Pharmacologic Substance|Hospital Course|5627,5637|false|false|false|C0028978|omeprazole|Omeprazole
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5644,5651|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|5644,5651|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|5644,5651|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Attribute|Clinical Attribute|Hospital Course|5653,5660|false|false|false|C1545665|Views delayed|Delayed
Drug|Biomedical or Dental Material|Hospital Course|5653,5668|false|false|false|C1707664|Delayed Release Dosage Form|Delayed Release
Event|Event|Hospital Course|5661,5668|false|false|false|||Release
Finding|Functional Concept|Hospital Course|5661,5668|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|5661,5668|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5661,5668|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Event|Event|Hospital Course|5675,5678|false|false|false|||Sig
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5689,5696|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|5689,5696|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|5689,5696|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Attribute|Clinical Attribute|Hospital Course|5698,5705|false|false|false|C1545665|Views delayed|Delayed
Drug|Biomedical or Dental Material|Hospital Course|5698,5713|false|false|false|C1707664|Delayed Release Dosage Form|Delayed Release
Event|Event|Hospital Course|5706,5713|false|false|false|||Release
Finding|Functional Concept|Hospital Course|5706,5713|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|5706,5713|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5706,5713|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|Hospital Course|5743,5752|false|false|false|C0030049|oxycodone|Oxycodone
Drug|Pharmacologic Substance|Hospital Course|5743,5752|false|false|false|C0030049|oxycodone|Oxycodone
Event|Event|Hospital Course|5743,5752|false|false|false|||Oxycodone
Procedure|Laboratory Procedure|Hospital Course|5743,5752|false|false|false|C0524222|Oxycodone measurement|Oxycodone
Drug|Pharmacologic Substance|Hospital Course|5743,5766|false|false|false|C0717368|acetaminophen / oxycodone|Oxycodone-Acetaminophen
Drug|Organic Chemical|Hospital Course|5753,5766|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Hospital Course|5753,5766|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|Hospital Course|5753,5766|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|Hospital Course|5753,5766|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Drug|Biomedical or Dental Material|Hospital Course|5774,5780|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|5790,5797|false|false|false|C0039225|Tablet Dosage Form|Tablets
Event|Event|Hospital Course|5790,5797|false|false|false|||Tablets
Event|Event|Hospital Course|5825,5831|false|false|false|||needed
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5838,5845|false|false|false|C1314782|Levemir|Levemir
Drug|Hormone|Hospital Course|5838,5845|false|false|false|C1314782|Levemir|Levemir
Drug|Pharmacologic Substance|Hospital Course|5838,5845|false|false|false|C1314782|Levemir|Levemir
Drug|Biomedical or Dental Material|Hospital Course|5858,5866|false|false|false|C0037633;C0525069;C1382100|Pharmaceutical Solutions;Solution Dosage Form;Solutions|Solution
Drug|Substance|Hospital Course|5858,5866|false|false|false|C0037633;C0525069;C1382100|Pharmaceutical Solutions;Solution Dosage Form;Solutions|Solution
Event|Event|Hospital Course|5858,5866|false|false|false|||Solution
Finding|Conceptual Entity|Hospital Course|5858,5866|false|false|false|C2699488|Resolution|Solution
Event|Event|Hospital Course|5867,5870|false|false|false|||Sig
Finding|Functional Concept|Hospital Course|5881,5893|false|false|false|C1522438|Subcutaneous Route of Administration|Subcutaneous
Finding|Idea or Concept|Hospital Course|5903,5906|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|5903,5906|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Hospital Course|5916,5919|false|false|false|||qAM
Drug|Organic Chemical|Hospital Course|5934,5943|false|false|false|C0025598|metformin|Metformin
Drug|Pharmacologic Substance|Hospital Course|5934,5943|false|false|false|C0025598|metformin|Metformin
Drug|Biomedical or Dental Material|Hospital Course|5951,5957|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|5971,5977|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|5971,5977|false|false|false|||Tablet
Disorder|Disease or Syndrome|Hospital Course|5987,5992|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|Hospital Course|5996,5999|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|5996,5999|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Biologically Active Substance|Hospital Course|6007,6016|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Element, Ion, or Isotope|Hospital Course|6007,6016|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Food|Hospital Course|6007,6016|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Inorganic Chemical|Hospital Course|6007,6016|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Pharmacologic Substance|Hospital Course|6007,6016|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Event|Event|Hospital Course|6007,6016|false|false|false|||Potassium
Finding|Physiologic Function|Hospital Course|6007,6016|false|false|false|C4553027|Potassium metabolic function|Potassium
Procedure|Laboratory Procedure|Hospital Course|6007,6016|false|false|false|C0202194|Potassium measurement|Potassium
Drug|Inorganic Chemical|Hospital Course|6007,6025|false|false|false|C0032825|potassium chloride|Potassium Chloride
Drug|Pharmacologic Substance|Hospital Course|6007,6025|false|false|false|C0032825|potassium chloride|Potassium Chloride
Drug|Element, Ion, or Isotope|Hospital Course|6017,6025|false|false|false|C0008203;C0596019|Chlorides;chloride ion|Chloride
Event|Event|Hospital Course|6017,6025|false|false|false|||Chloride
Finding|Physiologic Function|Hospital Course|6017,6025|false|false|false|C4553021|Chloride metabolic function|Chloride
Procedure|Laboratory Procedure|Hospital Course|6017,6025|false|false|false|C0201952|Chloride measurement|Chloride
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6033,6040|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|6033,6040|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|6033,6040|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Finding|Functional Concept|Hospital Course|6042,6051|false|false|false|C0443318|Sustained|Sustained
Drug|Biomedical or Dental Material|Hospital Course|6042,6059|false|false|false|C1710261|Sustained Release Dosage Form|Sustained Release
Event|Event|Hospital Course|6052,6059|false|false|false|||Release
Finding|Functional Concept|Hospital Course|6052,6059|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|6052,6059|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6052,6059|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6074,6081|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|6074,6081|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|6074,6081|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Event|Event|Hospital Course|6093,6100|false|false|false|||Release
Finding|Functional Concept|Hospital Course|6093,6100|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|6093,6100|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6093,6100|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Finding|Intellectual Product|Hospital Course|6104,6108|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|Hospital Course|6104,6114|false|false|false|C3537736|Once A Day|once a day
Finding|Idea or Concept|Hospital Course|6111,6114|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|6111,6114|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|Hospital Course|6122,6135|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Drug|Pharmacologic Substance|Hospital Course|6122,6135|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Drug|Biomedical or Dental Material|Hospital Course|6143,6149|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|6143,6149|false|false|false|||Tablet
Drug|Biomedical or Dental Material|Hospital Course|6143,6161|false|false|false|C0991582|Sublingual Tablet|Tablet, Sublingual
Finding|Finding|Hospital Course|6151,6161|false|false|false|C0001565;C4521982|Sublingual (intended site);Sublingual Route of Administration|Sublingual
Finding|Functional Concept|Hospital Course|6151,6161|false|false|false|C0001565;C4521982|Sublingual (intended site);Sublingual Route of Administration|Sublingual
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6162,6165|false|false|false|C0262329|Short insular gyrus|Sig
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6162,6165|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Drug|Immunologic Factor|Hospital Course|6162,6165|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Finding|Receptor|Hospital Course|6162,6165|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Drug|Biomedical or Dental Material|Hospital Course|6175,6181|false|false|false|C0039225|Tablet Dosage Form|tablet
Event|Event|Hospital Course|6175,6181|false|false|false|||tablet
Finding|Finding|Hospital Course|6183,6193|false|false|false|C0001565;C4521982|Sublingual (intended site);Sublingual Route of Administration|Sublingual
Finding|Functional Concept|Hospital Course|6183,6193|false|false|false|C0001565;C4521982|Sublingual (intended site);Sublingual Route of Administration|Sublingual
Event|Event|Hospital Course|6203,6209|false|false|false|||needed
Anatomy|Body Location or Region|Hospital Course|6214,6219|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Hospital Course|6214,6219|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Hospital Course|6214,6224|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|Hospital Course|6214,6224|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Hospital Course|6220,6224|false|false|false|C2598155||pain
Event|Event|Hospital Course|6220,6224|false|false|false|||pain
Finding|Functional Concept|Hospital Course|6220,6224|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|6220,6224|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|6226,6229|false|false|false|||Sit
Finding|Finding|Hospital Course|6226,6229|false|false|false|C0277814;C0728713;C1539668;C1539774|Does sit;HHAT gene;SIT1 gene;Sitting position|Sit
Finding|Gene or Genome|Hospital Course|6226,6229|false|false|false|C0277814;C0728713;C1539668;C1539774|Does sit;HHAT gene;SIT1 gene;Sitting position|Sit
Event|Event|Hospital Course|6245,6251|false|false|false|||taking
Event|Event|Hospital Course|6253,6257|false|false|false|||Take
Drug|Biomedical or Dental Material|Hospital Course|6262,6265|false|false|false|C0039225|Tablet Dosage Form|tab
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6272,6281|false|false|false|C0886384|5 minutes Office visit|5 minutes
Event|Event|Hospital Course|6274,6281|false|false|false|||minutes
Anatomy|Body Location or Region|Hospital Course|6288,6293|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Hospital Course|6288,6293|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Hospital Course|6288,6298|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|Hospital Course|6288,6298|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Hospital Course|6294,6298|false|false|false|C2598155||pain
Event|Event|Hospital Course|6294,6298|false|false|false|||pain
Finding|Functional Concept|Hospital Course|6294,6298|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|6294,6298|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|6299,6307|false|false|false|||resolves
Attribute|Clinical Attribute|Hospital Course|6313,6317|true|false|false|C2598155||pain
Event|Event|Hospital Course|6313,6317|true|false|false|||pain
Finding|Functional Concept|Hospital Course|6313,6317|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|6313,6317|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|6322,6330|true|false|false|||resolved
Event|Event|Hospital Course|6339,6343|true|false|false|||call
Drug|Hazardous or Poisonous Substance|Hospital Course|6344,6347|true|false|false|C0015063|Ethyl Methanesulfonate|EMS
Drug|Organic Chemical|Hospital Course|6344,6347|true|false|false|C0015063|Ethyl Methanesulfonate|EMS
Drug|Pharmacologic Substance|Hospital Course|6344,6347|true|false|false|C0015063|Ethyl Methanesulfonate|EMS
Event|Event|Hospital Course|6344,6347|true|false|false|||EMS
Finding|Gene or Genome|Hospital Course|6344,6347|true|false|false|C5203240|EMSLR gene|EMS
Procedure|Health Care Activity|Hospital Course|6344,6347|true|false|false|C0013961|Emergency Medical Services|EMS
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6355,6365|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Pharmacologic Substance|Hospital Course|6355,6365|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Biomedical or Dental Material|Hospital Course|6371,6377|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|6391,6397|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|6391,6397|false|false|false|||Tablet
Drug|Biomedical or Dental Material|Hospital Course|6425,6431|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|6436,6443|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|6436,6443|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|6452,6462|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|Hospital Course|6452,6462|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Organic Chemical|Hospital Course|6452,6471|false|false|false|C0700548|metoprolol tartrate|Metoprolol Tartrate
Drug|Pharmacologic Substance|Hospital Course|6452,6471|false|false|false|C0700548|metoprolol tartrate|Metoprolol Tartrate
Drug|Organic Chemical|Hospital Course|6463,6471|false|false|false|C0039328;C0144544|Tartrates;tartrate|Tartrate
Drug|Pharmacologic Substance|Hospital Course|6463,6471|false|false|false|C0039328;C0144544|Tartrates;tartrate|Tartrate
Event|Event|Hospital Course|6463,6471|false|false|false|||Tartrate
Drug|Biomedical or Dental Material|Hospital Course|6478,6484|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|6494,6501|false|false|false|C0039225|Tablet Dosage Form|Tablets
Disorder|Mental or Behavioral Dysfunction|Hospital Course|6505,6508|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6505,6508|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|6505,6508|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|6505,6508|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|6505,6508|false|false|false|C1332410|BID gene|BID
Disorder|Disease or Syndrome|Hospital Course|6513,6518|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|Hospital Course|6521,6524|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|6521,6524|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Biomedical or Dental Material|Hospital Course|6536,6542|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|6547,6554|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|6547,6554|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|6563,6573|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Pharmacologic Substance|Hospital Course|6563,6573|false|false|false|C0022251|isosorbide|Isosorbide
Event|Event|Hospital Course|6563,6573|false|false|false|||Isosorbide
Drug|Organic Chemical|Hospital Course|6563,6585|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Drug|Pharmacologic Substance|Hospital Course|6563,6585|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Event|Event|Hospital Course|6574,6585|false|false|false|||Mononitrate
Drug|Biomedical or Dental Material|Hospital Course|6592,6598|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|6609,6616|false|false|false|||Release
Finding|Functional Concept|Hospital Course|6609,6616|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|6609,6616|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6609,6616|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Event|Event|Hospital Course|6624,6627|false|false|false|||Sig
Drug|Biomedical or Dental Material|Hospital Course|6637,6643|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|6637,6643|false|false|false|||Tablet
Event|Event|Hospital Course|6654,6661|false|false|false|||Release
Finding|Functional Concept|Hospital Course|6654,6661|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|6654,6661|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6654,6661|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Biomedical or Dental Material|Hospital Course|6695,6701|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|6712,6719|false|false|false|||Release
Finding|Functional Concept|Hospital Course|6712,6719|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|6712,6719|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6712,6719|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Finding|Idea or Concept|Hospital Course|6730,6737|false|false|false|C0807726|refill|Refills
Event|Event|Hospital Course|6745,6754|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|6745,6754|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|6745,6754|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|6745,6754|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|6745,6754|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|6745,6766|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|6745,6766|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|6755,6766|false|false|false|C2926604||Disposition
Event|Event|Hospital Course|6755,6766|false|false|false|||Disposition
Procedure|Health Care Activity|Hospital Course|6755,6766|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|Hospital Course|6768,6772|false|false|false|||Home
Finding|Idea or Concept|Hospital Course|6768,6772|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|6768,6772|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|6768,6772|false|false|false|C1553498|home health encounter|Home
Event|Event|Hospital Course|6775,6784|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|6775,6784|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|6775,6784|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|6775,6784|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|6775,6784|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|6775,6794|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|6785,6794|false|false|false|C0945731||Diagnosis
Event|Event|Hospital Course|6785,6794|false|false|false|||Diagnosis
Finding|Classification|Hospital Course|6785,6794|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|6785,6794|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|6785,6794|false|false|false|C0011900|Diagnosis|Diagnosis
Finding|Finding|Hospital Course|6806,6814|false|false|false|C0741302|atypia morphology|Atypical
Finding|Sign or Symptom|Hospital Course|6806,6825|false|false|false|C0262384|Atypical chest pain|Atypical Chest pain
Anatomy|Body Location or Region|Hospital Course|6815,6820|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|Hospital Course|6815,6820|false|false|false|C0741025|Chest problem|Chest
Attribute|Clinical Attribute|Hospital Course|6815,6825|false|false|false|C2926613||Chest pain
Finding|Sign or Symptom|Hospital Course|6815,6825|false|false|false|C0008031|Chest Pain|Chest pain
Attribute|Clinical Attribute|Hospital Course|6821,6825|false|true|false|C2598155||pain
Event|Event|Hospital Course|6821,6825|false|false|false|||pain
Finding|Functional Concept|Hospital Course|6821,6825|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|6821,6825|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6828,6836|false|false|false|C0018787|Heart|Coronary
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6828,6843|false|false|false|C0205042|Coronary artery|Coronary artery
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6837,6843|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|Hospital Course|6837,6843|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Event|Event|Hospital Course|6844,6850|false|false|false|||disase
Disorder|Neoplastic Process|Hospital Course|6851,6860|false|false|false|C0027627|Neoplasm Metastasis|Secondary
Event|Event|Hospital Course|6851,6860|false|false|false|||Secondary
Finding|Functional Concept|Hospital Course|6851,6860|false|false|false|C1522484|metastatic qualifier|Secondary
Disorder|Disease or Syndrome|Hospital Course|6863,6875|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|Hospital Course|6863,6875|false|false|false|||Hypertension
Disorder|Disease or Syndrome|Hospital Course|6878,6886|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|Diabetes
Event|Event|Hospital Course|6878,6886|false|false|false|||Diabetes
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6888,6895|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|Hospital Course|6888,6895|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|Hospital Course|6888,6895|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|Hospital Course|6888,6895|false|false|false|||insulin
Finding|Gene or Genome|Hospital Course|6888,6895|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|Hospital Course|6888,6895|false|false|false|C0202098|Insulin measurement|insulin
Event|Event|Hospital Course|6896,6905|false|false|false|||dependent
Finding|Functional Concept|Hospital Course|6896,6905|false|false|false|C3244310|dependent|dependent
Event|Event|Discharge Condition|6930,6938|false|false|false|||Afebrile
Finding|Finding|Discharge Condition|6930,6938|false|false|false|C0277797|Apyrexial|Afebrile
Anatomy|Body Location or Region|Discharge Condition|6940,6945|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|Discharge Condition|6940,6945|false|false|false|C0741025|Chest problem|Chest
Attribute|Clinical Attribute|Discharge Condition|6940,6950|false|false|false|C2926613||Chest pain
Finding|Sign or Symptom|Discharge Condition|6940,6950|false|false|false|C0008031|Chest Pain|Chest pain
Attribute|Clinical Attribute|Discharge Condition|6946,6950|false|false|false|C2598155||pain
Event|Event|Discharge Condition|6946,6950|false|false|false|||pain
Finding|Functional Concept|Discharge Condition|6946,6950|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Condition|6946,6950|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|Discharge Condition|6946,6955|false|false|false|C0908489|Pain-Free|pain free
Event|Event|Discharge Condition|6951,6955|false|false|false|||free
Finding|Functional Concept|Discharge Condition|6951,6955|false|false|false|C0332296|Free of (attribute)|free
Event|Event|Discharge Condition|6957,6963|false|false|false|||stable
Finding|Intellectual Product|Discharge Condition|6957,6963|false|false|false|C1547311|Patient Condition Code - Stable|stable
Event|Event|Discharge Instructions|7003,7015|false|false|false|||hospitalized
Anatomy|Body Location or Region|Discharge Instructions|7032,7037|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Discharge Instructions|7032,7037|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Discharge Instructions|7032,7042|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|Discharge Instructions|7032,7042|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Discharge Instructions|7038,7042|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|7038,7042|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|7038,7042|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|7038,7042|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|7065,7070|true|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Discharge Instructions|7065,7070|true|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Discharge Instructions|7065,7070|true|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|Discharge Instructions|7065,7077|true|false|false|C0027051|Myocardial Infarction|heart attack
Event|Event|Discharge Instructions|7071,7077|true|false|false|||attack
Finding|Finding|Discharge Instructions|7071,7077|true|false|false|C1261512;C1304680|Attack (finding);Attack behavior|attack
Finding|Social Behavior|Discharge Instructions|7071,7077|true|false|false|C1261512;C1304680|Attack (finding);Attack behavior|attack
Anatomy|Body Location or Region|Discharge Instructions|7085,7090|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Discharge Instructions|7085,7090|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Discharge Instructions|7085,7095|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|Discharge Instructions|7085,7095|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Discharge Instructions|7091,7095|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|7091,7095|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|7091,7095|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|7091,7095|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Discharge Instructions|7096,7104|false|false|false|||resolved
Disorder|Disease or Syndrome|Discharge Instructions|7112,7117|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Discharge Instructions|7112,7117|false|false|false|||blood
Finding|Body Substance|Discharge Instructions|7112,7117|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Event|Event|Discharge Instructions|7119,7127|false|false|false|||pressure
Finding|Finding|Discharge Instructions|7119,7127|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|Discharge Instructions|7119,7127|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|Discharge Instructions|7119,7127|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|Discharge Instructions|7119,7127|false|false|false|C0033095||pressure
Finding|Finding|Discharge Instructions|7132,7140|false|false|false|C2984078;C3889124|A little bit;Only a Little|a little
Disorder|Disease or Syndrome|Discharge Instructions|7134,7140|false|false|false|C0023882|Little's Disease|little
Event|Event|Discharge Instructions|7134,7140|false|false|false|||little
Finding|Finding|Discharge Instructions|7134,7140|false|false|false|C3889124|Only a Little|little
Finding|Finding|Discharge Instructions|7141,7144|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|Discharge Instructions|7141,7144|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Event|Event|Discharge Instructions|7152,7159|false|false|false|||regimen
Finding|Intellectual Product|Discharge Instructions|7152,7159|false|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|7152,7159|false|false|false|C0040808|Treatment Protocols|regimen
Event|Event|Discharge Instructions|7185,7191|false|false|false|||taking
Finding|Finding|Discharge Instructions|7192,7199|false|false|false|C4534363|At home|at home
Event|Event|Discharge Instructions|7195,7199|false|false|false|||home
Finding|Idea or Concept|Discharge Instructions|7195,7199|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Discharge Instructions|7195,7199|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Discharge Instructions|7195,7199|false|false|false|C1553498|home health encounter|home
Event|Event|Discharge Instructions|7202,7209|false|false|false|||Several
Event|Event|Discharge Instructions|7234,7241|false|false|false|||changed
Event|Event|Discharge Instructions|7247,7251|false|false|false|||made
Event|Event|Discharge Instructions|7266,7273|false|false|false|||changes
Finding|Functional Concept|Discharge Instructions|7266,7273|false|false|false|C0392747|Changing|changes
Attribute|Clinical Attribute|Discharge Instructions|7282,7293|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|7282,7293|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Discharge Instructions|7282,7293|false|false|false|||medications
Finding|Intellectual Product|Discharge Instructions|7282,7293|false|false|false|C4284232|Medications|medications
Event|Event|Discharge Instructions|7301,7308|false|false|false|||changed
Drug|Organic Chemical|Discharge Instructions|7314,7319|false|false|false|C0590690|Imdur|imdur
Drug|Pharmacologic Substance|Discharge Instructions|7314,7319|false|false|false|C0590690|Imdur|imdur
Event|Event|Discharge Instructions|7314,7319|false|false|false|||imdur
Event|Event|Discharge Instructions|7340,7347|false|false|false|||changed
Drug|Amino Acid, Peptide, or Protein|Discharge Instructions|7353,7363|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|Discharge Instructions|7353,7363|false|false|false|C0065374|lisinopril|lisinopril
Event|Event|Discharge Instructions|7353,7363|false|false|false|||lisinopril
Event|Event|Discharge Instructions|7383,7395|false|false|false|||discontinued
Drug|Organic Chemical|Discharge Instructions|7401,7409|false|false|false|C0004147|atenolol|atenolol
Drug|Pharmacologic Substance|Discharge Instructions|7401,7409|false|false|false|C0004147|atenolol|atenolol
Event|Event|Discharge Instructions|7401,7409|false|false|false|||atenolol
Event|Event|Discharge Instructions|7417,7424|false|false|false|||started
Drug|Organic Chemical|Discharge Instructions|7425,7435|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|Discharge Instructions|7425,7435|false|false|false|C0025859|metoprolol|metoprolol
Event|Event|Discharge Instructions|7425,7435|false|false|false|||metoprolol
Attribute|Clinical Attribute|Discharge Instructions|7470,7476|false|false|false|C1718621|W stress|stress
Drug|Organic Chemical|Discharge Instructions|7470,7476|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|Discharge Instructions|7470,7476|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Finding|Finding|Discharge Instructions|7470,7476|false|false|false|C0038435|Stress|stress
Procedure|Diagnostic Procedure|Discharge Instructions|7470,7481|false|false|false|C0015260;C3494508|Exercise stress test;Stress Test|stress test
Anatomy|Body Location or Region|Discharge Instructions|7477,7481|false|false|false|C4318744|Test - temporal region|test
Event|Event|Discharge Instructions|7477,7481|false|false|false|||test
Finding|Functional Concept|Discharge Instructions|7477,7481|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Finding|Intellectual Product|Discharge Instructions|7477,7481|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Lab|Laboratory or Test Result|Discharge Instructions|7477,7481|false|false|false|C0456984|Test Result|test
Procedure|Laboratory Procedure|Discharge Instructions|7477,7481|false|false|false|C0022885|Laboratory Procedures|test
Event|Event|Discharge Instructions|7491,7497|false|false|false|||normal
Event|Event|Discharge Instructions|7507,7515|false|false|false|||continue
Phenomenon|Phenomenon or Process|Discharge Instructions|7520,7526|false|false|false|C3714578|Fix|adhere
Finding|Functional Concept|Discharge Instructions|7520,7529|false|false|false|C4281991|Follow|adhere to
Finding|Finding|Discharge Instructions|7532,7544|false|false|false|C0452415|Diet, Healthy|healthy diet
Drug|Food|Discharge Instructions|7540,7544|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|Discharge Instructions|7540,7544|false|false|false|||diet
Finding|Functional Concept|Discharge Instructions|7540,7544|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|Discharge Instructions|7540,7544|false|false|false|C0012159|Diet therapy|diet
Event|Event|Discharge Instructions|7549,7557|false|false|false|||exercise
Finding|Daily or Recreational Activity|Discharge Instructions|7549,7557|false|false|false|C0015259|Exercise|exercise
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|7549,7557|false|false|false|C1522704|Exercise Pain Management|exercise
Finding|Functional Concept|Discharge Instructions|7590,7600|true|false|false|C1524062|Additional|additional
Anatomy|Body Location or Region|Discharge Instructions|7601,7606|true|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Discharge Instructions|7601,7606|true|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Discharge Instructions|7601,7611|true|false|false|C2926613||chest pain
Finding|Sign or Symptom|Discharge Instructions|7601,7611|true|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Discharge Instructions|7607,7611|true|false|false|C2598155||pain
Event|Event|Discharge Instructions|7607,7611|true|false|false|||pain
Finding|Functional Concept|Discharge Instructions|7607,7611|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|7607,7611|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Discharge Instructions|7613,7622|true|false|false|||shortness
Finding|Body Substance|Discharge Instructions|7627,7633|false|false|false|C0225386|Breath|breath
Attribute|Clinical Attribute|Discharge Instructions|7635,7641|false|false|false|C4255480||nausea
Event|Event|Discharge Instructions|7635,7641|false|false|false|||nausea
Finding|Sign or Symptom|Discharge Instructions|7635,7641|false|false|false|C0027497|Nausea|nausea
Event|Event|Discharge Instructions|7643,7651|false|false|false|||vomiting
Finding|Sign or Symptom|Discharge Instructions|7643,7651|false|false|false|C0042963|Vomiting|vomiting
Event|Event|Discharge Instructions|7660,7664|false|false|false|||call
Disorder|Disease or Syndrome|Discharge Instructions|7670,7673|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|Discharge Instructions|7670,7673|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|Discharge Instructions|7670,7673|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|Discharge Instructions|7670,7673|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|Discharge Instructions|7670,7673|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|Discharge Instructions|7670,7673|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|Discharge Instructions|7670,7673|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|Discharge Instructions|7670,7673|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|Discharge Instructions|7670,7673|false|false|false|||PCP
Finding|Gene or Genome|Discharge Instructions|7670,7673|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|Discharge Instructions|7670,7673|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Event|Discharge Instructions|7677,7683|false|false|false|||return
Procedure|Health Care Activity|Discharge Instructions|7700,7708|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|7709,7721|false|false|false|C3263700||Instructions
Event|Event|Discharge Instructions|7709,7721|false|false|false|||Instructions
Finding|Intellectual Product|Discharge Instructions|7709,7721|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

