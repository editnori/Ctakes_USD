CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|true|false||Unit
null|Unit device|Device|true|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|true|false||Unit
null|Unit of Measure|LabModifier|true|false||Unit
null|Unit|LabModifier|true|false||Unit
null|Enzyme Unit|LabModifier|true|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Pharmaceutical Preparations|Drug|false|false||MEDICINEnull|Medicine|Title|false|false||MEDICINEnull|lisinopril|Drug|false|false||lisinopril
null|lisinopril|Drug|false|false||lisinoprilnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Chest Pain|Finding|false|false||Chest Painnull|null|Attribute|false|false||Chest Painnull|Chest problem|Finding|false|false||Chestnull|Chest|Anatomy|false|false||Chest
null|Anterior thoracic region|Anatomy|false|false||Chestnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Exercise|Finding|false|false||Exercisenull|Exercise Pain Management|Procedure|false|false||Exercisenull|echocardiography service|Procedure|false|false||Echocardiography
null|Echocardiography|Procedure|false|false||Echocardiographynull|PMH - past medical history|Finding|false|false||pmh
null|Medical History|Finding|false|false||pmhnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Known|Modifier|false|false||knownnull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Coronary Artery Bypass Surgery|Procedure|false|false||CABGnull|Numerous|LabModifier|false|false||multiplenull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Management procedure|Event|false|false||managednull|Angina Pectoris|Finding|false|false||angina
null|null|Finding|false|false||anginanull|null|Attribute|false|false||anginanull|Hypertensive disease|Disorder|false|false||HTNnull|Atypical chest pain|Finding|false|false||atypical chest painnull|atypia morphology|Finding|false|false||atypicalnull|Atypical|Modifier|false|false||atypicalnull|Chest Pain|Finding|false|false||chest painnull|null|Attribute|false|false||chest painnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Has patient|Finding|false|false||Patient hasnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Vessel Positions|Anatomy|false|false||vessel
null|Blood Vessel|Anatomy|false|false||vesselnull|Vessel (unit of presentation)|LabModifier|false|false||vesselnull|Coronary Artery Bypass Surgery|Procedure|false|false||CABGnull|Lima|Entity|false|false||LIMAnull|Leukocyte adhesion deficiency type 1|Disorder|false|false||LAD
null|Leukocyte adhesion deficiency|Disorder|false|false||LADnull|ITGB2 wt Allele|Finding|false|false||LAD
null|DLD gene|Finding|false|false||LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false||LADnull|Ladino Language|Entity|false|false||LADnull|Scalable Vector Graphics|Entity|false|false||SVGnull|Scalable Vector Graphics|Entity|false|false||SVGnull|null|Disorder|false|false||NSTEMInull|null|Finding|false|false||NSTEMInull|Catheterization|Procedure|false|false||cathnull|Occluded|Finding|false|false||occluded
null|Obstruction|Finding|false|false||occludednull|Graft Dosage Form|Drug|false|false||graft
null|Graft material|Drug|false|false||graftnull|Graft - Specimen Source Codes|Finding|false|false||graftnull|Graft Procedures on the Head|Procedure|false|false||graft
null|Grafting procedure|Procedure|false|false||graftnull|Transplanted tissue|Anatomy|false|false||graftnull|Small|LabModifier|false|false||smallnull|Diagonal|Modifier|false|false||diagonalnull|Macromolecular Branch|Drug|false|false||branchnull|Branch of|Modifier|false|false||branchnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Stenosis|Finding|false|false||stenosisnull|Stenosis <Pimeliinae>|Entity|false|false||stenosisnull|Stenosis Morphology|Modifier|false|false||stenosisnull|Leukocyte adhesion deficiency type 1|Disorder|false|false||LAD
null|Leukocyte adhesion deficiency|Disorder|false|false||LADnull|ITGB2 wt Allele|Finding|false|false||LAD
null|DLD gene|Finding|false|false||LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false||LADnull|Ladino Language|Entity|false|false||LADnull|null|Device|false|false||stentnull|Stenosis|Finding|false|false||stenosisnull|Stenosis <Pimeliinae>|Entity|false|false||stenosisnull|Stenosis Morphology|Modifier|false|false||stenosisnull|Methylcytosine Dioxygenase TET1|Drug|false|false||LCx
null|Methylcytosine Dioxygenase TET1|Drug|false|false||LCxnull|TET1 wt Allele|Finding|false|false||LCx
null|TET1 gene|Finding|false|false||LCxnull|Participation Type - origin|Finding|false|false||origin
null|National origin|Finding|false|false||originnull|Beginning|Time|false|false||originnull|Imdur|Drug|false|false||Imdur
null|Imdur|Drug|false|false||Imdurnull|Transcription Initiation|Finding|false|false||initiation
null|Initiation|Finding|false|false||initiation
null|null|Finding|false|false||initiationnull|AOD use initiation|Time|false|false||initiationnull|losartan|Drug|false|false||losartan
null|losartan|Drug|false|false||losartannull|Observation Interpretation - better|Finding|false|false||betternull|Better|Modifier|false|false||betternull|Control brand of phenylpropanolamine|Drug|false|false||control
null|CONTROL veterinary product|Drug|false|false||control
null|control substance|Drug|false|false||control
null|Control brand of phenylpropanolamine|Drug|false|false||controlnull|Control - Relationship modifier|Finding|false|false||control
null|Control function|Finding|false|false||control
null|Scientific Control|Finding|false|false||controlnull|Control Groups|Subject|false|false||controlnull|True Control Status|Modifier|false|false||control
null|control aspects|Modifier|false|false||controlnull|Often - answer to question|Finding|false|false||oftennull|Frequently|Time|false|false||oftennull|Angina, Unstable|Disorder|false|false||angina at rest
null|Angina decubitus|Disorder|false|false||angina at restnull|Angina Pectoris|Finding|false|false||angina
null|null|Finding|false|false||anginanull|null|Attribute|false|false||anginanull|At rest (qualifier value)|Finding|false|false||at restnull|REST protein, human|Drug|false|false||rest
null|REST protein, human|Drug|false|false||restnull|REST gene|Finding|false|false||rest
null|site-specific telomere resolvase activity|Finding|false|false||rest
null|Rest|Finding|false|false||restnull|Recent|Time|false|false||recentnull|BaseLine dental cement|Drug|false|false||baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|nitroglycerin|Drug|false|false||nitroglycerin
null|nitroglycerin|Drug|false|false||nitroglycerinnull|Approximate|Modifier|false|false||approximatelynull|Twice weekly|Time|false|false||twice weeklynull|Weekly|Time|false|false||weeklynull|Frequently|Time|false|false||frequentnull|Chest Pain|Finding|false|false||chest painsnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Pain|Finding|false|false||painsnull|Different|Modifier|false|false||differentnull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Angina Pectoris|Finding|false|false||angina
null|null|Finding|false|false||anginanull|null|Attribute|false|false||anginanull|Usually|Finding|false|false||usuallynull|Usual|Modifier|false|false||usuallynull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Current (present time)|Time|false|false||currentlynull|More|LabModifier|false|false||morenull|null|Finding|false|false||needlenull|Needle device|Device|false|false||needlenull|Needle Shape|Modifier|false|false||needlenull|Puncture wound|Disorder|false|false||pricksnull|Pricking sensation quality|Finding|false|false||pricksnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|More|LabModifier|false|false||morenull|Persistent|Time|false|false||persistentnull|Significant|Finding|true|false||significantnull|Event Seriousness - Significant|Modifier|true|false||significantnull|Relief brand of phenylephrine|Drug|true|false||relief
null|Relief brand of phenylephrine|Drug|true|false||reliefnull|Feeling relief|Finding|true|false||reliefnull|Observation Interpretation - worse|Finding|false|false||worse
null|Worse|Finding|false|false||worsenull|Worsening (qualifier value)|Modifier|false|false||worsenull|Breathing abnormally deep|Finding|false|false||deep breathing
null|Deep breathing|Finding|false|false||deep breathingnull|Deep Resection Margin|Attribute|false|false||deepnull|Deep (qualifier value)|Modifier|false|false||deepnull|outcomes otolaryngology breathing|Finding|false|false||breathing
null|Inspiration (function)|Finding|false|false||breathing
null|Respiration|Finding|false|false||breathingnull|null|Attribute|false|false||breathingnull|respiratory system process|Phenomenon|false|false||breathingnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|Anterior chest wall structure|Anatomy|false|false||anterior chestnull|Adenohypophyseal Diseases|Disorder|false|false||anteriornull|Anterior|Modifier|false|false||anteriornull|Chest problem|Finding|false|false||chestnull|Anterior thoracic region|Anatomy|false|false||chest
null|Chest|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|true|false||pain
null|Pain|Finding|true|false||painnull|null|Attribute|true|false||painnull|Coronary Artery Bypass Surgery|Procedure|false|false||CABGnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Dyspnea|Finding|false|false||SOBnull|Increased sweating|Finding|false|false||diaphoresisnull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|Palpitations|Finding|false|false||palpitationsnull|Paroxysmal|Time|true|false||paroxysmalnull|null|Finding|true|false||dyspnea
null|Dyspnea|Finding|true|false||dyspneanull|sleeping upright or using specific number of extra pillows (orthopnea)|Finding|true|false||orthopnea
null|Orthopnea|Finding|true|false||orthopneanull|Ankle edema (finding)|Finding|false|false||ankle edemanull|Lower extremity>Ankle|Anatomy|false|false||ankle
null|Ankle|Anatomy|false|false||ankle
null|Ankle joint structure|Anatomy|false|false||anklenull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Palpitations|Finding|false|false||palpitationsnull|Syncope|Finding|false|false||syncopenull|Syncope <Gastrophryninae>|Entity|false|false||syncopenull|Presyncope|Finding|false|false||presyncopenull|More|LabModifier|true|false||morenull|Cold brand of chlorpheniramine-phenylpropanolamine|Drug|true|false||cold
null|Cold brand of chlorpheniramine-phenylpropanolamine|Drug|true|false||coldnull|Common Cold|Disorder|true|false||cold
null|Chronic Obstructive Airway Disease|Disorder|true|false||coldnull|Cold Sensation|Finding|true|false||coldnull|Cold Therapy|Procedure|true|false||coldnull|Cold Temperature|Phenomenon|true|false||coldnull|Usual|Modifier|true|false||usualnull|Recent|Time|true|false||recentlynull|NUT Family Member 1, human|Drug|true|false||nut
null|NUT Family Member 1, human|Drug|true|false||nut
null|Nuts|Drug|true|false||nutnull|NUTM1 wt Allele|Finding|true|false||nut
null|NUTM1 gene|Finding|true|false||nutnull|Nut Device|Device|true|false||nutnull|Fever|Finding|true|false||feversnull|Chills|Finding|true|false||chillsnull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|Complaint (finding)|Finding|true|false||complaintsnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Current (present time)|Time|false|false||currentlynull|Loss (adaptation)|Finding|false|false||lossnull|Loss (quantitative)|LabModifier|false|false||lossnull|Impaired cognition|Disorder|false|false||cognitive impairmentnull|Cognitive|Finding|false|false||cognitivenull|Impaired health|Finding|false|false||impairment
null|Impaired|Finding|false|false||impairmentnull|Course|Time|false|false||Coursenull|Electrocardiogram image|Finding|false|false||EKG
null|Electrocardiogram|Finding|false|false||EKGnull|Electrocardiography|Procedure|false|false||EKGnull|Sinus brand of acetaminophen-pseudoephedrine|Drug|false|false||sinus
null|Sinus brand of acetaminophen-pseudoephedrine|Drug|false|false||sinusnull|pathologic fistula|Disorder|false|false||sinusnull|Sinus - general anatomical term|Anatomy|false|false||sinus
null|Nasal sinus|Anatomy|false|false||sinusnull|Lateral|Modifier|true|false||lateralnull|Mental Depression|Disorder|true|false||depressionsnull|Similarity|Modifier|true|false||similarnull|null|Time|true|false||priornull|Query Status Code - new|Finding|true|false||new
null|Act Status - new|Finding|true|false||newnull|Newar Language|Entity|true|false||newnull|New|Modifier|true|false||newnull|Ischemic|Finding|true|false||ischemicnull|Laboratory test finding|Lab|false|false||Labsnull|null|Modifier|false|false||unremarkablenull|Neg - answer|Finding|false|false||negnull|Negative - qualifier|Modifier|false|false||negnull|Plain chest X-ray|Procedure|false|false||CXRnull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|cardiac risk factors|Finding|false|false||CARDIAC RISK FACTORSnull|CARD.RISK|Finding|false|false||CARDIAC RISKnull|Cardiac attachment|Finding|false|false||CARDIACnull|Heart|Anatomy|false|false||CARDIACnull|Cardiac - anatomy qualifier|Modifier|false|false||CARDIACnull|risk factors - observation list|Finding|false|false||RISK FACTORS
null|risk factors|Finding|false|false||RISK FACTORS
null|History of - risk factor|Finding|false|false||RISK FACTORSnull|null|Attribute|false|false||RISK FACTORSnull|Risk|Finding|false|false||RISKnull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||Diabetes
null|Diabetes|Disorder|false|false||Diabetes
null|Diabetes Mellitus|Disorder|false|false||Diabetesnull|Dyslipidemias|Disorder|false|false||Dyslipidemianull|Hypertensive disease|Disorder|false|false||HTNnull|Cardiac attachment|Finding|false|false||CARDIACnull|Heart|Anatomy|false|false||CARDIACnull|Cardiac - anatomy qualifier|Modifier|false|false||CARDIACnull|Coronary Artery Disease|Disorder|false|false||Coronary artery disease
null|Coronary Arteriosclerosis|Disorder|false|false||Coronary artery diseasenull|Coronary artery|Anatomy|false|false||Coronary arterynull|Heart|Anatomy|false|false||Coronarynull|Coronary|Modifier|false|false||Coronarynull|Arteriopathic disease|Disorder|false|false||artery diseasenull|Arterial system|Anatomy|false|false||artery
null|Arteries|Anatomy|false|false||arterynull|Disease|Disorder|false|false||diseasenull|diastolic congestive heart failure|Disorder|false|false||Diastolic congestive heart failurenull|Diastole|Attribute|false|false||Diastolicnull|Congestive heart failure|Disorder|false|false||congestive heart failurenull|Congestive|Modifier|false|false||congestivenull|Congestive heart failure|Disorder|false|false||heart failure
null|Heart failure|Disorder|false|false||heart failurenull|Malignant neoplasm of heart|Disorder|false|false||heart
null|benign neoplasm of heart|Disorder|false|false||heartnull|HEART PROBLEM|Finding|false|false||heartnull|Chest>Heart|Anatomy|false|false||heart
null|Heart|Anatomy|false|false||heartnull|Failure (biologic function)|Finding|false|false||failure
null|Failure|Finding|false|false||failure
null|Personal failure|Finding|false|false||failurenull|Coronary Artery Bypass Surgery|Procedure|false|false||CABGnull|Coronary Artery Bypass Surgery|Procedure|false|false||CABGnull|Coronary Artery Bypass, Off-Pump|Procedure|false|false||Off pump coronary artery bypassnull|matrix metalloproteinase 7 activity|Finding|false|false||pumpnull|null|Device|false|false||pumpnull|Pump Dosing Unit|LabModifier|false|false||pumpnull|Coronary Artery Bypass Surgery|Procedure|false|false||coronary artery bypass graftnull|coronary artery graft device|Device|false|false||coronary artery bypass graftnull|Coronary Artery Bypass Surgery|Procedure|false|false||coronary artery bypassnull|Coronary artery|Anatomy|false|false||coronary arterynull|Heart|Anatomy|false|false||coronarynull|Coronary|Modifier|false|false||coronarynull|Arterial bypass graft|Procedure|false|false||artery bypass graftnull|Arterial system|Anatomy|false|false||artery
null|Arteries|Anatomy|false|false||arterynull|Bypass graft|Procedure|false|false||bypass graftnull|Creation of shunt|Procedure|false|false||bypassnull|Graft Dosage Form|Drug|false|false||graft
null|Graft material|Drug|false|false||graftnull|Graft - Specimen Source Codes|Finding|false|false||graftnull|Graft Procedures on the Head|Procedure|false|false||graft
null|Grafting procedure|Procedure|false|false||graftnull|Transplanted tissue|Anatomy|false|false||graftnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Structure of internal thoracic artery|Anatomy|false|false||internal mammary arterynull|Code System Type - Internal|Modifier|false|false||internal
null|Internal Surface|Modifier|false|false||internal
null|Internal|Modifier|false|false||internalnull|Mammary Arteries|Anatomy|false|false||mammary arterynull|Mammary gland|Anatomy|false|false||mammary
null|Breast|Anatomy|false|false||mammarynull|Arterial system|Anatomy|false|false||artery
null|Arteries|Anatomy|false|false||arterynull|Anterior descending branch of left coronary artery|Anatomy|false|false||left anterior descending artery
null|null|Anatomy|false|false||left anterior descending arterynull|Left anterior|Modifier|false|false||left anteriornull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Adenohypophyseal Diseases|Disorder|false|false||anteriornull|Anterior|Modifier|false|false||anteriornull|Sequencing - Descending|Finding|false|false||descendingnull|Descending|Modifier|false|false||descendingnull|Arterial system|Anatomy|false|false||artery
null|Arteries|Anatomy|false|false||arterynull|Great saphenous vein structure|Anatomy|false|false||saphenous vein
null|Saphenous Vein|Anatomy|false|false||saphenous veinnull|Veins|Anatomy|false|false||veinnull|Graft material|Drug|false|false||graftsnull|Transplanted tissue|Anatomy|false|false||graftsnull|grafting qualifier|Modifier|false|false||graftsnull|Diagonal|Modifier|false|false||diagonalnull|Obtuse|Modifier|false|false||obtusenull|Target Awareness - marginal|Finding|false|false||marginalnull|Marginal (quality)|Modifier|false|false||marginal
null|Marginal|Modifier|false|false||marginalnull|Procedure on artery|Procedure|false|false||arteriesnull|Arteries|Anatomy|false|false||arteries
null|Arterial system|Anatomy|false|false||arteriesnull|Percutaneous Coronary Intervention|Procedure|false|false||PERCUTANEOUS CORONARY INTERVENTIONSnull|Percutaneous Route of Drug Administration|Finding|false|false||PERCUTANEOUSnull|Percutaneous|Modifier|false|false||PERCUTANEOUSnull|Heart|Anatomy|false|false||CORONARYnull|Coronary|Modifier|false|false||CORONARYnull|Nursing interventions|Procedure|false|false||INTERVENTIONS
null|Intervention regimes|Procedure|false|false||INTERVENTIONSnull|null|Attribute|false|false||INTERVENTIONSnull|Burning Mouth Syndrome|Disorder|false|false||BMSnull|Proximal Resection Margin|Attribute|false|false||proximalnull|Proximal|Modifier|false|false||proximalnull|Leukocyte adhesion deficiency type 1|Disorder|false|false||LAD
null|Leukocyte adhesion deficiency|Disorder|false|false||LADnull|ITGB2 wt Allele|Finding|false|false||LAD
null|DLD gene|Finding|false|false||LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false||LADnull|Ladino Language|Entity|false|false||LADnull|DES protein, human|Drug|false|false||DES
null|Desmosine|Drug|false|false||DES
null|Desmosine|Drug|false|false||DES
null|DES protein, human|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DESnull|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|Disorder|false|false||DESnull|DES gene|Finding|false|false||DESnull|Middle|Modifier|false|false||midnull|Leukocyte adhesion deficiency type 1|Disorder|false|false||LAD
null|Leukocyte adhesion deficiency|Disorder|false|false||LADnull|ITGB2 wt Allele|Finding|false|false||LAD
null|DLD gene|Finding|false|false||LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false||LADnull|Ladino Language|Entity|false|false||LADnull|DES protein, human|Drug|false|false||DES
null|Desmosine|Drug|false|false||DES
null|Desmosine|Drug|false|false||DES
null|DES protein, human|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DESnull|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|Disorder|false|false||DESnull|DES gene|Finding|false|false||DESnull|Graph Edge|Finding|false|false||edgenull|Along edge (qualifier value)|Modifier|false|false||edgenull|Middle|Modifier|false|false||midnull|Leukocyte adhesion deficiency type 1|Disorder|false|false||LAD
null|Leukocyte adhesion deficiency|Disorder|false|false||LADnull|ITGB2 wt Allele|Finding|false|false||LAD
null|DLD gene|Finding|false|false||LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false||LADnull|Ladino Language|Entity|false|false||LADnull|DES protein, human|Drug|false|false||DES
null|Desmosine|Drug|false|false||DES
null|Desmosine|Drug|false|false||DES
null|DES protein, human|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DESnull|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|Disorder|false|false||DESnull|DES gene|Finding|false|false||DESnull|Stenosis|Finding|false|false||stenosisnull|Stenosis <Pimeliinae>|Entity|false|false||stenosisnull|Stenosis Morphology|Modifier|false|false||stenosisnull|Distal Resection Margin|Attribute|false|false||distalnull|Distal (qualifier value)|Modifier|false|false||distalnull|null|Device|false|false||stentnull|DES protein, human|Drug|false|false||DES
null|Desmosine|Drug|false|false||DES
null|Desmosine|Drug|false|false||DES
null|DES protein, human|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DESnull|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|Disorder|false|false||DESnull|DES gene|Finding|false|false||DESnull|Pacing up and down|Finding|false|false||PACINGnull|Disruptive, Impulse Control, and Conduct Disorders|Disorder|false|false||ICD
null|Type II Mucolipidosis|Disorder|false|false||ICDnull|International Classification of Diseases|Finding|false|false||ICD
null|GNPTAB wt Allele|Finding|false|false||ICDnull|Icd Regimen|Procedure|false|false||ICDnull|between lunch and dinner|Time|false|false||ICDnull|Morbid obesity|Disorder|true|false||Morbid obesitynull|Obesity|Disorder|true|false||obesitynull|BODY MASS INDEX QUANTITATIVE TRAIT LOCUS 20|Finding|true|false||obesitynull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|Gastroesophageal reflux disease|Disorder|false|false||GERDnull|Right tendinous cuff|Anatomy|false|false||Right rotator cuffnull|Table Cell Horizontal Align - right|Finding|false|false||Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|Rotator Cuff Injuries|Disorder|false|false||rotator cuff injurynull|Rotator Cuff|Anatomy|false|false||rotator cuffnull|null|Device|false|false||rotatornull|Cuffing (morphologic abnormality)|Finding|false|false||cuffnull|Cuff - body part|Anatomy|false|false||cuffnull|Cuff Device|Device|false|false||cuffnull|Traumatic AND/OR non-traumatic injury|Disorder|false|false||injury
null|Traumatic injury|Disorder|false|false||injurynull|Bursitis|Disorder|false|false||bursitisnull|Migraine Disorders|Disorder|false|false||Migrainesnull|Cancer patients and suicide and depression|Disorder|false|false||Depression
null|Mental Depression|Disorder|false|false||Depression
null|Depressive disorder|Disorder|false|false||Depression
null|Depressed mood|Disorder|false|false||Depressionnull|Depression - motion|Finding|false|false||Depression
null|null|Finding|false|false||Depressionnull|Depression - recess|Modifier|false|false||Depressionnull|Degenerative polyarthritis|Disorder|false|false||DJDnull|Hemorrhoids|Disorder|false|false||Hemorrhoidsnull|Rosacea|Disorder|false|false||Rosaceanull|Rosacea <Prayinae>|Entity|false|false||Rosaceanull|Ward (environment)|Device|false|false||wardnull|Ward (person)|Subject|false|false||wardnull|Ward (environment)|Entity|false|false||wardnull|ErbB Receptors|Drug|true|false||her family
null|ErbB Receptors|Drug|true|false||her familynull|ErbB Receptors|Finding|true|false||her familynull|Entity Name Part Type - family|Finding|true|false||family
null|Last Name|Finding|true|false||family
null|Living Arrangement - Family|Finding|true|false||family
null|Family (taxonomic)|Finding|true|false||family
null|Family Collection|Finding|true|false||familynull|Family|Subject|true|false||familynull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|Exam|Finding|false|false||EXAMnull|Medical Examination|Procedure|false|false||EXAMnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||GENERALnull|General medical service|Procedure|false|false||GENERALnull|Generalized|Modifier|false|false||GENERALnull|Oriented to place|Finding|false|false||Orientednull|Orientation, Spatial|Modifier|false|false||Orientednull|Mood (psychological function)|Finding|false|false||Mood
null|mood (physical finding)|Finding|false|false||Mood
null|Mood (attribute)|Finding|false|false||Moodnull|null|Attribute|false|false||Moodnull|Appropriate|Modifier|false|false||appropriatenull|HEENT|Anatomy|false|false||HEENTnull|Scleral Diseases|Disorder|false|false||Scleranull|examination of sclera|Procedure|false|false||Scleranull|Sclera|Anatomy|false|false||Scleranull|Anicteric|Finding|false|false||anictericnull|Pupil equal round and reacting to light|Finding|false|false||PERRLnull|Malignant neoplasm of conjunctiva|Disorder|true|false||Conjunctiva
null|Benign neoplasm of conjunctiva|Disorder|true|false||Conjunctiva
null|Conjunctival Diseases|Disorder|true|false||Conjunctivanull|Specimen Type - Conjunctiva|Finding|true|false||Conjunctiva
null|null|Finding|true|false||Conjunctivanull|examination of conjunctiva|Procedure|true|false||Conjunctiva
null|Procedure on conjunctiva|Procedure|true|false||Conjunctivanull|Structure of palpebral conjunctiva|Anatomy|true|false||Conjunctiva
null|conjunctiva|Anatomy|true|false||Conjunctivanull|Pink color|Modifier|true|false||pinknull|Pallor of skin|Finding|true|false||pallornull|Cyanosis|Finding|true|false||cyanosisnull|Oral mucous membrane structure|Anatomy|true|false||oral mucosanull|Oral Dosage Form|Drug|true|false||oralnull|Oral Route of Administration|Finding|true|false||oral
null|Oral (intended site)|Finding|true|false||oralnull|Oral cavity|Anatomy|true|false||oralnull|Oral|Modifier|true|false||oralnull|null|Finding|true|false||mucosanull|Mucous Membrane|Anatomy|true|false||mucosanull|Eyelid Xanthoma|Disorder|true|false||xanthelasma
null|Xanthoma|Disorder|true|false||xanthelasmanull|Passive joint movement of neck (finding)|Finding|false|false||NECK
null|Neck problem|Finding|false|false||NECKnull|dendritic spine neck|Anatomy|false|false||NECK
null|Neck|Anatomy|false|false||NECKnull|Supple|Finding|false|false||Supplenull|Jugular venous pressure|Finding|false|false||JVPnull|Chest problem|Finding|false|false||Chestnull|Chest|Anatomy|false|false||Chest
null|Anterior thoracic region|Anatomy|false|false||Chestnull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|Diffuse|Modifier|false|false||diffusenull|thiamine triphosphorate|Drug|false|false||TTP
null|ZFP36 protein, human|Drug|false|false||TTP
null|ZFP36 protein, human|Drug|false|false||TTP
null|thiamine triphosphorate|Drug|false|false||TTPnull|Congenital Thrombotic Thrombocytopenic Purpura|Disorder|false|false||TTP
null|Purpura, Thrombotic Thrombocytopenic|Disorder|false|false||TTPnull|ZFP36 wt Allele|Finding|false|false||TTP
null|ZFP36 gene|Finding|false|false||TTP
null|ADAMTS13 gene|Finding|false|false||TTPnull|Time to Progression|Time|false|false||TTPnull|Anterior chest wall structure|Anatomy|false|false||anterior chest wall
null|null|Anatomy|false|false||anterior chest wallnull|Anterior chest wall structure|Anatomy|false|false||anterior chestnull|Adenohypophyseal Diseases|Disorder|false|false||anteriornull|Anterior|Modifier|false|false||anteriornull|Chest wall structure|Anatomy|false|false||chest wall
null|Chest>Chest wall|Anatomy|false|false||chest wallnull|Chest problem|Finding|false|false||chestnull|Anterior thoracic region|Anatomy|false|false||chest
null|Chest|Anatomy|false|false||chestnull|Walls of a building|Device|false|false||wallnull|Cardiac attachment|Finding|false|false||CARDIACnull|Heart|Anatomy|false|false||CARDIACnull|Cardiac - anatomy qualifier|Modifier|false|false||CARDIACnull|Coronary Artery Bypass Surgery|Procedure|true|false||CABGnull|Cardiac thrill (finding)|Finding|true|false||thrillsnull|hoist [device]|Device|true|false||liftsnull|Lung|Anatomy|false|false||LUNGSnull|Coarse|Modifier|false|false||coarsenull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Basilar|Modifier|false|false||basilarnull|Basilar Rales|Finding|false|false||crackles
null|Rales|Finding|false|false||cracklesnull|Consistent with|Finding|false|false||consistent withnull|Compatible|Modifier|false|false||consistent withnull|Consistent with|Finding|false|false||consistentnull|Pleural Diseases|Disorder|false|false||pleuralnull|Pleura|Anatomy|false|false||pleuralnull|Pleural|Modifier|false|false||pleuralnull|Process Pharmacologic Substance|Drug|false|false||processnull|Process (qualifier value)|Finding|false|false||processnull|bony process|Anatomy|false|false||processnull|Process|Phenomenon|false|false||processnull|Plain chest X-ray|Procedure|true|false||CXRnull|Language Ability Proficiency - Good|Finding|true|false||good
null|Language Proficiency - Good|Finding|true|false||goodnull|Specimen Quality - Good|Modifier|true|false||good
null|Good|Modifier|true|false||goodnull|Air Movements|Phenomenon|true|false||air movementnull|Air (substance)|Drug|true|false||air
null|air|Drug|true|false||air
null|air|Drug|true|false||airnull|ACUTE INSULIN RESPONSE|Finding|true|false||air
null|AIRN gene|Finding|true|false||air
null|AI/RHEUM|Finding|true|false||airnull|Movement|Finding|true|false||movementnull|Wheezing|Finding|true|false||wheezesnull|Rhonchi|Finding|true|false||rhonchinull|Malignant neoplasm of abdomen|Disorder|false|false||ABDOMENnull|Abdomen problem|Finding|false|false||ABDOMENnull|Abdomen|Anatomy|false|false||ABDOMEN
null|Abdominal Cavity|Anatomy|false|false||ABDOMENnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||Softnull|Soft|Modifier|false|false||Softnull|LRRC4B gene|Finding|true|false||HSMnull|Emotional tenderness|Finding|true|false||tenderness
null|Sore to touch|Finding|true|false||tendernessnull|Absence of Biallelic TCRgamma Deletion|Disorder|true|false||Abdnull|ABD (body structure)|Anatomy|true|false||Abd
null|Abdomen|Anatomy|true|false||Abdnull|Procedure on aorta|Procedure|true|false||aortanull|Chest+Abdomen>Aorta|Anatomy|true|false||aorta
null|Aorta|Anatomy|true|false||aortanull|Palpation|Procedure|true|false||palpationnull|Abdominal bruit|Finding|true|false||abdominal bruitsnull|Abdomen|Anatomy|true|false||abdominalnull|Abdominal (qualifier value)|Modifier|true|false||abdominalnull|Bruit|Finding|true|false||bruitsnull|All extremities|Anatomy|false|false||EXTREMITIES
null|Limb structure|Anatomy|false|false||EXTREMITIESnull|Femur|Anatomy|true|false||femoralnull|Bruit|Finding|true|false||bruitsnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false||SKIN
null|Skin and subcutaneous tissue disorders|Disorder|false|false||SKINnull|Skin Specimen Source Code|Finding|false|false||SKIN
null|Skin Specimen|Finding|false|false||SKINnull|Skin, Human|Anatomy|false|false||SKIN
null|Skin|Anatomy|false|false||SKINnull|Stasis dermatitis|Disorder|true|false||stasis dermatitisnull|Stasis|Finding|true|false||stasisnull|Dermatitis|Disorder|true|false||dermatitisnull|Ulcer|Finding|true|false||ulcersnull|Scar Tissue|Finding|true|false||scars
null|Cicatrix|Finding|true|false||scarsnull|Xanthoma|Disorder|true|false||xanthomasnull|null|Drug|false|false||PULSESnull|Physiologic pulse|Finding|false|false||PULSESnull|Pulse taking|Procedure|false|false||PULSESnull|Neurology speciality|Title|false|false||Neuronull|Neurologic (qualifier value)|Modifier|false|false||Neuronull|Gross (qualifier value)|Modifier|true|false||grossnull|Deficit|Modifier|true|false||deficitsnull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|Exam|Finding|false|false||EXAMnull|Medical Examination|Procedure|false|false||EXAMnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||GENERALnull|General medical service|Procedure|false|false||GENERALnull|Generalized|Modifier|false|false||GENERALnull|Oriented to place|Finding|false|false||Orientednull|Orientation, Spatial|Modifier|false|false||Orientednull|Mood (psychological function)|Finding|false|false||Mood
null|mood (physical finding)|Finding|false|false||Mood
null|Mood (attribute)|Finding|false|false||Moodnull|null|Attribute|false|false||Moodnull|Appropriate|Modifier|false|false||appropriatenull|Flat affect|Finding|false|false||flat affectnull|Residential flat|Device|false|false||flatnull|Flat shape|Modifier|false|false||flatnull|Affect (mental function)|Finding|false|false||affectnull|assessment of affect|Procedure|false|false||affectnull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|HEENT|Anatomy|false|false||HEENTnull|Scleral Diseases|Disorder|false|false||Scleranull|examination of sclera|Procedure|false|false||Scleranull|Sclera|Anatomy|false|false||Scleranull|Anicteric|Finding|false|false||anictericnull|Pupil equal round and reacting to light|Finding|false|false||PERRLnull|Malignant neoplasm of conjunctiva|Disorder|true|false||Conjunctiva
null|Benign neoplasm of conjunctiva|Disorder|true|false||Conjunctiva
null|Conjunctival Diseases|Disorder|true|false||Conjunctivanull|Specimen Type - Conjunctiva|Finding|true|false||Conjunctiva
null|null|Finding|true|false||Conjunctivanull|examination of conjunctiva|Procedure|true|false||Conjunctiva
null|Procedure on conjunctiva|Procedure|true|false||Conjunctivanull|Structure of palpebral conjunctiva|Anatomy|true|false||Conjunctiva
null|conjunctiva|Anatomy|true|false||Conjunctivanull|Pink color|Modifier|true|false||pinknull|Pallor of skin|Finding|true|false||pallornull|Cyanosis|Finding|true|false||cyanosisnull|Oral mucous membrane structure|Anatomy|true|false||oral mucosanull|Oral Dosage Form|Drug|true|false||oralnull|Oral Route of Administration|Finding|true|false||oral
null|Oral (intended site)|Finding|true|false||oralnull|Oral cavity|Anatomy|true|false||oralnull|Oral|Modifier|true|false||oralnull|null|Finding|true|false||mucosanull|Mucous Membrane|Anatomy|true|false||mucosanull|Eyelid Xanthoma|Disorder|true|false||xanthelasma
null|Xanthoma|Disorder|true|false||xanthelasmanull|Structure of cornea of left eye|Anatomy|false|false||Left corneanull|Table Cell Horizontal Align - left|Finding|false|false||Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|Malignant neoplasm of cornea|Disorder|false|false||cornea
null|Corneal Diseases|Disorder|false|false||cornea
null|Benign neoplasm of cornea|Disorder|false|false||corneanull|SpecimenType - Cornea|Finding|false|false||corneanull|Cornea|Anatomy|false|false||corneanull|Scar Tissue|Finding|false|false||scar tissue
null|Cicatrix|Finding|false|false||scar tissuenull|Scar Tissue|Finding|false|false||scar
null|Cicatrix|Finding|false|false||scar
null|RPS4X gene|Finding|false|false||scarnull|Tissue Specimen Code|Finding|false|false||tissuenull|Body tissue|Anatomy|false|false||tissuenull|Medial|Modifier|false|false||medialnull|Passive joint movement of neck (finding)|Finding|false|false||NECK
null|Neck problem|Finding|false|false||NECKnull|dendritic spine neck|Anatomy|false|false||NECK
null|Neck|Anatomy|false|false||NECKnull|Supple|Finding|false|false||Supplenull|Residential flat|Device|false|false||flatnull|Flat shape|Modifier|false|false||flatnull|Jugular venous pressure|Finding|false|false||JVPnull|Goiter|Disorder|true|false||thyromegalynull|Chest problem|Finding|false|false||CHESTnull|Chest|Anatomy|false|false||CHEST
null|Anterior thoracic region|Anatomy|false|false||CHESTnull|thiamine triphosphorate|Drug|false|false||TTP
null|ZFP36 protein, human|Drug|false|false||TTP
null|ZFP36 protein, human|Drug|false|false||TTP
null|thiamine triphosphorate|Drug|false|false||TTPnull|Congenital Thrombotic Thrombocytopenic Purpura|Disorder|false|false||TTP
null|Purpura, Thrombotic Thrombocytopenic|Disorder|false|false||TTPnull|ZFP36 wt Allele|Finding|false|false||TTP
null|ZFP36 gene|Finding|false|false||TTP
null|ADAMTS13 gene|Finding|false|false||TTPnull|Time to Progression|Time|false|false||TTPnull|Sternum|Anatomy|false|false||sternumnull|Cardiac attachment|Finding|false|false||CARDIACnull|Heart|Anatomy|false|false||CARDIACnull|Cardiac - anatomy qualifier|Modifier|false|false||CARDIACnull|distant heart sounds|Finding|false|false||Distant heart soundsnull|Distant Metastasis|Finding|false|false||Distantnull|Distant|Modifier|false|false||Distantnull|Heart Sounds|Finding|false|false||heart soundsnull|auscultation of heart sounds|Procedure|false|false||heart soundsnull|null|Attribute|false|false||heart soundsnull|Malignant neoplasm of heart|Disorder|false|false||heart
null|benign neoplasm of heart|Disorder|false|false||heartnull|HEART PROBLEM|Finding|false|false||heartnull|Chest>Heart|Anatomy|false|false||heart
null|Heart|Anatomy|false|false||heartnull|null|Device|false|false||soundsnull|null|Phenomenon|false|false||soundsnull|Cardiac thrill (finding)|Finding|true|false||thrillsnull|hoist [device]|Device|true|false||liftsnull|Lung|Anatomy|false|false||LUNGSnull|cetrimonium bromide|Drug|true|false||CTABnull|Wheezing|Finding|true|false||wheezingnull|Basilar Rales|Finding|true|false||rales
null|Rales|Finding|true|false||ralesnull|Rhonchi|Finding|true|false||rhonchinull|Malignant neoplasm of abdomen|Disorder|true|false||ABDOMENnull|Abdomen problem|Finding|true|false||ABDOMENnull|Abdomen|Anatomy|true|false||ABDOMEN
null|Abdominal Cavity|Anatomy|true|false||ABDOMENnull|Obesity|Disorder|false|false||Obesenull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||softnull|Soft|Modifier|false|false||softnull|LRRC4B gene|Finding|true|false||HSMnull|Emotional tenderness|Finding|true|false||tenderness
null|Sore to touch|Finding|true|false||tendernessnull|Absence of Biallelic TCRgamma Deletion|Disorder|true|false||Abdnull|ABD (body structure)|Anatomy|true|false||Abd
null|Abdomen|Anatomy|true|false||Abdnull|Procedure on aorta|Procedure|true|false||aortanull|Chest+Abdomen>Aorta|Anatomy|true|false||aorta
null|Aorta|Anatomy|true|false||aortanull|Palpation|Procedure|true|false||palpationnull|Abdominal bruit|Finding|true|false||abdominal bruitsnull|Abdomen|Anatomy|true|false||abdominalnull|Abdominal (qualifier value)|Modifier|true|false||abdominalnull|Bruit|Finding|true|false||bruitsnull|All extremities|Anatomy|false|false||EXTREMITIES
null|Limb structure|Anatomy|false|false||EXTREMITIESnull|Femur|Anatomy|true|false||femoralnull|Bruit|Finding|true|false||bruitsnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false||SKIN
null|Skin and subcutaneous tissue disorders|Disorder|false|false||SKINnull|Skin Specimen Source Code|Finding|false|false||SKIN
null|Skin Specimen|Finding|false|false||SKINnull|Skin, Human|Anatomy|false|false||SKIN
null|Skin|Anatomy|false|false||SKINnull|Stasis dermatitis|Disorder|true|false||stasis dermatitisnull|Stasis|Finding|true|false||stasisnull|Dermatitis|Disorder|true|false||dermatitisnull|Ulcer|Finding|true|false||ulcersnull|Scar Tissue|Finding|true|false||scars
null|Cicatrix|Finding|true|false||scarsnull|Xanthoma|Disorder|true|false||xanthomasnull|null|Drug|false|false||PULSESnull|Physiologic pulse|Finding|false|false||PULSESnull|Pulse taking|Procedure|false|false||PULSESnull|Radial|Finding|false|false||radial
null|Circumpennate|Finding|false|false||radialnull|DSPP wt Allele|Finding|false|false||DPP
null|DSPP gene|Finding|false|false||DPPnull|Neurology speciality|Title|false|false||Neuronull|Neurologic (qualifier value)|Modifier|false|false||Neuronull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|Laboratory test finding|Lab|false|false||LABSnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Alanine Transaminase|Drug|false|false||ALT
null|Alanine Transaminase|Drug|false|false||ALTnull|Liposarcoma, well differentiated|Disorder|false|false||ALT
null|Atypical Lipoma|Disorder|false|false||ALTnull|null|Finding|false|false||ALT
null|Alternative Billing Concepts|Finding|false|false||ALT
null|GPT gene|Finding|false|false||ALTnull|Antibiotic Lock Therapy|Procedure|false|false||ALTnull|Southern Altai Language|Entity|false|false||ALTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||ASTnull|Atypical Spitz Nevus|Disorder|false|false||ASTnull|SLC17A5 wt Allele|Finding|false|false||AST
null|SLC17A5 gene|Finding|false|false||AST
null|GOT1 gene|Finding|false|false||ASTnull|Asterion|Anatomy|false|false||ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|Alkaline Phosphatase|Drug|false|false||AlkPhos
null|Alkaline Phosphatase|Drug|false|false||AlkPhosnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|lipase|Drug|false|false||Lipase
null|lipase|Drug|false|false||Lipase
null|lipase|Drug|false|false||Lipasenull|Lipase measurement|Procedure|false|false||Lipasenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MB
null|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MBnull|creatine kinase activity|Finding|false|false||CK-MBnull|Serum creatine phosphokinase MB isoenzyme measurement|Procedure|false|false||CK-MB
null|Creatine kinase MB measurement|Procedure|false|false||CK-MBnull|CD79A wt Allele|Finding|false|false||MB-1
null|CD79A gene|Finding|false|false||MB-1null|Blood calcium measurement|Procedure|false|false||BLOOD Calciumnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Plain chest X-ray|Procedure|false|false||CXRnull|Coronal (qualifier value)|Modifier|false|false||Frontalnull|Lateral|Modifier|false|false||lateralnull|View|Modifier|false|false||viewsnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Persistent|Time|false|false||persistentnull|Left costodiaphragmatic recess|Anatomy|false|false||left costophrenic anglenull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Costophrenic angle|Anatomy|false|false||costophrenic anglenull|Angular|Modifier|false|false||anglenull|Suggestive of|Finding|false|false||suggestive ofnull|Suggestive of|Finding|false|false||suggestivenull|Cicatrization|Finding|false|false||scarring
null|Cicatrix|Finding|false|false||scarringnull|Thickening of pleura|Disorder|false|false||pleural thickeningnull|Pleural Diseases|Disorder|false|false||pleuralnull|Pleura|Anatomy|false|false||pleuralnull|Pleural|Modifier|false|false||pleuralnull|Thickened|Finding|false|false||thickeningnull|Lung|Anatomy|false|false||lungsnull|Remote control command - Clear|Finding|false|false||clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|Limited (extensiveness)|Finding|false|false||limitsnull|Median Sternotomy|Procedure|false|false||Median sternotomynull|Median (qualifier value)|Modifier|false|false||Median
null|Midline (qualifier value)|Modifier|false|false||Mediannull|Statistical Median|LabModifier|false|false||Median
null|Population Median|LabModifier|false|false||Median
null|Sample Median|LabModifier|false|false||Mediannull|Sternotomy (procedure)|Procedure|false|false||sternotomynull|Bone Wires|Device|false|false||wiresnull|Mediastinum|Anatomy|false|false||mediastinalnull|Mediastinal|Modifier|false|false||mediastinalnull|Clip|Device|false|false||clipsnull|Admission Level of Care Code - Acute|Finding|true|false||acute
null|Acute - Triage Code|Finding|true|false||acutenull|acute|Time|true|false||acutenull|Cardiovascular disease+Pulmonary disease|Disorder|true|false||cardiopulmonarynull|Cardiopulmonary|Anatomy|true|false||cardiopulmonarynull|Process Pharmacologic Substance|Drug|true|false||processnull|Process (qualifier value)|Finding|true|false||processnull|bony process|Anatomy|true|false||processnull|Process|Phenomenon|true|false||processnull|Exercise|Finding|false|false||Exercisenull|Exercise Pain Management|Procedure|false|false||Exercisenull|Stress bismuth subsalicylate|Drug|false|false||Stress
null|Stress bismuth subsalicylate|Drug|false|false||Stressnull|Stress|Finding|false|false||Stressnull|W stress|Attribute|false|false||Stressnull|impression (attitude)|Finding|false|false||IMPRESSION
null|EKG impression|Finding|false|false||IMPRESSIONnull|atypia morphology|Finding|false|false||Atypicalnull|Atypical|Modifier|false|false||Atypicalnull|Sudden onset (contextual qualifier) (qualifier value)|Finding|false|false||sudden onset ofnull|Sudden onset (contextual qualifier) (qualifier value)|Finding|false|false||sudden onsetnull|Sudden onset (attribute)|Time|false|false||sudden onsetnull|Sudden (qualifier value)|Modifier|false|false||suddennull|Onset of (contextual qualifier)|Modifier|false|false||onset ofnull|Onset of (contextual qualifier)|Modifier|false|false||onsetnull|Age of Onset|LabModifier|false|false||onsetnull|Chest tightness|Finding|false|false||chest tightnessnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Tightness sensation quality|Modifier|false|false||tightnessnull|ST segment|Finding|false|false||ST segmentnull|Anatomical segmentation|Modifier|false|false||segmentnull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|IPSS-R Risk Category Low|Finding|false|false||low
null|IPSS Risk Category Low|Finding|false|false||low
null|low confidentiality|Finding|false|false||lownull|Low - MessageWaitingPriority|Modifier|false|false||low
null|low|Modifier|false|false||low
null|low exposure|Modifier|false|false||lownull|null|LabModifier|false|false||lownull|Workload|LabModifier|false|false||workloadnull|Rest|Finding|false|false||Restingnull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Systolic Hypertension|Disorder|false|false||systolic hypertensionnull|Systole|Finding|false|false||systolicnull|Hypertensive disease|Disorder|false|false||hypertensionnull|Blunted|Modifier|false|false||bluntednull|Hemodynamics|Finding|false|false||hemodynamicnull|hemodynamics (procedure)|Procedure|false|false||hemodynamicnull|response to exercise|Finding|false|false||response to exercisenull|Communication Response|Finding|false|false||response
null|Disease Response|Finding|false|false||response
null|Answer (statement)|Finding|false|false||responsenull|Response process|Subject|false|false||responsenull|Exercise|Finding|false|false||exercisenull|Exercise Pain Management|Procedure|false|false||exercisenull|ECHO protocol|Procedure|false|false||Echo
null|Extension for Community Healthcare Outcomes|Procedure|false|false||Echonull|Echo <Calopterygidae>|Entity|false|false||Echonull|Report (document)|Finding|false|false||reportnull|Reporting|Procedure|false|false||reportnull|null|Attribute|false|false||reportnull|Exercise|Finding|false|false||Exercisenull|Exercise Pain Management|Procedure|false|false||Exercisenull|ECHO protocol|Procedure|false|false||Echo
null|Extension for Community Healthcare Outcomes|Procedure|false|false||Echonull|Echo <Calopterygidae>|Entity|false|false||Echonull|impression (attitude)|Finding|false|false||IMPRESSION
null|EKG impression|Finding|false|false||IMPRESSIONnull|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group|Finding|false|false||Poor
null|Patient Condition Code - Poor|Finding|false|false||Poornull|Poverty|Subject|false|false||Poornull|Language Proficiency - Poor|Modifier|false|false||Poor
null|Specimen Quality - Poor|Modifier|false|false||Poor
null|Poor - grade|Modifier|false|false||Poor
null|Poor - qualifier|Modifier|false|false||Poornull|Functional Relationship|Finding|false|false||functional
null|Function (attribute)|Finding|false|false||functional
null|Functional|Finding|false|false||functionalnull|Exercise capacity|LabModifier|false|false||exercise capacitynull|Exercise|Finding|false|false||exercisenull|Exercise Pain Management|Procedure|false|false||exercisenull|Capacity|LabModifier|false|false||capacitynull|Equine Gonadotropins|Drug|false|false||ECG
null|Equine Gonadotropins|Drug|false|false||ECG
null|Equine Gonadotropins|Drug|false|false||ECGnull|Electrocardiogram image|Finding|false|false||ECG
null|Electrocardiogram|Finding|false|false||ECGnull|Electrocardiography|Procedure|false|false||ECGnull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|Absent|Finding|false|false||absence ofnull|Absence (morphologic abnormality)|Disorder|false|false||absencenull|Absent|Finding|false|false||absencenull|Evidence of (contextual qualifier)|Finding|false|false||evidence ofnull|Evidence|Finding|false|false||evidencenull|Induce (action)|Finding|false|false||induciblenull|Ischemia|Finding|false|false||ischemianull|Ischemia Procedure|Procedure|false|false||ischemianull|IPSS-R Risk Category Low|Finding|false|false||low
null|IPSS Risk Category Low|Finding|false|false||low
null|low confidentiality|Finding|false|false||lownull|Low - MessageWaitingPriority|Modifier|false|false||low
null|low|Modifier|false|false||low
null|low exposure|Modifier|false|false||lownull|null|LabModifier|false|false||lownull|Workload|LabModifier|false|false||workloadnull|Rest|Finding|false|false||Restingnull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Systolic Hypertension|Disorder|false|false||systolic hypertensionnull|Systole|Finding|false|false||systolicnull|Hypertensive disease|Disorder|false|false||hypertensionnull|Blunted|Modifier|false|false||bluntednull|Hemodynamics|Finding|false|false||hemodynamicnull|hemodynamics (procedure)|Procedure|false|false||hemodynamicnull|Communication Response|Finding|false|false||response
null|Disease Response|Finding|false|false||response
null|Answer (statement)|Finding|false|false||responsenull|Response process|Subject|false|false||responsenull|Physiological|Finding|false|false||physiologicnull|Stress bismuth subsalicylate|Drug|false|false||stress
null|Stress bismuth subsalicylate|Drug|false|false||stressnull|Stress|Finding|false|false||stressnull|W stress|Attribute|false|false||stressnull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|Laboratory test finding|Lab|false|false||LABSnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Phos <Photinae>|Entity|false|false||Phosnull|Infantile Neuroaxonal Dystrophy|Disorder|false|false||PLANnull|Treatment Plan|Finding|false|false||PLAN
null|Planned|Finding|false|false||PLAN
null|null|Finding|false|false||PLANnull|PMH - past medical history|Finding|false|false||pmh
null|Medical History|Finding|false|false||pmhnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Known|Modifier|false|false||knownnull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Coronary Artery Bypass Surgery|Procedure|false|false||CABGnull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Angina Pectoris|Finding|false|false||angina
null|null|Finding|false|false||anginanull|null|Attribute|false|false||anginanull|Hypertensive disease|Disorder|false|false||HTNnull|Chest Pain|Finding|false|false||chest painnull|null|Attribute|false|false||chest painnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Angina, Unstable|Disorder|false|false||crescendo anginanull|Crescendo|Drug|false|false||crescendo
null|Crescendo|Drug|false|false||crescendonull|Angina Pectoris|Finding|false|false||angina
null|null|Finding|false|false||anginanull|null|Attribute|false|false||anginanull|Chest Pain|Finding|false|false||Chest painnull|null|Attribute|false|false||Chest painnull|Chest problem|Finding|false|false||Chestnull|Chest|Anatomy|false|false||Chest
null|Anterior thoracic region|Anatomy|false|false||Chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|IPSS-R Risk Category High|Finding|false|false||high
null|Message Waiting Priority - High|Finding|false|false||high
null|high - ActExposureLevelCode|Finding|false|false||high
null|IPSS Risk Category High|Finding|false|false||high
null|High (finding)|Finding|false|false||highnull|Observation Value - High|Modifier|false|false||high
null|High|Modifier|false|false||high
null|Abnormally high|Modifier|false|false||highnull|Heart|Anatomy|false|false||coronarynull|Coronary|Modifier|false|false||coronarynull|Risk|Finding|false|false||risknull|Recent|Time|true|false||recentnull|CAT protein, human|Drug|true|false||cat
null|CAT protein, human|Drug|true|false||cat
null|Cat hair antigen|Drug|true|false||cat
null|Cat hair antigen|Drug|true|false||cat
null|Chloramphenicol O-Acetyltransferase|Drug|true|false||cat
null|Chloramphenicol O-Acetyltransferase|Drug|true|false||catnull|Truncus Arteriosus, Persistent|Disorder|true|false||catnull|CAT gene|Finding|true|false||cat
null|Cutaneous Assessment Tool|Finding|true|false||cat
null|Chloramphenicol Acetyl Transferase Gene|Finding|true|false||cat
null|catalase activity|Finding|true|false||cat
null|Chronic Obstructive Pulmonary Disease Assessment Test scale|Finding|true|false||catnull|allergy testing cat|Procedure|true|false||cat
null|X-Ray Computed Tomography|Procedure|true|false||cat
null|cytarabine/thioguanine protocol|Procedure|true|false||catnull|Cat (organism)|Entity|true|false||cat
null|Family Felidae|Entity|true|false||cat
null|Catalan language|Entity|true|false||cat
null|Felis catus|Entity|true|false||catnull|6 months|Time|true|false||6 monthsnull|month|Time|true|false||monthsnull|FBXW7 wt Allele|Finding|true|false||ago
null|FBXW7 gene|Finding|true|false||agonull|Disease|Disorder|true|false||diseasenull|FACT Complex|Drug|false|false||Fact
null|FACT Complex|Drug|false|false||Factnull|SSRP1 wt Allele|Finding|false|false||Fact
null|SUPT16H gene|Finding|false|false||Factnull|Foundation for the Accreditation of Cellular Therapy|Subject|false|false||Factnull|physical examination (physical finding)|Finding|false|false||physical examnull|Physical Examination|Procedure|false|false||physical examnull|physical examination (physical finding)|Finding|false|false||physical
null|Physical|Finding|false|false||physicalnull|Physical Examination|Procedure|false|false||physicalnull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Cardiac attachment|Finding|false|false||cardiacnull|Heart|Anatomy|false|false||cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||cardiacnull|Science of Etiology|Finding|false|false||cause
null|Etiology aspects|Finding|false|false||causenull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Impaired cognition|Disorder|false|false||cognitive impairmentnull|Cognitive|Finding|false|false||cognitivenull|Impaired health|Finding|false|false||impairment
null|Impaired|Finding|false|false||impairmentnull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Stenosis|Finding|false|false||stenosisnull|Stenosis <Pimeliinae>|Entity|false|false||stenosisnull|Stenosis Morphology|Modifier|false|false||stenosisnull|Echocardiography, Stress|Procedure|false|false||stress echonull|Stress bismuth subsalicylate|Drug|false|false||stress
null|Stress bismuth subsalicylate|Drug|false|false||stressnull|Stress|Finding|false|false||stressnull|W stress|Attribute|false|false||stressnull|Extension for Community Healthcare Outcomes|Procedure|false|false||echo
null|ECHO protocol|Procedure|false|false||echonull|Echo <Calopterygidae>|Entity|false|false||echonull|Functional Relationship|Finding|false|false||functional
null|Function (attribute)|Finding|false|false||functional
null|Functional|Finding|false|false||functionalnull|Congenital Abnormality|Disorder|false|false||abnormalitynull|Abnormality|Finding|false|false||abnormalitynull|Exertion|Finding|false|false||exertionnull|ECHO protocol|Procedure|true|false||ECHO
null|Extension for Community Healthcare Outcomes|Procedure|true|false||ECHOnull|Echo <Calopterygidae>|Entity|true|false||ECHOnull|Congenital Abnormality|Disorder|true|false||abnormalitiesnull|teratologic|Finding|true|false||abnormalitiesnull|Atypical chest pain|Finding|false|false||atypical chest painnull|atypia morphology|Finding|false|false||atypicalnull|Atypical|Modifier|false|false||atypicalnull|Chest Pain|Finding|false|false||chest painnull|null|Attribute|false|false||chest painnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Stress bismuth subsalicylate|Drug|false|false||stress
null|Stress bismuth subsalicylate|Drug|false|false||stressnull|Stress|Finding|false|false||stressnull|W stress|Attribute|false|false||stressnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Arylsulfatase A, human|Drug|false|false||ASA
null|Arylsulfatase A, human|Drug|false|false||ASA
null|aspirin|Drug|false|false||ASA
null|aspirin|Drug|false|false||ASAnull|ARSA gene|Finding|false|false||ASAnull|Plavix|Drug|false|false||plavix
null|Plavix|Drug|false|false||plavixnull|Hydroxymethylglutaryl-CoA Reductase Inhibitors|Drug|false|false||statin
null|Hydroxymethylglutaryl-CoA Reductase Inhibitors|Drug|false|false||statinnull|EEF1A2 gene|Finding|false|false||statinnull|3-hydroxy-3-methylglutaryl-coenzyme A reductase inhibitor (disposition)|Modifier|false|false||statinnull|nitrate ion|Drug|false|false||nitrate
null|nitrate ion|Drug|false|false||nitrate
null|Nitrate|Drug|false|false||nitrate
null|Nitrates|Drug|false|false||nitratenull|metoprolol|Drug|false|false||metoprolol
null|metoprolol|Drug|false|false||metoprololnull|In-House|Finding|false|false||in-housenull|House (environment)|Device|false|false||housenull|Home environment|Modifier|false|false||housenull|Telephone Number|Finding|true|false||tele
null|TCAP gene|Finding|true|false||telenull|Alarms (package insert)|Finding|true|false||alarmsnull|Alarm device|Device|true|false||alarmsnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Stress bismuth subsalicylate|Drug|false|false||stress
null|Stress bismuth subsalicylate|Drug|false|false||stressnull|Stress|Finding|false|false||stressnull|W stress|Attribute|false|false||stressnull|Follow-up status|Finding|false|false||follow-upnull|follow-up|Procedure|false|false||follow-upnull|Follow - dosing instruction imperative|Finding|false|false||follow
null|Follow|Finding|false|false||follownull|Followed by|Time|false|false||follownull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|Chronic - Admission Level of Care Code|Finding|false|false||CHRONICnull|Provision of recurring care for chronic illness|Procedure|false|false||CHRONICnull|chronic|Time|false|false||CHRONICnull|diastolic congestive heart failure|Disorder|false|false||Diastolic CHFnull|Diastole|Attribute|false|false||Diastolicnull|Congestive heart failure|Disorder|false|false||CHFnull|Choroidal fissure|Anatomy|false|false||CHFnull|Aspects of signs|Finding|true|false||signs
null|Physical findings|Finding|true|false||signsnull|Manufactured sign|Device|true|false||signsnull|Fluid Overload|Finding|true|false||fluid overload
null|Hypervolemia (finding)|Finding|true|false||fluid overloadnull|fluid - substance|Drug|true|false||fluid
null|Liquid substance|Drug|true|false||fluidnull|Fluid Specimen Code|Finding|true|false||fluidnull|Fluid behavior|Modifier|true|false||fluidnull|Current (present time)|Time|true|false||currentlynull|BaseLine dental cement|Drug|true|false||baselinenull|baseline - TableCellVerticalAlign|Finding|true|false||baselinenull|Baseline|LabModifier|true|false||baselinenull|Diuresis|Finding|true|false||diuresisnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Daily|Time|true|false||dailynull|Aspects of signs|Finding|true|false||signs
null|Physical findings|Finding|true|false||signsnull|Manufactured sign|Device|true|false||signsnull|Decompensation|Finding|true|false||decompensationnull|Diuresis|Finding|true|false||diuresisnull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||Diabetes
null|Diabetes|Disorder|false|false||Diabetes
null|Diabetes Mellitus|Disorder|false|false||Diabetesnull|Hospital Information Systems|Finding|false|false||HISSnull|In-House|Finding|false|false||in-housenull|House (environment)|Device|false|false||housenull|Home environment|Modifier|false|false||housenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|insulin, regular, human|Drug|false|false||insulin
null|Insulin [EPC]|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulinnull|INS gene|Finding|false|false||insulinnull|Insulin measurement|Procedure|false|false||insulinnull|GDC Regimen Terminology|Finding|false|false||regimennull|Treatment Protocols|Procedure|false|false||regimennull|Lantus|Drug|false|false||lantus
null|Lantus|Drug|false|false||lantusnull|Once a day, at bedtime|Time|false|false||QHSnull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|MEDICATION LIST|Finding|false|false||Medication listnull|Pharmaceutical Preparations|Drug|false|false||Medicationnull|medication - HL7 publishing domain|Finding|false|false||Medication
null|Medications|Finding|false|false||Medicationnull|List|Finding|false|false||list
null|Sequence Data Type|Finding|false|false||listnull|Accurate (qualifier value)|Modifier|false|false||accuratenull|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||completenull|Completion Status for valid values - Complete|Finding|false|false||complete
null|Data operation - complete|Finding|false|false||complete
null|Finish - dosing instruction imperative|Finding|false|false||completenull|Complete|Modifier|false|false||completenull|losartan potassium|Drug|false|false||Losartan Potassium
null|losartan potassium|Drug|false|false||Losartan Potassiumnull|losartan|Drug|false|false||Losartan
null|losartan|Drug|false|false||Losartannull|Potassium Drug Class|Drug|false|false||Potassium
null|Dietary Potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassiumnull|Potassium metabolic function|Finding|false|false||Potassiumnull|Potassium measurement|Procedure|false|false||Potassiumnull|Daily|Time|false|false||DAILYnull|aspirin|Drug|false|false||Aspirin
null|aspirin|Drug|false|false||Aspirinnull|Daily|Time|false|false||DAILYnull|carisoprodol|Drug|false|false||carisoprodol
null|carisoprodol|Drug|false|false||carisoprodolnull|Oral Dosage Form|Drug|false|false||Oralnull|Oral Route of Administration|Finding|false|false||Oral
null|Oral (intended site)|Finding|false|false||Oralnull|Oral cavity|Anatomy|false|false||Oralnull|Oral|Modifier|false|false||Oralnull|Once a day, at bedtime|Time|false|false||qhsnull|Spasm|Finding|false|false||spasm
null|KANTR gene|Finding|false|false||spasmnull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Once a day, at bedtime|Time|false|false||at bedtimenull|Once a day, at bedtime|Time|false|false||bedtime
null|Bedtime (qualifier value)|Time|false|false||bedtimenull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Spasm|Finding|false|false||muscle spasmnull|Muscle (organ)|Anatomy|false|false||muscle
null|Muscle Tissue|Anatomy|false|false||musclenull|Spasm|Finding|false|false||spasm
null|KANTR gene|Finding|false|false||spasmnull|pantoprazole|Drug|false|false||Pantoprazole
null|pantoprazole|Drug|false|false||Pantoprazolenull|Every twenty four hours|Time|false|false||Q24Hnull|trazodone|Drug|false|false||traZODONE
null|trazodone|Drug|false|false||traZODONEnull|acetaminophen / oxycodone|Drug|false|false||Oxycodone-Acetaminophennull|oxycodone|Drug|false|false||Oxycodone
null|oxycodone|Drug|false|false||Oxycodonenull|Oxycodone measurement|Procedure|false|false||Oxycodonenull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Tablet Dosage Form|Drug|false|false||TABnull|Tablet Dosing Unit|LabModifier|false|false||TABnull|Every eight hours|Time|false|false||Q8Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|atorvastatin|Drug|false|false||Atorvastatin
null|atorvastatin|Drug|false|false||Atorvastatinnull|Daily|Time|false|false||DAILYnull|nitroglycerin|Drug|false|false||Nitroglycerin
null|nitroglycerin|Drug|false|false||Nitroglycerinnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Chest Pain|Finding|false|false||chest painnull|null|Attribute|false|false||chest painnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|metoprolol succinate|Drug|false|false||Metoprolol Succinate
null|metoprolol succinate|Drug|false|false||Metoprolol Succinatenull|metoprolol|Drug|false|false||Metoprolol
null|metoprolol|Drug|false|false||Metoprololnull|succinate|Drug|false|false||Succinate
null|Succinates|Drug|false|false||Succinatenull|Daily|Time|false|false||DAILYnull|isosorbide mononitrate|Drug|false|false||Isosorbide Mononitrate
null|isosorbide mononitrate|Drug|false|false||Isosorbide Mononitratenull|isosorbide|Drug|false|false||Isosorbide
null|isosorbide|Drug|false|false||Isosorbidenull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Daily|Time|false|false||DAILYnull|clopidogrel|Drug|false|false||Clopidogrel
null|clopidogrel|Drug|false|false||Clopidogrelnull|Daily|Time|false|false||DAILYnull|fluticasone propionate|Drug|false|false||Fluticasone Propionate
null|fluticasone propionate|Drug|false|false||Fluticasone Propionatenull|fluticasone|Drug|false|false||Fluticasone
null|fluticasone|Drug|false|false||Fluticasonenull|propionate|Drug|false|false||Propionate
null|Propionates|Drug|false|false||Propionatenull|Puff Dosing Unit|LabModifier|false|false||PUFF
null|Picofarad|LabModifier|false|false||PUFFnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Units
null|Unit of Measure|LabModifier|false|false||Units
null|Unit|LabModifier|false|false||Unitsnull|Bedtime (qualifier value)|Time|false|false||Bedtime
null|Once a day, at bedtime|Time|false|false||Bedtimenull|insulin, regular, human|Drug|false|false||Insulin
null|Insulin [EPC]|Drug|false|false||Insulin
null|INS protein, human|Drug|false|false||Insulin
null|INS protein, human|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Insulin Drug Class|Drug|false|false||Insulin
null|Insulin Drug Class|Drug|false|false||Insulin
null|insulin, regular, human|Drug|false|false||Insulin
null|insulin, regular, human|Drug|false|false||Insulinnull|INS gene|Finding|false|false||Insulinnull|Insulin measurement|Procedure|false|false||Insulinnull|sliding scale|Procedure|false|false||Sliding Scalenull|Sliding|Finding|false|false||Slidingnull|Scale, LOINC Axis 5|Finding|false|false||Scale
null|Base Number|Finding|false|false||Scale
null|Scale - rank|Finding|false|false||Scalenull|Integumentary scale|Anatomy|false|false||Scalenull|Weight measurement scales|Device|false|false||Scalenull|Scaling|Event|false|false||Scalenull|Unit dose|LabModifier|false|false||Dose
null|Dosage|LabModifier|false|false||Dosenull|Override|Finding|false|false||Overridenull|Indication of (contextual qualifier)|Finding|false|false||Reasonnull|Levemir|Drug|false|false||Levemir
null|Levemir|Drug|false|false||Levemir
null|Levemir|Drug|false|false||Levemirnull|Once a day, at bedtime|Time|false|false||QHSnull|Diagnostic Service Section ID - Pharmacy|Finding|false|false||pharmacy
null|Pharmacy domain|Finding|false|false||pharmacynull|Pharmaceutical Services|Procedure|false|false||pharmacynull|Pharmacy facility|Device|false|false||pharmacynull|Pharmacy (field)|Title|false|false||pharmacynull|Pharmacy facility|Entity|false|false||pharmacynull|List|Finding|false|false||list
null|Sequence Data Type|Finding|false|false||listnull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|aspirin|Drug|false|false||Aspirin
null|aspirin|Drug|false|false||Aspirinnull|Daily|Time|false|false||DAILYnull|atorvastatin|Drug|false|false||Atorvastatin
null|atorvastatin|Drug|false|false||Atorvastatinnull|Daily|Time|false|false||DAILYnull|clopidogrel|Drug|false|false||Clopidogrel
null|clopidogrel|Drug|false|false||Clopidogrelnull|Daily|Time|false|false||DAILYnull|fluticasone propionate|Drug|false|false||Fluticasone Propionate
null|fluticasone propionate|Drug|false|false||Fluticasone Propionatenull|fluticasone|Drug|false|false||Fluticasone
null|fluticasone|Drug|false|false||Fluticasonenull|propionate|Drug|false|false||Propionate
null|Propionates|Drug|false|false||Propionatenull|Puff Dosing Unit|LabModifier|false|false||PUFF
null|Picofarad|LabModifier|false|false||PUFFnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Units
null|Unit of Measure|LabModifier|false|false||Units
null|Unit|LabModifier|false|false||Unitsnull|Bedtime (qualifier value)|Time|false|false||Bedtime
null|Once a day, at bedtime|Time|false|false||Bedtimenull|insulin, regular, human|Drug|false|false||Insulin
null|Insulin [EPC]|Drug|false|false||Insulin
null|INS protein, human|Drug|false|false||Insulin
null|INS protein, human|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Insulin Drug Class|Drug|false|false||Insulin
null|Insulin Drug Class|Drug|false|false||Insulin
null|insulin, regular, human|Drug|false|false||Insulin
null|insulin, regular, human|Drug|false|false||Insulinnull|INS gene|Finding|false|false||Insulinnull|Insulin measurement|Procedure|false|false||Insulinnull|sliding scale|Procedure|false|false||Sliding Scalenull|Sliding|Finding|false|false||Slidingnull|Scale, LOINC Axis 5|Finding|false|false||Scale
null|Base Number|Finding|false|false||Scale
null|Scale - rank|Finding|false|false||Scalenull|Integumentary scale|Anatomy|false|false||Scalenull|Weight measurement scales|Device|false|false||Scalenull|Scaling|Event|false|false||Scalenull|Unit dose|LabModifier|false|false||Dose
null|Dosage|LabModifier|false|false||Dosenull|Override|Finding|false|false||Overridenull|Indication of (contextual qualifier)|Finding|false|false||Reasonnull|Levemir|Drug|false|false||Levemir
null|Levemir|Drug|false|false||Levemir
null|Levemir|Drug|false|false||Levemirnull|Once a day, at bedtime|Time|false|false||QHSnull|Diagnostic Service Section ID - Pharmacy|Finding|false|false||pharmacy
null|Pharmacy domain|Finding|false|false||pharmacynull|Pharmaceutical Services|Procedure|false|false||pharmacynull|Pharmacy facility|Device|false|false||pharmacynull|Pharmacy (field)|Title|false|false||pharmacynull|Pharmacy facility|Entity|false|false||pharmacynull|List|Finding|false|false||list
null|Sequence Data Type|Finding|false|false||listnull|losartan potassium|Drug|false|false||Losartan Potassium
null|losartan potassium|Drug|false|false||Losartan Potassiumnull|losartan|Drug|false|false||Losartan
null|losartan|Drug|false|false||Losartannull|Potassium Drug Class|Drug|false|false||Potassium
null|Dietary Potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassiumnull|Potassium metabolic function|Finding|false|false||Potassiumnull|Potassium measurement|Procedure|false|false||Potassiumnull|Daily|Time|false|false||DAILYnull|nitroglycerin|Drug|false|false||Nitroglycerin
null|nitroglycerin|Drug|false|false||Nitroglycerinnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Chest Pain|Finding|false|false||chest painnull|null|Attribute|false|false||chest painnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|pantoprazole|Drug|false|false||Pantoprazole
null|pantoprazole|Drug|false|false||Pantoprazolenull|Every twenty four hours|Time|false|false||Q24Hnull|trazodone|Drug|false|false||traZODONE
null|trazodone|Drug|false|false||traZODONEnull|carisoprodol|Drug|false|false||carisoprodol
null|carisoprodol|Drug|false|false||carisoprodolnull|Oral Dosage Form|Drug|false|false||Oralnull|Oral Route of Administration|Finding|false|false||Oral
null|Oral (intended site)|Finding|false|false||Oralnull|Oral cavity|Anatomy|false|false||Oralnull|Oral|Modifier|false|false||Oralnull|Once a day, at bedtime|Time|false|false||qhsnull|Spasm|Finding|false|false||spasm
null|KANTR gene|Finding|false|false||spasmnull|metoprolol succinate|Drug|false|false||Metoprolol Succinate
null|metoprolol succinate|Drug|false|false||Metoprolol Succinatenull|metoprolol|Drug|false|false||Metoprolol
null|metoprolol|Drug|false|false||Metoprololnull|succinate|Drug|false|false||Succinate
null|Succinates|Drug|false|false||Succinatenull|Daily|Time|false|false||DAILYnull|acetaminophen / oxycodone|Drug|false|false||Oxycodone-Acetaminophennull|oxycodone|Drug|false|false||Oxycodone
null|oxycodone|Drug|false|false||Oxycodonenull|Oxycodone measurement|Procedure|false|false||Oxycodonenull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Tablet Dosage Form|Drug|false|false||TABnull|Tablet Dosing Unit|LabModifier|false|false||TABnull|Every eight hours|Time|false|false||Q8Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|isosorbide mononitrate|Drug|false|false||Isosorbide Mononitrate
null|isosorbide mononitrate|Drug|false|false||Isosorbide Mononitratenull|isosorbide|Drug|false|false||Isosorbide
null|isosorbide|Drug|false|false||Isosorbidenull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Daily|Time|false|false||DAILYnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Atypical chest pain|Finding|false|false||Atypical Chest Painnull|atypia morphology|Finding|false|false||Atypicalnull|Atypical|Modifier|false|false||Atypicalnull|Chest Pain|Finding|false|false||Chest Painnull|null|Attribute|false|false||Chest Painnull|Chest problem|Finding|false|false||Chestnull|Chest|Anatomy|false|false||Chest
null|Anterior thoracic region|Anatomy|false|false||Chestnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Confusion|Disorder|false|false||Confusednull|Precaution Code - Confused|Finding|false|false||Confused
null|Clouded consciousness|Finding|false|false||Confusednull|Sometimes|Time|false|false||sometimesnull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Coordination of Benefits - Independent|Finding|false|false||Independent
null|Religious Affiliation - Independent|Finding|false|false||Independent
null|Independence|Finding|false|false||Independent
null|Independently able|Finding|false|false||Independentnull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Chest Pain|Finding|false|false||chest painnull|null|Attribute|false|false||chest painnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|AML Lab Table|Finding|false|false||lab
null|LAT2 gene|Finding|false|false||lab
null|EWS Lab Table|Finding|false|false||labnull|Laboratory|Device|false|false||labnull|Labrador retriever|Entity|false|false||lab
null|Laboratory|Entity|false|false||labnull|Chest|Anatomy|false|false||chestsnull|Electrocardiogram image|Finding|false|false||EKG
null|Electrocardiogram|Finding|false|false||EKGnull|Electrocardiography|Procedure|false|false||EKGnull|Malignant neoplasm of heart|Disorder|true|false||heart
null|benign neoplasm of heart|Disorder|true|false||heartnull|HEART PROBLEM|Finding|true|false||heartnull|Chest>Heart|Anatomy|true|false||heart
null|Heart|Anatomy|true|false||heartnull|Attack (finding)|Finding|true|false||attack
null|Attack behavior|Finding|true|false||attacknull|Attack device|Device|true|false||attacknull|Exercise stress test|Procedure|false|false||stress test
null|Stress Test|Procedure|false|false||stress testnull|Stress bismuth subsalicylate|Drug|false|false||stress
null|Stress bismuth subsalicylate|Drug|false|false||stressnull|Stress|Finding|false|false||stressnull|W stress|Attribute|false|false||stressnull|Tests (qualifier value)|Finding|false|false||test
null|Testing|Finding|false|false||testnull|Laboratory Procedures|Procedure|false|false||testnull|Test - temporal region|Anatomy|false|false||testnull|Test Result|Lab|false|false||testnull|Test Dosing Unit|LabModifier|false|false||testnull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Patient Outcome - Worsening|Finding|true|false||worseningnull|Worsening (qualifier value)|Modifier|true|false||worseningnull|Coronary Artery Disease|Disorder|true|false||coronary artery disease
null|Coronary Arteriosclerosis|Disorder|true|false||coronary artery diseasenull|Coronary artery|Anatomy|true|false||coronary arterynull|Heart|Anatomy|true|false||coronarynull|Coronary|Modifier|true|false||coronarynull|Arteriopathic disease|Disorder|true|false||artery diseasenull|Arterial system|Anatomy|true|false||artery
null|Arteries|Anatomy|true|false||arterynull|Disease|Disorder|true|false||diseasenull|Chest Pain|Finding|false|false||chest painnull|null|Attribute|false|false||chest painnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Touching|Finding|false|false||touchingnull|Tactile|Modifier|false|false||touchingnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Usual|Modifier|true|false||typicalnull|Coronary Artery Disease|Disorder|true|false||coronary artery disease
null|Coronary Arteriosclerosis|Disorder|true|false||coronary artery diseasenull|Coronary artery|Anatomy|true|false||coronary arterynull|Heart|Anatomy|true|false||coronarynull|Coronary|Modifier|true|false||coronarynull|Arteriopathic disease|Disorder|true|false||artery diseasenull|Arterial system|Anatomy|true|false||artery
null|Arteries|Anatomy|true|false||arterynull|Disease|Disorder|true|false||diseasenull|Administration Method - Pain|Finding|true|false||pain
null|Pain|Finding|true|false||painnull|null|Attribute|true|false||painnull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Relate - vinyl resin|Drug|false|false||relatednull|Role Link Type - related|Finding|false|false||related
null|Related (finding)|Finding|false|false||relatednull|Definitely Related to Intervention|Modifier|false|false||related
null|Relationships|Modifier|false|false||relatednull|Musculoskeletal Pain|Finding|false|false||musculoskeletal painnull|Musculoskeletal|Finding|false|false||musculoskeletalnull|null|Attribute|false|false||musculoskeletalnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|MEDICATION LIST|Finding|false|false||medication listnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|List|Finding|false|false||list
null|Sequence Data Type|Finding|false|false||listnull|follow-up|Procedure|false|false||followupnull|Cardiologists|Subject|false|false||cardiologistnull|Further|Modifier|false|false||furthernull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions