CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Neurology speciality|Title|false|false||NEUROLOGYnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|amoxicillin|Drug|false|false||amoxicillin
null|amoxicillin|Drug|false|false||amoxicillinnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Chief complaint (finding)|Finding|false|false||Chief Complaintnull|Complaint (finding)|Finding|false|false||Complaintnull|null|Attribute|false|false||Complaintnull|Weakness|Finding|false|false||Weakness
null|Asthenia|Finding|false|false||Weaknessnull|Lethargy|Finding|false|false||lethargynull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|History of present illness (finding)|Finding|false|false||History of Present Illnessnull|null|Attribute|false|false||History of Present Illnessnull|Medical History|Finding|false|false||History ofnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Present illness|Finding|false|false||Present Illnessnull|Present|Finding|false|false||Present
null|Presentation|Finding|false|false||Presentnull|Illness (finding)|Finding|false|false||Illnessnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Transaction counts and value totals - year|Finding|false|false||year
null|Precision - year|Finding|false|false||yearnull|year|Time|false|false||yearnull|Old|Time|false|false||oldnull|Females|Subject|false|false||female
null|Woman|Subject|false|false||femalenull|Female, Self-Report|Modifier|false|false||female
null|Female Phenotype|Modifier|false|false||femalenull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Abdominal Pain|Finding|false|false|C0000726|abdominal painnull|Abdomen|Anatomy|false|false|C0000737;C1549543;C0030193|abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Administration Method - Pain|Finding|false|false|C0000726|pain
null|Pain|Finding|false|false|C0000726|painnull|null|Attribute|false|false||painnull|Anemia|Disorder|false|false||anemianull|Anemia <Anemiaceae>|Entity|false|false||anemianull|Recent|Time|false|false||recentnull|Saccharum officinale, sucrose, cane sugar, Homeopathic preparation|Drug|false|false||sucrose
null|Saccharum officinale, sucrose, cane sugar, Homeopathic preparation|Drug|false|false||sucrose
null|sucrose|Drug|false|false||sucrose
null|sucrose|Drug|false|false||sucrose
null|sucrose|Drug|false|false||sucrosenull|Infusion route|Finding|false|false||infusionnull|Infusion procedures|Procedure|false|false||infusionnull|Infusion reaction|Finding|false|false||infusion reactionnull|Infusion route|Finding|false|false||infusionnull|Infusion procedures|Procedure|false|false||infusionnull|Reaction|Finding|false|false||reactionnull|Mottling|Finding|false|false||mottlingnull|Abnormal color|Finding|false|false||discolorationnull|Foot|Anatomy|false|false||feetnull|Foot Unit of Length|LabModifier|false|false||feetnull|Steroids|Drug|false|false||steroids
null|Steroids|Drug|false|false||steroidsnull|Lethargy|Finding|false|false||lethargynull|Headache|Finding|false|false||headachenull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Quantity limited request - Records|Finding|false|false||records
null|Records|Finding|false|false||recordsnull|Query Quantity Unit - Records|Modifier|false|false||recordsnull|Aunt|Subject|false|false||Auntnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Much|Finding|false|false||muchnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Aunt|Subject|false|false||auntnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Recent|Time|false|false||recentlynull|Illness (finding)|Finding|true|false||illnessnull|Behavioral change|Finding|false|false||behavioral changenull|Behavior|Finding|false|false||behavioralnull|Changing|Finding|false|false||changenull|Change - procedure|Procedure|false|false||changenull|Delta (difference)|LabModifier|false|false||change
null|Changed status|LabModifier|false|false||changenull|Cold brand of chlorpheniramine-phenylpropanolamine|Drug|false|false||cold
null|Cold brand of chlorpheniramine-phenylpropanolamine|Drug|false|false||coldnull|Common Cold|Disorder|false|false||cold
null|Chronic Obstructive Airway Disease|Disorder|false|false||coldnull|Cold Sensation|Finding|false|false||coldnull|Cold Therapy|Procedure|false|false||coldnull|Cold Temperature|Phenomenon|false|false||coldnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|null|Finding|false|false||transfusionnull|Transfusion (procedure)|Procedure|false|false||transfusion
null|Blood Transfusion|Procedure|false|false||transfusionnull|Mandibular right first molar prosthesis|Device|false|false||30Pnull|Aunt|Subject|false|false||auntnull|Visit|Finding|false|false||visitnull|Endoglin, human|Drug|false|false||end
null|Endoglin, human|Drug|false|false||endnull|end - ActRelationshipCheckpoint|Finding|false|false||end
null|ENG gene|Finding|false|false||end
null|ENG wt Allele|Finding|false|false||endnull|Stop (qualifier value)|Time|false|false||endnull|End|Modifier|false|false||endnull|Infusion route|Finding|false|false||infusionnull|Infusion procedures|Procedure|false|false||infusionnull|Purple|Modifier|false|false||purplenull|Lower Extremity|Anatomy|false|false||lower extremitiesnull|Body Site Modifier - Lower|Anatomy|false|false|C2003888|lowernull|Lower (action)|Event|false|false|C1548802|lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|All extremities|Anatomy|false|false||extremities
null|Limb structure|Anatomy|false|false||extremitiesnull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|Tachycardia|Finding|false|false|C4037974;C0018787|heart racingnull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787|heart
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787|heartnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|heartnull|Chest>Heart|Anatomy|false|false|C0039231;C1561444;C0153957;C0153500;C0795691|heart
null|Heart|Anatomy|false|false|C0039231;C1561444;C0153957;C0153500;C0795691|heartnull|Racing - Production Class Code|Finding|false|false|C4037974;C0018787|racingnull|Racing animals|Entity|false|false||racingnull|Androgen Binding Protein|Drug|false|false||SBP
null|Androgen Binding Protein|Drug|false|false||SBPnull|CCHCR1 wt Allele|Finding|false|false||SBP
null|SHBG wt Allele|Finding|false|false||SBPnull|Systolic blood pressure measurement|Procedure|false|false||SBPnull|Systolic Pressure|Attribute|false|false||SBPnull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Quantity limited request - Records|Finding|false|false||records
null|Records|Finding|false|false||recordsnull|Query Quantity Unit - Records|Modifier|false|false||recordsnull|Shivering|Finding|false|false||shiveringnull|Eye|Anatomy|false|false|C5848506|eyesnull|null|Attribute|false|false|C0015392|eyesnull|Mottling|Finding|false|false||mottlednull|Hand|Anatomy|false|false||handsnull|Foot|Anatomy|false|false||feetnull|Foot Unit of Length|LabModifier|false|false||feetnull|Concern|Finding|false|false||concernnull|Respiratory distress|Finding|false|false||respiratory distressnull|Respiratory attachment|Finding|false|false||respiratory
null|respiratory|Finding|false|false||respiratory
null|null|Finding|false|false||respiratory
null|Respiratory specimen|Finding|false|false||respiratorynull|Respiratory rate|Attribute|false|false||respiratorynull|Emotional distress|Finding|false|false||distress
null|Distress|Finding|false|false||distressnull|Benadryl|Drug|false|false||Benadryl
null|Benadryl|Drug|false|false||Benadrylnull|hydrocortisone|Drug|false|false||hydrocortisone
null|hydrocortisone|Drug|false|false||hydrocortisone
null|hydrocortisone|Drug|false|false||hydrocortisonenull|Cortisol Measurement|Procedure|false|false||hydrocortisonenull|5 Hours|Time|false|false||5 hoursnull|Hour|Time|false|false||hoursnull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Lethargy|Finding|false|false||lethargicnull|Frequently|Time|false|false||frequentlynull|Able to sit up|Finding|false|false||able to sit upnull|Able to sit|Finding|false|false||able to sitnull|Able (qualifier value)|Finding|false|false||ablenull|Ability|Subject|false|false||ablenull|Does sit up|Finding|false|false||sit upnull|Does sit|Finding|false|false||sit
null|Sitting position|Finding|false|false||sit
null|HHAT gene|Finding|false|false||sit
null|SIT1 gene|Finding|false|false||sitnull|Walking (function)|Finding|false|false||walknull|Issue (document)|Finding|false|false||issue
null|Problem|Finding|false|false||issuenull|Issue (action)|Event|false|false||issuenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|BORNHOLM EYE DISEASE|Disorder|false|false||bednull|Bachelor of Education|Finding|false|false||bednull|Beds|Device|false|false||bednull|Patient Location - Bed|Modifier|false|false||bednull|Aunt|Subject|false|false||auntnull|Still|Disorder|false|false||stillnull|Headache|Finding|false|false||headachenull|null|Finding|false|false||transfusionnull|Transfusion (procedure)|Procedure|false|false||transfusion
null|Blood Transfusion|Procedure|false|false||transfusionnull|Place - dosing instruction imperative|Finding|false|false||placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|Characteristics|Modifier|false|false||characteristicnull|Aunt|Subject|false|false||auntnull|Acetaminophen [EPC]|Drug|false|false||acetaminophen
null|acetaminophen|Drug|false|false||acetaminophen
null|acetaminophen|Drug|false|false||acetaminophennull|Acetaminophen measurement|Procedure|false|false||acetaminophennull|Water Specimen|Drug|false|false||water
null|water|Drug|false|false||water
null|water|Drug|false|false||waternull|Water - Specimen Source Codes|Finding|false|false||waternull|Hydrotherapy|Procedure|false|false||waternull|Sleep brand of diphenhydramine hydrochloride|Drug|false|false||sleep
null|Sleep brand of diphenhydramine hydrochloride|Drug|false|false||sleepnull|Sleep|Finding|false|false||sleepnull|next - HtmlLinkType|Finding|false|false||nextnull|Following|Time|false|false||next
null|Then|Time|false|false||nextnull|Adjacent|Modifier|false|false||nextnull|Few hours|Time|false|false||few hoursnull|Hour|Time|false|false||hoursnull|Awake (finding)|Finding|false|false||awakenull|Awakening (time frame)|Time|false|false||awakenull|Several|LabModifier|false|false||severalnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Bathroom|Device|false|false||bathroom
null|Toilet Facilities|Device|false|false||bathroomnull|Then - dosing instruction fragment|Finding|false|false||Thennull|Then|Time|false|false||Thennull|Late|Time|false|false||laternull|Late|Time|false|false||laternull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Aunt|Subject|false|false||auntnull|Worried|Finding|false|false||worriednull|Able (qualifier value)|Finding|false|false||ablenull|Ability|Subject|false|false||ablenull|Headache|Finding|false|false||headachenull|Drowsiness|Finding|false|false||sleepynull|Processing type - Evaluation|Finding|false|false||evaluationnull|Evaluation procedure|Procedure|false|false||evaluation
null|Evaluation|Procedure|false|false||evaluationnull|Drowsiness|Finding|false|false||drowsynull|Authorization Mode - Voice|Finding|false|false||voice
null|Voice G-code|Finding|false|false||voice
null|Voice|Finding|false|false||voicenull|TelecommunicationCapabilities - voice|Modifier|false|false||voicenull|Alert brand of caffeine|Drug|false|false||alert
null|Alert brand of caffeine|Drug|false|false||alertnull|Mentally alert|Finding|false|false||alert
null|Consciousness clear|Finding|false|false||alert
null|Alert note|Finding|false|false||alert
null|Alert|Finding|false|false||alertnull|null|Attribute|false|false||alertnull|Oriented to place|Finding|false|false||orientednull|Orientation, Spatial|Modifier|false|false||orientednull|Consistent with|Finding|false|false|C4266572;C0015392;C0700042|consistentnull|Carcinoma in situ of eye|Disorder|false|false|C4266572;C0015392;C0700042|eye
null|Disorder of eye|Disorder|false|false|C4266572;C0015392;C0700042|eyenull|Eye - Specimen Source Code|Finding|false|false|C4266572;C0015392;C0700042|eye
null|Eye problem|Finding|false|false|C4266572;C0015392;C0700042|eye
null|Eye Specimen|Finding|false|false|C4266572;C0015392;C0700042|eyenull|Head>Eye|Anatomy|false|false|C1550636;C1546630;C0262477;C0016385;C0154094;C0015397;C0332290|eye
null|Eye|Anatomy|false|false|C1550636;C1546630;C0262477;C0016385;C0154094;C0015397;C0332290|eye
null|Orbital region|Anatomy|false|false|C1550636;C1546630;C0262477;C0016385;C0154094;C0015397;C0332290|eyenull|Cardiac Flutter|Finding|false|false|C4266572;C0015392;C0700042|flutteringnull|Pupil|Anatomy|false|false|C4722408|pupilsnull|Reactive to light|Finding|false|false||reactive to lightnull|Reactive Therapy|Procedure|false|false|C0034121|reactivenull|Reactive|Modifier|false|false||reactivenull|TNFSF14 protein, human|Drug|false|false||light
null|TNFSF14 protein, human|Drug|false|false||lightnull|Light - subjective measurement|Finding|false|false||light
null|TNFSF14 wt Allele|Finding|false|false||light
null|TNFSF14 gene|Finding|false|false||light
null|Light color|Finding|false|false||lightnull|Phototherapy|Procedure|false|false||lightnull|Light|Phenomenon|false|false||lightnull|Light (qualifier)|Modifier|false|false||lightnull|Extraocular eye movement|Finding|false|false|C4266572;C0015392;C0700042|extraocular eye movementsnull|Extraocular|Finding|false|false|C4266572;C0015392;C0700042|extraocularnull|Eye Movements|Finding|false|false|C4266572;C0015392;C0700042|eye movementsnull|Carcinoma in situ of eye|Disorder|false|false|C4266572;C0015392;C0700042|eye
null|Disorder of eye|Disorder|false|false|C4266572;C0015392;C0700042|eyenull|Eye - Specimen Source Code|Finding|false|false|C4266572;C0015392;C0700042|eye
null|Eye problem|Finding|false|false|C4266572;C0015392;C0700042|eye
null|Eye Specimen|Finding|false|false|C4266572;C0015392;C0700042|eyenull|Head>Eye|Anatomy|false|false|C1550636;C1546630;C0262477;C0702182;C0241886;C0154094;C0015397;C0026649;C0015413|eye
null|Eye|Anatomy|false|false|C1550636;C1546630;C0262477;C0702182;C0241886;C0154094;C0015397;C0026649;C0015413|eye
null|Orbital region|Anatomy|false|false|C1550636;C1546630;C0262477;C0702182;C0241886;C0154094;C0015397;C0026649;C0015413|eyenull|Movement|Finding|false|false|C4266572;C0015392;C0700042|movementsnull|Full|Modifier|false|false||fullnull|Focal|Modifier|false|false||focalnull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|AML Lab Table|Finding|false|false||Lab
null|LAT2 gene|Finding|false|false||Lab
null|EWS Lab Table|Finding|false|false||Labnull|Laboratory|Device|false|false||Labnull|Labrador retriever|Entity|false|false||Lab
null|Laboratory|Entity|false|false||Labnull|Work|Event|false|false||worknull|Leukocytes|Anatomy|false|false||WBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|sodium bicarbonate|Drug|false|false||bicarb
null|sodium bicarbonate|Drug|false|false||bicarbnull|Ferritin|Drug|false|false||Ferritin
null|Ferritin|Drug|false|false||Ferritin
null|Ferritin|Drug|false|false||Ferritinnull|Ferritin measurement|Procedure|false|false||Ferritinnull|Carbon dioxide measurement, partial pressure|Procedure|false|false||PCO2null|Carbon dioxide, partial pressure|Lab|false|false||PCO2null|Leukocytes|Anatomy|false|false||WBCnull|Monocytes|Anatomy|false|false|C1521746;C0863146;C0337438;C0202202|monocytesnull|glucose|Drug|false|false||glucose
null|glucose|Drug|false|false||glucose
null|glucose|Drug|false|false||glucosenull|Glucose measurement|Procedure|false|false|C0026473|glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||glucosenull|Proteins|Drug|false|false||protein
null|Proteins|Drug|false|false||proteinnull|Protein Info|Finding|false|false|C0026473|proteinnull|Protein measurement|Procedure|false|false|C0026473|proteinnull|Yellow color (finding)|Finding|true|false|C0026473|xanthochromianull|tocilizumab|Drug|false|false||MRA
null|tocilizumab|Drug|false|false||MRA
null|tocilizumab|Drug|false|false||MRAnull|Magnetic Resonance Angiography|Procedure|false|false||MRAnull|MRI-Based Angiogram|Lab|false|false||MRAnull|MRV|Drug|false|false||MRV
null|MRV|Drug|false|false||MRVnull|Thrombus|Finding|true|false||thrombus
null|Blood Clot|Finding|true|false||thrombusnull|Thrombus <Thrombidae>|Entity|true|false||thrombusnull|Thrombosis|Finding|false|false||thrombosisnull|Further|Modifier|false|false||furthernull|Disease Management|Procedure|false|false||managementnull|Management Occupations|Subject|false|false||managementnull|Management procedure|Event|false|false||management
null|Administration occupational activities|Event|false|false||managementnull|Published Interview|Finding|false|false||interviewnull|Interview|Event|false|false||interviewnull|Much|Finding|false|false||muchnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Feel Tired question|Finding|false|false||tired
null|Fatigue|Finding|false|false||tired
null|Feeling tired|Finding|false|false||tirednull|Eye|Anatomy|false|false|C5848506|eyesnull|null|Attribute|false|false|C0015392|eyesnull|Sexual Orientation - Questioning|Finding|false|false||questioningnull|Gender Questioning|Subject|false|false||questioningnull|Headache|Finding|false|false||headachenull|Photophobia|Finding|false|false||photophobianull|Unable|Finding|false|false||unablenull|Participate|Event|false|false||participatenull|Sexual Orientation - Questioning|Finding|false|false||questioningnull|Gender Questioning|Subject|false|false||questioningnull|Often - answer to question|Finding|false|false||oftennull|Frequently|Time|false|false||oftennull|Weepiness|Finding|false|false||tearfulnull|Hardness|Modifier|false|false||hardnull|Indirect exposure mechanism - Father|Finding|false|false||father
null|Relationship - Father|Finding|false|false||father
null|Father - courtesy title|Finding|false|false||fathernull|Father (person)|Subject|false|false||fathernull|Aunt|Subject|false|false||auntnull|Medical History|Finding|true|false||history ofnull|History of present illness (finding)|Finding|true|false||history
null|History of previous events|Finding|true|false||history
null|Historical aspects qualifier|Finding|true|false||history
null|Medical History|Finding|true|false||history
null|Concept History|Finding|true|false||historynull|History|Subject|false|false||historynull|Seizures|Finding|true|false||seizuresnull|Central Nervous System|Anatomy|false|false||CNSnull|Clinical Nurse Specialists|Subject|false|false||CNSnull|Certified Nurse Specialist|Title|false|false||CNSnull|Staphylococcus, coagulase negative (organism)|Entity|true|false||CNSnull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|Brain Concussion|Disorder|false|false||concussionnull|year|Time|false|false||yearsnull|Old|Time|false|false||oldnull|PMH - past medical history|Finding|false|false||Past Medical History
null|Medical History|Finding|false|false||Past Medical Historynull|Medical History|Finding|false|false||Medical Historynull|Medical referral type|Finding|false|false||Medical
null|Medical|Finding|false|false||Medical
null|Medical school type|Finding|false|false||Medicalnull|Medical service|Procedure|false|false||Medicalnull|Medical History|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|History of present illness (finding)|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Anemia|Disorder|false|false||Anemianull|Anemia <Anemiaceae>|Entity|false|false||Anemianull|Social and personal history|Finding|false|false||Social History
null|Social History|Finding|false|false||Social Historynull|Social|Finding|false|false||Socialnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Family Medical History|Finding|false|false||Family Historynull|Entity Name Part Type - family|Finding|false|false||Family
null|Last Name|Finding|false|false||Family
null|Living Arrangement - Family|Finding|false|false||Family
null|Family (taxonomic)|Finding|false|false||Family
null|Family Collection|Finding|false|false||Familynull|Family|Subject|false|false||Familynull|History of present illness (finding)|Finding|false|true||History
null|History of previous events|Finding|false|true||History
null|Historical aspects qualifier|Finding|false|true||History
null|Medical History|Finding|false|true||History
null|Concept History|Finding|false|true||Historynull|History|Subject|false|false||Historynull|Relationship - Mother|Finding|false|false||Mothernull|Mother (person)|Subject|false|false||Mothernull|Celiac Disease|Disorder|false|false||celiac diseasenull|CTLA4 gene|Finding|false|false||celiac diseasenull|Celiac Disease|Disorder|false|false||celiacnull|Disease|Disorder|false|false||diseasenull|Hypothyroidism, Autoimmune|Disorder|false|false||autoimmune hypothyroidismnull|Autoimmune reaction|Finding|false|false||autoimmune
null|Autoimmune|Finding|false|false||autoimmunenull|Hypothyroidism|Disorder|false|false||hypothyroidismnull|Diffuse alveolar damage|Disorder|false|false||Dadnull|Disability Assessment for Dementia Questionnaire|Finding|false|false||Dadnull|Healthy|Modifier|false|false||healthynull|Cousin|Subject|false|false||cousinnull|Seizures|Finding|false|false||seizuresnull|physical examination (physical finding)|Finding|false|false||Physical Examnull|Physical Examination|Procedure|false|false||Physical Examnull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||Generalnull|General medical service|Procedure|false|false||Generalnull|Generalized|Modifier|false|false||Generalnull|Infrequent|Time|false|false||occasionalnull|Eye lid|Anatomy|false|false|C0154094;C0015397|eye lidnull|Carcinoma in situ of eye|Disorder|false|false|C4266572;C0015392;C0700042;C2706046|eye
null|Disorder of eye|Disorder|false|false|C4266572;C0015392;C0700042;C2706046|eyenull|Eye - Specimen Source Code|Finding|false|false|C4266572;C0015392;C0700042|eye
null|Eye problem|Finding|false|false|C4266572;C0015392;C0700042|eye
null|Eye Specimen|Finding|false|false|C4266572;C0015392;C0700042|eyenull|Head>Eye|Anatomy|false|false|C1550636;C1546630;C0262477;C0154094;C0015397;C0016385|eye
null|Eye|Anatomy|false|false|C1550636;C1546630;C0262477;C0154094;C0015397;C0016385|eye
null|Orbital region|Anatomy|false|false|C1550636;C1546630;C0262477;C0154094;C0015397;C0016385|eyenull|Cardiac Flutter|Finding|false|false|C4266572;C0015392;C0700042|flutteringnull|Benign neoplasm of the lip|Disorder|false|false|C0023759|lip
null|Lymphoid interstitial pneumonia|Disorder|false|false|C0023759|lipnull|SMG1 wt Allele|Finding|false|false|C0023759|lip
null|SMG1 gene|Finding|false|false|C0023759|lipnull|Lip structure|Anatomy|false|false|C0153932;C0264511;C1846919;C3889123;C0362076|lipnull|Movement|Finding|false|false||movementsnull|Infrequent|Time|false|false||occasionalnull|Bradykinesia|Finding|false|false||slow movementsnull|Slow|Modifier|false|false||slownull|Movement|Finding|false|false|C0018670;C0152336|movementsnull|Problems with head|Disorder|false|false|C0018670;C0152336;C0023759|headnull|Procedure on head|Procedure|false|false|C0018670;C0152336|headnull|Structure of head of caudate nucleus|Anatomy|false|false|C0876917;C0362076;C0026649|head
null|Head|Anatomy|false|false|C0876917;C0362076;C0026649|headnull|Head Device|Device|false|false||headnull|Side|Modifier|false|false||sidenull|Side|Modifier|false|false||sidenull|HEENT|Anatomy|false|false||HEENTnull|Physical trauma|Disorder|true|false||trauma
null|Traumatic injury|Disorder|true|false||trauma
null|Trauma|Disorder|true|false||traumanull|Trauma assessment and care|Procedure|true|false||traumanull|Trauma, nursing specialty|Title|false|false||traumanull|trauma qualifier|Modifier|false|false||traumanull|jaundice|Finding|true|false||jaundice
null|Icterus|Finding|true|false||jaundice
null|yellow skin or eyes (symptom)|Finding|true|false||jaundicenull|Lesion|Finding|true|false|C0521367|lesionsnull|Oropharyngeal|Anatomy|false|false|C0221198|oropharynxnull|Pulmonary ventilator management|Procedure|false|false||Pulmnull|Hereditary Multiple Exostoses|Disorder|false|false||Extnull|EXT1 wt Allele|Finding|false|false||Ext
null|EXT1 gene|Finding|false|false||Extnull|Clammy skin|Finding|false|false||clammynull|Feels warm|Finding|false|false||warmnull|warming process|Phenomenon|false|false||warmnull|Eruption of skin (disorder)|Disorder|true|false||rashnull|Skin rash|Finding|true|false||rash
null|Eruptions|Finding|true|false||rash
null|Exanthema|Finding|true|false||rashnull|Neurologic (qualifier value)|Modifier|false|false||Neurologicnull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Frequently|Time|false|false||frequentlynull|Feeling upset|Finding|false|false||upsetnull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Weepiness|Finding|false|false||tearfulnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Ablepharon|Disorder|false|false|C0015392|Eyes opennull|Eye|Anatomy|false|false|C0266574;C5848506|Eyesnull|null|Attribute|false|false|C0015392|Eyesnull|Open|Modifier|false|false||opennull|Authorization Mode - Voice|Finding|false|false||voice
null|Voice G-code|Finding|false|false||voice
null|Voice|Finding|false|false||voicenull|TelecommunicationCapabilities - voice|Modifier|false|false||voicenull|Full|Modifier|false|false||fullnull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|MDF Attribute Type - Name|Finding|true|false||name
null|Person Name|Finding|true|false||name
null|Name|Finding|true|false||namenull|Name (property) (qualifier value)|Modifier|false|false||namenull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Feel Tired question|Finding|false|false||tired
null|Fatigue|Finding|false|false||tired
null|Feeling tired|Finding|false|false||tirednull|Unable|Finding|false|false||unablenull|Provide (product)|Drug|false|false||providenull|Providing (action)|Event|false|false||providenull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Speech|Finding|false|false||Speechnull|Speech assessment|Procedure|false|false||Speechnull|Spontaneous|Finding|true|false||spontaneousnull|Speech|Finding|false|false||speechnull|Speech assessment|Procedure|false|false||speechnull|system output|Finding|true|false||outputnull|Measurement of fluid output|Procedure|true|false||outputnull|LITAF gene|Finding|false|false||simplenull|Simple|Modifier|false|false||simplenull|Open|Modifier|false|false||opennull|Eye|Anatomy|false|false|C5848506|eyesnull|null|Attribute|false|false|C0015392|eyesnull|hoist [device]|Device|false|false||liftnull|Lifting|Event|false|false|C1140621|liftnull|Leg|Anatomy|false|false|C0206244;C5781420|legsnull|null|Attribute|false|false|C1140621|legsnull|Able (qualifier value)|Finding|false|false||ablenull|Ability|Subject|false|false||ablenull|MDF Attribute Type - Name|Finding|false|false||name
null|Person Name|Finding|false|false||name
null|Name|Finding|false|false||namenull|Name (property) (qualifier value)|Modifier|false|false||namenull|Key - HL7UpdateMode|Finding|false|false||key
null|Key - value|Finding|false|false||keynull|Feathers (allergen)|Drug|false|false|C0015731;C1744713|feathernull|null|Anatomy|false|false|C3486460|feather
null|Feathers|Anatomy|false|false|C3486460|feathernull|Cerebrovascular accident|Disorder|false|false|C2340164|strokenull|Stroke (heart beat)|Finding|false|false|C2340164|strokenull|Heart Diseases|Disorder|false|false|C2340164|cardnull|Card (document)|Finding|false|false|C2340164|cardnull|CaRD Regimen|Procedure|false|false|C2340164|cardnull|Stratum radiatum|Anatomy|false|false|C1720594;C5202809;C0018799;C0038454;C5977286;C3275277|cardnull|Card - Blister Pack|Device|false|false||cardnull|cardiology (field)|Title|false|false||cardnull|Then - dosing instruction fragment|Finding|false|false|C2340164|thennull|Then|Time|false|false||thennull|Eye|Anatomy|false|false|C5848506|eyesnull|null|Attribute|false|false|C0015392|eyesnull|Firstly|Modifier|false|false||firstnull|First (number)|LabModifier|false|false||firstnull|Sentence|Finding|false|false||sentencenull|Cerebrovascular accident|Disorder|false|false|C2340164|strokenull|Stroke (heart beat)|Finding|false|false|C2340164|strokenull|Heart Diseases|Disorder|false|false|C2340164|cardnull|Card (document)|Finding|false|false|C2340164|cardnull|CaRD Regimen|Procedure|false|false|C2340164|cardnull|Stratum radiatum|Anatomy|false|false|C0038454;C3275277;C1720594;C5977286;C0018799;C5202809|cardnull|Card - Blister Pack|Device|false|false||cardnull|cardiology (field)|Title|false|false||cardnull|Then - dosing instruction fragment|Finding|false|false|C2340164|thennull|Then|Time|false|false||thennull|More|LabModifier|false|false||morenull|Eye|Anatomy|false|false|C5848506|eyesnull|null|Attribute|false|false|C0015392|eyesnull|Cerebrovascular accident|Disorder|false|false|C2340164|strokenull|Stroke (heart beat)|Finding|false|false|C2340164|strokenull|Heart Diseases|Disorder|false|false|C2340164|cardnull|Card (document)|Finding|false|false|C2340164|cardnull|CaRD Regimen|Procedure|false|false|C2340164|cardnull|Stratum radiatum|Anatomy|false|false|C3275277;C0018799;C0038454;C5977286;C5202809|cardnull|Card - Blister Pack|Device|false|false||cardnull|cardiology (field)|Title|false|false||cardnull|Picture|Device|false|false||picture
null|photograph|Device|false|false||picturenull|Further|Modifier|false|false||furthernull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Neoplasm of uncertain or unknown behavior of cranial nerves|Disorder|false|false|C0010268;C0037303;C0027740|Cranial Nerves
null|Benign neoplasm of cranial nerves|Disorder|false|false|C0010268;C0037303;C0027740|Cranial Nervesnull|Cranial Nerves|Anatomy|false|false|C0004992;C0496937|Cranial Nervesnull|Bone structure of cranium|Anatomy|false|false|C0004992;C0496937|Cranialnull|Cranial|Modifier|false|false||Cranialnull|Nerve|Anatomy|false|false|C0004992;C0496937|Nervesnull|Pupil|Anatomy|false|false||Pupilsnull|Nystagmus|Disorder|false|false||nystagmusnull|Social confrontation skill|Finding|false|false||confrontationnull|Confrontation visual field test|Procedure|false|false||confrontation
null|Confrontation|Procedure|false|false||confrontationnull|Ophthalmoscopy|Procedure|false|false||Fundoscopic examnull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Papilledema|Disorder|true|false||papilledemanull|Exudate|Finding|false|false||exudatesnull|Hemorrhage|Finding|false|false||hemorrhagesnull|Roman numeral VII|Finding|false|false|C2338708;C3496273;C3496274|VIInull|Lamina VII of gray matter of spinal cord|Anatomy|false|false|C0445385|VII
null|lobule VII|Anatomy|false|false|C0445385|VII
null|layer VII (Cajal)|Anatomy|false|false|C0445385|VIInull|Facial Paresis|Disorder|true|false|C0015450|facial droopnull|Unilateral facial palsy|Finding|true|false|C0015450|facial droopnull|Face|Anatomy|false|false|C0427055;C4022719|facialnull|Facial|Modifier|false|false||facialnull|Face|Anatomy|false|false||facialnull|Facial|Modifier|false|false||facialnull|Set of muscles|Anatomy|false|false||musculaturenull|Symmetric Relationship|Finding|false|false||symmetric
null|Symmetrical|Finding|false|false||symmetricnull|Grimaces|Finding|false|false||grimacenull|Roman numeral VIII|Finding|false|false|C2327388;C0228488|VIII
null|COX8A gene|Finding|false|false|C2327388;C0228488|VIIInull|Lamina VIII of gray matter of spinal cord|Anatomy|false|false|C0445599;C1413661|VIII
null|Cerebellar pyramis|Anatomy|false|false|C0445599;C1413661|VIIInull|outcomes otolaryngology hearing|Finding|false|false||Hearing
null|Hearing finding|Finding|false|false||Hearing
null|Hearing|Finding|false|false||Hearingnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Palate|Anatomy|false|false||Palatenull|Benign neoplasm of tongue|Disorder|false|false|C1660780;C0040408|Tonguenull|Procedure on tongue|Procedure|false|false|C0040408;C1660780|Tonguenull|Tongue|Anatomy|false|false|C0872394;C0153933|Tonguenull|midline cell component|Anatomy|false|false|C0153933;C0872394|midlinenull|Midline (qualifier value)|Modifier|false|false||midlinenull|motor movement|Finding|false|false||Motornull|Motor Device|Device|false|false||Motornull|Bulk (conceptual)|Drug|false|false||bulk
null|Dietary Fiber|Drug|false|false||bulknull|Alveolar rhabdomyosarcoma|Disorder|false|false|C0446516|armsnull|Adherence to Refills and Medications Scale|Finding|false|false|C0446516|arms
null|KIDINS220 gene|Finding|false|false|C0446516|armsnull|Upper arm|Anatomy|false|false|C5575339;C2681631;C0206655;C5782111|armsnull|null|Attribute|false|false|C0446516|armsnull|Alveolar rhabdomyosarcoma|Disorder|false|false|C0446516|armsnull|Adherence to Refills and Medications Scale|Finding|false|false|C0446516|arms
null|KIDINS220 gene|Finding|false|false|C0446516|armsnull|Upper arm|Anatomy|false|false|C0206655;C5575339;C2681631;C5782111;C0362076|armsnull|null|Attribute|false|false|C0446516|armsnull|Problems with head|Disorder|false|false|C0018670;C0152336;C0446516|headnull|Procedure on head|Procedure|false|false|C0018670;C0152336|headnull|Structure of head of caudate nucleus|Anatomy|false|false|C0362076;C5575339;C2681631;C0206655;C0876917|head
null|Head|Anatomy|false|false|C0362076;C5575339;C2681631;C0206655;C0876917|headnull|Head Device|Device|false|false||headnull|Alveolar rhabdomyosarcoma|Disorder|false|false|C0018670;C0152336;C0446516|armsnull|Adherence to Refills and Medications Scale|Finding|false|false|C0446516;C0018670;C0152336|arms
null|KIDINS220 gene|Finding|false|false|C0446516;C0018670;C0152336|armsnull|Upper arm|Anatomy|false|false|C5575339;C2681631;C0206655;C5782111|armsnull|null|Attribute|false|false|C0446516|armsnull|Slow|Modifier|false|false||slowlynull|FANCONI ANEMIA, COMPLEMENTATION GROUP E|Disorder|false|false|C0015450;C4266571|facenull|FANCE wt Allele|Finding|false|false|C0015450;C4266571|face
null|FANCE gene|Finding|false|false|C0015450;C4266571|face
null|ELOVL6 gene|Finding|false|false|C0015450;C4266571|facenull|Head>Face|Anatomy|false|false|C1423759;C2828055;C1414531;C3159311;C2346952;C3160739|face
null|Face|Anatomy|false|false|C1423759;C2828055;C1414531;C3159311;C2346952;C3160739|facenull|Face (spatial concept)|Modifier|false|false||facenull|Slow|Modifier|false|false||slowlynull|Drops - Drug Form|Drug|false|false||dropsnull|Drop Dosing Unit|LabModifier|false|false||dropsnull|BORNHOLM EYE DISEASE|Disorder|false|false|C0015450;C4266571|bednull|Bachelor of Education|Finding|false|false|C0015450;C4266571|bednull|Beds|Device|false|false||bednull|Patient Location - Bed|Modifier|false|false||bednull|Disease Controlled|Finding|false|false||controlled
null|Control function|Finding|false|false||controlled
null|Controlled mark|Finding|false|false||controllednull|Alveolar rhabdomyosarcoma|Disorder|false|false|C0446516|armsnull|Adherence to Refills and Medications Scale|Finding|false|false|C0446516|arms
null|KIDINS220 gene|Finding|false|false|C0446516|armsnull|Upper arm|Anatomy|false|false|C5782111;C5575339;C2681631;C0206655|armsnull|null|Attribute|false|false|C0446516|armsnull|Side|Modifier|false|false||sidenull|Rails (medical device)|Device|false|false||railsnull|BORNHOLM EYE DISEASE|Disorder|false|false||bednull|Bachelor of Education|Finding|false|false||bednull|Beds|Device|false|false||bednull|Patient Location - Bed|Modifier|false|false||bednull|Leg|Anatomy|false|false|C5781420|legsnull|null|Attribute|false|false|C1140621|legsnull|Sensory (qualifier value)|Modifier|false|false||Sensorynull|Slightly (qualifier value)|Modifier|false|false||slightly
null|Slight (qualifier value)|Modifier|false|false||slightlynull|Upper Extremity|Anatomy|false|false||upper extremitiesnull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|All extremities|Anatomy|false|false||extremities
null|Limb structure|Anatomy|false|false||extremitiesnull|Lower Extremity|Anatomy|false|false|C2003888|lower extremitiesnull|Body Site Modifier - Lower|Anatomy|false|false|C2003888|lowernull|Lower (action)|Event|false|false|C0278454;C0015385;C0023216;C1548802|lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|All extremities|Anatomy|false|false|C2003888|extremities
null|Limb structure|Anatomy|false|false|C2003888|extremitiesnull|Stimulus|Phenomenon|false|false||stimulinull|TRI-AAT9-1 gene|Finding|false|false||Tri
null|Temptation and Restraint Inventory|Finding|false|false||Trinull|Fenamole|Drug|false|false||Pat
null|Fenamole|Drug|false|false||Patnull|Paroxysmal atrial tachycardia|Disorder|false|false||Patnull|glutamate-prephenate aminotransferase activity|Finding|false|false||Pat
null|aspartate-prephenate aminotransferase activity|Finding|false|false||Pat
null|protein acetyltransferase activity|Finding|false|false||Patnull|Thermoacoustic Computed Tomography|Procedure|false|false||Patnull|acetylcholine|Drug|false|false||Ach
null|acetylcholine|Drug|false|false||Ach
null|acetylcholine|Drug|false|false||Achnull|Achondroplasia|Disorder|false|false||Achnull|FGFR3 wt Allele|Finding|false|false||Ach
null|FGFR3 gene|Finding|false|false||Ach
null|Ache|Finding|false|false||Achnull|Acoli Language|Entity|false|false||Achnull|Plantar (qualifier value)|Anatomy|false|false||Plantar
null|Sole of Foot|Anatomy|false|false||Plantarnull|Communication Response|Finding|false|false||response
null|Disease Response|Finding|false|false||response
null|Answer (statement)|Finding|false|false||responsenull|Response process|Subject|false|false||responsenull|Flexor (Anatomical coordinate)|Anatomy|false|false||flexornull|Flexor <Diplocrepinae>|Entity|false|false||flexornull|Coordination of Benefits - Coordination|Finding|false|false||Coordination
null|Coordinated|Finding|false|false||Coordination
null|Physiologic Coordination|Finding|false|false||Coordinationnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Gait|Finding|false|false||Gaitnull|Relationship modifier - Patient|Finding|true|false||patient
null|Specimen Type - Patient|Finding|true|false||patient
null|Mail Claim Party - Patient|Finding|true|false||patient
null|Report source - Patient|Finding|true|false||patient
null|null|Finding|true|false||patient
null|Disabled Person Code - Patient|Finding|true|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|true|false||patientnull|BORNHOLM EYE DISEASE|Disorder|false|false||bednull|Bachelor of Education|Finding|false|false||bednull|Beds|Device|false|false||bednull|Patient Location - Bed|Modifier|false|false||bednull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||Generalnull|General medical service|Procedure|false|false||Generalnull|Generalized|Modifier|false|false||Generalnull|Chairs|Device|false|false||chairnull|Chairperson|Subject|false|false||chairnull|Eye|Anatomy|false|false|C5848506|eyesnull|null|Attribute|false|false|C0015392|eyesnull|HEENT|Anatomy|false|false||HEENTnull|Physical trauma|Disorder|true|false||trauma
null|Traumatic injury|Disorder|true|false||trauma
null|Trauma|Disorder|true|false||traumanull|Trauma assessment and care|Procedure|true|false||traumanull|Trauma, nursing specialty|Title|false|false||traumanull|trauma qualifier|Modifier|false|false||traumanull|jaundice|Finding|true|false||jaundice
null|Icterus|Finding|true|false||jaundice
null|yellow skin or eyes (symptom)|Finding|true|false||jaundicenull|Lesion|Finding|true|false|C0521367|lesionsnull|Oropharyngeal|Anatomy|false|false|C0221198|oropharynxnull|continuous electrocardiogram sinus bradycardia|Finding|false|false|C1305231;C0030471|sinus bradycardia
null|Sinus Bradycardia by ECG Finding|Finding|false|false|C1305231;C0030471|sinus bradycardia
null|Sinus bradycardia|Finding|false|false|C1305231;C0030471|sinus bradycardianull|Sinus brand of acetaminophen-pseudoephedrine|Drug|false|false|C1305231;C0030471|sinus
null|Sinus brand of acetaminophen-pseudoephedrine|Drug|false|false|C1305231;C0030471|sinusnull|pathologic fistula|Disorder|false|false|C1305231;C0030471|sinusnull|Sinus - general anatomical term|Anatomy|false|false|C0723346;C0085610;C5235162;C2108107;C0016169|sinus
null|Nasal sinus|Anatomy|false|false|C0723346;C0085610;C5235162;C2108107;C0016169|sinusnull|Bradycardia by ECG Finding|Finding|false|false||bradycardia
null|Bradycardia|Finding|false|false||bradycardianull|Pulmonary ventilator management|Procedure|false|false||Pulmnull|Hereditary Multiple Exostoses|Disorder|false|false||Extnull|EXT1 wt Allele|Finding|false|false||Ext
null|EXT1 gene|Finding|false|false||Extnull|Feels warm|Finding|false|false||Warmnull|warming process|Phenomenon|false|false||Warmnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Eruption of skin (disorder)|Disorder|true|false||rashnull|Skin rash|Finding|true|false||rash
null|Eruptions|Finding|true|false||rash
null|Exanthema|Finding|true|false||rashnull|Mottling|Finding|false|false||mottlingnull|Neurologic (qualifier value)|Modifier|false|false||Neurologicnull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Slow|Modifier|false|false||slownull|Shortened|Modifier|false|false||shortnull|Short Value|LabModifier|false|false||short
null|Short|LabModifier|false|false||shortnull|Sentence|Finding|false|false||sentencenull|More|LabModifier|false|false||Morenull|Humor|Finding|false|false||humornull|Humor therapy|Procedure|false|false||humornull|complex (molecular entity)|Drug|false|false||complexnull|Complex|Modifier|false|false||complexnull|Sentence|Finding|false|false||sentencesnull|Eye|Anatomy|false|false|C5848506;C3810854;C0587267|Eyesnull|null|Attribute|false|false|C0015392|Eyesnull|Close|Finding|false|false|C0015392|close
null|Closed|Finding|false|false|C0015392|closenull|Speech|Finding|false|false||Speechnull|Speech assessment|Procedure|false|false||Speechnull|Spontaneous|Finding|true|false||spontaneousnull|Speech|Finding|true|false||speechnull|Speech assessment|Procedure|true|false||speechnull|system output|Finding|true|false||outputnull|Measurement of fluid output|Procedure|true|false||outputnull|LITAF gene|Finding|false|false||simplenull|Simple|Modifier|false|false||simplenull|Neoplasm of uncertain or unknown behavior of cranial nerves|Disorder|false|false|C0010268;C0037303;C0027740|Cranial Nerves
null|Benign neoplasm of cranial nerves|Disorder|false|false|C0010268;C0037303;C0027740|Cranial Nervesnull|Cranial Nerves|Anatomy|false|false|C0004992;C0496937|Cranial Nervesnull|Bone structure of cranium|Anatomy|false|false|C0004992;C0496937|Cranialnull|Cranial|Modifier|false|false||Cranialnull|Nerve|Anatomy|false|false|C0004992;C0496937|Nervesnull|Pupil|Anatomy|false|false||Pupilsnull|Nystagmus|Disorder|false|false||nystagmusnull|facial sensation|Finding|false|false|C0015450|facial sensationnull|Face|Anatomy|false|false|C2229507;C0517999;C1554187;C0036658;C0542538|facialnull|Facial|Modifier|false|false||facialnull|Observation of Sensation|Finding|false|false|C0015450|sensation
null|Sensory perception|Finding|false|false|C0015450|sensationnull|sensory exam|Procedure|false|false|C0015450|sensationnull|Sensation quality|Modifier|false|false||sensationnull|Gender Status - Intact|Finding|false|false|C0015450|intactnull|Intact|Modifier|false|false||intactnull|Roman numeral VII|Finding|false|false|C2338708;C3496273;C3496274|VIInull|Lamina VII of gray matter of spinal cord|Anatomy|false|false|C0445385|VII
null|lobule VII|Anatomy|false|false|C0445385|VII
null|layer VII (Cajal)|Anatomy|false|false|C0445385|VIInull|Facial Paresis|Disorder|true|false|C0015450|facial droopnull|Unilateral facial palsy|Finding|true|false|C0015450|facial droopnull|Face|Anatomy|false|false|C4022719;C0427055|facialnull|Facial|Modifier|false|false||facialnull|Face|Anatomy|false|false|C0332516;C2699744|facialnull|Facial|Modifier|false|false||facialnull|Set of muscles|Anatomy|false|false||musculaturenull|Symmetric Relationship|Finding|false|false|C0015450|symmetric
null|Symmetrical|Finding|false|false|C0015450|symmetricnull|Grimaces|Finding|false|false||grimacenull|Limited component (foundation metadata concept)|Finding|false|false||limited
null|Limited (extensiveness)|Finding|false|false||limitednull|Face|Anatomy|false|false||facialnull|Facial|Modifier|false|false||facialnull|Movement|Finding|false|false||movementsnull|Palate|Anatomy|false|false|C0153933;C0872394|palatenull|tongue midline|Finding|false|false|C1660780;C0040408|tongue midlinenull|Benign neoplasm of tongue|Disorder|false|false|C1660780;C0040408;C0700374|tonguenull|Procedure on tongue|Procedure|false|false|C0040408;C0700374;C1660780|tonguenull|Tongue|Anatomy|false|false|C0872394;C0153933;C3693372|tonguenull|midline cell component|Anatomy|false|false|C0153933;C3693372;C0872394|midlinenull|Midline (qualifier value)|Modifier|false|false||midlinenull|motor movement|Finding|false|false||Motornull|Motor Device|Device|false|false||Motornull|Bulk (conceptual)|Drug|false|false||bulk
null|Dietary Fiber|Drug|false|false||bulknull|Lifting|Event|false|false|C0015385|Liftingnull|Limb structure|Anatomy|false|false|C0206655;C0206244;C5575339;C2681631|arms and legsnull|Alveolar rhabdomyosarcoma|Disorder|false|false|C0446516;C1140621;C0015385|armsnull|Adherence to Refills and Medications Scale|Finding|false|false|C0446516;C0015385|arms
null|KIDINS220 gene|Finding|false|false|C0446516;C0015385|armsnull|Upper arm|Anatomy|false|false|C5782111;C0206655;C5575339;C2681631|armsnull|null|Attribute|false|false|C0446516|armsnull|Leg|Anatomy|false|false|C0206655;C5781420|legsnull|null|Attribute|false|false|C1140621|legsnull|Gravity (physical force)|Phenomenon|true|false||gravitynull|Gravity - Unit of Force|LabModifier|false|false||gravitynull|Resistance (Psychotherapeutic)|Finding|true|false||resistance
null|social resistance|Finding|true|false||resistance
null|Resistance Process|Finding|true|false||resistancenull|Resistance|Attribute|true|false||resistancenull|Sensory (qualifier value)|Modifier|false|false||Sensorynull|Observation of Sensation|Finding|false|false||Sensation
null|Sensory perception|Finding|false|false||Sensationnull|sensory exam|Procedure|false|false||Sensationnull|Sensation quality|Modifier|false|false||Sensationnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Touch sensation|Finding|false|false||touch
null|Touch Perception|Finding|false|false||touchnull|Therapeutic Touch|Procedure|false|false||touchnull|Tactile|Modifier|false|false||touchnull|Body temperature measurement|Procedure|false|false||temperaturenull|Body Temperature|Subject|false|false||temperaturenull|Temperature|LabModifier|false|false||temperaturenull|Patella|Anatomy|false|false||patellarnull|Biceps brachii muscle structure|Anatomy|false|false||bicepsnull|Structure of brachioradialis muscle|Anatomy|false|false||brachioradialisnull|Coordination of Benefits - Coordination|Finding|false|false||Coordination
null|Coordinated|Finding|false|false||Coordination
null|Physiologic Coordination|Finding|false|false||Coordinationnull|Cerebellar Dysmetria|Finding|true|false||dysmetrianull|Tremor|Finding|true|false||tremornull|Gait|Finding|false|false||Gaitnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|Laboratory test finding|Lab|false|false||labsnull|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSEnull|Glucose measurement|Procedure|false|false||GLUCOSEnull|Glucose^1.5H post dose glucagon|Lab|false|false||GLUCOSEnull|urea|Drug|false|false||UREA
null|urea|Drug|false|false||UREA
null|urea|Drug|false|false||UREAnull|Urea measurement|Procedure|false|false||UREAnull|Sodium supplements|Drug|false|false||SODIUM
null|sodium|Drug|false|false||SODIUM
null|sodium|Drug|false|false||SODIUM
null|Sodium Drug Class|Drug|false|false||SODIUMnull|Sodium metabolic function|Finding|false|false||SODIUMnull|Sodium measurement|Procedure|false|false||SODIUMnull|Potassium Drug Class|Drug|false|false||POTASSIUM
null|Dietary Potassium|Drug|false|false||POTASSIUM
null|potassium|Drug|false|false||POTASSIUM
null|potassium|Drug|false|false||POTASSIUM
null|potassium|Drug|false|false||POTASSIUM
null|Potassium supplement|Drug|false|false||POTASSIUM
null|Potassium supplement|Drug|false|false||POTASSIUMnull|Potassium metabolic function|Finding|false|false||POTASSIUMnull|Potassium measurement|Procedure|false|false||POTASSIUMnull|chloride ion|Drug|false|false||CHLORIDE
null|Chlorides|Drug|false|false||CHLORIDEnull|Chloride metabolic function|Finding|false|false||CHLORIDEnull|Chloride measurement|Procedure|false|false||CHLORIDEnull|Total|Modifier|false|false||TOTALnull|carbon dioxide|Drug|false|false||CO2
null|carbon dioxide|Drug|false|false||CO2null|MT-CO2 gene|Finding|false|false||CO2
null|null|Finding|false|false||CO2
null|C2 wt Allele|Finding|false|false||CO2null|blood anion gap (lab test)|Procedure|false|false||ANION GAP
null|Anion gap measurement|Procedure|false|false||ANION GAPnull|Anion Gap|Attribute|false|false||ANION GAPnull|Anion gap result|Lab|false|false||ANION GAPnull|Anions|Drug|false|false||ANIONnull|Ras GTPase-Activating Protein 1, Human|Drug|false|false||GAP
null|Ras GTPase-Activating Protein 1, Human|Drug|false|false||GAP
null|GTPase-Activating Proteins|Drug|false|false||GAP
null|GTPase-Activating Proteins|Drug|false|false||GAPnull|RASA1 wt Allele|Finding|false|false||GAP
null|RASA1 gene|Finding|false|false||GAPnull|Gap (space)|Modifier|false|false||GAPnull|Alanine Transaminase|Drug|false|false||ALT
null|Alanine Transaminase|Drug|false|false||ALTnull|Liposarcoma, well differentiated|Disorder|false|false||ALT
null|Atypical Lipoma|Disorder|false|false||ALTnull|null|Finding|false|false||ALT
null|Alternative Billing Concepts|Finding|false|false||ALT
null|GPT gene|Finding|false|false||ALTnull|Antibiotic Lock Therapy|Procedure|false|false||ALTnull|Southern Altai Language|Entity|false|false||ALTnull|SGPT - Glutamate pyruvate transaminase|Drug|false|false||SGPT
null|SGPT - Glutamate pyruvate transaminase|Drug|false|false||SGPTnull|GPT gene|Finding|false|false||SGPTnull|Serum Alanine Transaminase Test|Procedure|false|false||SGPTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false|C1185650|AST
null|Aspartate Transaminase|Drug|false|false|C1185650|AST
null|Aspartate Transaminase|Drug|false|false|C1185650|AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false|C1185650|AST
null|SLC17A5 protein, human|Drug|false|false|C1185650|AST
null|SLC17A5 protein, human|Drug|false|false|C1185650|ASTnull|Atypical Spitz Nevus|Disorder|false|false|C1185650|ASTnull|SLC17A5 wt Allele|Finding|false|false|C1185650|AST
null|SLC17A5 gene|Finding|false|false|C1185650|AST
null|GOT1 gene|Finding|false|false|C1185650|ASTnull|Asterion|Anatomy|false|false|C0201899;C4522245;C1415181;C0004002;C0242192;C1121182;C1415181;C1420113;C5960784|ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||SGOT
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||SGOTnull|GOT1 gene|Finding|false|false|C1185650|SGOTnull|Aspartate aminotransferase measurement|Procedure|false|false|C1185650|SGOTnull|Alkaline Phosphatase|Drug|false|false||ALK PHOS
null|Alkaline Phosphatase|Drug|false|false||ALK PHOSnull|Alkaline phosphatase measurement|Procedure|false|false||ALK PHOSnull|ALK protein, human|Drug|false|false||ALK
null|ALK protein, human|Drug|false|false||ALKnull|ALK protein, human|Finding|false|false||ALK
null|ALK gene|Finding|false|false||ALK
null|ALK wt Allele|Finding|false|false||ALKnull|Phos <Photinae>|Entity|false|false||PHOSnull|CALCIUM SUPPLEMENTS|Drug|false|false||CALCIUM
null|calcium|Drug|false|false||CALCIUM
null|calcium|Drug|false|false||CALCIUM
null|calcium|Drug|false|false||CALCIUM
null|CALCIUM SUPPLEMENTS|Drug|false|false||CALCIUM
null|Calcium, Dietary|Drug|false|false||CALCIUM
null|Calcium [EPC]|Drug|false|false||CALCIUM
null|Calcium Drug Class|Drug|false|false||CALCIUMnull|Calcium metabolic function|Finding|false|false||CALCIUMnull|Calcium measurement|Procedure|false|false||CALCIUMnull|phosphate ion|Drug|false|false||PHOSPHATE
null|Phosphates|Drug|false|false||PHOSPHATE
null|phosphate ion|Drug|false|false||PHOSPHATEnull|Phosphate measurement|Procedure|false|false||PHOSPHATEnull|Magnesium supplements, alimentary tract and metabolism|Drug|false|false||MAGNESIUM
null|magnesium|Drug|false|false||MAGNESIUM
null|magnesium|Drug|false|false||MAGNESIUM
null|Magnesium Drug Class|Drug|false|false||MAGNESIUM
null|Magnesium supplements, alimentary tract and metabolism|Drug|false|false||MAGNESIUMnull|Magnesium measurement|Procedure|false|false||MAGNESIUMnull|TGM2 protein, human|Drug|false|false||tTG
null|TGM2 protein, human|Drug|false|false||tTG
null|TGM2 protein, human|Drug|false|false||tTGnull|TGM2 wt Allele|Finding|false|false||tTGnull|immunoglobulin A, human|Drug|false|false||IgA
null|immunoglobulin A|Drug|false|false||IgA
null|immunoglobulin A|Drug|false|false||IgA
null|immunoglobulin A, human|Drug|false|false||IgAnull|CD79A wt Allele|Finding|false|false||IgA
null|CD79A gene|Finding|false|false||IgAnull|Immunoglobulin A measurement|Procedure|false|false||IgAnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C0014792;C1114281|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||HGB
null|Hemoglobin|Drug|false|false||HGBnull|CYGB gene|Finding|false|false||HGBnull|Hemoglobin concentration|Lab|false|false||HGBnull|Hemopoietic stem cell transplant|Procedure|false|false||HCT
null|Hematocrit Measurement|Procedure|false|false||HCTnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||PLTnull|Count Dosing Unit|LabModifier|false|false||COUNT
null|Count|LabModifier|false|false||COUNTnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Hour|Time|false|false||HOURSnull|Random|Modifier|false|false||RANDOMnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Rh Negative Blood Group|Finding|false|false||NEGATIVE
null|Negative|Finding|false|false||NEGATIVE
null|Negative Finding|Finding|false|false||NEGATIVEnull|Expression Negative|Lab|false|false||NEGATIVEnull|Negative - qualifier|Modifier|false|false||NEGATIVE
null|Negative Charge|Modifier|false|false||NEGATIVEnull|Negative Number|LabModifier|false|false||NEGATIVEnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Opiates|Drug|false|false||opiates
null|Opiates|Drug|false|false||opiates
null|Opiates|Drug|false|false||opiates
null|Opiate Alkaloids|Drug|false|false||opiates
null|Opiate Alkaloids|Drug|false|false||opiates
null|Opiate Alkaloids|Drug|false|false||opiatesnull|Opiate Measurement|Procedure|false|false||opiatesnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|cocaine|Drug|false|false||cocaine
null|cocaine|Drug|false|false||cocaine
null|cocaine|Drug|false|false||cocaine
null|cocaine|Drug|false|false||cocainenull|Poisoning by cocaine|Disorder|false|false||cocainenull|Cocaine measurement|Procedure|false|false||cocainenull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Color of urine|Finding|false|false||URINE  COLORnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|color additive|Drug|false|false||COLOR
null|Coloring Excipient|Drug|false|false||COLORnull|color - solid dosage form|Modifier|false|false||COLOR
null|Color|Modifier|false|false||COLORnull|Color quantity|LabModifier|false|false||COLORnull|Cereal plant straw|Drug|false|false||Strawnull|Straw package type|Device|false|false||Strawnull|Straw Color|Modifier|false|false||Strawnull|Straw (unit of presentation)|LabModifier|false|false||Strawnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Hematuria|Disorder|false|false||URINE  BLOODnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|nitrite ion|Drug|false|false||NITRITE
null|Nitrites|Drug|false|false||NITRITE
null|Nitrites|Drug|false|false||NITRITE
null|Nitrites|Drug|false|false||NITRITE
null|nitrite ion|Drug|false|false||NITRITE
null|nitrite ion|Drug|false|false||NITRITEnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Proteins|Drug|false|false||PROTEIN
null|Proteins|Drug|false|false||PROTEINnull|Protein Info|Finding|false|false||PROTEINnull|Protein measurement|Procedure|false|false||PROTEINnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSEnull|Glucose measurement|Procedure|false|false||GLUCOSEnull|Glucose^1.5H post dose glucagon|Lab|false|false||GLUCOSEnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Ketones|Drug|false|false||KETONEnull|bilirubin preparation|Drug|false|false||BILIRUBIN
null|bilirubin preparation|Drug|false|false||BILIRUBIN
null|Bilirubin|Drug|false|false||BILIRUBIN
null|Bilirubin|Drug|false|false||BILIRUBINnull|Bilirubin, total measurement|Procedure|false|false||BILIRUBIN
null|blood bilirubin level test|Procedure|false|false||BILIRUBINnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|null|Lab|false|false|C0014792|URINE  RBC
null|Red blood cells urine positive|Lab|false|false|C0014792|URINE  RBCnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C0014792;C0221752;C2188659;C1114281|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Leukocytes|Anatomy|false|false||WBCnull|bacteria aspects|Finding|false|false||BACTERIAnull|Bacteria <walking sticks>|Entity|false|false||BACTERIA
null|Bacteria|Entity|false|false||BACTERIAnull|Yeast, Dried|Drug|false|false||YEAST
null|Candida albicans allergenic extract|Drug|false|false||YEAST
null|Candida albicans allergenic extract|Drug|false|false||YEAST
null|Candida albicans allergenic extract|Drug|false|false||YEASTnull|Saccharomyces cerevisiae|Entity|false|false||YEAST
null|Yeasts|Entity|false|false||YEASTnull|Tissue Factor Pathway Inhibitor, human|Drug|false|false||EPI
null|epinephrine|Drug|false|false||EPI
null|epinephrine|Drug|false|false||EPI
null|epinephrine|Drug|false|false||EPI
null|Tissue Factor Pathway Inhibitor, human|Drug|false|false||EPInull|Exocrine pancreatic insufficiency|Disorder|false|false||EPInull|Eysenck personality inventory|Finding|false|false||EPI
null|TFPI wt Allele|Finding|false|false||EPI
null|TFPI gene|Finding|false|false||EPInull|Electronic Portal Imaging|Procedure|false|false||EPI
null|Echo-Planar Imaging|Procedure|false|false||EPInull|Mucus in urine (finding)|Finding|false|false||URINE  MUCOUSnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Mucus (substance)|Finding|false|false||MUCOUS
null|mucus layer|Finding|false|false||MUCOUSnull|Mucous appearance|Modifier|false|false||MUCOUSnull|Retinoic Acid Response Element|Finding|false|false||RAREnull|Infrequent|Time|false|false||RAREnull|Rare|Modifier|false|false||RAREnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C0014792;C1114281|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||HGB
null|Hemoglobin|Drug|false|false||HGBnull|CYGB gene|Finding|false|false||HGBnull|Hemoglobin concentration|Lab|false|false||HGBnull|Hemopoietic stem cell transplant|Procedure|false|false||HCT
null|Hematocrit Measurement|Procedure|false|false||HCTnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Monos|Drug|false|false||MONOS
null|Mono-S|Drug|false|false||MONOS
null|Monos|Drug|false|false||MONOSnull|SARCOIDOSIS, EARLY-ONSET|Disorder|false|false||EOS
null|Familial eosinophilia|Disorder|false|false||EOSnull|PRSS33 gene|Finding|false|false||EOS
null|IKZF4 gene|Finding|false|false||EOSnull|Eos <Loriini>|Entity|false|false||EOSnull|Primed lymphocyte test|Procedure|false|false||PLTnull|Count Dosing Unit|LabModifier|false|false||COUNT
null|Count|LabModifier|false|false||COUNTnull|Partial pressure of Oxygen|Finding|false|false||PO2
null|US Military enlisted E5|Finding|false|false||PO2null|PO2 measurement|Procedure|false|false||PO2null|Carbon dioxide measurement, partial pressure|Procedure|false|false||PCO2null|Carbon dioxide, partial pressure|Lab|false|false||PCO2null|Total|Modifier|false|false||TOTALnull|carbon dioxide|Drug|false|false||CO2
null|carbon dioxide|Drug|false|false||CO2null|MT-CO2 gene|Finding|false|false|C2987514|CO2
null|null|Finding|false|false|C2987514|CO2
null|C2 wt Allele|Finding|false|false|C2987514|CO2null|nitrogenous base|Drug|false|false|C2987514|BASE
null|Base|Drug|false|false|C2987514|BASE
null|Dental Base|Drug|false|false|C2987514|BASE
null|base - RoleClass|Drug|false|false|C2987514|BASEnull|Base - General Qualifier|Finding|false|false|C2987514|BASE
null|BPIFA4P gene|Finding|false|false|C2987514|BASE
null|Base - RX Component Type|Finding|false|false|C2987514|BASEnull|Anatomical base|Anatomy|false|false|C4284286;C1537986;C0860710;C0947611;C0282411;C1704464;C0178499;C1550601;C1880279;C1549548;C1705938;C1843354|BASEnull|Base - unit of product usage|LabModifier|false|false||BASEnull|Published Comment|Finding|false|false|C2987514|COMMENTS
null|Comment|Finding|false|false|C2987514|COMMENTSnull|Green color|Modifier|false|false||GREENnull|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSEnull|Glucose measurement|Procedure|false|false||GLUCOSEnull|Glucose^1.5H post dose glucagon|Lab|false|false||GLUCOSEnull|urea|Drug|false|false||UREA
null|urea|Drug|false|false||UREA
null|urea|Drug|false|false||UREAnull|Urea measurement|Procedure|false|false||UREAnull|Sodium supplements|Drug|false|false||SODIUM
null|sodium|Drug|false|false||SODIUM
null|sodium|Drug|false|false||SODIUM
null|Sodium Drug Class|Drug|false|false||SODIUMnull|Sodium metabolic function|Finding|false|false||SODIUMnull|Sodium measurement|Procedure|false|false||SODIUMnull|Potassium Drug Class|Drug|false|false||POTASSIUM
null|Dietary Potassium|Drug|false|false||POTASSIUM
null|potassium|Drug|false|false||POTASSIUM
null|potassium|Drug|false|false||POTASSIUM
null|potassium|Drug|false|false||POTASSIUM
null|Potassium supplement|Drug|false|false||POTASSIUM
null|Potassium supplement|Drug|false|false||POTASSIUMnull|Potassium metabolic function|Finding|false|false||POTASSIUMnull|Potassium measurement|Procedure|false|false||POTASSIUMnull|chloride ion|Drug|false|false||CHLORIDE
null|Chlorides|Drug|false|false||CHLORIDEnull|Chloride metabolic function|Finding|false|false||CHLORIDEnull|Chloride measurement|Procedure|false|false||CHLORIDEnull|Total|Modifier|false|false||TOTALnull|carbon dioxide|Drug|false|false||CO2
null|carbon dioxide|Drug|false|false||CO2null|MT-CO2 gene|Finding|false|false||CO2
null|null|Finding|false|false||CO2
null|C2 wt Allele|Finding|false|false||CO2null|blood anion gap (lab test)|Procedure|false|false||ANION GAP
null|Anion gap measurement|Procedure|false|false||ANION GAPnull|Anion Gap|Attribute|false|false||ANION GAPnull|Anion gap result|Lab|false|false||ANION GAPnull|Anions|Drug|false|false||ANIONnull|Ras GTPase-Activating Protein 1, Human|Drug|false|false||GAP
null|Ras GTPase-Activating Protein 1, Human|Drug|false|false||GAP
null|GTPase-Activating Proteins|Drug|false|false||GAP
null|GTPase-Activating Proteins|Drug|false|false||GAPnull|RASA1 wt Allele|Finding|false|false||GAP
null|RASA1 gene|Finding|false|false||GAPnull|Gap (space)|Modifier|false|false||GAPnull|Alanine Transaminase|Drug|false|false||ALT
null|Alanine Transaminase|Drug|false|false||ALTnull|Liposarcoma, well differentiated|Disorder|false|false||ALT
null|Atypical Lipoma|Disorder|false|false||ALTnull|null|Finding|false|false||ALT
null|Alternative Billing Concepts|Finding|false|false||ALT
null|GPT gene|Finding|false|false||ALTnull|Antibiotic Lock Therapy|Procedure|false|false||ALTnull|Southern Altai Language|Entity|false|false||ALTnull|SGPT - Glutamate pyruvate transaminase|Drug|false|false||SGPT
null|SGPT - Glutamate pyruvate transaminase|Drug|false|false||SGPTnull|GPT gene|Finding|false|false||SGPTnull|Serum Alanine Transaminase Test|Procedure|false|false||SGPTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false|C1185650|AST
null|Aspartate Transaminase|Drug|false|false|C1185650|AST
null|Aspartate Transaminase|Drug|false|false|C1185650|AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false|C1185650|AST
null|SLC17A5 protein, human|Drug|false|false|C1185650|AST
null|SLC17A5 protein, human|Drug|false|false|C1185650|ASTnull|Atypical Spitz Nevus|Disorder|false|false|C1185650|ASTnull|SLC17A5 wt Allele|Finding|false|false|C1185650|AST
null|SLC17A5 gene|Finding|false|false|C1185650|AST
null|GOT1 gene|Finding|false|false|C1185650|ASTnull|Asterion|Anatomy|false|false|C1415181;C1420113;C5960784;C0201899;C1415181;C4522245;C0004002;C0242192;C1121182|ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||SGOT
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||SGOTnull|GOT1 gene|Finding|false|false|C1185650|SGOTnull|Aspartate aminotransferase measurement|Procedure|false|false|C1185650|SGOTnull|Creatine Kinase|Drug|false|false||CPK
null|Creatine Kinase|Drug|false|false||CPKnull|PIK3C2A gene|Finding|false|false||CPKnull|Creatine kinase measurement|Procedure|false|false||CPKnull|ALK protein, human|Drug|false|false||ALK
null|ALK protein, human|Drug|false|false||ALKnull|ALK protein, human|Finding|false|false||ALK
null|ALK gene|Finding|false|false||ALK
null|ALK wt Allele|Finding|false|false||ALKnull|Phos <Photinae>|Entity|false|false||PHOSnull|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MB
null|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MBnull|creatine kinase activity|Finding|false|false||CK-MBnull|Serum creatine phosphokinase MB isoenzyme measurement|Procedure|false|false||CK-MB
null|Creatine kinase MB measurement|Procedure|false|false||CK-MBnull|Albumin|Drug|false|false||ALBUMIN
null|Albumins|Drug|false|false||ALBUMIN
null|Albumins|Drug|false|false||ALBUMIN
null|Albumin|Drug|false|false||ALBUMINnull|Albumin metabolic function|Finding|false|false||ALBUMIN
null|ALB gene|Finding|false|false||ALBUMINnull|Albumin measurement|Procedure|false|false||ALBUMINnull|CALCIUM SUPPLEMENTS|Drug|false|false||CALCIUM
null|calcium|Drug|false|false||CALCIUM
null|calcium|Drug|false|false||CALCIUM
null|calcium|Drug|false|false||CALCIUM
null|CALCIUM SUPPLEMENTS|Drug|false|false||CALCIUM
null|Calcium, Dietary|Drug|false|false||CALCIUM
null|Calcium [EPC]|Drug|false|false||CALCIUM
null|Calcium Drug Class|Drug|false|false||CALCIUMnull|Calcium metabolic function|Finding|false|false||CALCIUMnull|Calcium measurement|Procedure|false|false||CALCIUMnull|phosphate ion|Drug|false|false||PHOSPHATE
null|Phosphates|Drug|false|false||PHOSPHATE
null|phosphate ion|Drug|false|false||PHOSPHATEnull|Phosphate measurement|Procedure|false|false||PHOSPHATEnull|Magnesium supplements, alimentary tract and metabolism|Drug|false|false||MAGNESIUM
null|magnesium|Drug|false|false||MAGNESIUM
null|magnesium|Drug|false|false||MAGNESIUM
null|Magnesium Drug Class|Drug|false|false||MAGNESIUM
null|Magnesium supplements, alimentary tract and metabolism|Drug|false|false||MAGNESIUMnull|Magnesium measurement|Procedure|false|false||MAGNESIUMnull|vitamin B12|Drug|false|false||VIT B12
null|cobalamins|Drug|false|false||VIT B12
null|cobalamins|Drug|false|false||VIT B12
null|vitamin B12|Drug|false|false||VIT B12
null|vitamin B12|Drug|false|false||VIT B12null|VIT gene|Finding|false|false||VIT
null|EWS Vitals Table|Finding|false|false||VIT
null|AML Vitals Table|Finding|false|false||VITnull|VIT Regimen|Procedure|false|false||VITnull|TNFAIP1 wt Allele|Finding|false|false||B12
null|NDUFB3 gene|Finding|false|false||B12
null|TNFAIP1 gene|Finding|false|false||B12null|thyrotropin|Drug|false|false||TSH
null|thyrotropin|Drug|false|false||TSH
null|thyrotropin|Drug|false|false||TSHnull|Thyroid stimulating hormone measurement|Procedure|false|false||TSHnull|null|Attribute|false|false||TSHnull|thyrotropin|Drug|false|false||TSH
null|thyrotropin|Drug|false|false||TSH
null|thyrotropin|Drug|false|false||TSHnull|Thyroid stimulating hormone measurement|Procedure|false|false||TSHnull|null|Attribute|false|false||TSHnull|Titer|LabModifier|false|false||TITERnull|C-Reactive Protein, human|Drug|false|false||CRP
null|C-reactive protein|Drug|false|false||CRP
null|C-reactive protein|Drug|false|false||CRP
null|C-Reactive Protein, human|Drug|false|false||CRPnull|CRP wt Allele|Finding|false|false||CRP
null|CRP gene|Finding|false|false||CRP
null|CSRP1 gene|Finding|false|false||CRP
null|PPIAP10 gene|Finding|false|false||CRPnull|Pidgin and Creole language|Entity|false|false||CRPnull|Rh Negative Blood Group|Finding|false|false||NEGATIVE
null|Negative|Finding|false|false||NEGATIVE
null|Negative Finding|Finding|false|false||NEGATIVEnull|Expression Negative|Lab|false|false||NEGATIVEnull|Negative - qualifier|Modifier|false|false||NEGATIVE
null|Negative Charge|Modifier|false|false||NEGATIVEnull|Negative Number|LabModifier|false|false||NEGATIVEnull|Arylsulfatase A, human|Drug|false|false||ASA
null|Arylsulfatase A, human|Drug|false|false||ASA
null|aspirin|Drug|false|false||ASA
null|aspirin|Drug|false|false||ASAnull|ARSA gene|Finding|false|false||ASAnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|CNS depressants ethanol|Drug|false|false||ETHANOL
null|CNS depressants ethanol|Drug|false|false||ETHANOL
null|antiseptics ethanol|Drug|false|false||ETHANOL
null|antiseptics ethanol|Drug|false|false||ETHANOL
null|ethanol|Drug|false|false||ETHANOL
null|ethanol|Drug|false|false||ETHANOLnull|Toxic effect of ethyl alcohol|Disorder|false|false||ETHANOLnull|Ethanol measurement|Procedure|false|false||ETHANOLnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Electroencephalography|Procedure|false|false||EEGnull|impression (attitude)|Finding|false|false||IMPRESSION
null|EKG impression|Finding|false|false||IMPRESSIONnull|Telemetry|Procedure|false|false||telemetrynull|Background|Finding|false|false||backgroundnull|Waking|Finding|false|false||wakingnull|Upon Awakening - schedule frequency|Time|false|false||wakingnull|Sleep brand of diphenhydramine hydrochloride|Drug|false|false||sleep
null|Sleep brand of diphenhydramine hydrochloride|Drug|false|false||sleepnull|Sleep|Finding|false|false||sleepnull|Patterns|Modifier|false|false||patternsnull|Focal|Modifier|false|false||focalnull|Congenital Abnormality|Disorder|true|false||abnormalitiesnull|teratologic|Finding|true|false||abnormalitiesnull|Seizures|Finding|false|false||seizuresnull|Bradycardia by ECG Finding|Finding|false|false||bradycardia
null|Bradycardia|Finding|false|false||bradycardianull|Imaging problem|Finding|false|false||IMAGINGnull|Diagnostic Imaging|Procedure|false|false||IMAGING
null|Imaging Techniques|Procedure|false|false||IMAGINGnull|Imaging Technology|Title|false|false||IMAGINGnull|Nuclear magnetic resonance imaging brain|Procedure|false|false|C4266577;C0006104|MRI BRAINnull|CYREN gene|Finding|false|false|C4266577;C0006104|MRInull|Magnetic resonance imaging service|Procedure|false|false|C4266577;C0006104|MRI
null|Magnetic Resonance Imaging|Procedure|false|false|C4266577;C0006104|MRInull|Maori Language|Entity|false|false||MRInull|Brain Diseases|Disorder|false|false|C4266577;C0006104|BRAINnull|Head>Brain|Anatomy|false|false|C4028269;C0024485;C0587658;C1824234;C0006111|BRAIN
null|Brain|Anatomy|false|false|C4028269;C0024485;C0587658;C1824234;C0006111|BRAINnull|Contrast Media|Drug|true|false||CONTRASTnull|Contrast|Modifier|false|false||CONTRASTnull|findings aspects|Finding|false|false||FINDINGSnull|null|Attribute|false|false||FINDINGSnull|FLAIR (product)|Drug|false|false||FLAIR
null|FLAIR (product)|Drug|false|false||FLAIRnull|Fluid Attenuated Inversion Recovery|Procedure|false|false||FLAIRnull|Isointense|Finding|false|false||isointensenull|Lesion|Finding|false|false|C1660780|lesion
null|null|Finding|false|false|C1660780|lesionnull|midline cell component|Anatomy|false|false|C1546698;C0221198|midlinenull|Midline (qualifier value)|Modifier|false|false||midlinenull|Adenohypophyseal Diseases|Disorder|false|false||anteriornull|Anterior|Modifier|false|false||anteriornull|Posterior Pituitary Hormone Drug Class|Drug|false|false|C0447640;C0032009;C0032005|posterior pituitary
null|posterior pituitary hormones|Drug|false|false|C0447640;C0032009;C0032005|posterior pituitary
null|posterior pituitary hormones|Drug|false|false|C0447640;C0032009;C0032005|posterior pituitary
null|posterior pituitary hormones|Drug|false|false|C0447640;C0032009;C0032005|posterior pituitary
null|Posterior Pituitary Hormone Drug Class|Drug|false|false|C0447640;C0032009;C0032005|posterior pituitarynull|Pituitary Gland, Posterior|Anatomy|false|false|C3714635;C0032017;C0304812;C0032002;C0751438|posterior pituitary
null|pars nervosa of hypophysis|Anatomy|false|false|C3714635;C0032017;C0304812;C0032002;C0751438|posterior pituitarynull|Posterior pituitary disease|Disorder|false|false|C0032005;C0447640;C0032009|posteriornull|Dorsal|Modifier|false|false||posteriornull|Pituitary hormone preparation|Drug|false|false|C0447640;C0032009;C0032005|pituitary
null|Pituitary hormone preparation|Drug|false|false|C0447640;C0032009;C0032005|pituitary
null|Pituitary hormone preparation|Drug|false|false|C0447640;C0032009;C0032005|pituitarynull|Pituitary Diseases|Disorder|false|false|C0032005;C0447640;C0032009|pituitarynull|Pituitary Gland|Anatomy|false|false|C3714635;C0032017;C0751438;C0032002;C0304812|pituitarynull|Evidence|Finding|true|false||evidencenull|Hemorrhage|Finding|false|false||hemorrhagenull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Mass Effect|Finding|false|false||mass effectnull|Mass of body structure|Finding|false|false||mass
null|Morphology, Attenuation, Size, and Structure Criteria|Finding|false|false||mass
null|null|Finding|false|false||mass
null|FBN1 wt Allele|Finding|false|false||mass
null|FBN1 gene|Finding|false|false||mass
null|Mass of body region|Finding|false|false||massnull|Mass, a measure of quantity of matter|LabModifier|false|false||mass
null|Molecular Mass|LabModifier|false|false||massnull|Effect, Appearance|Modifier|false|false||effect
null|Effect|Modifier|false|false||effectnull|Midline Shift|Finding|false|false|C1660780|midline shiftnull|midline cell component|Anatomy|false|false|C0021308;C2347509;C4086580;C0333051|midlinenull|Midline (qualifier value)|Modifier|false|false||midlinenull|shift displacement|Finding|false|false|C1660780|shiftnull|Physical Shift|Phenomenon|false|false|C1660780|shiftnull|Infarction|Finding|false|false|C1660780|infarctionnull|Heart Ventricle|Anatomy|false|false|C2827597|ventriclesnull|Diameter (qualifier value)|LabModifier|false|false||calibernull|Computer Configuration|Finding|false|false|C0018827|configurationnull|With configuration|Modifier|false|false||configurationnull|Observation Interpretation - Abnormal|Finding|true|false||abnormal
null|Abnormal|Finding|true|false||abnormalnull|Refractive surgery enhancement|Procedure|true|false||enhancementnull|Enhance (action)|Event|true|false||enhancementnull|Contrast Media|Drug|false|false||contrastnull|Contrast|Modifier|false|false||contrastnull|Administration (procedure)|Procedure|false|false||administrationnull|Administration occupational activities|Event|false|false||administrationnull|impression (attitude)|Finding|false|false||IMPRESSION
null|EKG impression|Finding|false|false||IMPRESSIONnull|FLAIR (product)|Drug|false|false||FLAIR
null|FLAIR (product)|Drug|false|false||FLAIRnull|Fluid Attenuated Inversion Recovery|Procedure|false|false||FLAIRnull|Isointense|Finding|false|false||isointensenull|Lesion|Finding|false|false|C1660780|lesion
null|null|Finding|false|false|C1660780|lesionnull|midline cell component|Anatomy|false|false|C1546698;C0221198|midlinenull|Midline (qualifier value)|Modifier|false|false||midlinenull|Adenohypophyseal Diseases|Disorder|false|false||anteriornull|Anterior|Modifier|false|false||anteriornull|Posterior Pituitary Hormone Drug Class|Drug|false|false|C0447640;C0032009;C0032005|posterior pituitary
null|posterior pituitary hormones|Drug|false|false|C0447640;C0032009;C0032005|posterior pituitary
null|posterior pituitary hormones|Drug|false|false|C0447640;C0032009;C0032005|posterior pituitary
null|posterior pituitary hormones|Drug|false|false|C0447640;C0032009;C0032005|posterior pituitary
null|Posterior Pituitary Hormone Drug Class|Drug|false|false|C0447640;C0032009;C0032005|posterior pituitarynull|Pituitary Gland, Posterior|Anatomy|false|false|C0332148;C0750492;C3714635;C0032017;C0751438;C0032002|posterior pituitary
null|pars nervosa of hypophysis|Anatomy|false|false|C0332148;C0750492;C3714635;C0032017;C0751438;C0032002|posterior pituitarynull|Posterior pituitary disease|Disorder|false|false|C0447640;C0032009;C0032005|posteriornull|Dorsal|Modifier|false|false||posteriornull|Pituitary hormone preparation|Drug|false|false|C0032005|pituitary
null|Pituitary hormone preparation|Drug|false|false|C0032005|pituitary
null|Pituitary hormone preparation|Drug|false|false|C0032005|pituitarynull|Pituitary Diseases|Disorder|false|false|C0447640;C0032009;C0032005|pituitarynull|Pituitary Gland|Anatomy|false|false|C3714635;C0032017;C0032002;C0332148;C0750492;C0304812;C0751438|pituitarynull|Probable diagnosis|Finding|false|false|C0447640;C0032009;C0032005|likely
null|Probably|Finding|false|false|C0447640;C0032009;C0032005|likelynull|Cleaved|Modifier|false|false||cleftnull|Cyst|Disorder|false|false||cystnull|SpecimenType - Cyst|Finding|false|false||cyst
null|null|Finding|false|false||cystnull|Cyst form of protozoa|Entity|false|false||cystnull|Further|Modifier|false|false||Furthernull|Processing type - Evaluation|Finding|false|false||evaluationnull|Evaluation procedure|Procedure|false|false||evaluation
null|Evaluation|Procedure|false|false||evaluationnull|Pituitary hormone preparation|Drug|false|false|C0032005|pituitary
null|Pituitary hormone preparation|Drug|false|false|C0032005|pituitary
null|Pituitary hormone preparation|Drug|false|false|C0032005|pituitarynull|Pituitary Diseases|Disorder|false|false|C0032005|pituitarynull|Pituitary Gland|Anatomy|false|false|C0304812;C0032002|pituitarynull|BRIEF Health Literacy Screening Tool|Finding|false|false||Brief
null|Behavior Rating Inventory of Executive Function|Finding|false|false||Briefnull|Brief|Time|false|false||Briefnull|Shortened|Modifier|false|false||Briefnull|Hospital course|Finding|false|false||Hospital Coursenull|null|Attribute|false|false||Hospital Coursenull|Organization unit type - Hospital|Finding|false|false||Hospitalnull|Hospitals|Device|false|false||Hospitalnull|Hospitals|Entity|false|false||Hospitalnull|Hospital environment|Modifier|false|false||Hospitalnull|Course|Time|false|false||Coursenull|Worksheet|Finding|false|false||worksheetnull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|famotidine|Drug|false|false||famotidine
null|famotidine|Drug|false|false||famotidinenull|Daily|Time|false|false||dailynull|Contraceptive methods|Procedure|false|false||birth controlnull|Entity Name Part Qualifier - birth|Finding|false|false||birth
null|Childbirth|Finding|false|false||birth
null|birth (history)|Finding|false|false||birth
null|Name Given at Birth|Finding|false|false||birth
null|Birth|Finding|false|false||birthnull|Control brand of phenylpropanolamine|Drug|false|false||control
null|CONTROL veterinary product|Drug|false|false||control
null|control substance|Drug|false|false||control
null|Control brand of phenylpropanolamine|Drug|false|false||controlnull|Control - Relationship modifier|Finding|false|false||control
null|Control function|Finding|false|false||control
null|Scientific Control|Finding|false|false||controlnull|Control Groups|Subject|false|false||controlnull|True Control Status|Modifier|false|false||control
null|control aspects|Modifier|false|false||controlnull|Aunt|Subject|false|false||auntnull|microgram|LabModifier|false|false||mcgnull|Daily|Time|false|false||DAILYnull|famotidine|Drug|false|false||Famotidine
null|famotidine|Drug|false|false||Famotidinenull|Daily|Time|false|false||DAILYnull|metoprolol tartrate|Drug|false|false||Metoprolol Tartrate
null|metoprolol tartrate|Drug|false|false||Metoprolol Tartratenull|metoprolol|Drug|false|false||Metoprolol
null|metoprolol|Drug|false|false||Metoprololnull|tartrate|Drug|false|false||Tartrate
null|Tartrates|Drug|false|false||Tartrate
null|tartrate|Drug|false|false||Tartratenull|Daily|Time|false|false||DAILYnull|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin Drug Class|Drug|false|false||Multivitamins
null|Multivitamin Drug Class|Drug|false|false||Multivitaminsnull|Minerals|Drug|false|false||mineralsnull|Tablet Dosage Form|Drug|false|false||TABnull|Tablet Dosing Unit|LabModifier|false|false||TABnull|Daily|Time|false|false||DAILYnull|Once a day, at bedtime|Time|false|false||QHSnull|Entity|Entity|false|false||itemnull|Miscellaneous|Modifier|false|false||miscellaneousnull|Once - dosing instruction fragment|Finding|false|false||ONCEnull|Once (schedule frequency)|Time|false|false||ONCEnull|Forecast of outcome|Procedure|false|false||Prognosisnull|null|Attribute|false|false||Prognosisnull|Language Ability Proficiency - Good|Finding|false|false||Good
null|Language Proficiency - Good|Finding|false|false||Goodnull|Specimen Quality - Good|Modifier|false|false||Good
null|Good|Modifier|false|false||Goodnull|month|Time|false|false||monthsnull|PRSS30P gene|Finding|false|false||Dispnull|Dispense (activity)|Event|false|false||Dispnull|refill|Finding|false|false||Refillsnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|long-term care|Procedure|false|false||Extended Carenull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|In care (finding)|Finding|false|false||Care
null|Continuity Assessment Record and Evaluation|Finding|false|false||Carenull|care activity|Event|false|false||Carenull|ADMIN.FACILITY|Finding|false|false||Facilitynull|Facility (object)|Device|false|false||Facilitynull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Functional Relationship|Finding|false|false||Functional
null|Function (attribute)|Finding|false|false||Functional
null|Functional|Finding|false|false||Functionalnull|Neurologic (qualifier value)|Modifier|false|false||neurologicalnull|Syndrome|Disorder|false|false||syndromenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Disease|Disorder|false|false||Conditionnull|Logical Condition|Finding|false|false||Conditionnull|null|Attribute|false|false||Conditionnull|Condition|Modifier|false|false||Conditionnull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Lethargy|Finding|false|false||Lethargicnull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Coordination of Benefits - Independent|Finding|false|false||Independent
null|Religious Affiliation - Independent|Finding|false|false||Independent
null|Independence|Finding|false|false||Independent
null|Independently able|Finding|false|false||Independentnull|Discharge instructions|Finding|false|false||Discharge Instructionsnull|hospital discharge instructions (treatment)|Procedure|false|false||Discharge Instructionsnull|null|Attribute|false|false||Discharge Instructionsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructionsnull|FBXW7-AS1 gene|Finding|false|false||Dearnull|Production Class Code - Pleasure|Finding|false|false||pleasure
null|pleasurable emotion|Finding|false|false||pleasurenull|Pleasure - Animals raised for recreation|Entity|false|false||pleasurenull|care of - AddressPartType|Finding|false|false||care ofnull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Headache|Finding|false|false||headachenull|Lethargy|Finding|false|false||lethargynull|Weakness|Finding|false|false||weakness
null|Asthenia|Finding|false|false||weaknessnull|Iron Drug Class|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|Ferrum metallicum, Homeopathic preparation|Drug|false|false||ironnull|Iron measurement|Procedure|false|false||ironnull|Infusion route|Finding|false|false||infusionnull|Infusion procedures|Procedure|false|false||infusionnull|MDF AttributeType - Number|Finding|false|false||numbernull|Count of entities|LabModifier|false|false||number
null|Numbers|LabModifier|false|false||numbernull|Tests (qualifier value)|Finding|false|false||testsnull|Laboratory Procedures|Procedure|false|false||testsnull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Reassuring (procedure)|Procedure|false|false||reassuringnull|CYREN gene|Finding|false|false|C4266577;C0006104|MRInull|Magnetic resonance imaging service|Procedure|false|false|C4266577;C0006104|MRI
null|Magnetic Resonance Imaging|Procedure|false|false|C4266577;C0006104|MRInull|Maori Language|Entity|false|false||MRInull|Brain Diseases|Disorder|false|false|C4266577;C0006104|brainnull|Head>Brain|Anatomy|false|false|C0024485;C0587658;C1824234;C0006111|brain
null|Brain|Anatomy|false|false|C0024485;C0587658;C1824234;C0006111|brainnull|Evidence|Finding|true|false||evidencenull|Cerebrovascular accident|Disorder|false|false||strokenull|Stroke (heart beat)|Finding|false|false||strokenull|Inflammation|Finding|false|false||inflammationnull|Electroencephalography|Procedure|false|false|C4266577;C0006104|EEGnull|Brain Waves|Finding|false|false|C4266577;C0006104|brain wavesnull|Brain Diseases|Disorder|false|false|C4266577;C0006104|brainnull|Head>Brain|Anatomy|false|false|C0678909;C0006111;C0013819|brain
null|Brain|Anatomy|false|false|C0678909;C0006111;C0013819|brainnull|null|Phenomenon|false|false||wavesnull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Seizures|Finding|true|false||seizurenull|Weakness|Finding|false|false||weakness
null|Asthenia|Finding|false|false||weaknessnull|Course|Time|false|false||coursenull|Hospitalization|Procedure|false|false||hospitalizationnull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Strength (attribute)|Finding|false|false||strengthnull|Pharmaceutical Strength|LabModifier|false|false||strength
null|Physical Strength|LabModifier|false|false||strengthnull|Long Variable|Modifier|false|false||long
null|Long|Modifier|false|false||longnull|Hardness|Modifier|false|false||hardnull|Vitelliform Macular Dystrophy|Disorder|false|false||bestnull|BEST1 wt Allele|Finding|false|false||best
null|BEST1 gene|Finding|false|false||bestnull|best (quality)|Modifier|false|false||bestnull|Care team|Finding|false|false||Care Teamnull|null|Attribute|false|false||Care Teamnull|In care (finding)|Finding|false|false||Care
null|Continuity Assessment Record and Evaluation|Finding|false|false||Carenull|care activity|Event|false|false||Carenull|Team|Subject|false|false||Teamnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions