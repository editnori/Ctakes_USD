CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Pharmaceutical Preparations|Drug|false|false||MEDICINEnull|Medicine|Title|false|false||MEDICINEnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|sulfa|Drug|false|false||Sulfanull|Sulfonamide Anti-Infective Agents|Drug|false|false||Sulfonamide
null|Sulfonamide Anti-Infective Agents|Drug|false|false||Sulfonamide
null|Sulfonamides|Drug|false|false||Sulfonamide
null|Sulfonamides|Drug|false|false||Sulfonamide
null|Sulfonamide [EPC]|Drug|false|false||Sulfonamidenull|Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE|Drug|false|false||Antibiotics
null|Antibiotics|Drug|false|false||Antibiotics
null|Antibiotics, ophthalmologic|Drug|false|false||Antibiotics
null|Antibiotics, Gynecological|Drug|false|false||Antibiotics
null|antibiotics, intestinal|Drug|false|false||Antibiotics
null|Antibiotic throat preparations|Drug|false|false||Antibiotics
null|Antibiotics, Antitubercular|Drug|false|false||Antibiotics
null|Antibiotics for systemic use|Drug|false|false||Antibiotics
null|Antifungal Antibiotics, Topical|Drug|false|false||Antibioticsnull|codeine|Drug|false|false||Codeine
null|codeine|Drug|false|false||Codeinenull|Bactrim|Drug|false|false||Bactrim
null|Bactrim|Drug|false|false||Bactrimnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Chief complaint (finding)|Finding|false|false||Chief Complaintnull|Complaint (finding)|Finding|false|false||Complaintnull|null|Attribute|false|false||Complaintnull|Weakness|Finding|false|false||Weakness
null|Asthenia|Finding|false|false||Weaknessnull|Nausea and vomiting|Finding|false|false||nausea/vomitingnull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|Vomiting|Finding|false|false||vomitingnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|History of present illness (finding)|Finding|false|false||History of Present Illnessnull|null|Attribute|false|false||History of Present Illnessnull|Medical History|Finding|false|false||History ofnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Present illness|Finding|false|false||Present Illnessnull|Present|Finding|false|false||Present
null|Presentation|Finding|false|false||Presentnull|Illness (finding)|Finding|false|false||Illnessnull|Recent|Time|false|false||recentlynull|Metastatic malignant neoplasm|Disorder|false|false||metastatic cancer
null|Disseminated Malignant Neoplasm|Disorder|false|false||metastatic cancer
null|Neoplasm Metastasis|Disorder|false|false||metastatic cancernull|metastatic qualifier|Finding|false|false||metastatic
null|Metastatic to|Finding|false|false||metastaticnull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|unknown vaccine or immune globulin|Drug|false|false||unknown
null|Unknown - Vaccines administered|Drug|false|false||unknown
null|Unknown - Vaccines administered|Drug|false|false||unknown
null|unknown vaccine or immune globulin|Drug|false|false||unknownnull|Unknown - Patient_s Relationship to Insured|Finding|false|false||unknown
null|Unknown - Special Program Code|Finding|false|false||unknown
null|Unknown - Production Class Code|Finding|false|false||unknown
null|Unknown - Patient Outcome|Finding|false|false||unknown
null|Unknown - Recreational Drug Use Code|Finding|false|false||unknown
null|Unknown - Escort Required|Finding|false|false||unknown
null|Unknown - Transport Arranged|Finding|false|false||unknown
null|Unknown - Living Arrangement|Finding|false|false||unknown
null|Unknown - Employment Status|Finding|false|false||unknown
null|Unknown - Relationship|Finding|false|false||unknown
null|Unknown - publishing section|Finding|false|false||unknown
null|Unknown Publicity Code|Finding|false|false||unknown
null|Unknown - Event reason|Finding|false|false||unknown
null|Unknown - Religion|Finding|false|false||unknown
null|Unknown - Organ Donor Code|Finding|false|false||unknown
null|unknown - NullFlavor|Finding|false|false||unknown
null|Unknown - Notify Clergy Code|Finding|false|false||unknown
null|Unknown - Administrative Gender|Finding|false|false||unknown
null|Unknown - Patient Condition Code|Finding|false|false||unknown
null|Unknown - Living Will Code|Finding|false|false||unknown
null|Marital Status - Unknown|Finding|false|false||unknown
null|Unknown - mode of arrival code|Finding|false|false||unknown
null|Unknown - Patient Class|Finding|false|false||unknown
null|Unknown - Event Expected|Finding|false|false||unknown
null|Unknown - Expanded yes/no indicator|Finding|false|false||unknown
null|Unknown - Immunization Registry Status|Finding|false|false||unknown
null|Unknown - Container status|Finding|false|false||unknown
null|Unknown - CWE statuses|Finding|false|false||unknown
null|Unknown - Job Status|Finding|false|false||unknown
null|Unknown - Precaution Code|Finding|false|false||unknown
null|Unknown - Contact Role|Finding|false|false||unknown
null|Unknown - Living Dependency|Finding|false|false||unknownnull|Ethnic group unknown|Subject|false|false||unknownnull|Unknown - Allergy Severity|Modifier|false|false||unknown
null|Unknown - HL7 update mode|Modifier|false|false||unknown
null|Unknown|Modifier|false|false||unknownnull|null|Time|false|false||priornull|Presentation|Finding|false|false||presentingnull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|Vomiting|Finding|false|false||vomitingnull|Fever symptoms (finding)|Finding|false|false||fever
null|Fever|Finding|false|false||fevernull|Has patient|Finding|false|false||Patient hasnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Vomiting|Finding|false|false||vomitingnull|week|Time|false|false||weeksnull|Metastatic malignant neoplasm|Disorder|false|false||metastatic cancer
null|Disseminated Malignant Neoplasm|Disorder|false|false||metastatic cancer
null|Neoplasm Metastasis|Disorder|false|false||metastatic cancernull|metastatic qualifier|Finding|false|false||metastatic
null|Metastatic to|Finding|false|false||metastaticnull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Upper abdomen (surface region)|Anatomy|false|false|C0153662;C1512806;C4723750;C1547310;C0941288;C4521161;C3251814;C3641766|upper abdomen
null|Upper abdomen structure|Anatomy|false|false|C0153662;C1512806;C4723750;C1547310;C0941288;C4521161;C3251814;C3641766|upper abdomennull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|Abdomen|Anatomy|false|false|C4723750;C1547310;C0153662;C0941288;C3641766;C4521161;C3251814|abdomen andnull|Malignant neoplasm of abdomen|Disorder|false|false|C2937240;C0230165;C0000726;C0230168;C0000726|abdomennull|Abdomen problem|Finding|false|false|C0230168;C0000726;C0000726;C2937240;C0230165|abdomennull|Abdomen|Anatomy|false|false|C0941288;C4521161;C3251814;C0153662;C4723750;C1547310;C3641766|abdomen
null|Abdominal Cavity|Anatomy|false|false|C0941288;C4521161;C3251814;C0153662;C4723750;C1547310;C3641766|abdomennull|Very Poor|Finding|false|false|C0000726;C2937240;C0230165;C0230168;C0000726|very poornull|Very|Modifier|false|false||verynull|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group|Finding|false|false|C0000726;C2937240;C0230165;C0230168;C0000726|poor
null|Patient Condition Code - Poor|Finding|false|false|C0000726;C2937240;C0230165;C0230168;C0000726|poornull|Poverty|Subject|false|false||poornull|Language Proficiency - Poor|Modifier|false|false||poor
null|Specimen Quality - Poor|Modifier|false|false||poor
null|Poor - grade|Modifier|false|false||poor
null|Poor - qualifier|Modifier|false|false||poornull|Intake|Finding|false|false|C2937240;C0230165|intakenull|Measurement of fluid intake|Procedure|false|false|C0230168;C0000726;C2937240;C0230165;C0000726|intake
null|Intake (treatment)|Procedure|false|false|C0230168;C0000726;C2937240;C0230165;C0000726|intakenull|Feel Weak (question)|Finding|false|false||weak
null|Weakness|Finding|false|false||weaknull|Weak|Modifier|false|false||weaknull|Time periods|Time|false|false||time periodnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Menstruation|Finding|false|false||periodnull|Clinical Trial Period|Procedure|false|false||periodnull|per period (qualifier value)|Time|false|false||period
null|Time periods|Time|false|false||periodnull|Transaction counts and value totals - Period|LabModifier|false|false||periodnull|Vomiting|Finding|false|false||vomitingnull|Abdominal Pain|Finding|false|false|C0000726|abdominal painnull|Abdomen|Anatomy|false|false|C0000737;C1549543;C0030193|abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Administration Method - Pain|Finding|false|false|C0000726|pain
null|Pain|Finding|false|false|C0000726|painnull|null|Attribute|false|false||painnull|week|Time|false|false||weeksnull|More|LabModifier|false|false||morenull|Fatigue|Finding|false|false||fatiguednull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Upper Respiratory Infections|Disorder|false|false||URInull|Uniform Resource Identifier|Finding|false|false||URI
null|URI1 gene|Finding|false|false||URI
null|URI1 wt Allele|Finding|false|false||URInull|Symptoms aspect|Finding|true|false||symptoms
null|Symptoms|Finding|true|false||symptomsnull|Urinary tract|Anatomy|false|false||urinarynull|urinary|Modifier|false|false||urinarynull|Complaint (finding)|Finding|false|false||complaintsnull|Constipation|Finding|false|false||constipatednull|Antiemetics|Drug|false|false||anti-emeticsnull|Last|Modifier|false|false||Lastnull|Defecation|Finding|false|false|C0021853|bowel movementnull|Intestines|Anatomy|false|false|C0011135|bowelnull|Movement|Finding|false|false||movementnull|Gas - SpecimenType|Drug|false|false||gas
null|Gases|Drug|false|false||gas
null|Gas Dosage Form|Drug|false|false||gasnull|Gas - Specimen Source Codes|Finding|false|false||gas
null|gastrointestinal gas|Finding|false|false||gas
null|PAGR1 wt Allele|Finding|false|false||gas
null|GALNS wt Allele|Finding|false|false||gas
null|GALNS gene|Finding|false|false||gas
null|GAST wt Allele|Finding|false|false||gas
null|GAST gene|Finding|false|false||gas
null|germacrene-A synthase activity|Finding|false|false||gas
null|PAGR1 gene|Finding|false|false||gasnull|Edema of lower extremity|Finding|false|false|C0023216;C1548802;C0015385|lower extremity edemanull|Lower Extremity|Anatomy|false|false|C0239340;C0085649;C0013604|lower extremitynull|Body Site Modifier - Lower|Anatomy|false|false|C0085649;C0239340;C2003888|lowernull|Lower (action)|Event|false|false|C1548802|lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Peripheral edema|Finding|false|false|C1548802;C0023216;C0015385|extremity edemanull|Limb structure|Anatomy|false|false|C0013604;C0085649;C0239340|extremitynull|Edema|Finding|false|false|C0023216;C0015385|edemanull|null|Attribute|false|false||edemanull|Present|Finding|false|false||present
null|Presentation|Finding|false|false||presentnull|Several|LabModifier|false|false||severalnull|week|Time|false|false||weeksnull|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|liver
null|liver extract|Drug|false|false|C4037986;C1278929;C0023884|liver
null|liver extract|Drug|false|false|C4037986;C1278929;C0023884|liver
null|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|liver
null|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|livernull|Benign neoplasm of liver|Disorder|false|false|C4037986;C1278929;C0023884|liver
null|Liver diseases|Disorder|false|false|C4037986;C1278929;C0023884|livernull|Liver problem|Finding|false|false|C4037986;C1278929;C0023884|livernull|Procedures on liver|Procedure|false|false|C4037986;C1278929;C0023884|livernull|Abdomen>Liver|Anatomy|false|false|C0023895;C0496870;C0577060;C0721399;C0023899;C0872387;C1705694;C0812270|liver
null|null|Anatomy|false|false|C0023895;C0496870;C0577060;C0721399;C0023899;C0872387;C1705694;C0812270|liver
null|Liver|Anatomy|false|false|C0023895;C0496870;C0577060;C0721399;C0023899;C0872387;C1705694;C0812270|livernull|ETV3 wt Allele|Finding|false|false|C4037986;C1278929;C0023884|mets
null|ETV3 gene|Finding|false|false|C4037986;C1278929;C0023884|metsnull|Several|LabModifier|false|false||severalnull|week|Time|false|false||weeksnull|ibuprofen|Drug|false|false||ibuprofen
null|ibuprofen|Drug|false|false||ibuprofennull|biopsy characteristics|Finding|false|false||biopsy
null|null|Finding|false|false||biopsynull|Biopsy Procedures on the Pharynx, Adenoids, and Tonsils|Procedure|false|false||biopsy
null|Biopsy|Procedure|false|false||biopsy
null|Consent Type - biopsy|Procedure|false|false||biopsynull|Initial (abbreviation)|Finding|false|false||initialnull|Initially|Time|false|false||initialnull|Firstly|Modifier|false|false||initialnull|Laboratory test finding|Lab|false|false||Labsnull|Significant|Finding|false|false|C0023516|significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|Leukocytes|Anatomy|false|false|C0750502|WBCnull|5'-Inosinic acid, 2'-deoxy-2'-fluoro-, homopolymer|Drug|false|false||polys
null|Poly A|Drug|false|false||polysnull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|Ketones|Drug|false|false||ketonesnull|Toxic effect of ketones|Disorder|false|false||ketonesnull|Ketone bodies measurement, quantitative|Procedure|false|false||ketones
null|Urine ketone test|Procedure|false|false||ketonesnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Zofran|Drug|false|false||zofran
null|Zofran|Drug|false|false||zofrannull|Plain chest X-ray|Procedure|false|false||CXRnull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|Left sided|Modifier|false|false||left sided
null|Left|Modifier|false|false||left sidednull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Abnormally opaque structure (morphologic abnormality)|Finding|false|false||opacity
null|Decreased translucency|Finding|false|false||opacitynull|Peptide Nucleic Acids|Drug|false|false||PNAnull|metastatic qualifier|Finding|false|false||metastatic
null|Metastatic to|Finding|false|false||metastaticnull|diseae|Entity|false|false||diseaenull|Smear - instruction imperative|Event|false|false||spreadnull|Spreading (qualifier value)|Modifier|false|false||spreadnull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|cefepime|Drug|false|false||cefepime
null|cefepime|Drug|false|false||cefepimenull|Pneumonia|Disorder|false|false||pneumonianull|Transfer - product ownership|Finding|false|false||transfer
null|Transfer Technique|Finding|false|false||transfer
null|ActClass - transfer|Finding|false|false||transfer
null|null|Finding|false|false||transfernull|Transfer (immobility management)|Procedure|false|false||transfernull|Current (present time)|Time|false|false||Currentlynull|Feel Weak (question)|Finding|false|false||feel weak
null|Weakness|Finding|false|false||feel weaknull|Feel Weak (question)|Finding|false|false||weak
null|Weakness|Finding|false|false||weaknull|Weak|Modifier|false|false||weaknull|Nausea|Finding|false|false||nauseousnull|C22orf39 gene|Finding|false|false||pantsnull|Underpants|Device|false|false||pants
null|Trousers|Device|false|false||pantsnull|Feel Weak (question)|Finding|false|false||weak
null|Weakness|Finding|false|false||weaknull|Weak|Modifier|false|false||weaknull|Feel Tired question|Finding|false|false||tired
null|Fatigue|Finding|false|false||tired
null|Feeling tired|Finding|false|false||tirednull|Review of systems (procedure)|Procedure|false|false||REVIEW OF SYSTEMSnull|null|Attribute|false|false||REVIEW OF SYSTEMS
null|null|Attribute|false|false||REVIEW OF SYSTEMSnull|Review of|Finding|false|false||REVIEW OFnull|Review (Publication Type)|Finding|false|false||REVIEW
null|Act Class - review|Finding|false|false||REVIEWnull|System|Finding|false|false||SYSTEMSnull|Proline dehydrogenase deficiency|Disorder|false|false||HPInull|History of present illness (finding)|Finding|false|false||HPI
null|allene oxide synthase activity|Finding|false|false||HPInull|Night sweats|Finding|false|false||night sweatsnull|Night time|Time|false|false||nightnull|Sweating|Finding|false|false||sweats
null|Sweat|Finding|false|false||sweatsnull|Headache|Finding|false|false||headachenull|Vision|Finding|false|false||visionnull|null|Attribute|false|false||visionnull|Specialized Stand Alone Plan - Vision|Entity|false|false||visionnull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|Rhinorrhea|Finding|false|false||rhinorrheanull|Congestion|Finding|false|false||congestionnull|Sore Throat brand of benzocaine & menthol|Drug|false|false|C0230069;C3665375;C0031354|sore throat
null|Sore Throat brand of Phenol|Drug|false|false|C0230069;C3665375;C0031354|sore throat
null|Sore Throat brand of Phenol|Drug|false|false|C0230069;C3665375;C0031354|sore throat
null|Sore Throat brand of benzocaine & menthol|Drug|false|false|C0230069;C3665375;C0031354|sore throatnull|Pharyngitis|Disorder|false|false|C0230069;C3665375;C0031354|sore throatnull|Sore Throat|Finding|false|false|C0230069;C3665375;C0031354|sore throatnull|Sore to touch|Finding|false|false||sore
null|Sore skin|Finding|false|false||sorenull|Sore sensation quality|Modifier|false|false||sorenull|Throat Homeopathic Medication|Drug|false|false|C0230069;C3665375;C0031354|throatnull|Specimen Type - Throat|Finding|false|false|C0230069;C3665375;C0031354|throat
null|null|Finding|false|false|C0230069;C3665375;C0031354|throatnull|Throat|Anatomy|false|false|C0018932;C1550663;C1547926;C3244654;C0723402;C1950455;C0031350;C0242429|throat
null|Anterior portion of neck|Anatomy|false|false|C0018932;C1550663;C1547926;C3244654;C0723402;C1950455;C0031350;C0242429|throat
null|Pharyngeal structure|Anatomy|false|false|C0018932;C1550663;C1547926;C3244654;C0723402;C1950455;C0031350;C0242429|throatnull|Hematochezia|Disorder|false|false|C0230069;C3665375;C0031354|BRBPRnull|Melena|Finding|false|false||melenanull|Hematochezia|Disorder|false|false||hematochezianull|Blood in stool|Finding|false|false||hematochezianull|Dysuria|Finding|false|false||dysurianull|Hematuria|Disorder|false|false||hematurianull|PMH - past medical history|Finding|false|false||Past Medical History
null|Medical History|Finding|false|false||Past Medical Historynull|Medical History|Finding|false|false||Medical Historynull|Medical referral type|Finding|false|false||Medical
null|Medical|Finding|false|false||Medical
null|Medical school type|Finding|false|false||Medicalnull|Medical service|Procedure|false|false||Medicalnull|Medical History|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|History of present illness (finding)|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|PMH - past medical history|Finding|false|false||PMH
null|Medical History|Finding|false|false||PMHnull|Enneking High Surgical Grade|Finding|false|false||high grade
null|Severe (severity modifier)|Finding|false|false||high gradenull|Message Waiting Priority - High|Finding|false|false||high
null|high - ActExposureLevelCode|Finding|false|false||high
null|IPSS Risk Category High|Finding|false|false||high
null|IPSS-R Risk Category High|Finding|false|false||high
null|High (finding)|Finding|false|false||highnull|Observation Value - High|Modifier|false|false||high
null|High|Modifier|false|false||high
null|Abnormally high|Modifier|false|false||highnull|Histopathologic Grade|Finding|false|false||grade
null|Grade|Finding|false|false||grade
null|School Grade|Finding|false|false||gradenull|Exploratory laparotomy|Procedure|false|false||exploratory laparotomynull|Laparotomy|Procedure|false|false||laparotomynull|Lysis|Finding|false|false||lysis
null|pathologic cytolysis|Finding|false|false||lysisnull|Tissue Adhesions|Finding|false|false||adhesionsnull|Small intestine excision|Procedure|false|false|C4319010;C0021852;C0021853|small bowel resectionnull|Abdomen>Small bowel|Anatomy|false|false|C0741614;C0015252;C0728940;C0192601|small bowel
null|Intestines, Small|Anatomy|false|false|C0741614;C0015252;C0728940;C0192601|small bowelnull|Small|LabModifier|false|false||smallnull|Bowel resection|Procedure|false|false|C0021853;C4319010;C0021852|bowel resectionnull|Intestines|Anatomy|false|false|C0741614;C0192601|bowelnull|removal technique|Procedure|false|false|C4319010;C0021852|resection
null|Excision|Procedure|false|false|C4319010;C0021852|resectionnull|Anastomosis of small intestine to small intestine|Procedure|false|false||enteroenterostomy
null|Anastomosis of intestine|Procedure|false|false||enteroenterostomynull|Carcinoid Tumor|Disorder|false|false||carcinoidnull|Hyperlipidemia|Disorder|false|false||hyperlipidemia
null|Hyperlipoproteinemias|Disorder|false|false||hyperlipidemianull|Serum lipids high (finding)|Finding|false|false||hyperlipidemianull|Vitamin B 12 Deficiency|Disorder|false|false||vitamin B12 deficiencynull|Decreased circulating vitamin B12 concentration|Finding|false|false||vitamin B12 deficiencynull|Vitamin B12 [EPC]|Drug|false|false||vitamin B12
null|cobalamins|Drug|false|false||vitamin B12
null|cobalamins|Drug|false|false||vitamin B12
null|vitamin B12|Drug|false|false||vitamin B12
null|vitamin B12|Drug|false|false||vitamin B12
null|vitamin B12|Drug|false|false||vitamin B12null|VITAMIN B12 MEASUREMENT|Procedure|false|false||vitamin B12null|Vitamins|Drug|false|false||vitamin
null|Vitamins|Drug|false|false||vitamin
null|Vitamins|Drug|false|false||vitaminnull|TNFAIP1 wt Allele|Finding|false|false||B12
null|NDUFB3 gene|Finding|false|false||B12
null|TNFAIP1 gene|Finding|false|false||B12null|Malnutrition|Disorder|false|false||deficiencynull|Deficiency|Finding|false|false||deficiencynull|deficiency aspects|Modifier|false|false||deficiencynull|Neck|Anatomy|false|false|C0029408|cervicalnull|Cervical|Modifier|false|false||cervicalnull|Degenerative polyarthritis|Disorder|false|false|C0027530|DJDnull|Degenerative polyarthritis|Disorder|false|false||osteoarthritisnull|Lung excision|Procedure|false|false|C4037972;C0024109|lung resectionnull|Lung diseases|Disorder|false|false|C4037972;C0024109|lungnull|Lung Problem|Finding|false|false|C4037972;C0024109|lungnull|Chest>Lung|Anatomy|false|false|C0024115;C0396565;C0740941|lung
null|Lung|Anatomy|false|false|C0024115;C0396565;C0740941|lungnull|removal technique|Procedure|false|false||resection
null|Excision|Procedure|false|false||resectionnull|Consent Type - Hysterectomy|Finding|false|false||hysterectomynull|Hysterectomy|Procedure|false|false||hysterectomynull|Right arm|Anatomy|false|false|C1522541;C5400986;C4761640;C1824218;C3715044;C0543467;C3495676;C0038895;C1457907;C1547138|R armnull|Anorectal Malformations|Disorder|false|false|C0446516;C1140618;C1269078;C4048756|armnull|AKR1A1 wt Allele|Finding|false|false|C0446516;C1140618;C1269078;C4048756|arm
null|ARMC9 gene|Finding|false|false|C0446516;C1140618;C1269078;C4048756|armnull|Protocol Treatment Arm|Procedure|false|false|C4048756;C0446516;C1140618;C1269078|arm
null|Axillary Reverse Mapping|Procedure|false|false|C4048756;C0446516;C1140618;C1269078|arm
null|Study Arm|Procedure|false|false|C4048756;C0446516;C1140618;C1269078|armnull|Upper arm|Anatomy|false|false|C1824218;C3715044;C3495676;C1522541;C5400986;C4761640|arm
null|null|Anatomy|false|false|C1824218;C3715044;C3495676;C1522541;C5400986;C4761640|arm
null|Upper Extremity|Anatomy|false|false|C1824218;C3715044;C3495676;C1522541;C5400986;C4761640|armnull|Level of Care - Surgery|Finding|false|false|C4048756|surgery
null|Surgical procedure finding|Finding|false|false|C4048756|surgery
null|Surgical aspects|Finding|false|false|C4048756|surgerynull|Operative Surgical Procedures|Procedure|false|false|C4048756|surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Social and personal history|Finding|false|false||Social History
null|Social History|Finding|false|false||Social Historynull|Social|Finding|false|false||Socialnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Family Medical History|Finding|false|false||Family Historynull|Entity Name Part Type - family|Finding|false|false||Family
null|Last Name|Finding|false|false||Family
null|Living Arrangement - Family|Finding|false|false||Family
null|Family (taxonomic)|Finding|false|false||Family
null|Family Collection|Finding|false|false||Familynull|Family|Subject|false|false||Familynull|History of present illness (finding)|Finding|false|true||History
null|History of previous events|Finding|false|true||History
null|Historical aspects qualifier|Finding|false|true||History
null|Medical History|Finding|false|true||History
null|Concept History|Finding|false|true||Historynull|History|Subject|false|false||Historynull|Relationship - Mother|Finding|false|false||Mothernull|Mother (person)|Subject|false|false||Mothernull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Youngest|Modifier|false|false||Youngestnull|In Touch|Device|false|false||in touchnull|Touch Perception|Finding|false|false||touch
null|Touch sensation|Finding|false|false||touchnull|Therapeutic Touch|Procedure|false|false||touchnull|Tactile|Modifier|false|false||touchnull|Sibling|Subject|false|false||siblingsnull|Indirect exposure mechanism - Father|Finding|false|false||Father
null|Relationship - Father|Finding|false|false||Father
null|Father - courtesy title|Finding|false|false||Fathernull|Father (person)|Subject|false|false||Fathernull|physical examination (physical finding)|Finding|false|false||Physical Examnull|Physical Examination|Procedure|false|false||Physical Examnull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|physical examination (physical finding)|Finding|false|false||Physical Examnull|Physical Examination|Procedure|false|false||Physical Examnull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||GENERALnull|General medical service|Procedure|false|false||GENERALnull|Generalized|Modifier|false|false||GENERALnull|Obesity|Disorder|false|false||Obesenull|Woman|Subject|false|false||woman
null|Human, Female adult|Subject|false|false||womannull|Feeling comfortable|Finding|false|false||comfortablenull|patient appears in no acute distress (physical finding)|Finding|false|false||in no acute distressnull|Admission Level of Care Code - Acute|Finding|true|false||acute
null|Acute - Triage Code|Finding|true|false||acutenull|acute|Time|false|false||acutenull|Emotional distress|Finding|true|false||distress
null|Distress|Finding|true|false||distressnull|HEENT|Anatomy|false|false||HEENTnull|PERRLA|Finding|false|false||PERRLAnull|Anicteric|Finding|false|false||anictericnull|Slightly (qualifier value)|Modifier|false|false||slightly
null|Slight (qualifier value)|Modifier|false|false||slightlynull|Mucus (substance)|Finding|false|false||mucus
null|mucus layer|Finding|false|false||mucus
null|null|Finding|false|false||mucusnull|Membrane Tissue|Anatomy|false|false||membranesnull|Passive joint movement of neck (finding)|Finding|false|false|C0027530;C3159206|NECK
null|Neck problem|Finding|false|false|C0027530;C3159206|NECKnull|dendritic spine neck|Anatomy|false|false|C0812434;C0684335|NECK
null|Neck|Anatomy|false|false|C0812434;C0684335|NECKnull|Supple|Finding|false|false||supplenull|Obesity|Disorder|false|false||obesenull|Lung|Anatomy|false|false||LUNGSnull|Distant Metastasis|Finding|false|false||Distantnull|Distant|Modifier|false|false||Distantnull|null|Attribute|false|false||breath sounds
null|Respiratory Sounds|Attribute|false|false||breath soundsnull|Breath|Finding|false|false||breathnull|null|Device|false|false||soundsnull|null|Phenomenon|false|false||soundsnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Basilar Rales|Finding|false|false||crackles
null|Rales|Finding|false|false||cracklesnull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787|HEART
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787|HEARTnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|HEARTnull|Chest>Heart|Anatomy|false|false|C0795691;C0153957;C0153500|HEART
null|Heart|Anatomy|false|false|C0795691;C0153957;C0153500|HEARTnull|MAS1L gene|Finding|true|false||MRGnull|Malignant neoplasm of abdomen|Disorder|false|false|C0230168;C0000726|ABDOMENnull|Abdomen problem|Finding|false|false|C0230168;C0000726|ABDOMENnull|Abdomen|Anatomy|false|false|C0153662;C0941288|ABDOMEN
null|Abdominal Cavity|Anatomy|false|false|C0153662;C0941288|ABDOMENnull|Bowel sounds|Finding|false|false|C0021853|bowel soundsnull|Intestines|Anatomy|false|false|C0232693|bowelnull|null|Device|false|false||soundsnull|null|Phenomenon|false|false||soundsnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||softnull|Soft|Modifier|false|false||softnull|Epigastric|Anatomy|false|false||epigastricnull|Structure of right upper quadrant of abdomen|Anatomy|false|false|C0684239;C0234233|RUQnull|RUQ - Right upper quadrant|Modifier|false|false||RUQnull|Emotional tenderness|Finding|false|false|C0230177|tenderness
null|Sore to touch|Finding|false|false|C0230177|tendernessnull|Palpation|Procedure|false|false||palpationnull|Massive|Modifier|false|false||markedlynull|Hepatomegaly|Finding|false|false|C4037986;C1278929;C0023884|enlarged livernull|Enlargement procedure|Procedure|false|false||enlargednull|Enlarged|Modifier|false|false||enlargednull|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|liver
null|liver extract|Drug|false|false|C4037986;C1278929;C0023884|liver
null|liver extract|Drug|false|false|C4037986;C1278929;C0023884|liver
null|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|liver
null|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|livernull|Benign neoplasm of liver|Disorder|false|false|C4037986;C1278929;C0023884|liver
null|Liver diseases|Disorder|false|false|C4037986;C1278929;C0023884|livernull|Liver problem|Finding|false|false|C4037986;C1278929;C0023884|livernull|Procedures on liver|Procedure|false|false|C4037986;C1278929;C0023884|livernull|Abdomen>Liver|Anatomy|false|false|C0019209;C0872387;C0577060;C0721399;C0023899;C0023895;C0496870|liver
null|null|Anatomy|false|false|C0019209;C0872387;C0577060;C0721399;C0023899;C0023895;C0496870|liver
null|Liver|Anatomy|false|false|C0019209;C0872387;C0577060;C0721399;C0023899;C0023895;C0496870|livernull|Liver edge palpable|Finding|false|false|C4037986;C1278929;C0023884|liver edge palpablenull|Liver edge|Finding|false|false|C4037986;C1278929;C0023884|liver edgenull|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|liver
null|liver extract|Drug|false|false|C4037986;C1278929;C0023884|liver
null|liver extract|Drug|false|false|C4037986;C1278929;C0023884|liver
null|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|liver
null|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|livernull|Benign neoplasm of liver|Disorder|false|false|C4037986;C1278929;C0023884|liver
null|Liver diseases|Disorder|false|false|C4037986;C1278929;C0023884|livernull|Liver problem|Finding|false|false|C4037986;C1278929;C0023884|livernull|Procedures on liver|Procedure|false|false|C4037986;C1278929;C0023884|livernull|Abdomen>Liver|Anatomy|false|false|C0721399;C0023899;C0023895;C0496870;C0577060;C0426690;C0426689;C0872387|liver
null|null|Anatomy|false|false|C0721399;C0023899;C0023895;C0496870;C0577060;C0426690;C0426689;C0872387|liver
null|Liver|Anatomy|false|false|C0721399;C0023899;C0023895;C0496870;C0577060;C0426690;C0426689;C0872387|livernull|Graph Edge|Finding|false|false||edgenull|Along edge (qualifier value)|Modifier|false|false||edgenull|Palpable|Modifier|false|false||palpablenull|Rib Cage|Anatomy|false|false|C4555210;C5552712;C1426669|rib cagenull|Bone structure of rib|Anatomy|false|false|C1426669;C5552712|ribnull|CAGE Antibody|Drug|false|false|C0222762|cage
null|CAGE Antibody|Drug|false|false|C0222762|cage
null|CAGE Antibody|Drug|false|false|C0222762|cagenull|DDX53 gene|Finding|false|false|C0222762;C0035561|cagenull|CAP Analysis of Gene Expression|Procedure|false|false|C0222762;C0035561|cagenull|Spinal cage|Device|false|false||cage
null|null|Device|false|false||cagenull|Protective muscle spasm|Finding|true|false||guardingnull|All extremities|Anatomy|false|false||EXTREMITIES
null|Limb structure|Anatomy|false|false||EXTREMITIESnull|Edema of lower extremity|Finding|false|false|C1548802;C0015385;C0023216|lower extremity edemanull|Lower Extremity|Anatomy|false|false|C0085649;C0013604;C0239340|lower extremitynull|Body Site Modifier - Lower|Anatomy|false|false|C0239340;C2003888;C0013604;C0085649|lowernull|Lower (action)|Event|false|false|C1548802|lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Peripheral edema|Finding|false|false|C0015385;C0023216;C1548802|extremity edemanull|Limb structure|Anatomy|false|false|C0085649;C0239340;C0013604|extremitynull|Edema|Finding|false|false|C1548802;C0015385;C0023216|edemanull|null|Attribute|false|false||edemanull|null|Finding|false|false||pulses radialnull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false||pulsesnull|Radial|Finding|false|false||radial
null|Circumpennate|Finding|false|false||radialnull|Neurology speciality|Title|false|false||NEUROnull|Neurologic (qualifier value)|Modifier|false|false||NEUROnull|Awake (finding)|Finding|false|false||awakenull|Awakening (time frame)|Time|false|false||awakenull|Central Nervous System|Anatomy|false|false||CNsnull|Clinical Nurse Specialists|Subject|false|false||CNsnull|Certified Nurse Specialist|Title|false|false||CNsnull|Staphylococcus, coagulase negative (organism)|Entity|false|false||CNsnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Muscle Strength|Finding|false|false|C4083049;C0026845|muscle strengthnull|null|Attribute|false|false|C4083049;C0026845|muscle strengthnull|Muscle (organ)|Anatomy|false|false|C0808080;C0517349;C4050373|muscle
null|Muscle Tissue|Anatomy|false|false|C0808080;C0517349;C4050373|musclenull|Strength (attribute)|Finding|false|false|C4083049;C0026845|strengthnull|Pharmaceutical Strength|LabModifier|false|false||strength
null|Physical Strength|LabModifier|false|false||strengthnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|physical examination (physical finding)|Finding|false|false||Physical Examnull|Physical Examination|Procedure|false|false||Physical Examnull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||Generalnull|General medical service|Procedure|false|false||Generalnull|Generalized|Modifier|false|false||Generalnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Admission Level of Care Code - Acute|Finding|true|false||acute
null|Acute - Triage Code|Finding|true|false||acutenull|acute|Time|false|false||acutenull|Emotional distress|Finding|true|false||distress
null|Distress|Finding|true|false||distressnull|Obesity|Disorder|false|false||obesenull|Woman|Subject|false|false||woman
null|Human, Female adult|Subject|false|false||womannull|HEENT|Anatomy|false|false|C2228481;C0036412|HEENTnull|Scleral Diseases|Disorder|false|false|C0036410;C1512338|Scleranull|examination of sclera|Procedure|false|false|C0036410;C1512338|Scleranull|Sclera|Anatomy|false|false|C2228481;C0036412;C0205180|Scleranull|Anicteric|Finding|false|false|C0036410|anictericnull|Myelofibrosis|Disorder|false|false|C0694605|MMMnull|Medial part of medial mammillary nucleus|Anatomy|false|false|C0026987|MMMnull|Oropharyngeal|Anatomy|false|false|C1550016|oropharynxnull|Remote control command - Clear|Finding|false|false|C0521367|clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|Passive joint movement of neck (finding)|Finding|false|false|C0027530;C3159206|Neck
null|Neck problem|Finding|false|false|C0027530;C3159206|Necknull|dendritic spine neck|Anatomy|false|false|C5550999;C0398738;C0428897;C0332254;C0812434;C0684335;C1414063;C1706333|Neck
null|Neck|Anatomy|false|false|C5550999;C0398738;C0428897;C0332254;C0812434;C0684335;C1414063;C1706333|Necknull|Supple|Finding|false|false|C0027530;C3159206|supplenull|Jugular venous pressure|Finding|false|false|C0027530;C3159206|JVPnull|Elevated|Modifier|false|false||elevated
null|High|Modifier|false|false||elevatednull|Leukocyte adhesion deficiency type 1|Disorder|true|false|C0027530;C3159206;C0226032|LAD
null|Leukocyte adhesion deficiency|Disorder|true|false|C0027530;C3159206;C0226032|LADnull|ITGB2 wt Allele|Finding|true|false|C0226032;C0027530;C3159206|LAD
null|DLD gene|Finding|true|false|C0226032;C0027530;C3159206|LADnull|Anterior descending branch of left coronary artery|Anatomy|true|false|C1414063;C1706333;C5550999;C0398738|LADnull|Ladino Language|Entity|true|false||LADnull|Lung|Anatomy|false|false|C1550016|Lungsnull|Remote control command - Clear|Finding|false|false|C0024109|Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Auscultation|Procedure|false|false||auscultationnull|Breath|Finding|false|false||breathnull|null|Device|false|false||soundnull|null|Phenomenon|false|false||soundnull|Left posterior|Modifier|false|false||left posteriornull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Posterior pituitary disease|Disorder|false|false||posteriornull|Dorsal|Modifier|false|false||posteriornull|Basilar|Modifier|false|false||basilarnull|Lung field|Anatomy|false|false|C1553496;C2349184;C2346620;C1521738;C0024115;C0740941|lung fieldnull|Lung diseases|Disorder|false|false|C4037972;C0024109;C0225759|lungnull|Lung Problem|Finding|false|false|C4037972;C0024109;C0225759|lungnull|Chest>Lung|Anatomy|false|false|C0024115;C0740941|lung
null|Lung|Anatomy|false|false|C0024115;C0740941|lungnull|Knowledge Field|Finding|false|false|C0225759|field
null|Force Field|Finding|false|false|C0225759|field
null|Field|Finding|false|false|C0225759|fieldnull|field - patient encounter|Procedure|false|false|C0225759|fieldnull|Wheezing|Finding|true|false||wheezesnull|Basilar Rales|Finding|true|false||rales
null|Rales|Finding|true|false||ralesnull|Regular|Modifier|false|false||Regularnull|Amount type - Rate|Finding|false|false||ratenull|Rating (action)|Event|false|false||ratenull|Rate|LabModifier|false|false||ratenull|Rhythm|Finding|false|false||rhythm
null|rhythmic process (biological)|Finding|false|false||rhythmnull|Heart murmur|Finding|true|false||murmursnull|Pericardial friction rub|Finding|true|false||rubsnull|Malignant neoplasm of abdomen|Disorder|false|false|C0230168;C0000726|Abdomennull|Abdomen problem|Finding|false|false|C0230168;C0000726|Abdomennull|Abdomen|Anatomy|false|false|C0153662;C0941288;C3542022;C0028754|Abdomen
null|Abdominal Cavity|Anatomy|false|false|C0153662;C0941288;C3542022;C0028754|Abdomennull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false|C0230168;C0000726|softnull|Soft|Modifier|false|false||softnull|Obesity|Disorder|false|false|C0230168;C0000726|obesenull|Tender|Modifier|false|false||tendernull|Intestines|Anatomy|false|false||bowelnull|null|Device|false|false||soundsnull|null|Phenomenon|false|false||soundsnull|Present|Finding|false|false||present
null|Presentation|Finding|false|false||presentnull|Rebound tenderness|Finding|true|false||rebound tendernessnull|Emotional tenderness|Finding|true|false||tenderness
null|Sore to touch|Finding|true|false||tendernessnull|Protective muscle spasm|Finding|true|false||guardingnull|Organomegaly|Finding|false|false||organomegalynull|Hereditary Multiple Exostoses|Disorder|false|false||Extnull|EXT1 wt Allele|Finding|false|false||Ext
null|EXT1 gene|Finding|false|false||Extnull|Feels warm|Finding|false|false||warmnull|warming process|Phenomenon|false|false||warmnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false||pulsesnull|Clubbing|Disorder|true|false||clubbingnull|Cyanosis|Finding|true|false||cyanosisnull|Pitting edema|Finding|false|false||pitting edemanull|Pitting|Finding|false|false||pittingnull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Neurology speciality|Title|false|false||Neuronull|Neurologic (qualifier value)|Modifier|false|false||Neuronull|CNS 2|Finding|false|false||CNs2null|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Motor function (finding)|Finding|false|false||motor functionnull|Motor function (observable entity)|Phenomenon|false|false||motor functionnull|motor movement|Finding|false|false||motornull|Motor Device|Device|false|false||motornull|Function (attribute)|Finding|false|false||function
null|physiological aspects|Finding|false|false||function
null|Mathematical Operator|Finding|false|false||function
null|Functional Status|Finding|false|false||functionnull|Function Axis|Subject|false|false||functionnull|Laboratory test finding|Lab|false|false||Labsnull|Admission activity|Procedure|false|false||ADMIT
null|Hospital admission|Procedure|false|false||ADMITnull|Laboratory test finding|Lab|false|false||LABSnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0851353;C0005768;C0229664;C0005767|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C1114281;C0014792|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Lymph|Finding|false|false||Lymphsnull|Monos|Drug|false|false||Monos
null|Mono-S|Drug|false|false||Monos
null|Monos|Drug|false|false||Monosnull|SARCOIDOSIS, EARLY-ONSET|Disorder|false|false||Eos
null|Familial eosinophilia|Disorder|false|false||Eosnull|PRSS33 gene|Finding|false|false||Eos
null|IKZF4 gene|Finding|false|false||Eosnull|Eos <Loriini>|Entity|false|false||Eosnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Alanine Transaminase|Drug|false|false||ALT
null|Alanine Transaminase|Drug|false|false||ALTnull|Liposarcoma, well differentiated|Disorder|false|false|C1185650|ALT
null|Atypical Lipoma|Disorder|false|false|C1185650|ALTnull|null|Finding|false|false|C1185650|ALT
null|Alternative Billing Concepts|Finding|false|false|C1185650|ALT
null|GPT gene|Finding|false|false|C1185650|ALTnull|Antibiotic Lock Therapy|Procedure|false|false|C1185650|ALTnull|Southern Altai Language|Entity|false|false||ALTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false|C1185650|AST
null|Aspartate Transaminase|Drug|false|false|C1185650|AST
null|Aspartate Transaminase|Drug|false|false|C1185650|AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false|C1185650|AST
null|SLC17A5 protein, human|Drug|false|false|C1185650|AST
null|SLC17A5 protein, human|Drug|false|false|C1185650|ASTnull|Atypical Spitz Nevus|Disorder|false|false|C1185650|ASTnull|SLC17A5 wt Allele|Finding|false|false|C1185650|AST
null|SLC17A5 gene|Finding|false|false|C1185650|AST
null|GOT1 gene|Finding|false|false|C1185650|ASTnull|Asterion|Anatomy|false|false|C4553172;C0004002;C0242192;C1121182;C2257651;C1415274;C1140170;C4522245;C1266129;C1370889;C1415181;C1420113;C5960784|ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|Alkaline Phosphatase|Drug|false|false||AlkPhos
null|Alkaline Phosphatase|Drug|false|false||AlkPhosnull|Blood calcium measurement|Procedure|false|false||BLOOD Calciumnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Blood albumin|Procedure|false|false||BLOOD Albuminnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Albumin|Drug|false|false||Albumin
null|Albumins|Drug|false|false||Albumin
null|Albumins|Drug|false|false||Albumin
null|Albumin|Drug|false|false||Albuminnull|Albumin metabolic function|Finding|false|false||Albumin
null|ALB gene|Finding|false|false||Albuminnull|Albumin measurement|Procedure|false|false||Albuminnull|lactate in blood (lab test)|Procedure|false|false||BLOOD Lactatenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|lactate|Drug|false|false||Lactate
null|lactate|Drug|false|false||Lactate
null|Lactates|Drug|false|false||Lactatenull|Lactic acid measurement|Procedure|false|false||Lactatenull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|Laboratory test finding|Lab|false|false||LABSnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0851353;C0005768;C0229664;C0005767|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C0014792;C1114281|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Alanine Transaminase|Drug|false|false||ALT
null|Alanine Transaminase|Drug|false|false||ALTnull|Liposarcoma, well differentiated|Disorder|false|false||ALT
null|Atypical Lipoma|Disorder|false|false||ALTnull|null|Finding|false|false||ALT
null|Alternative Billing Concepts|Finding|false|false||ALT
null|GPT gene|Finding|false|false||ALTnull|Antibiotic Lock Therapy|Procedure|false|false||ALTnull|Southern Altai Language|Entity|false|false||ALTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false|C1185650|AST
null|Aspartate Transaminase|Drug|false|false|C1185650|AST
null|Aspartate Transaminase|Drug|false|false|C1185650|AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false|C1185650|AST
null|SLC17A5 protein, human|Drug|false|false|C1185650|AST
null|SLC17A5 protein, human|Drug|false|false|C1185650|ASTnull|Atypical Spitz Nevus|Disorder|false|false|C1185650|ASTnull|SLC17A5 wt Allele|Finding|false|false|C1185650|AST
null|SLC17A5 gene|Finding|false|false|C1185650|AST
null|GOT1 gene|Finding|false|false|C1185650|ASTnull|Asterion|Anatomy|false|false|C0004002;C0242192;C1121182;C0851148;C1415181;C1420113;C5960784;C0202113;C4522245|ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|Lactate Dehydrogenase|Drug|false|false||LDH
null|Lactate Dehydrogenase|Drug|false|false||LDHnull|Lifetime Drinking History|Finding|false|false|C1185650|LDHnull|Lactate dehydrogenase measurement|Procedure|false|false|C1185650|LDHnull|Alkaline Phosphatase|Drug|false|false||AlkPhos
null|Alkaline Phosphatase|Drug|false|false||AlkPhosnull|Blood calcium measurement|Procedure|false|false||BLOOD Calciumnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Imaging problem|Finding|false|false||IMAGINGnull|Diagnostic Imaging|Procedure|false|false||IMAGING
null|Imaging Techniques|Procedure|false|false||IMAGINGnull|Imaging Technology|Title|false|false||IMAGINGnull|Final report|Finding|false|false||Final Reportnull|Diagnosis Type - Final|Finding|false|false||Finalnull|Final|Time|false|false||Finalnull|End-stage|Modifier|false|false||Finalnull|Report (document)|Finding|false|false||Reportnull|Reporting|Procedure|false|false||Reportnull|null|Attribute|false|false||Reportnull|History of present illness (finding)|Finding|false|false||HISTORY
null|History of previous events|Finding|false|false||HISTORY
null|Historical aspects qualifier|Finding|false|false||HISTORY
null|Medical History|Finding|false|false||HISTORY
null|Concept History|Finding|false|false||HISTORYnull|History|Subject|false|false||HISTORYnull|New diagnosis (finding)|Finding|false|false||New diagnosisnull|New Diagnosis Procedure|Procedure|false|false||New diagnosisnull|Query Status Code - new|Finding|false|false||New
null|Act Status - new|Finding|false|false||Newnull|Newar Language|Entity|false|false||Newnull|New|Modifier|false|false||Newnull|Diagnosis Classification - Diagnosis|Finding|false|false||diagnosis
null|diagnosis aspects|Finding|false|false||diagnosisnull|Diagnosis|Procedure|false|false||diagnosisnull|null|Attribute|false|false||diagnosisnull|Metastatic malignant neoplasm|Disorder|false|false||metastatic cancer
null|Disseminated Malignant Neoplasm|Disorder|false|false||metastatic cancer
null|Neoplasm Metastasis|Disorder|false|false||metastatic cancernull|metastatic qualifier|Finding|false|false||metastatic
null|Metastatic to|Finding|false|false||metastaticnull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|unknown vaccine or immune globulin|Drug|false|false||unknown
null|Unknown - Vaccines administered|Drug|false|false||unknown
null|Unknown - Vaccines administered|Drug|false|false||unknown
null|unknown vaccine or immune globulin|Drug|false|false||unknownnull|Unknown - mode of arrival code|Finding|false|false||unknown
null|Unknown - Special Program Code|Finding|false|false||unknown
null|Unknown - Production Class Code|Finding|false|false||unknown
null|Unknown - Patient Outcome|Finding|false|false||unknown
null|Unknown - Recreational Drug Use Code|Finding|false|false||unknown
null|Unknown - Escort Required|Finding|false|false||unknown
null|Unknown - Transport Arranged|Finding|false|false||unknown
null|Unknown - Living Arrangement|Finding|false|false||unknown
null|Unknown - Employment Status|Finding|false|false||unknown
null|Unknown - Relationship|Finding|false|false||unknown
null|Unknown - publishing section|Finding|false|false||unknown
null|Unknown Publicity Code|Finding|false|false||unknown
null|Unknown - Event reason|Finding|false|false||unknown
null|Unknown - Religion|Finding|false|false||unknown
null|Unknown - Organ Donor Code|Finding|false|false||unknown
null|unknown - NullFlavor|Finding|false|false||unknown
null|Unknown - Notify Clergy Code|Finding|false|false||unknown
null|Unknown - Administrative Gender|Finding|false|false||unknown
null|Unknown - Patient Condition Code|Finding|false|false||unknown
null|Unknown - Living Will Code|Finding|false|false||unknown
null|Marital Status - Unknown|Finding|false|false||unknown
null|Unknown - Patient Class|Finding|false|false||unknown
null|Unknown - Event Expected|Finding|false|false||unknown
null|Unknown - Expanded yes/no indicator|Finding|false|false||unknown
null|Unknown - Immunization Registry Status|Finding|false|false||unknown
null|Unknown - Container status|Finding|false|false||unknown
null|Unknown - CWE statuses|Finding|false|false||unknown
null|Unknown - Patient_s Relationship to Insured|Finding|false|false||unknown
null|Unknown - Job Status|Finding|false|false||unknown
null|Unknown - Precaution Code|Finding|false|false||unknown
null|Unknown - Contact Role|Finding|false|false||unknown
null|Unknown - Living Dependency|Finding|false|false||unknownnull|Ethnic group unknown|Subject|false|false||unknownnull|Unknown - Allergy Severity|Modifier|false|false||unknown
null|Unknown - HL7 update mode|Modifier|false|false||unknown
null|Unknown|Modifier|false|false||unknownnull|True primary (qualifier value)|Time|false|false||primarynull|Primary|Modifier|false|false||primarynull|Extent|Modifier|false|false||extent ofnull|Extent|Modifier|false|false||extentnull|Lesion|Finding|false|false||lesionsnull|Comparison|Event|false|false||COMPARISONnull|null|Attribute|false|false|C1508499;C4266535;C0030797;C0559769;C0000726|CT abdomen and pelvisnull|CT of abdomen|Procedure|false|false|C0000726;C4266535;C0030797;C0559769;C1508499;C0230168;C0000726|CT abdomennull|null|Attribute|false|false|C0230168;C0000726|CT abdomennull|Abdominopelvic structure|Anatomy|false|false|C0153662;C1715387;C0153663;C0941288;C0412620|abdomen and pelvisnull|Abdomen|Anatomy|false|false|C0412620;C0153662;C1715387|abdomen andnull|Malignant neoplasm of abdomen|Disorder|false|false|C1508499;C0000726;C0230168;C0000726|abdomennull|Abdomen problem|Finding|false|false|C1508499;C0230168;C0000726|abdomennull|Abdomen|Anatomy|false|false|C1644645;C0153662;C0412620;C0941288|abdomen
null|Abdominal Cavity|Anatomy|false|false|C1644645;C0153662;C0412620;C0941288|abdomennull|Malignant neoplasm of pelvis|Disorder|false|false|C1508499;C4266535;C0030797;C0559769|pelvisnull|Pelvis problem|Finding|false|false|C4266535;C0030797;C0559769|pelvisnull|Pelvis+|Anatomy|false|false|C1715387;C0412620;C0812455;C0153663|pelvis
null|Pelvic cavity structure|Anatomy|false|false|C1715387;C0412620;C0812455;C0153663|pelvis
null|Pelvis|Anatomy|false|false|C1715387;C0412620;C0812455;C0153663|pelvisnull|Techniques|Finding|false|false||TECHNIQUEnull|Multidetector Computed Tomography|Procedure|false|false|C0460005|Multidetector CTnull|Trunk structure|Anatomy|false|false|C3179130|torsonull|Intravenous Route of Administration|Finding|false|false||intravenousnull|Intravenous|Modifier|false|false||intravenousnull|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C1272919;C1527415;C4521986|oralnull|Oral|Modifier|false|false||oralnull|Contrast Media|Drug|false|false||contrastnull|Contrast|Modifier|false|false||contrastnull|Coronal (qualifier value)|Modifier|false|false||Coronal
null|Coronal plane|Modifier|false|false||Coronalnull|Sagittal plane|Anatomy|false|false||sagittalnull|Sagittal|Modifier|false|false||sagittalnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Assessment of body build|Procedure|false|false|C0460148;C0444584;C4082212;C1268086;C0152338|body habitusnull|Document Body|Finding|false|false|C0460148;C0444584;C4082212;C1268086;C0152338|bodynull|Structure of body of caudate nucleus|Anatomy|false|false|C1318474;C1551342|body
null|Human body structure|Anatomy|false|false|C1318474;C1551342|body
null|Body structure|Anatomy|false|false|C1318474;C1551342|body
null|Adult human body|Anatomy|false|false|C1318474;C1551342|body
null|Whole body|Anatomy|false|false|C1318474;C1551342|bodynull|Human body|Subject|false|false||bodynull|findings aspects|Finding|false|false||FINDINGSnull|null|Attribute|false|false||FINDINGSnull|Chest problem|Finding|false|false|C1527391;C0817096|CHESTnull|Chest|Anatomy|false|false|C0741025|CHEST
null|Anterior thoracic region|Anatomy|false|false|C0741025|CHESTnull|Multiple Pulmonary Nodules|Finding|false|false|C0024109|pulmonary nodulesnull|Pulmonary (intended site)|Finding|false|false|C0024109|pulmonarynull|Lung|Anatomy|false|false|C4522268;C2707265;C0748164|pulmonarynull|null|Attribute|false|false|C0024109|pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|AKT1S1 wt Allele|Finding|false|false|C0796494|lobe
null|AKT1S1 gene|Finding|false|false|C0796494|lobenull|lobe|Anatomy|false|false|C3539671;C1428707|lobenull|Structure of left upper lobe of lung|Anatomy|false|false|C1552822;C3539671;C1428707|left upper lobenull|Table Cell Horizontal Align - left|Finding|false|false|C1261076;C0225756;C0796494|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Structure of upper lobe of lung|Anatomy|false|false|C1552822;C3539671;C1428707|upper lobenull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|AKT1S1 wt Allele|Finding|false|false|C0796494;C0225756;C1261076|lobe
null|AKT1S1 gene|Finding|false|false|C0796494;C0225756;C1261076|lobenull|lobe|Anatomy|false|false|C3539671;C1428707;C1552822|lobenull|Largest|LabModifier|false|false||largestnull|Diameter (qualifier value)|LabModifier|false|false||diameternull|Sequence - TransmissionRelationshipTypeCode|Finding|false|false||sequence
null|DNA Sequence|Finding|false|false||sequence
null|RNA Sequence|Finding|false|false||sequence
null|Sequence|Finding|false|false||sequence
null|Base Sequence|Finding|false|false||sequence
null|Sequence - ParameterizedDataType|Finding|false|false||sequencenull|Intrauterine growth restriction, metaphyseal dysplasia, adrenal hypoplasia congenita, and genital anomaly syndrome|Disorder|false|false||imagenull|Image (foundation metadata concept)|Finding|false|false||image
null|Image|Finding|false|false||image
null|Medical Image|Finding|false|false||image
null|image - dosage form|Finding|false|false||imagenull|Integrated Molecular Analysis of Genomes and their Expression Consortium|Entity|false|false||imagenull|Physiologic calcification|Finding|false|false||Calcification
null|Calcification|Finding|false|false||Calcification
null|Calcinosis|Finding|false|false||Calcificationnull|Calcified (qualifier value)|Modifier|false|false||Calcificationnull|Structure of right pleural cavity|Anatomy|false|false|C1510420;C0011334;C0162326;C0004793;C1519249;C1547787;C3853789;C0162327;C3542466;C1704254;C1704922;C1696103;C1846009;C0032226;C1552823|right pleural cavitynull|Table Cell Horizontal Align - right|Finding|false|false|C0178802;C0225782|rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Pleural cavity|Anatomy|false|false|C0162326;C0004793;C1519249;C1547787;C3853789;C0162327;C1552823;C1510420;C0011334;C0032226;C3542466;C1704254;C1704922;C1696103;C1846009|pleural cavitynull|Pleural Diseases|Disorder|false|false|C0333343;C0178802;C0225782;C0032225|pleuralnull|Pleura|Anatomy|false|false|C0162326;C0004793;C1519249;C1547787;C3853789;C0162327;C1510420;C0011334;C0032226|pleuralnull|Pleural|Modifier|false|false||pleuralnull|Dental caries|Disorder|false|false|C0225782;C0178802;C0032225;C0333343|cavity
null|Cavitation|Disorder|false|false|C0225782;C0178802;C0032225;C0333343|cavitynull|Body cavities|Anatomy|false|false|C0032226;C3542466;C1704254;C1704922;C1696103;C0162326;C0004793;C1519249;C1547787;C3853789;C0162327;C1510420;C0011334;C1846009|cavitynull|Sequence - TransmissionRelationshipTypeCode|Finding|false|false|C0178802;C0225782;C0032225;C0333343|sequence
null|DNA Sequence|Finding|false|false|C0178802;C0225782;C0032225;C0333343|sequence
null|RNA Sequence|Finding|false|false|C0178802;C0225782;C0032225;C0333343|sequence
null|Sequence|Finding|false|false|C0178802;C0225782;C0032225;C0333343|sequence
null|Base Sequence|Finding|false|false|C0178802;C0225782;C0032225;C0333343|sequence
null|Sequence - ParameterizedDataType|Finding|false|false|C0178802;C0225782;C0032225;C0333343|sequencenull|Intrauterine growth restriction, metaphyseal dysplasia, adrenal hypoplasia congenita, and genital anomaly syndrome|Disorder|false|false|C0225782;C0333343;C0178802|imagenull|Image (foundation metadata concept)|Finding|false|false|C0225782;C0333343;C0178802|image
null|Image|Finding|false|false|C0225782;C0333343;C0178802|image
null|Medical Image|Finding|false|false|C0225782;C0333343;C0178802|image
null|image - dosage form|Finding|false|false|C0225782;C0333343;C0178802|imagenull|Integrated Molecular Analysis of Genomes and their Expression Consortium|Entity|false|false||imagenull|Adverse Event Probably Related to Intervention|Modifier|false|false||likely relatednull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Relate - vinyl resin|Drug|false|false||relatednull|Role Link Type - related|Finding|false|false||related
null|Related (finding)|Finding|false|false||relatednull|Definitely Related to Intervention|Modifier|false|false||related
null|Relationships|Modifier|false|false||relatednull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Medical History|Finding|false|false||history ofnull|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|History of present illness (finding)|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Act Relationship Subset - previous|Time|false|false||previous
null|Previous|Time|false|false||previousnull|Right lung|Anatomy|false|false|C0024115;C0740941;C0543467;C0038895;C1457907;C1547138;C1552823;C0038903|right lungnull|Table Cell Horizontal Align - right|Finding|false|false|C0225706|rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Pulmonary Surgical Procedures|Procedure|false|false|C4037972;C0024109;C0225706|lung surgerynull|Lung diseases|Disorder|false|false|C0225706;C4037972;C0024109|lungnull|Lung Problem|Finding|false|false|C0225706;C4037972;C0024109|lungnull|Chest>Lung|Anatomy|false|false|C0543467;C0740941;C0024115;C0038903;C0038895;C1457907;C1547138|lung
null|Lung|Anatomy|false|false|C0543467;C0740941;C0024115;C0038903;C0038895;C1457907;C1547138|lungnull|Level of Care - Surgery|Finding|false|false|C0225706;C4037972;C0024109|surgery
null|Surgical procedure finding|Finding|false|false|C0225706;C4037972;C0024109|surgery
null|Surgical aspects|Finding|false|false|C0225706;C4037972;C0024109|surgerynull|Operative Surgical Procedures|Procedure|false|false|C4037972;C0024109;C0225706|surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Pleural effusion (disorder)|Finding|true|false|C0032225|pleural effusion
null|Pleural effusion fluid|Finding|true|false|C0032225|pleural effusion
null|null|Finding|true|false|C0032225|pleural effusionnull|Pleural Diseases|Disorder|false|false|C0032225|pleuralnull|Pleura|Anatomy|false|false|C2073625;C1253943;C0032227;C0032226;C2317432;C1546613;C0013687|pleuralnull|Pleural|Modifier|false|false||pleuralnull|Effusion (substance)|Finding|true|false|C0032225|effusion
null|null|Finding|true|false|C0032225|effusion
null|effusion|Finding|true|false|C0032225|effusionnull|Pneumothorax|Disorder|true|false||pneumothoraxnull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|Mediastinum|Anatomy|false|false||mediastinalnull|Mediastinal|Modifier|false|false||mediastinalnull|Axilla|Anatomy|false|false|C4282165;C0497156|axillarynull|Hilar lymphadenopathy|Disorder|true|false||hilar adenopathynull|Hilar|Modifier|false|false||hilarnull|Lymphadenopathy|Disorder|false|false|C0004454|adenopathynull|Swollen Lymph Node|Finding|false|false|C0004454|adenopathynull|Cardiac attachment|Finding|false|false|C0018787|Cardiacnull|Heart|Anatomy|false|false|C1314974|Cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||Cardiacnull|size|Modifier|false|false||sizenull|size - solid dosage form|LabModifier|false|false||sizenull|Pericardial effusion|Disorder|true|false|C0031050;C0442031|pericardial effusionnull|Pericardial effusion body substance|Finding|true|false|C0031050;C0442031|pericardial effusionnull|Pericardial (qualifier value)|Anatomy|false|false|C0031039;C2317432;C1546613;C0013687;C1253937|pericardial
null|Pericardial sac structure|Anatomy|false|false|C0031039;C2317432;C1546613;C0013687;C1253937|pericardialnull|Effusion (substance)|Finding|true|false|C0031050;C0442031|effusion
null|null|Finding|true|false|C0031050;C0442031|effusion
null|effusion|Finding|true|false|C0031050;C0442031|effusionnull|Malignant neoplasm of abdomen|Disorder|false|false|C0230168;C0000726|ABDOMENnull|Abdomen problem|Finding|false|false|C0230168;C0000726|ABDOMENnull|Abdomen|Anatomy|false|false|C0941288;C0153662|ABDOMEN
null|Abdominal Cavity|Anatomy|false|false|C0941288;C0153662|ABDOMENnull|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|liver
null|liver extract|Drug|false|false|C4037986;C1278929;C0023884|liver
null|liver extract|Drug|false|false|C4037986;C1278929;C0023884|liver
null|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|liver
null|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|livernull|Benign neoplasm of liver|Disorder|false|false|C4037986;C1278929;C0023884|liver
null|Liver diseases|Disorder|false|false|C4037986;C1278929;C0023884|livernull|Liver problem|Finding|false|false|C4037986;C1278929;C0023884|livernull|Procedures on liver|Procedure|false|false|C4037986;C1278929;C0023884|livernull|Abdomen>Liver|Anatomy|false|false|C0721399;C0023899;C0023895;C0496870;C0577060;C1293134;C0872387|liver
null|null|Anatomy|false|false|C0721399;C0023899;C0023895;C0496870;C0577060;C1293134;C0872387|liver
null|Liver|Anatomy|false|false|C0721399;C0023899;C0023895;C0496870;C0577060;C1293134;C0872387|livernull|Enlargement procedure|Procedure|false|false|C4037986;C1278929;C0023884|enlargednull|Enlarged|Modifier|false|false||enlargednull|density|LabModifier|false|false||densitynull|Lesion|Finding|false|false|C0796494;C4037986;C1278929;C0023884|lesionsnull|lobe|Anatomy|false|false|C0872387;C0721399;C0023899;C0023895;C0496870;C0221198;C0577060|lobesnull|Liver brand of Vitamin B 12|Drug|true|false|C0796494;C4037986;C1278929;C0023884|liver
null|liver extract|Drug|true|false|C0796494;C4037986;C1278929;C0023884|liver
null|liver extract|Drug|true|false|C0796494;C4037986;C1278929;C0023884|liver
null|Liver brand of Vitamin B 12|Drug|true|false|C0796494;C4037986;C1278929;C0023884|liver
null|Liver brand of Vitamin B 12|Drug|true|false|C0796494;C4037986;C1278929;C0023884|livernull|Benign neoplasm of liver|Disorder|true|false|C4037986;C1278929;C0023884;C0796494|liver
null|Liver diseases|Disorder|true|false|C4037986;C1278929;C0023884;C0796494|livernull|Liver problem|Finding|true|false|C4037986;C1278929;C0023884;C0796494|livernull|Procedures on liver|Procedure|true|false|C0796494;C4037986;C1278929;C0023884|livernull|Abdomen>Liver|Anatomy|false|false|C0577060;C0023895;C0496870;C0721399;C0023899;C0872387;C0221198|liver
null|null|Anatomy|false|false|C0577060;C0023895;C0496870;C0721399;C0023899;C0872387;C0221198|liver
null|Liver|Anatomy|false|false|C0577060;C0023895;C0496870;C0721399;C0023899;C0872387;C0221198|livernull|veterans alcoholism screening test (VAST)|Finding|false|false|C0933845;C0736268|vastnull|majority|Finding|false|false|C0205054;C0933845;C0736268|majoritynull|Liver parenchyma|Anatomy|false|false|C0814230;C0680220|hepatic parenchymanull|Hepatic|Anatomy|false|false|C0680220|hepaticnull|Parenchyma|Anatomy|false|false|C0814230;C0680220|parenchymanull|Portal vein structure|Anatomy|false|false||portal vein
null|Abdomen>Portal vein|Anatomy|false|false||portal vein
null|null|Anatomy|false|false||portal veinnull|Hepatic|Anatomy|false|false||portalnull|Veins|Anatomy|false|false||veinnull|Legal patent|Finding|false|false||patentnull|Open|Modifier|false|false||patentnull|During values|Time|false|false||intranull|Extrahepatic|Modifier|false|false||extrahepaticnull|Duct (organ) structure|Anatomy|false|false|C1322279|duct
null|canal [body parts]|Anatomy|false|false|C1322279|ductnull|Duct Device|Device|false|false||ductnull|Pathological Dilatation|Finding|true|false||dilatation
null|Dilated|Finding|true|false||dilatationnull|Dilate procedure|Procedure|true|false|C0687028;C1550227|dilatationnull|examination of gallbladder|Procedure|false|false|C4071903;C1524055;C0016976|gallbladdernull|Gallbladder (MMHCC)|Anatomy|false|false|C2032932|gallbladder
null|Gallbladder|Anatomy|false|false|C2032932|gallbladder
null|Abdomen>Gallbladder|Anatomy|false|false|C2032932|gallbladdernull|null|Modifier|false|false||unremarkablenull|Small amount|LabModifier|false|false||small amountnull|Small|LabModifier|false|false||smallnull|Amount class - Amount|Finding|false|false||amountnull|Quantity|LabModifier|false|false||amountnull|Ascites|Disorder|false|false||ascitesnull|Peritoneal Effusion|Finding|false|false||ascitesnull|Adjacent|Modifier|false|false||adjacent tonull|Adjacent|Modifier|false|false||adjacentnull|To the right (qualifier value)|Modifier|false|false||to the rightnull|Right lobe of liver|Anatomy|false|false|C0872387;C0023895;C0496870;C0721399;C0023899;C0577060;C3539671;C1428707;C1552823|right lobe of the livernull|Table Cell Horizontal Align - right|Finding|false|false|C0796494;C4037986;C1278929;C0023884;C0227481|rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|AKT1S1 wt Allele|Finding|false|false|C0227481;C4037986;C1278929;C0023884;C0796494|lobe
null|AKT1S1 gene|Finding|false|false|C0227481;C4037986;C1278929;C0023884;C0796494|lobenull|lobe|Anatomy|false|false|C0577060;C1552823;C0023895;C0496870;C3539671;C1428707;C0721399;C0023899;C0872387|lobenull|Liver brand of Vitamin B 12|Drug|false|false|C0227481;C4037986;C1278929;C0023884;C0796494|liver
null|liver extract|Drug|false|false|C0227481;C4037986;C1278929;C0023884;C0796494|liver
null|liver extract|Drug|false|false|C0227481;C4037986;C1278929;C0023884;C0796494|liver
null|Liver brand of Vitamin B 12|Drug|false|false|C0227481;C4037986;C1278929;C0023884;C0796494|liver
null|Liver brand of Vitamin B 12|Drug|false|false|C0227481;C4037986;C1278929;C0023884;C0796494|livernull|Benign neoplasm of liver|Disorder|false|false|C0796494;C0227481;C4037986;C1278929;C0023884|liver
null|Liver diseases|Disorder|false|false|C0796494;C0227481;C4037986;C1278929;C0023884|livernull|Liver problem|Finding|false|false|C0796494;C4037986;C1278929;C0023884;C0227481|livernull|Procedures on liver|Procedure|false|false|C0227481;C0796494;C4037986;C1278929;C0023884|livernull|Abdomen>Liver|Anatomy|false|false|C1552823;C0577060;C0023895;C0496870;C3539671;C1428707;C0721399;C0023899;C0872387|liver
null|null|Anatomy|false|false|C1552823;C0577060;C0023895;C0496870;C3539671;C1428707;C0721399;C0023899;C0872387|liver
null|Liver|Anatomy|false|false|C1552823;C0577060;C0023895;C0496870;C3539671;C1428707;C0721399;C0023899;C0872387|livernull|Right kidney|Anatomy|false|false|C0812426;C0496927;C0496892;C4554465;C0869841;C1552823|right kidneynull|Table Cell Horizontal Align - right|Finding|false|false|C0227665;C0022646;C0227613|rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Neoplasm of uncertain or unknown behavior of kidney|Disorder|false|false|C0227665;C0022646;C0227613|kidney
null|Benign neoplasm of kidney|Disorder|false|false|C0227665;C0022646;C0227613|kidneynull|Kidney problem|Finding|false|false|C0227613;C0227665;C0022646|kidneynull|examination of kidney|Procedure|false|false|C0227613;C0227665;C0022646|kidney
null|Procedures on Kidney|Procedure|false|false|C0227613;C0227665;C0022646|kidneynull|Kidney|Anatomy|false|false|C0496927;C0496892;C0812426;C1552823;C4554465;C0869841|kidney
null|Both kidneys|Anatomy|false|false|C0496927;C0496892;C0812426;C1552823;C4554465;C0869841|kidneynull|MILDLY|Modifier|false|false||mildly
null|Mild (qualifier value)|Modifier|false|false||mildlynull|Hepatomegaly|Finding|false|false|C4037986;C1278929;C0023884|enlarged livernull|Enlargement procedure|Procedure|false|false|C4037986;C1278929;C0023884|enlargednull|Enlarged|Modifier|false|false||enlargednull|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|liver
null|liver extract|Drug|false|false|C4037986;C1278929;C0023884|liver
null|liver extract|Drug|false|false|C4037986;C1278929;C0023884|liver
null|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|liver
null|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|livernull|Benign neoplasm of liver|Disorder|false|false|C4037986;C1278929;C0023884|liver
null|Liver diseases|Disorder|false|false|C4037986;C1278929;C0023884|livernull|Liver problem|Finding|false|false|C4037986;C1278929;C0023884|livernull|Procedures on liver|Procedure|false|false|C4037986;C1278929;C0023884|livernull|Abdomen>Liver|Anatomy|false|false|C0019209;C0721399;C0023899;C0023895;C0496870;C0577060;C1293134;C0872387|liver
null|null|Anatomy|false|false|C0019209;C0721399;C0023899;C0023895;C0496870;C0577060;C1293134;C0872387|liver
null|Liver|Anatomy|false|false|C0019209;C0721399;C0023899;C0023895;C0496870;C0577060;C1293134;C0872387|livernull|density|LabModifier|false|false||densitynull|Lesion|Finding|false|false||lesion
null|null|Finding|false|false||lesionnull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|DNA Polymerase Epsilon Catalytic Subunit A, Human|Drug|false|false|C0935623;C0227613;C0227665;C0022646|pole
null|DNA Polymerase Epsilon Catalytic Subunit A, Human|Drug|false|false|C0935623;C0227613;C0227665;C0022646|polenull|POLE gene|Finding|false|false|C0227613;C0227665;C0022646;C0935623|polenull|anatomical pole|Anatomy|false|false|C0496927;C0496892;C1552823;C0812426;C4554465;C0869841;C3811771;C1418729|polenull|Right kidney|Anatomy|false|false|C1418729;C4554465;C0869841;C0332148;C0750492;C0496927;C0496892;C3811771;C0812426;C1552823|right kidneynull|Table Cell Horizontal Align - right|Finding|false|false|C0935623;C0227665;C0022646;C0227613|rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Neoplasm of uncertain or unknown behavior of kidney|Disorder|false|false|C0935623;C0227665;C0022646;C0227613|kidney
null|Benign neoplasm of kidney|Disorder|false|false|C0935623;C0227665;C0022646;C0227613|kidneynull|Kidney problem|Finding|false|false|C0935623;C0227665;C0022646;C0227613|kidneynull|examination of kidney|Procedure|false|false|C0227665;C0022646;C0227613;C0935623|kidney
null|Procedures on Kidney|Procedure|false|false|C0227665;C0022646;C0227613;C0935623|kidneynull|Kidney|Anatomy|false|false|C0496927;C0496892;C4554465;C0869841;C1552823;C1418729;C0812426;C3811771|kidney
null|Both kidneys|Anatomy|false|false|C0496927;C0496892;C4554465;C0869841;C1552823;C1418729;C0812426;C3811771|kidneynull|Probable diagnosis|Finding|false|false|C0227613|likely
null|Probably|Finding|false|false|C0227613|likelynull|Cyst|Disorder|false|false||cystnull|SpecimenType - Cyst|Finding|false|false||cyst
null|null|Finding|false|false||cystnull|Cyst form of protozoa|Entity|false|false||cystnull|Sequence - TransmissionRelationshipTypeCode|Finding|false|false||sequence
null|DNA Sequence|Finding|false|false||sequence
null|RNA Sequence|Finding|false|false||sequence
null|Sequence|Finding|false|false||sequence
null|Base Sequence|Finding|false|false||sequence
null|Sequence - ParameterizedDataType|Finding|false|false||sequencenull|Intrauterine growth restriction, metaphyseal dysplasia, adrenal hypoplasia congenita, and genital anomaly syndrome|Disorder|false|false||imagenull|Image (foundation metadata concept)|Finding|false|false||image
null|Image|Finding|false|false||image
null|Medical Image|Finding|false|false||image
null|image - dosage form|Finding|false|false||imagenull|Integrated Molecular Analysis of Genomes and their Expression Consortium|Entity|false|false||imagenull|Right kidney|Anatomy|false|false|C0812426;C4554465;C0869841;C0496927;C0496892;C1552823|right kidneynull|Table Cell Horizontal Align - right|Finding|false|false|C0227665;C0022646;C0227613|rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Neoplasm of uncertain or unknown behavior of kidney|Disorder|false|false|C0227665;C0022646;C0227613|kidney
null|Benign neoplasm of kidney|Disorder|false|false|C0227665;C0022646;C0227613|kidneynull|Kidney problem|Finding|false|false|C0227613;C0227665;C0022646|kidneynull|examination of kidney|Procedure|false|false|C0227613;C0227665;C0022646|kidney
null|Procedures on Kidney|Procedure|false|false|C0227613;C0227665;C0022646|kidneynull|Kidney|Anatomy|false|false|C0812426;C0496927;C0496892;C1552823;C4554465;C0869841|kidney
null|Both kidneys|Anatomy|false|false|C0812426;C0496927;C0496892;C1552823;C4554465;C0869841|kidneynull|null|Modifier|false|false||unremarkablenull|Left kidney|Anatomy|false|false|C4554465;C0869841;C1552822;C0496927;C0496892;C0812426|left kidneynull|Table Cell Horizontal Align - left|Finding|false|false|C0227614;C0227665;C0022646|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Neoplasm of uncertain or unknown behavior of kidney|Disorder|false|false|C0227665;C0022646;C0227614|kidney
null|Benign neoplasm of kidney|Disorder|false|false|C0227665;C0022646;C0227614|kidneynull|Kidney problem|Finding|false|false|C0227614;C0227665;C0022646|kidneynull|examination of kidney|Procedure|false|false|C0227614;C0227665;C0022646|kidney
null|Procedures on Kidney|Procedure|false|false|C0227614;C0227665;C0022646|kidneynull|Kidney|Anatomy|false|false|C0496927;C0496892;C4554465;C0869841;C0812426;C1552822|kidney
null|Both kidneys|Anatomy|false|false|C0496927;C0496892;C4554465;C0869841;C0812426;C1552822|kidneynull|Limited (extensiveness)|Finding|false|false||limitsnull|Adrenal Glands|Anatomy|false|false|C0812414;C0153470;C0869677|adrenalsnull|Malignant neoplasm of spleen|Disorder|false|false|C4037984;C0037993;C0001625|spleennull|Spleen problem|Finding|false|false|C4037984;C0037993;C0001625|spleennull|Procedures on Spleen|Procedure|false|false|C0001625;C4037984;C0037993|spleennull|Abdomen>Spleen|Anatomy|false|false|C0812414;C0153470;C0869677|spleen
null|Spleen|Anatomy|false|false|C0812414;C0153470;C0869677|spleennull|null|Modifier|false|false||unremarkablenull|pancreas extract|Drug|false|false|C4037927;C0030274|pancreas
null|pancreas extract|Drug|false|false|C4037927;C0030274|pancreasnull|Benign tumor of pancreas|Disorder|false|false|C4037927;C0030274|pancreas
null|Pancreatic Diseases|Disorder|false|false|C4037927;C0030274|pancreasnull|Pancreas problem|Finding|false|false|C4037927;C0030274|pancreasnull|Procedures on Pancreas|Procedure|false|false|C4037927;C0030274|pancreasnull|Abdomen>Pancreas|Anatomy|false|false|C0869826;C0347284;C0030286;C0813176;C0771711|pancreas
null|Pancreas|Anatomy|false|false|C0869826;C0347284;C0030286;C0813176;C0771711|pancreasnull|null|Finding|false|false||within normal limitsnull|Limited (extensiveness)|Finding|false|false||limitsnull|Small|LabModifier|false|false||smallnull|Large Intestine|Anatomy|false|false|C5890938;C1416798|large bowelnull|LARGE1 wt Allele|Finding|false|false|C0021851|large
null|LARGE1 gene|Finding|false|false|C0021851|largenull|Large|LabModifier|false|false||largenull|Intestines|Anatomy|false|false||bowelnull|null|Modifier|false|false||unremarkablenull|Retroperitoneal Space|Anatomy|false|false|C0497156|retroperitonealnull|Mesentery|Anatomy|false|false|C4282165;C0497156|mesentericnull|Lymphadenopathy|Disorder|true|false|C0035359;C0025474|adenopathynull|Swollen Lymph Node|Finding|true|false|C0025474|adenopathynull|Malignant neoplasm of pelvis|Disorder|false|false|C4266535;C0030797;C0559769|PELVISnull|Pelvis problem|Finding|false|false|C4266535;C0030797;C0559769|PELVISnull|Pelvis+|Anatomy|false|false|C0153663;C0812455|PELVIS
null|Pelvic cavity structure|Anatomy|false|false|C0153663;C0812455|PELVIS
null|Pelvis|Anatomy|false|false|C0153663;C0812455|PELVISnull|Malignant neoplasm of pelvis|Disorder|false|false|C4266535;C0030797;C0559769|pelvisnull|Pelvis problem|Finding|false|false|C4266535;C0030797;C0559769|pelvisnull|Pelvis+|Anatomy|false|false|C0812455;C0153663|pelvis
null|Pelvic cavity structure|Anatomy|false|false|C0812455;C0153663|pelvis
null|Pelvis|Anatomy|false|false|C0812455;C0153663|pelvisnull|Secondary to|Modifier|false|false||secondary tonull|Neoplasm Metastasis|Disorder|false|false||secondarynull|metastatic qualifier|Finding|false|false||secondarynull|Secondary to|Modifier|false|false||secondarynull|second (number)|LabModifier|false|false||secondarynull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Assessment of body build|Procedure|false|false|C0460148;C0444584;C4082212;C1268086;C0152338|body habitusnull|Document Body|Finding|false|false|C0460148;C0444584;C4082212;C1268086;C0152338|bodynull|Structure of body of caudate nucleus|Anatomy|false|false|C1551342;C1318474|body
null|Human body structure|Anatomy|false|false|C1551342;C1318474|body
null|Body structure|Anatomy|false|false|C1551342;C1318474|body
null|Adult human body|Anatomy|false|false|C1551342;C1318474|body
null|Whole body|Anatomy|false|false|C1551342;C1318474|bodynull|Human body|Subject|false|false||bodynull|Pelvis|Anatomy|false|false||pelvicnull|Neoplasm of uncertain or unknown behavior of bladder|Disorder|false|false|C0005682|bladder
null|Benign neoplasm of bladder|Disorder|false|false|C0005682|bladder
null|Carcinoma in situ of bladder|Disorder|false|false|C0005682|bladdernull|Procedures on bladder|Procedure|false|false|C0005682|bladdernull|Urinary Bladder|Anatomy|false|false|C0496930;C0154017;C0154091;C0872388|bladdernull|null|Modifier|false|false||unremarkablenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Status post|Time|false|false||status post
null|Post|Time|false|false||status postnull|What subject filter - Status|Finding|false|false||statusnull|null|Attribute|false|false||statusnull|Social status|Modifier|false|false||status
null|Status|Modifier|false|false||statusnull|SLC35G1 gene|Finding|false|false||post
null|DESI1 gene|Finding|false|false||postnull|Post Device|Device|false|false||postnull|Post|Time|false|false||postnull|Supracervical hysterectomy|Procedure|false|false||supracervical hysterectomy
null|Partial hysterectomy|Procedure|false|false||supracervical hysterectomynull|Consent Type - Hysterectomy|Finding|false|false||hysterectomynull|Hysterectomy|Procedure|false|false||hysterectomynull|Pelvis|Anatomy|false|false|C0497156;C4282165|pelvicnull|Lymphadenopathy|Disorder|true|false|C0030797|adenopathynull|Swollen Lymph Node|Finding|true|false|C0030797|adenopathynull|effusion|Finding|true|false||free fluidnull|Free of (attribute)|Finding|true|false||freenull|Empty (qualifier)|Modifier|false|false||freenull|fluid - substance|Drug|true|false||fluid
null|Liquid substance|Drug|true|false||fluidnull|Fluid Specimen Code|Finding|true|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Malignant neoplasm of pelvis|Disorder|false|false|C4266535;C0030797;C0559769|pelvisnull|Pelvis problem|Finding|false|false|C4266535;C0030797;C0559769|pelvisnull|Pelvis+|Anatomy|false|false|C0812455;C0153663|pelvis
null|Pelvic cavity structure|Anatomy|false|false|C0812455;C0153663|pelvis
null|Pelvis|Anatomy|false|false|C0812455;C0153663|pelvisnull|Bone Tissue, Human|Anatomy|false|false||OSSEOUS
null|Skeletal bone|Anatomy|false|false||OSSEOUSnull|Structure|Modifier|false|false||STRUCTURESnull|Bilateral|Modifier|false|false||Bilateralnull|Symmetrical|Finding|false|false||symmetricalnull|Sclerosis|Finding|false|false|C0020889|sclerosisnull|Bone structure of ilium|Anatomy|false|false|C0036429|iliacnull|Side|Modifier|false|false||sidenull|Sacroiliac joint structure|Anatomy|false|false|C0343261;C0029400;C0332290;C0152263;C0332290|sacroiliac jointsnull|sacroiliac|Anatomy|false|false|C0029400;C0343261;C0332290;C0152263|sacroiliacnull|Joints|Anatomy|false|false|C0332290;C0152263;C0343261;C0029400|joints
null|Articular system|Anatomy|false|false|C0332290;C0152263;C0343261;C0029400|jointsnull|Consistent with|Finding|false|false|C0036036|consistent withnull|Compatible|Modifier|false|false||consistent withnull|Consistent with|Finding|false|false|C0392905;C0022417;C0036036;C0555898|consistentnull|Osteitis condensans ilii|Disorder|false|false|C0036036;C0555898;C0392905;C0022417|osteitis condensans iliinull|Osteitis condensans|Disorder|false|false|C0392905;C0022417;C0036036;C0555898|osteitis condensansnull|Osteitis|Disorder|false|false|C0555898;C0036036;C0392905;C0022417|osteitisnull|Severe - Severity of Illness Code|Finding|false|false|C1285116;C0524470;C0019558;C0392905;C1269611;C0022417;C0022122;C0228391;C0019552;C4299095|severe
null|Intensity and Distress 5|Finding|false|false|C1285116;C0524470;C0019558;C0392905;C1269611;C0022417;C0022122;C0228391;C0019552;C4299095|severe
null|Severe - Triage Code|Finding|false|false|C1285116;C0524470;C0019558;C0392905;C1269611;C0022417;C0022122;C0228391;C0019552;C4299095|severe
null|Severe (severity modifier)|Finding|false|false|C1285116;C0524470;C0019558;C0392905;C1269611;C0022417;C0022122;C0228391;C0019552;C4299095|severe
null|Allergy Severity - Severe|Finding|false|false|C1285116;C0524470;C0019558;C0392905;C1269611;C0022417;C0022122;C0228391;C0019552;C4299095|severenull|Abnormal degeneration|Finding|false|false|C0019558;C0524470;C1285116|degenerative changenull|biologic degeneration|Finding|false|false|C0022122;C0228391;C0019552;C4299095;C0392905;C1269611;C0022417;C1285116;C0524470;C0019558|degenerative
null|Abnormal degeneration|Finding|false|false|C0022122;C0228391;C0019552;C4299095;C0392905;C1269611;C0022417;C1285116;C0524470;C0019558|degenerativenull|Changing|Finding|false|false|C0022122;C0228391;C0019552;C4299095;C0019558;C1285116;C0524470;C0392905;C1269611;C0022417|changenull|Change - procedure|Procedure|false|false|C0022122;C0228391;C0019552;C4299095;C0019558;C1285116;C0392905;C1269611;C0022417;C0524470|changenull|Delta (difference)|LabModifier|false|false||change
null|Changed status|LabModifier|false|false||changenull|Right hip joint structure|Anatomy|false|false|C5203119;C1547231;C0205082;C1547227;C1561581;C0392747;C1430701;C0529134;C1505163;C1654726;C0011164;C1880269;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C1292890;C0575044;C0011164;C4319952;C1552823|right hip jointnull|Right hip region structure|Anatomy|false|false|C0575044;C5203119;C1547231;C0205082;C1547227;C1561581;C1292890;C0392747;C1552823;C0011164;C1430701;C0529134;C1505163;C1654726;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C0011164;C1880269;C4319952|right hipnull|Table Cell Horizontal Align - right|Finding|false|false|C0392905;C1269611;C0022417;C0524470;C0019558;C0022122;C0228391;C0019552;C4299095;C1285116|rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Hip Joint|Anatomy|false|false|C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C0392747;C1292890;C0011164;C5203119;C1547231;C0205082;C1547227;C1561581;C0575044;C4319952;C1552823;C1430701;C0529134;C1505163;C1654726;C0011164;C1880269|hip jointnull|heme iron polypeptide|Drug|false|false|C0022122;C0228391;C0019552;C4299095;C0392905;C1269611;C0022417;C1285116;C0524470;C0019558|hip
null|ST13 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095;C0392905;C1269611;C0022417;C1285116;C0524470;C0019558|hip
null|ST13 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095;C0392905;C1269611;C0022417;C1285116;C0524470;C0019558|hip
null|RPL29 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095;C0392905;C1269611;C0022417;C1285116;C0524470;C0019558|hip
null|RPL29 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095;C0392905;C1269611;C0022417;C1285116;C0524470;C0019558|hip
null|HHIP protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095;C0392905;C1269611;C0022417;C1285116;C0524470;C0019558|hip
null|HHIP protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095;C0392905;C1269611;C0022417;C1285116;C0524470;C0019558|hip
null|heme iron polypeptide|Drug|false|false|C0022122;C0228391;C0019552;C4299095;C0392905;C1269611;C0022417;C1285116;C0524470;C0019558|hipnull|RPL29 wt Allele|Finding|false|false|C0019558;C0392905;C1269611;C0022417;C0022122;C0228391;C0019552;C4299095;C0524470;C1285116|hip
null|REG3A gene|Finding|false|false|C0019558;C0392905;C1269611;C0022417;C0022122;C0228391;C0019552;C4299095;C0524470;C1285116|hip
null|RPL29 gene|Finding|false|false|C0019558;C0392905;C1269611;C0022417;C0022122;C0228391;C0019552;C4299095;C0524470;C1285116|hip
null|ST13 wt Allele|Finding|false|false|C0019558;C0392905;C1269611;C0022417;C0022122;C0228391;C0019552;C4299095;C0524470;C1285116|hip
null|ST13 gene|Finding|false|false|C0019558;C0392905;C1269611;C0022417;C0022122;C0228391;C0019552;C4299095;C0524470;C1285116|hip
null|HHIP gene|Finding|false|false|C0019558;C0392905;C1269611;C0022417;C0022122;C0228391;C0019552;C4299095;C0524470;C1285116|hip
null|HHIP wt Allele|Finding|false|false|C0019558;C0392905;C1269611;C0022417;C0022122;C0228391;C0019552;C4299095;C0524470;C1285116|hip
null|REG3A wt Allele|Finding|false|false|C0019558;C0392905;C1269611;C0022417;C0022122;C0228391;C0019552;C4299095;C0524470;C1285116|hipnull|Procedure on hip|Procedure|false|false|C0392905;C1269611;C0022417;C0524470;C0019558;C1285116;C0022122;C0228391;C0019552;C4299095|hipnull|Lower extremity>Hip|Anatomy|false|false|C1430701;C0529134;C1505163;C1654726;C0392747;C0011164;C1880269;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C4319952;C5203119;C1547231;C0205082;C1547227;C1561581;C1292890;C1552823;C0575044|hip
null|Hip structure|Anatomy|false|false|C1430701;C0529134;C1505163;C1654726;C0392747;C0011164;C1880269;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C4319952;C5203119;C1547231;C0205082;C1547227;C1561581;C1292890;C1552823;C0575044|hip
null|Structure of habenulopeduncular tract|Anatomy|false|false|C1430701;C0529134;C1505163;C1654726;C0392747;C0011164;C1880269;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C4319952;C5203119;C1547231;C0205082;C1547227;C1561581;C1292890;C1552823;C0575044|hip
null|Bone structure of ischium|Anatomy|false|false|C1430701;C0529134;C1505163;C1654726;C0392747;C0011164;C1880269;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C4319952;C5203119;C1547231;C0205082;C1547227;C1561581;C1292890;C1552823;C0575044|hipnull|Joint problem|Finding|false|false|C0524470;C0392905;C1269611;C0022417;C0019558;C1285116;C0022122;C0228391;C0019552;C4299095|jointnull|null|Anatomy|false|false|C1552823;C0575044;C1430701;C0529134;C1505163;C1654726;C1292890;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C0392747;C0011164;C1880269;C5203119;C1547231;C0205082;C1547227;C1561581;C4319952|joint
null|Joints|Anatomy|false|false|C1552823;C0575044;C1430701;C0529134;C1505163;C1654726;C1292890;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C0392747;C0011164;C1880269;C5203119;C1547231;C0205082;C1547227;C1561581;C4319952|joint
null|Articular system|Anatomy|false|false|C1552823;C0575044;C1430701;C0529134;C1505163;C1654726;C1292890;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C0392747;C0011164;C1880269;C5203119;C1547231;C0205082;C1547227;C1561581;C4319952|jointnull|Joint Device|Device|false|false||jointnull|Articular space|Anatomy|false|false|C0575044|joint spacenull|Joint problem|Finding|false|false|C0392905;C1269611;C0022417;C0224497|jointnull|null|Anatomy|false|false|C0575044;C0015302;C1956089;C5442360|joint
null|Joints|Anatomy|false|false|C0575044;C0015302;C1956089;C5442360|joint
null|Articular system|Anatomy|false|false|C0575044;C0015302;C1956089;C5442360|jointnull|Joint Device|Device|false|false||jointnull|Space (Astronomy)|Phenomenon|false|false||spacenull|Space - property|Modifier|false|false||spacenull|Loss (adaptation)|Finding|false|false||lossnull|Loss (quantitative)|LabModifier|false|false||lossnull|Osteophyte formation|Finding|false|false|C0392905;C1269611;C0022417|osteophyte formationnull|Osteophyte|Disorder|false|false|C0392905;C1269611;C0022417|osteophyte
null|External hyperostosis|Disorder|false|false|C0392905;C1269611;C0022417|osteophytenull|Formation|Finding|false|false||formationnull|Anabolism|Phenomenon|false|false||formationnull|Formations|Modifier|false|false||formationnull|Destructive behavior|Finding|true|false||destructivenull|Bone Tissue, Human|Anatomy|false|false|C0221198|osseous
null|Skeletal bone|Anatomy|false|false|C0221198|osseousnull|Lesion|Finding|false|false|C4520924;C0262950|lesionsnull|impression (attitude)|Finding|false|false||IMPRESSION
null|EKG impression|Finding|false|false||IMPRESSIONnull|Numerous|LabModifier|false|false||Multiplenull|Pulmonary (intended site)|Finding|false|false|C0024109|pulmonarynull|Lung|Anatomy|false|false|C1513183;C0494165;C2707265;C2939419;C0027627;C4522268|pulmonarynull|null|Attribute|false|false|C0024109|pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Metastatic malignant neoplasm to liver|Disorder|false|false|C0205054;C0024109|hepatic metastasesnull|Hepatic|Anatomy|false|false|C2939419;C0027627;C0494165;C1513183|hepaticnull|Metastatic malignant neoplasm|Disorder|false|false|C0205054;C0024109|metastases
null|Neoplasm Metastasis|Disorder|false|false|C0205054;C0024109|metastasesnull|Metastatic Lesion|Finding|false|false|C0024109;C0205054|metastasesnull|Separate|Modifier|false|false||separatenull|True primary (qualifier value)|Time|false|false||primarynull|Primary|Modifier|false|false||primarynull|Lesion|Finding|false|false||lesion
null|null|Finding|false|false||lesionnull|BRIEF Health Literacy Screening Tool|Finding|false|false||Brief
null|Behavior Rating Inventory of Executive Function|Finding|false|false||Briefnull|Brief|Time|false|false||Briefnull|Shortened|Modifier|false|false||Briefnull|Hospital course|Finding|false|false||Hospital Coursenull|null|Attribute|false|false||Hospital Coursenull|Organization unit type - Hospital|Finding|false|false||Hospitalnull|Hospitals|Device|false|false||Hospitalnull|Hospitals|Entity|false|false||Hospitalnull|Hospital environment|Modifier|false|false||Hospitalnull|Course|Time|false|false||Coursenull|Recent|Time|false|false||recentlynull|Metastatic malignant neoplasm|Disorder|false|false||metastatic cancer
null|Disseminated Malignant Neoplasm|Disorder|false|false||metastatic cancer
null|Neoplasm Metastasis|Disorder|false|false||metastatic cancernull|metastatic qualifier|Finding|false|false||metastatic
null|Metastatic to|Finding|false|false||metastaticnull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|unknown vaccine or immune globulin|Drug|false|false||unknown
null|Unknown - Vaccines administered|Drug|false|false||unknown
null|Unknown - Vaccines administered|Drug|false|false||unknown
null|unknown vaccine or immune globulin|Drug|false|false||unknownnull|Unknown - mode of arrival code|Finding|false|false||unknown
null|Unknown - Special Program Code|Finding|false|false||unknown
null|Unknown - Production Class Code|Finding|false|false||unknown
null|Unknown - Patient Outcome|Finding|false|false||unknown
null|Unknown - Recreational Drug Use Code|Finding|false|false||unknown
null|Unknown - Escort Required|Finding|false|false||unknown
null|Unknown - Transport Arranged|Finding|false|false||unknown
null|Unknown - Living Arrangement|Finding|false|false||unknown
null|Unknown - Employment Status|Finding|false|false||unknown
null|Unknown - Relationship|Finding|false|false||unknown
null|Unknown - publishing section|Finding|false|false||unknown
null|Unknown Publicity Code|Finding|false|false||unknown
null|Unknown - Event reason|Finding|false|false||unknown
null|Unknown - Religion|Finding|false|false||unknown
null|Unknown - Organ Donor Code|Finding|false|false||unknown
null|unknown - NullFlavor|Finding|false|false||unknown
null|Unknown - Notify Clergy Code|Finding|false|false||unknown
null|Unknown - Administrative Gender|Finding|false|false||unknown
null|Unknown - Patient Condition Code|Finding|false|false||unknown
null|Unknown - Living Will Code|Finding|false|false||unknown
null|Marital Status - Unknown|Finding|false|false||unknown
null|Unknown - Patient Class|Finding|false|false||unknown
null|Unknown - Event Expected|Finding|false|false||unknown
null|Unknown - Expanded yes/no indicator|Finding|false|false||unknown
null|Unknown - Immunization Registry Status|Finding|false|false||unknown
null|Unknown - Container status|Finding|false|false||unknown
null|Unknown - CWE statuses|Finding|false|false||unknown
null|Unknown - Patient_s Relationship to Insured|Finding|false|false||unknown
null|Unknown - Job Status|Finding|false|false||unknown
null|Unknown - Precaution Code|Finding|false|false||unknown
null|Unknown - Contact Role|Finding|false|false||unknown
null|Unknown - Living Dependency|Finding|false|false||unknownnull|Ethnic group unknown|Subject|false|false||unknownnull|Unknown - Allergy Severity|Modifier|false|false||unknown
null|Unknown - HL7 update mode|Modifier|false|false||unknown
null|Unknown|Modifier|false|false||unknownnull|True primary (qualifier value)|Time|false|false||primarynull|Primary|Modifier|false|false||primarynull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|Vomiting|Finding|false|false||vomitingnull|Fever symptoms (finding)|Finding|false|false||fever
null|Fever|Finding|false|false||fevernull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Fever symptoms (finding)|Finding|false|false||Fever
null|Fever|Finding|false|false||Fevernull|Leukocytosis|Disorder|false|false||leukocytosisnull|Blood leukocyte number above reference range|Finding|false|false||leukocytosisnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Fever symptoms (finding)|Finding|false|false||fever
null|Fever|Finding|false|false||fevernull|Leukocytosis|Disorder|false|false||leukocytosisnull|Blood leukocyte number above reference range|Finding|false|false||leukocytosisnull|Initially|Time|false|false||initiallynull|SLC35G1 gene|Finding|false|false||post
null|DESI1 gene|Finding|false|false||postnull|Post Device|Device|false|false||postnull|Post|Time|false|false||postnull|Obstructed|Finding|false|false||obstructivenull|Peptide Nucleic Acids|Drug|false|false||PNAnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|cefepime|Drug|false|false||cefepime
null|cefepime|Drug|false|false||cefepimenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Trunk structure|Anatomy|false|false||torsonull|Continuous|Finding|false|false||ongoingnull|Primary malignant neoplasm|Disorder|false|false||malignancy
null|Malignant Neoplasms|Disorder|false|false||malignancynull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Primary Neoplasm|Disorder|true|false||primary tumornull|True primary (qualifier value)|Time|false|false||primarynull|Primary|Modifier|false|false||primarynull|Neoplasms|Disorder|true|false||tumornull|Tumor Mass|Finding|true|false||tumor
null|null|Finding|true|false||tumornull|Concern|Finding|true|false||concernnull|Pneumonia|Disorder|false|false||pneumonianull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Feel Weak (question)|Finding|false|false||weak
null|Weakness|Finding|false|false||weaknull|Weak|Modifier|false|false||weaknull|Unable|Finding|false|false||unablenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Living Alone|Finding|false|false||alonenull|alone - group size|Subject|false|false||alonenull|Singular|LabModifier|false|false||alonenull|Diagnostic Service Section ID - Physical Therapy|Finding|false|false||physical therapynull|Physical therapy|Procedure|false|false||physical therapynull|Physical therapy (field)|Title|false|false||physical therapynull|physical examination (physical finding)|Finding|false|false||physical
null|Physical|Finding|false|false||physicalnull|Physical Examination|Procedure|false|false||physicalnull|Therapy Object (animal model)|Finding|false|false||therapy
null|therapeutic aspects|Finding|false|false||therapynull|Therapeutic procedure|Procedure|false|false||therapynull|Rehab facility|Device|false|false||rehab facilitynull|Rehab facility|Entity|false|false||rehab facilitynull|Rehabilitation therapy|Procedure|false|false||rehabnull|ADMIN.FACILITY|Finding|false|false||facilitynull|Facility (object)|Device|false|false||facilitynull|Pediatric failure to thrive|Disorder|false|false||Failure to thrive
null|Failure to Thrive|Disorder|false|false||Failure to thrivenull|Failure (biologic function)|Finding|false|false||Failure
null|Failure|Finding|false|false||Failure
null|Personal failure|Finding|false|false||Failurenull|Thrive|Drug|false|false||thrive
null|Thrive|Drug|false|false||thrivenull|Transnasal humidified rapid-insufflation ventilatory exchange|Procedure|false|false||thrivenull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|6 weeks|Time|false|false||6 weeksnull|week|Time|false|false||weeksnull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|Vomiting|Finding|false|false||vomitingnull|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group|Finding|false|false||poor
null|Patient Condition Code - Poor|Finding|false|false||poornull|Poverty|Subject|false|false||poornull|Language Proficiency - Poor|Modifier|false|false||poor
null|Specimen Quality - Poor|Modifier|false|false||poor
null|Poor - grade|Modifier|false|false||poor
null|Poor - qualifier|Modifier|false|false||poornull|Intake|Finding|false|false||intakenull|Measurement of fluid intake|Procedure|false|false||intake
null|Intake (treatment)|Procedure|false|false||intakenull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Hepatomegaly|Finding|false|false|C4037986;C1278929;C0023884|enlarged livernull|Enlargement procedure|Procedure|false|false|C4037986;C1278929;C0023884|enlargednull|Enlarged|Modifier|false|false||enlargednull|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|liver
null|liver extract|Drug|false|false|C4037986;C1278929;C0023884|liver
null|liver extract|Drug|false|false|C4037986;C1278929;C0023884|liver
null|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|liver
null|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|livernull|Benign neoplasm of liver|Disorder|false|false|C4037986;C1278929;C0023884|liver
null|Liver diseases|Disorder|false|false|C4037986;C1278929;C0023884|livernull|Liver problem|Finding|false|false|C4037986;C1278929;C0023884|livernull|Procedures on liver|Procedure|false|false|C4037986;C1278929;C0023884|livernull|Abdomen>Liver|Anatomy|false|false|C0577060;C0872387;C0023895;C0496870;C0019209;C0721399;C0023899;C1293134|liver
null|null|Anatomy|false|false|C0577060;C0872387;C0023895;C0496870;C0019209;C0721399;C0023899;C1293134|liver
null|Liver|Anatomy|false|false|C0577060;C0872387;C0023895;C0496870;C0019209;C0721399;C0023899;C1293134|livernull|Defecation|Finding|false|false|C0021853|bowel movementsnull|Intestines|Anatomy|false|false|C0011135|bowelnull|Movement|Finding|false|false||movementsnull|Pass (indicator)|Finding|false|false||passnull|Gas - SpecimenType|Drug|false|false||gas
null|Gases|Drug|false|false||gas
null|Gas Dosage Form|Drug|false|false||gasnull|Gas - Specimen Source Codes|Finding|false|false||gas
null|gastrointestinal gas|Finding|false|false||gas
null|PAGR1 wt Allele|Finding|false|false||gas
null|GALNS wt Allele|Finding|false|false||gas
null|GALNS gene|Finding|false|false||gas
null|GAST wt Allele|Finding|false|false||gas
null|GAST gene|Finding|false|false||gas
null|germacrene-A synthase activity|Finding|false|false||gas
null|PAGR1 gene|Finding|false|false||gasnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Albumin|Drug|false|false||albumin
null|Albumins|Drug|false|false||albumin
null|Albumins|Drug|false|false||albumin
null|Albumin|Drug|false|false||albuminnull|Albumin metabolic function|Finding|false|false||albumin
null|ALB gene|Finding|false|false||albuminnull|Albumin measurement|Procedure|false|false||albuminnull|Ketones|Drug|false|false||ketonesnull|Toxic effect of ketones|Disorder|false|false||ketonesnull|Urine ketone test|Procedure|false|false||ketones
null|Ketone bodies measurement, quantitative|Procedure|false|false||ketonesnull|Portion of urine|Finding|false|false||urine
null|null|Finding|false|false||urine
null|Urine|Finding|false|false||urine
null|In Urine|Finding|false|false||urine
null|Urine specimen|Finding|false|false||urinenull|Weight Loss|Finding|false|false||weight loss
null|Losing Weight (question)|Finding|false|false||weight lossnull|Measured weight loss (observable entity)|LabModifier|false|false||weight lossnull|infant weight for previous delivery (history)|Finding|false|false||weight
null|Weight symptom (finding)|Finding|false|false||weightnull|Weighing patient|Procedure|false|false||weightnull|null|Attribute|false|false||weightnull|Body Weight|Subject|false|false||weightnull|Importance Weight|Modifier|false|false||weightnull|Weight|LabModifier|false|false||weightnull|Loss (adaptation)|Finding|false|false||lossnull|Loss (quantitative)|LabModifier|false|false||lossnull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|Peripheral edema|Finding|false|false||peripheral edemanull|Peripheral|Modifier|false|false||peripheralnull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Malnutrition|Disorder|false|false||poor nutritionnull|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group|Finding|false|false||poor
null|Patient Condition Code - Poor|Finding|false|false||poornull|Poverty|Subject|false|false||poornull|Language Proficiency - Poor|Modifier|false|false||poor
null|Specimen Quality - Poor|Modifier|false|false||poor
null|Poor - grade|Modifier|false|false||poor
null|Poor - qualifier|Modifier|false|false||poornull|Nutrition (function)|Finding|false|false||nutrition
null|Nutritional status|Finding|false|false||nutrition
null|Nutrition outcomes|Finding|false|false||nutritionnull|Feeding and dietary regimes|Procedure|false|false||nutrition
null|Nutritional Study|Procedure|false|false||nutritionnull|Science of nutrition|Title|false|false||nutritionnull|Starvation|Finding|false|false||starvationnull|Ketosis|Disorder|false|false||ketosis
null|Ketoacidosis|Disorder|false|false||ketosisnull|Nutrition (function)|Finding|false|false||Nutrition
null|Nutritional status|Finding|false|false||Nutrition
null|Nutrition outcomes|Finding|false|false||Nutritionnull|Feeding and dietary regimes|Procedure|false|false||Nutrition
null|Nutritional Study|Procedure|false|false||Nutritionnull|Science of nutrition|Title|false|false||Nutritionnull|Consultation|Procedure|false|false||consultnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Hospital Stay|Time|false|false||hospital staynull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Platelet Glycoprotein 4, human|Drug|false|false|C0001527|fat
null|FAT1 protein, human|Drug|false|false|C0001527|fat
null|FAT1 protein, human|Drug|false|false|C0001527|fat
null|Fatty acid glycerol esters|Drug|false|false|C0001527|fat
null|Fatty acid glycerol esters|Drug|false|false|C0001527|fatnull|Platelet Glycoprotein 4, human|Finding|false|false|C0001527|fat
null|CD36 gene|Finding|false|false|C0001527|fat
null|FAT1 gene|Finding|false|false|C0001527|fat
null|CD36 wt Allele|Finding|false|false|C0001527|fat
null|FAT1 wt Allele|Finding|false|false|C0001527|fatnull|doxorubicin/fluorouracil/triazinate protocol|Procedure|false|false|C0001527|fatnull|Adipose tissue|Anatomy|false|false|C0279453;C1435181;C0015677;C3887682;C3887682;C0812278;C1705088;C1708004;C1366645|fatnull|Obese build|Subject|false|false||fatnull|Fantse Language|Entity|false|false||fatnull|CARNATION INSTANT|Drug|false|false||Carnation Instantnull|Carnation|Entity|false|false||Carnationnull|Breakfast|Finding|false|false||Breakfastnull|With breakfast|Time|false|false||Breakfastnull|Chronic back pain|Finding|false|false||Chronic back painnull|Chronic - Admission Level of Care Code|Finding|false|false||Chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||Chronicnull|chronic|Time|false|false||Chronicnull|Back Pain|Finding|false|false||back painnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|gabapentin|Drug|false|false||gabapentin
null|gabapentin|Drug|false|false||gabapentinnull|Cancer patients and suicide and depression|Disorder|false|false||Depression
null|Mental Depression|Disorder|false|false||Depression
null|Depressive disorder|Disorder|false|false||Depression
null|Depressed mood|Disorder|false|false||Depressionnull|Depression - motion|Finding|false|false||Depression
null|null|Finding|false|false||Depressionnull|Depression - recess|Modifier|false|false||Depressionnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|bupropion|Drug|false|false||bupropion
null|bupropion|Drug|false|false||bupropionnull|sertraline|Drug|false|false||sertraline
null|sertraline|Drug|false|false||sertralinenull|hydrochlorothiazide|Drug|false|false||HCTZ
null|hydrochlorothiazide|Drug|false|false||HCTZnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|hydrochlorothiazide|Drug|false|false||hctz
null|hydrochlorothiazide|Drug|false|false||hctznull|Hospitalization|Procedure|false|false||hospitalizationnull|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group|Finding|false|false||poor
null|Patient Condition Code - Poor|Finding|false|false||poornull|Poverty|Subject|false|false||poornull|Language Proficiency - Poor|Modifier|false|false||poor
null|Specimen Quality - Poor|Modifier|false|false||poor
null|Poor - grade|Modifier|false|false||poor
null|Poor - qualifier|Modifier|false|false||poornull|Intake|Finding|false|false||intakenull|Measurement of fluid intake|Procedure|false|false||intake
null|Intake (treatment)|Procedure|false|false||intakenull|Concern|Finding|false|false||concernnull|dehydration (Na, H2O)|Disorder|false|false||dehydration
null|Dehydration|Disorder|false|false||dehydrationnull|Dehydration procedure|Procedure|false|false||dehydrationnull|Systemic arterial pressure|Finding|false|false||Blood pressuresnull|Blood and lymphatic system disorders|Disorder|false|false||Bloodnull|peripheral blood|Finding|false|false||Blood
null|Blood|Finding|false|false||Blood
null|In Blood|Finding|false|false||Bloodnull|Pressure (finding)|Finding|false|false||pressuresnull|null|Phenomenon|false|false||pressuresnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|hydrochlorothiazide|Drug|false|false||HCTZ
null|hydrochlorothiazide|Drug|false|false||HCTZnull|Issue (document)|Finding|false|false||issue
null|Problem|Finding|false|false||issuenull|Issue (action)|Event|false|false||issuenull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|Hyperlipidemia|Disorder|false|false||Hyperlipidemia
null|Hyperlipoproteinemias|Disorder|false|false||Hyperlipidemianull|Serum lipids high (finding)|Finding|false|false||Hyperlipidemianull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|metastatic qualifier|Finding|false|false|C1184743|metastatic
null|Metastatic to|Finding|false|false|C1184743|metastaticnull|Process Pharmacologic Substance|Drug|false|false|C1184743|processnull|Process (qualifier value)|Finding|false|false|C1184743|processnull|bony process|Anatomy|false|false|C1522484;C0036525;C1951340;C4521054;C1522240|processnull|Process|Phenomenon|false|false|C1184743|processnull|Hydroxymethylglutaryl-CoA Reductase Inhibitors|Drug|false|false||statin
null|Hydroxymethylglutaryl-CoA Reductase Inhibitors|Drug|false|false||statinnull|EEF1A2 gene|Finding|false|false||statinnull|3-hydroxy-3-methylglutaryl-coenzyme A reductase inhibitor (disposition)|Modifier|false|false||statinnull|during hospitalization|Time|false|false||during hospitalizationnull|Hospitalization|Procedure|false|false||hospitalizationnull|Medical referral type|Finding|false|false||medical
null|Medical|Finding|false|false||medical
null|Medical school type|Finding|false|false||medicalnull|Medical service|Procedure|false|false||medicalnull|GDC Regimen Terminology|Finding|false|false||regimennull|Treatment Protocols|Procedure|false|false||regimennull|Insomnia homeopathic medication|Drug|false|false||Insomnianull|Sleeplessness|Finding|false|false||Insomnianull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|trazodone|Drug|false|false||trazodone
null|trazodone|Drug|false|false||trazodonenull|Transition Mutation|Disorder|false|false||TRANSITIONnull|Transition (action)|Event|false|false||TRANSITIONnull|MDF Attribute Type - Code|Finding|false|false||CODE
null|A Codes|Finding|false|false||CODE
null|Code|Finding|false|false||CODEnull|Coding|Event|false|false||CODEnull|Full|Modifier|false|false||FULLnull|Confirmation|Finding|false|false||Confirmednull|Confirmed by|Modifier|false|false||Confirmednull|Contact - HL7 Attribution|Finding|false|false||CONTACT
null|Contact with|Finding|false|false||CONTACT
null|Communication Contact|Finding|false|false||CONTACTnull|contact person|Subject|false|false||CONTACTnull|Physical contact|Phenomenon|false|false||CONTACTnull|Personal Contact|Event|false|false||CONTACTnull|Relationship - Friend|Finding|false|false||friendnull|friend|Subject|false|false||friendnull|hydrochlorothiazide|Drug|false|false||HCTZ
null|hydrochlorothiazide|Drug|false|false||HCTZnull|On admission|Time|false|false||on admissionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|consider|Finding|false|false||considernull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|Platelet Glycoprotein 4, human|Drug|false|false|C0001527|fat
null|FAT1 protein, human|Drug|false|false|C0001527|fat
null|FAT1 protein, human|Drug|false|false|C0001527|fat
null|Fatty acid glycerol esters|Drug|false|false|C0001527|fat
null|Fatty acid glycerol esters|Drug|false|false|C0001527|fatnull|Platelet Glycoprotein 4, human|Finding|false|false|C0001527|fat
null|CD36 gene|Finding|false|false|C0001527|fat
null|FAT1 gene|Finding|false|false|C0001527|fat
null|CD36 wt Allele|Finding|false|false|C0001527|fat
null|FAT1 wt Allele|Finding|false|false|C0001527|fatnull|doxorubicin/fluorouracil/triazinate protocol|Procedure|false|false|C0001527|fatnull|Adipose tissue|Anatomy|false|false|C3887682;C0812278;C1705088;C1708004;C1366645;C2698559;C0279453;C1435181;C0015677;C3887682|fatnull|Obese build|Subject|false|false||fatnull|Fantse Language|Entity|false|false||fatnull|CARNATION INSTANT|Drug|false|false||Carnation Instantnull|Carnation|Entity|false|false||Carnationnull|Breakfast|Finding|false|false|C0001527|Breakfastnull|With breakfast|Time|false|false||Breakfastnull|Meal (occasion for eating)|Finding|false|false||mealsnull|With meals|Time|false|false||mealsnull|Neoplasms|Disorder|false|false||oncologynull|oncology services|Procedure|false|false||oncologynull|oncology (field)|Title|false|false||oncologynull|Further|Modifier|false|false||furthernull|Diagnosis Classification - Diagnosis|Finding|false|false||diagnosis
null|diagnosis aspects|Finding|false|false||diagnosisnull|Diagnosis|Procedure|false|false||diagnosisnull|null|Attribute|false|false||diagnosisnull|Disease Management|Procedure|false|false||managementnull|Management Occupations|Subject|false|false||managementnull|Management procedure|Event|false|false||management
null|Administration occupational activities|Event|false|false||managementnull|Primary malignant neoplasm|Disorder|false|false||malignancy
null|Malignant Neoplasms|Disorder|false|false||malignancynull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|MEDICATION LIST|Finding|false|false||Medication listnull|Pharmaceutical Preparations|Drug|false|false||Medicationnull|medication - HL7 publishing domain|Finding|false|false||Medication
null|Medications|Finding|false|false||Medicationnull|List|Finding|false|false||list
null|Sequence Data Type|Finding|false|false||listnull|Accurate (qualifier value)|Modifier|false|false||accuratenull|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||completenull|Completion Status for valid values - Complete|Finding|false|false||complete
null|Data operation - complete|Finding|false|false||complete
null|Finish - dosing instruction imperative|Finding|false|false||completenull|Complete|Modifier|false|false||completenull|albuterol|Drug|false|false||Albuterol
null|albuterol|Drug|false|false||Albuterolnull|Inhaler (unit of presentation)|Finding|false|false||Inhalernull|Inhaler|Device|false|false||Inhalernull|Inhaler Dosing Unit|LabModifier|false|false||Inhalernull|Puff Dosing Unit|LabModifier|false|false||PUFF
null|Picofarad|LabModifier|false|false||PUFFnull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Dyspnea|Finding|false|false||SOBnull|bupropion|Drug|false|false||BuPROPion
null|bupropion|Drug|false|false||BuPROPionnull|Daily|Time|false|false||DAILYnull|gabapentin|Drug|false|false||Gabapentin
null|gabapentin|Drug|false|false||Gabapentinnull|sertraline|Drug|false|false||Sertraline
null|sertraline|Drug|false|false||Sertralinenull|Daily|Time|false|false||DAILYnull|simvastatin|Drug|false|false||Simvastatin
null|simvastatin|Drug|false|false||Simvastatinnull|Daily|Time|false|false||DAILYnull|trazodone|Drug|false|false||traZODONE
null|trazodone|Drug|false|false||traZODONEnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Sleep brand of diphenhydramine hydrochloride|Drug|false|false||sleep
null|Sleep brand of diphenhydramine hydrochloride|Drug|false|false||sleepnull|Sleep|Finding|false|false||sleepnull|ibuprofen|Drug|false|false||Ibuprofen
null|ibuprofen|Drug|false|false||Ibuprofennull|Every twelve hours|Time|false|false||Q12Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|hydrochlorothiazide|Drug|false|false||Hydrochlorothiazide
null|hydrochlorothiazide|Drug|false|false||Hydrochlorothiazidenull|Daily|Time|false|false||DAILYnull|ondansetron|Drug|false|false||Ondansetron
null|ondansetron|Drug|false|false||Ondansetronnull|Every eight hours|Time|false|false||Q8Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|albuterol|Drug|false|false||Albuterol
null|albuterol|Drug|false|false||Albuterolnull|Inhaler (unit of presentation)|Finding|false|false||Inhalernull|Inhaler|Device|false|false||Inhalernull|Inhaler Dosing Unit|LabModifier|false|false||Inhalernull|Puff Dosing Unit|LabModifier|false|false||PUFF
null|Picofarad|LabModifier|false|false||PUFFnull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Dyspnea|Finding|false|false||SOBnull|bupropion|Drug|false|false||BuPROPion
null|bupropion|Drug|false|false||BuPROPionnull|Daily|Time|false|false||DAILYnull|gabapentin|Drug|false|false||Gabapentin
null|gabapentin|Drug|false|false||Gabapentinnull|sertraline|Drug|false|false||Sertraline
null|sertraline|Drug|false|false||Sertralinenull|Daily|Time|false|false||DAILYnull|trazodone|Drug|false|false||traZODONE
null|trazodone|Drug|false|false||traZODONEnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Sleep brand of diphenhydramine hydrochloride|Drug|false|false||sleep
null|Sleep brand of diphenhydramine hydrochloride|Drug|false|false||sleepnull|Sleep|Finding|false|false||sleepnull|ondansetron|Drug|false|false||Ondansetron
null|ondansetron|Drug|false|false||Ondansetronnull|Every eight hours|Time|false|false||Q8Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|bisacodyl|Drug|false|false||Bisacodyl
null|bisacodyl|Drug|false|false||Bisacodylnull|Daily|Time|false|false||DAILYnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Constipation|Finding|false|false||constipationnull|oxycodone|Drug|false|false||OxycoDONE
null|oxycodone|Drug|false|false||OxycoDONEnull|Oxycodone measurement|Procedure|false|false||OxycoDONEnull|Immediate Release Dosage Form|Drug|false|false||Immediate Releasenull|Query Priority - Immediate|Finding|false|false||Immediate
null|immediate - ResponseCode|Finding|false|false||Immediatenull|Immediate|Time|false|false||Immediate
null|Stat (do immediately)|Time|false|false||Immediatenull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Sedation|Finding|false|false||sedation
null|Sedated state|Finding|false|false||sedationnull|Sedation procedure|Procedure|false|false||sedationnull|oxycodone|Drug|false|false||oxycodone
null|oxycodone|Drug|false|false||oxycodonenull|Oxycodone measurement|Procedure|false|false||oxycodonenull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false|C0230028;C0226896|by mouthnull|Oral cavity|Anatomy|false|false|C1527415|mouth
null|Oral region|Anatomy|false|false|C1527415|mouthnull|6 Hours|Time|false|false||6 hoursnull|Hour|Time|false|false||hoursnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|enoxaparin sodium|Drug|false|false||Enoxaparin Sodium
null|enoxaparin sodium|Drug|false|false||Enoxaparin Sodiumnull|enoxaparin|Drug|false|false||Enoxaparin
null|enoxaparin|Drug|false|false||Enoxaparinnull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|Daily|Time|false|false||DAILYnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|long-term care|Procedure|false|false||Extended Carenull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|In care (finding)|Finding|false|false||Care
null|Continuity Assessment Record and Evaluation|Finding|false|false||Carenull|care activity|Event|false|false||Carenull|ADMIN.FACILITY|Finding|false|false||Facilitynull|Facility (object)|Device|false|false||Facilitynull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Metastatic malignant neoplasm|Disorder|false|false||Metastatic disease
null|Metastatic Neoplasm|Disorder|false|false||Metastatic disease
null|Neoplasm Metastasis|Disorder|false|false||Metastatic diseasenull|Metastatic Lesion|Finding|false|false||Metastatic diseasenull|metastatic qualifier|Finding|false|false||Metastatic
null|Metastatic to|Finding|false|false||Metastaticnull|Disease|Disorder|false|false||diseasenull|unknown vaccine or immune globulin|Drug|false|false||unknown
null|Unknown - Vaccines administered|Drug|false|false||unknown
null|Unknown - Vaccines administered|Drug|false|false||unknown
null|unknown vaccine or immune globulin|Drug|false|false||unknownnull|Unknown - mode of arrival code|Finding|false|false||unknown
null|Unknown - Special Program Code|Finding|false|false||unknown
null|Unknown - Production Class Code|Finding|false|false||unknown
null|Unknown - Patient Outcome|Finding|false|false||unknown
null|Unknown - Recreational Drug Use Code|Finding|false|false||unknown
null|Unknown - Escort Required|Finding|false|false||unknown
null|Unknown - Transport Arranged|Finding|false|false||unknown
null|Unknown - Living Arrangement|Finding|false|false||unknown
null|Unknown - Employment Status|Finding|false|false||unknown
null|Unknown - Relationship|Finding|false|false||unknown
null|Unknown - publishing section|Finding|false|false||unknown
null|Unknown Publicity Code|Finding|false|false||unknown
null|Unknown - Event reason|Finding|false|false||unknown
null|Unknown - Religion|Finding|false|false||unknown
null|Unknown - Organ Donor Code|Finding|false|false||unknown
null|unknown - NullFlavor|Finding|false|false||unknown
null|Unknown - Notify Clergy Code|Finding|false|false||unknown
null|Unknown - Administrative Gender|Finding|false|false||unknown
null|Unknown - Patient Condition Code|Finding|false|false||unknown
null|Unknown - Living Will Code|Finding|false|false||unknown
null|Marital Status - Unknown|Finding|false|false||unknown
null|Unknown - Patient Class|Finding|false|false||unknown
null|Unknown - Event Expected|Finding|false|false||unknown
null|Unknown - Expanded yes/no indicator|Finding|false|false||unknown
null|Unknown - Immunization Registry Status|Finding|false|false||unknown
null|Unknown - Container status|Finding|false|false||unknown
null|Unknown - CWE statuses|Finding|false|false||unknown
null|Unknown - Patient_s Relationship to Insured|Finding|false|false||unknown
null|Unknown - Job Status|Finding|false|false||unknown
null|Unknown - Precaution Code|Finding|false|false||unknown
null|Unknown - Contact Role|Finding|false|false||unknown
null|Unknown - Living Dependency|Finding|false|false||unknownnull|Ethnic group unknown|Subject|false|false||unknownnull|Unknown - Allergy Severity|Modifier|false|false||unknown
null|Unknown - HL7 update mode|Modifier|false|false||unknown
null|Unknown|Modifier|false|false||unknownnull|True primary (qualifier value)|Time|false|false||primarynull|Primary|Modifier|false|false||primarynull|Weakness|Finding|false|false||Weakness
null|Asthenia|Finding|false|false||Weaknessnull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Tumor Burden|Procedure|false|false||tumor burdennull|Neoplasms|Disorder|false|false||tumornull|Tumor Mass|Finding|false|false||tumor
null|null|Finding|false|false||tumornull|Burden|Finding|false|false||burdennull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Disease|Disorder|false|false||Conditionnull|Logical Condition|Finding|false|false||Conditionnull|null|Attribute|false|false||Conditionnull|Condition|Modifier|false|false||Conditionnull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Coordination of Benefits - Independent|Finding|false|false||Independent
null|Religious Affiliation - Independent|Finding|false|false||Independent
null|Independence|Finding|false|false||Independent
null|Independently able|Finding|false|false||Independentnull|Discharge instructions|Finding|false|false||Discharge Instructionsnull|hospital discharge instructions (treatment)|Procedure|false|false||Discharge Instructionsnull|null|Attribute|false|false||Discharge Instructionsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructionsnull|FBXW7-AS1 gene|Finding|false|false||Dearnull|Processing type - Evaluation|Finding|false|false||evaluationnull|Evaluation procedure|Procedure|false|false||evaluation
null|Evaluation|Procedure|false|false||evaluationnull|Several|LabModifier|false|false||severalnull|week|Time|false|false||weeksnull|Weakness|Finding|false|false||weakness
null|Asthenia|Finding|false|false||weaknessnull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|Marker Device|Device|false|false||markersnull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|Initially|Time|false|false||initiallynull|Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE|Drug|false|false||antibiotics
null|Antibiotics|Drug|false|false||antibiotics
null|Antibiotics, ophthalmologic|Drug|false|false||antibiotics
null|Antibiotics, Gynecological|Drug|false|false||antibiotics
null|antibiotics, intestinal|Drug|false|false||antibiotics
null|Antibiotic throat preparations|Drug|false|false||antibiotics
null|Antibiotics, Antitubercular|Drug|false|false||antibiotics
null|Antibiotics for systemic use|Drug|false|false||antibiotics
null|Antifungal Antibiotics, Topical|Drug|false|false||antibioticsnull|Radionuclide Imaging|Procedure|false|false|C0460005|scan
null|Scanning|Procedure|false|false|C0460005|scannull|Trunk structure|Anatomy|false|false|C0034606;C0441633|torsonull|Metastatic malignant neoplasm|Disorder|false|false||metastatic disease
null|Metastatic Neoplasm|Disorder|false|false||metastatic disease
null|Neoplasm Metastasis|Disorder|false|false||metastatic diseasenull|Metastatic Lesion|Finding|false|false||metastatic diseasenull|metastatic qualifier|Finding|false|false||metastatic
null|Metastatic to|Finding|false|false||metastaticnull|Disease|Disorder|false|false||diseasenull|Carcinoma of unknown primary|Disorder|false|false||cancer of unknown originnull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Unknown (origin) (qualifier value)|Finding|false|false||unknown originnull|unknown vaccine or immune globulin|Drug|false|false||unknown
null|Unknown - Vaccines administered|Drug|false|false||unknown
null|Unknown - Vaccines administered|Drug|false|false||unknown
null|unknown vaccine or immune globulin|Drug|false|false||unknownnull|Unknown - mode of arrival code|Finding|false|false||unknown
null|Unknown - Special Program Code|Finding|false|false||unknown
null|Unknown - Production Class Code|Finding|false|false||unknown
null|Unknown - Patient Outcome|Finding|false|false||unknown
null|Unknown - Recreational Drug Use Code|Finding|false|false||unknown
null|Unknown - Escort Required|Finding|false|false||unknown
null|Unknown - Transport Arranged|Finding|false|false||unknown
null|Unknown - Living Arrangement|Finding|false|false||unknown
null|Unknown - Employment Status|Finding|false|false||unknown
null|Unknown - Relationship|Finding|false|false||unknown
null|Unknown - publishing section|Finding|false|false||unknown
null|Unknown Publicity Code|Finding|false|false||unknown
null|Unknown - Event reason|Finding|false|false||unknown
null|Unknown - Religion|Finding|false|false||unknown
null|Unknown - Organ Donor Code|Finding|false|false||unknown
null|unknown - NullFlavor|Finding|false|false||unknown
null|Unknown - Notify Clergy Code|Finding|false|false||unknown
null|Unknown - Administrative Gender|Finding|false|false||unknown
null|Unknown - Patient Condition Code|Finding|false|false||unknown
null|Unknown - Living Will Code|Finding|false|false||unknown
null|Marital Status - Unknown|Finding|false|false||unknown
null|Unknown - Patient Class|Finding|false|false||unknown
null|Unknown - Event Expected|Finding|false|false||unknown
null|Unknown - Expanded yes/no indicator|Finding|false|false||unknown
null|Unknown - Immunization Registry Status|Finding|false|false||unknown
null|Unknown - Container status|Finding|false|false||unknown
null|Unknown - CWE statuses|Finding|false|false||unknown
null|Unknown - Patient_s Relationship to Insured|Finding|false|false||unknown
null|Unknown - Job Status|Finding|false|false||unknown
null|Unknown - Precaution Code|Finding|false|false||unknown
null|Unknown - Contact Role|Finding|false|false||unknown
null|Unknown - Living Dependency|Finding|false|false||unknownnull|Ethnic group unknown|Subject|false|false||unknownnull|Unknown - Allergy Severity|Modifier|false|false||unknown
null|Unknown - HL7 update mode|Modifier|false|false||unknown
null|Unknown|Modifier|false|false||unknownnull|Participation Type - origin|Finding|false|false||origin
null|National origin|Finding|false|false||originnull|Beginning|Time|false|false||originnull|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|liver
null|liver extract|Drug|false|false|C4037986;C1278929;C0023884|liver
null|liver extract|Drug|false|false|C4037986;C1278929;C0023884|liver
null|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|liver
null|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|livernull|Benign neoplasm of liver|Disorder|false|false|C4037986;C1278929;C0023884;C0024109|liver
null|Liver diseases|Disorder|false|false|C4037986;C1278929;C0023884;C0024109|livernull|Liver problem|Finding|false|false|C4037986;C1278929;C0023884;C0024109|livernull|Procedures on liver|Procedure|false|false|C4037986;C1278929;C0023884;C0024109|livernull|Abdomen>Liver|Anatomy|false|false|C0023895;C0496870;C0872387;C0721399;C0023899;C0577060|liver
null|null|Anatomy|false|false|C0023895;C0496870;C0872387;C0721399;C0023899;C0577060|liver
null|Liver|Anatomy|false|false|C0023895;C0496870;C0872387;C0721399;C0023899;C0577060|livernull|Lung|Anatomy|false|false|C0872387;C0023895;C0496870;C0577060|lungsnull|Weakness|Finding|false|false||weakness
null|Asthenia|Finding|false|false||weaknessnull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|most likely|Finding|false|false||most likelynull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Hepatomegaly|Finding|false|false|C4037986;C1278929;C0023884|enlarged livernull|Enlargement procedure|Procedure|false|false|C4037986;C1278929;C0023884|enlargednull|Enlarged|Modifier|false|false||enlargednull|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|liver
null|liver extract|Drug|false|false|C4037986;C1278929;C0023884|liver
null|liver extract|Drug|false|false|C4037986;C1278929;C0023884|liver
null|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|liver
null|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|livernull|Benign neoplasm of liver|Disorder|false|false|C4037986;C1278929;C0023884|liver
null|Liver diseases|Disorder|false|false|C4037986;C1278929;C0023884|livernull|Liver problem|Finding|false|false|C4037986;C1278929;C0023884|livernull|Procedures on liver|Procedure|false|false|C4037986;C1278929;C0023884|livernull|Abdomen>Liver|Anatomy|false|false|C0023895;C0496870;C1293134;C0721399;C0023899;C0019209;C0577060;C0872387|liver
null|null|Anatomy|false|false|C0023895;C0496870;C1293134;C0721399;C0023899;C0019209;C0577060;C0872387|liver
null|Liver|Anatomy|false|false|C0023895;C0496870;C1293134;C0721399;C0023899;C0019209;C0577060;C0872387|livernull|Oncologists|Subject|false|false||oncologistnull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|Further|Modifier|false|false||furthernull|Diagnosis Classification - Diagnosis|Finding|false|false||diagnosis
null|diagnosis aspects|Finding|false|false||diagnosisnull|Diagnosis|Procedure|false|false||diagnosisnull|null|Attribute|false|false||diagnosisnull|Biomaterial Treatment|Finding|false|false||treatment
null|Treating|Finding|false|false||treatment
null|therapeutic aspects|Finding|false|false||treatmentnull|treatment - ActInformationManagementReason|Procedure|false|false||treatment
null|Administration (procedure)|Procedure|false|false||treatment
null|Therapeutic procedure|Procedure|false|false||treatmentnull|Primary malignant neoplasm|Disorder|false|false||malignancy
null|Malignant Neoplasms|Disorder|false|false||malignancynull|Rehabilitation Centers|Device|false|false||rehabilitation facilitynull|Rehabilitation Centers|Entity|false|false||rehabilitation facilitynull|Encounter due to care involving use of rehabilitation procedures|Finding|false|false||rehabilitation
null|Rehabilitation aspects|Finding|false|false||rehabilitationnull|Rehabilitation therapy|Procedure|false|false||rehabilitationnull|null|Title|false|false||rehabilitationnull|ADMIN.FACILITY|Finding|false|false||facilitynull|Facility (object)|Device|false|false||facilitynull|Help document|Finding|false|false||helpnull|Assisted (qualifier value)|Modifier|false|false||helpnull|REGAIN|Drug|false|false||regainnull|Strength (attribute)|Finding|false|false||strengthnull|Pharmaceutical Strength|LabModifier|false|false||strength
null|Physical Strength|LabModifier|false|false||strengthnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Anticipated|Finding|false|false||anticipatednull|Length of Stay|Time|false|false||length of staynull|Length|LabModifier|false|false||lengthnull|Less Than|LabModifier|false|false||LESS THANnull|Smaller|Modifier|false|false||LESSnull|Less Than|LabModifier|false|false||LESSnull|30 days|Time|false|false||30 DAYSnull|day|Time|false|false||DAYSnull|Fix|Phenomenon|false|false||attachednull|MEDICATION LIST|Finding|false|false||medication listnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|List|Finding|false|false||list
null|Sequence Data Type|Finding|false|false||listnull|Production Class Code - Pleasure|Finding|false|false||pleasure
null|pleasurable emotion|Finding|false|false||pleasurenull|Pleasure - Animals raised for recreation|Entity|false|false||pleasurenull|care of - AddressPartType|Finding|false|false||care ofnull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|NCK-Interacting Protein with SH3 Domain|Drug|false|false||wishnull|NCKIPSD wt Allele|Finding|false|false||wish
null|NCKIPSD gene|Finding|false|false||wishnull|Vitelliform Macular Dystrophy|Disorder|false|false||bestnull|BEST1 wt Allele|Finding|false|false||best
null|BEST1 gene|Finding|false|false||bestnull|best (quality)|Modifier|false|false||bestnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions