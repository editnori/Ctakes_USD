 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|26,30
No|31,33
:|33,34
_|37,38
_|38,39
_|39,40
<EOL>|40,41
<EOL>|42,43
Admission|43,52
Date|53,57
:|57,58
_|60,61
_|61,62
_|62,63
Discharge|77,86
Date|87,91
:|91,92
_|95,96
_|96,97
_|97,98
<EOL>|98,99
<EOL>|100,101
Date|101,105
of|106,108
Birth|109,114
:|114,115
_|117,118
_|118,119
_|119,120
Sex|133,136
:|136,137
F|140,141
<EOL>|141,142
<EOL>|143,144
Service|144,151
:|151,152
UROLOGY|153,160
<EOL>|160,161
<EOL>|162,163
Allergies|163,172
:|172,173
<EOL>|174,175
No|175,177
Known|178,183
Allergies|184,193
/|194,195
Adverse|196,203
Drug|204,208
Reactions|209,218
<EOL>|218,219
<EOL>|220,221
Attending|221,230
:|230,231
_|232,233
_|233,234
_|234,235
.|235,236
<EOL>|236,237
<EOL>|238,239
Chief|239,244
Complaint|245,254
:|254,255
<EOL>|255,256
Bladder|256,263
cancer|264,270
<EOL>|270,271
<EOL>|272,273
Major|273,278
Surgical|279,287
or|288,290
Invasive|291,299
Procedure|300,309
:|309,310
<EOL>|310,311
robotic|311,318
anterior|319,327
exenteration|328,340
and|341,344
open|345,349
ileal|350,355
conduit|356,363
<EOL>|363,364
<EOL>|364,365
<EOL>|366,367
History|367,374
of|375,377
Present|378,385
Illness|386,393
:|393,394
<EOL>|394,395
_|395,396
_|396,397
_|397,398
with|399,403
invasive|404,412
bladder|413,420
cancer|421,427
,|427,428
pelvic|429,435
MRI|436,439
concerning|440,450
for|451,454
<EOL>|455,456
invasion|456,464
into|465,469
anterior|470,478
vaginal|479,486
wall|487,491
,|491,492
now|493,496
s|497,498
/|498,499
p|499,500
robotic|501,508
anterior|509,517
<EOL>|518,519
exent|519,524
(|525,526
Dr|526,528
_|529,530
_|530,531
_|531,532
and|533,536
open|537,541
ileal|542,547
conduit|548,555
(|556,557
Dr|557,559
_|560,561
_|561,562
_|562,563
.|563,564
<EOL>|564,565
<EOL>|566,567
Past|567,571
Medical|572,579
History|580,587
:|587,588
<EOL>|588,589
Hypertension|589,601
,|601,602
laparoscopic|603,615
cholecystectomy|616,631
<EOL>|631,632
six|632,635
months|636,642
ago|643,646
,|646,647
left|648,652
knee|653,657
replacement|658,669
six|670,673
to|674,676
_|677,678
_|678,679
_|679,680
years|681,686
ago|687,690
,|690,691
<EOL>|691,692
laminectomy|692,703
of|704,706
L5|707,709
-|709,710
S1|710,712
at|713,715
age|716,719
_|720,721
_|721,722
_|722,723
,|723,724
two|725,728
vaginal|729,736
deliveries|737,747
.|747,748
<EOL>|748,749
<EOL>|749,750
<EOL>|751,752
Social|752,758
History|759,766
:|766,767
<EOL>|767,768
_|768,769
_|769,770
_|770,771
<EOL>|771,772
Family|772,778
History|779,786
:|786,787
<EOL>|787,788
Negative|788,796
for|797,800
bladder|801,808
CA|809,811
.|811,812
<EOL>|812,813
<EOL>|813,814
<EOL>|815,816
Physical|816,824
Exam|825,829
:|829,830
<EOL>|830,831
A|831,832
&|832,833
Ox3|833,836
<EOL>|836,837
Breathing|837,846
comfortably|847,858
on|859,861
RA|862,864
<EOL>|864,865
WWP|865,868
<EOL>|868,869
Abd|869,872
S|873,874
/|874,875
ND|875,877
/|877,878
appropriate|878,889
postsurgical|890,902
tenderness|903,913
to|914,916
palpation|917,926
<EOL>|926,927
Urostomy|927,935
pink|936,940
,|940,941
viable|942,948
<EOL>|948,949
<EOL>|950,951
Pertinent|951,960
Results|961,968
:|968,969
<EOL>|969,970
_|970,971
_|971,972
_|972,973
06|974,976
:|976,977
50AM|977,981
BLOOD|982,987
WBC|988,991
-|991,992
7.6|992,995
RBC|996,999
-|999,1000
3|1000,1001
.|1001,1002
41|1002,1004
*|1004,1005
Hgb|1006,1009
-|1009,1010
10|1010,1012
.|1012,1013
6|1013,1014
*|1014,1015
Hct|1016,1019
-|1019,1020
32|1020,1022
.|1022,1023
5|1023,1024
*|1024,1025
<EOL>|1026,1027
MCV|1027,1030
-|1030,1031
95|1031,1033
MCH|1034,1037
-|1037,1038
31.1|1038,1042
MCHC|1043,1047
-|1047,1048
32.6|1048,1052
RDW|1053,1056
-|1056,1057
14.4|1057,1061
RDWSD|1062,1067
-|1067,1068
50|1068,1070
.|1070,1071
2|1071,1072
*|1072,1073
Plt|1074,1077
_|1078,1079
_|1079,1080
_|1080,1081
<EOL>|1081,1082
_|1082,1083
_|1083,1084
_|1084,1085
06|1086,1088
:|1088,1089
50AM|1089,1093
BLOOD|1094,1099
Plt|1100,1103
_|1104,1105
_|1105,1106
_|1106,1107
<EOL>|1107,1108
_|1108,1109
_|1109,1110
_|1110,1111
06|1112,1114
:|1114,1115
45AM|1115,1119
BLOOD|1120,1125
Glucose|1126,1133
-|1133,1134
117|1134,1137
*|1137,1138
UreaN|1139,1144
-|1144,1145
23|1145,1147
*|1147,1148
Creat|1149,1154
-|1154,1155
0.6|1155,1158
Na|1159,1161
-|1161,1162
136|1162,1165
<EOL>|1166,1167
K|1167,1168
-|1168,1169
4.4|1169,1172
Cl|1173,1175
-|1175,1176
104|1176,1179
HCO3|1180,1184
-|1184,1185
23|1185,1187
AnGap|1188,1193
-|1193,1194
13|1194,1196
<EOL>|1196,1197
_|1197,1198
_|1198,1199
_|1199,1200
06|1201,1203
:|1203,1204
45AM|1204,1208
BLOOD|1209,1214
Calcium|1215,1222
-|1222,1223
7|1223,1224
.|1224,1225
9|1225,1226
*|1226,1227
Phos|1228,1232
-|1232,1233
3.4|1233,1236
Mg|1237,1239
-|1239,1240
2.0|1240,1243
<EOL>|1243,1244
<EOL>|1245,1246
Brief|1246,1251
Hospital|1252,1260
Course|1261,1267
:|1267,1268
<EOL>|1268,1269
Ms.|1269,1272
_|1273,1274
_|1274,1275
_|1275,1276
was|1277,1280
admitted|1281,1289
to|1290,1292
the|1293,1296
Urology|1297,1304
service|1305,1312
after|1313,1318
<EOL>|1319,1320
undergoing|1320,1330
[|1331,1332
robotic|1332,1339
anterior|1340,1348
exenteration|1349,1361
with|1362,1366
ileal|1367,1372
conduit|1373,1380
]|1380,1381
.|1381,1382
<EOL>|1383,1384
No|1384,1386
concerning|1387,1397
intrao|1398,1404
-|1404,1405
perative|1405,1413
events|1414,1420
occurred|1421,1429
;|1429,1430
please|1431,1437
see|1438,1441
<EOL>|1442,1443
dictated|1443,1451
operative|1452,1461
note|1462,1466
for|1467,1470
details|1471,1478
.|1478,1479
Patient|1480,1487
received|1488,1496
<EOL>|1497,1498
_|1498,1499
_|1499,1500
_|1500,1501
intravenous|1502,1513
antibiotic|1514,1524
prophylaxis|1525,1536
and|1537,1540
deep|1541,1545
vein|1546,1550
<EOL>|1551,1552
thrombosis|1552,1562
prophylaxis|1563,1574
with|1575,1579
subcutaneous|1580,1592
heparin|1593,1600
.|1600,1601
The|1602,1605
<EOL>|1606,1607
post-operative|1607,1621
course|1622,1628
was|1629,1632
notable|1633,1640
for|1641,1644
several|1645,1652
episodes|1653,1661
of|1662,1664
emesis|1665,1671
<EOL>|1672,1673
prompting|1673,1682
NGT|1683,1686
placement|1687,1696
on|1697,1699
_|1700,1701
_|1701,1702
_|1702,1703
.|1703,1704
Pt|1706,1708
self|1709,1713
removed|1714,1721
the|1722,1725
NGT|1726,1729
on|1730,1732
_|1733,1734
_|1734,1735
_|1735,1736
,|1736,1737
<EOL>|1738,1739
but|1739,1742
nausea|1743,1749
/|1749,1750
emesis|1750,1756
resolved|1757,1765
thereafter|1766,1776
and|1777,1780
pt|1781,1783
was|1784,1787
gradually|1788,1797
<EOL>|1798,1799
advanced|1799,1807
to|1808,1810
a|1811,1812
regular|1813,1820
diet|1821,1825
with|1826,1830
passage|1831,1838
of|1839,1841
flatus|1842,1848
without|1849,1856
issue|1857,1862
.|1862,1863
<EOL>|1864,1865
With|1866,1870
advacement|1871,1881
of|1882,1884
diet|1885,1889
,|1889,1890
patient|1891,1898
was|1899,1902
transitioned|1903,1915
from|1916,1920
IV|1921,1923
pain|1924,1928
<EOL>|1929,1930
medication|1930,1940
to|1941,1943
oral|1944,1948
pain|1949,1953
medications|1954,1965
.|1965,1966
The|1967,1970
ostomy|1971,1977
nurse|1978,1983
<EOL>|1983,1984
saw|1984,1987
the|1988,1991
patient|1992,1999
for|2000,2003
ostomy|2004,2010
teaching|2011,2019
.|2019,2020
At|2021,2023
the|2024,2027
time|2028,2032
of|2033,2035
discharge|2036,2045
<EOL>|2046,2047
the|2047,2050
wound|2051,2056
was|2057,2060
healing|2061,2068
well|2069,2073
with|2074,2078
no|2079,2081
evidence|2082,2090
of|2091,2093
erythema|2094,2102
,|2102,2103
<EOL>|2104,2105
swelling|2105,2113
,|2113,2114
or|2115,2117
purulent|2118,2126
drainage|2127,2135
.|2135,2136
Her|2137,2140
drain|2141,2146
was|2147,2150
removed|2151,2158
.|2158,2159
The|2160,2163
<EOL>|2164,2165
ostomy|2165,2171
was|2172,2175
perfused|2176,2184
and|2185,2188
patent|2189,2195
,|2195,2196
and|2197,2200
one|2201,2204
ureteral|2205,2213
stent|2214,2219
had|2220,2223
<EOL>|2224,2225
fallen|2225,2231
out|2232,2235
spontaneously|2236,2249
.|2249,2250
_|2252,2253
_|2253,2254
_|2254,2255
was|2256,2259
consulted|2260,2269
and|2270,2273
recommended|2274,2285
<EOL>|2286,2287
disposition|2287,2298
to|2299,2301
rehab|2302,2307
.|2307,2308
Post-operative|2310,2324
follow|2325,2331
up|2332,2334
appointments|2335,2347
<EOL>|2348,2349
were|2349,2353
arranged|2354,2362
/|2362,2363
discussed|2363,2372
and|2373,2376
the|2377,2380
patient|2381,2388
was|2389,2392
discharged|2393,2403
to|2404,2406
rehab|2407,2412
<EOL>|2413,2414
for|2414,2417
further|2418,2425
recovery|2426,2434
.|2434,2435
<EOL>|2435,2436
<EOL>|2436,2437
<EOL>|2438,2439
Medications|2439,2450
on|2451,2453
Admission|2454,2463
:|2463,2464
<EOL>|2464,2465
The|2465,2468
Preadmission|2469,2481
Medication|2482,2492
list|2493,2497
is|2498,2500
accurate|2501,2509
and|2510,2513
complete|2514,2522
.|2522,2523
<EOL>|2523,2524
1.|2524,2526
Heparin|2527,2534
5000|2535,2539
UNIT|2540,2544
SC|2545,2547
ONCE|2548,2552
<EOL>|2553,2554
Start|2554,2559
:|2559,2560
in|2561,2563
O.R.|2564,2568
Holding|2569,2576
Area|2577,2581
<EOL>|2582,2583
2.|2583,2585
Losartan|2586,2594
Potassium|2595,2604
50|2605,2607
mg|2608,2610
PO|2611,2613
DAILY|2614,2619
<EOL>|2620,2621
3.|2621,2623
Atorvastatin|2624,2636
10|2637,2639
mg|2640,2642
PO|2643,2645
QPM|2646,2649
<EOL>|2650,2651
4.|2651,2653
Levothyroxine|2654,2667
Sodium|2668,2674
175|2675,2678
mcg|2679,2682
PO|2683,2685
DAILY|2686,2691
<EOL>|2692,2693
<EOL>|2693,2694
<EOL>|2695,2696
Discharge|2696,2705
Medications|2706,2717
:|2717,2718
<EOL>|2718,2719
1.|2719,2721
Acetaminophen|2723,2736
650|2737,2740
mg|2741,2743
PO|2744,2746
Q6H|2747,2750
<EOL>|2752,2753
2.|2753,2755
Docusate|2757,2765
Sodium|2766,2772
100|2773,2776
mg|2777,2779
PO|2780,2782
BID|2783,2786
<EOL>|2787,2788
take|2788,2792
while|2793,2798
taking|2799,2805
narcotic|2806,2814
pain|2815,2819
meds|2820,2824
<EOL>|2825,2826
RX|2826,2828
*|2829,2830
docusate|2830,2838
sodium|2839,2845
[|2846,2847
Colace|2847,2853
]|2853,2854
100|2855,2858
mg|2859,2861
1|2862,2863
capsule|2864,2871
(|2871,2872
s|2872,2873
)|2873,2874
by|2875,2877
mouth|2878,2883
twice|2884,2889
<EOL>|2890,2891
a|2891,2892
day|2893,2896
Disp|2897,2901
#|2902,2903
*|2903,2904
50|2904,2906
Capsule|2907,2914
Refills|2915,2922
:|2922,2923
*|2923,2924
0|2924,2925
<EOL>|2926,2927
3.|2927,2929
Enoxaparin|2931,2941
Sodium|2942,2948
40|2949,2951
mg|2952,2954
SC|2955,2957
DAILY|2958,2963
<EOL>|2964,2965
Start|2965,2970
:|2970,2971
_|2972,2973
_|2973,2974
_|2974,2975
,|2975,2976
First|2977,2982
Dose|2983,2987
:|2987,2988
Next|2989,2993
Routine|2994,3001
Administration|3002,3016
Time|3017,3021
<EOL>|3022,3023
RX|3023,3025
*|3026,3027
enoxaparin|3027,3037
40|3038,3040
mg|3041,3043
/|3043,3044
0.4|3044,3047
mL|3048,3050
40|3051,3053
mg|3054,3056
sc|3057,3059
daily|3060,3065
Disp|3066,3070
#|3071,3072
*|3072,3073
28|3073,3075
Syringe|3076,3083
<EOL>|3084,3085
Refills|3085,3092
:|3092,3093
*|3093,3094
0|3094,3095
<EOL>|3096,3097
4.|3097,3099
Nitrofurantoin|3101,3115
Monohyd|3116,3123
(|3124,3125
MacroBID|3125,3133
)|3133,3134
100|3135,3138
mg|3139,3141
PO|3142,3144
DAILY|3145,3150
<EOL>|3151,3152
take|3152,3156
while|3157,3162
ureteral|3163,3171
stents|3172,3178
are|3179,3182
in|3183,3185
place|3186,3191
<EOL>|3192,3193
RX|3193,3195
*|3196,3197
nitrofurantoin|3197,3211
monohyd|3212,3219
/|3219,3220
m|3220,3221
-|3221,3222
cryst|3222,3227
[|3228,3229
Macrobid|3229,3237
]|3237,3238
100|3239,3242
mg|3243,3245
1|3246,3247
<EOL>|3248,3249
capsule|3249,3256
(|3256,3257
s|3257,3258
)|3258,3259
by|3260,3262
mouth|3263,3268
daily|3269,3274
Disp|3275,3279
#|3280,3281
*|3281,3282
14|3282,3284
Capsule|3285,3292
Refills|3293,3300
:|3300,3301
*|3301,3302
0|3302,3303
<EOL>|3304,3305
5.|3305,3307
OxyCODONE|3309,3318
(|3319,3320
Immediate|3320,3329
Release|3330,3337
)|3337,3338
5|3339,3340
mg|3341,3343
PO|3344,3346
Q4H|3347,3350
:|3350,3351
PRN|3351,3354
Pain|3355,3359
-|3360,3361
<EOL>|3362,3363
Moderate|3363,3371
<EOL>|3372,3373
RX|3373,3375
*|3376,3377
oxycodone|3377,3386
5|3387,3388
mg|3389,3391
1|3392,3393
tablet|3394,3400
(|3400,3401
s|3401,3402
)|3402,3403
by|3404,3406
mouth|3407,3412
q4h|3413,3416
prn|3417,3420
Disp|3421,3425
#|3426,3427
*|3427,3428
30|3428,3430
Tablet|3431,3437
<EOL>|3438,3439
Refills|3439,3446
:|3446,3447
*|3447,3448
0|3448,3449
<EOL>|3450,3451
6.|3451,3453
Atorvastatin|3455,3467
10|3468,3470
mg|3471,3473
PO|3474,3476
QPM|3477,3480
<EOL>|3482,3483
7.|3483,3485
Levothyroxine|3487,3500
Sodium|3501,3507
175|3508,3511
mcg|3512,3515
PO|3516,3518
DAILY|3519,3524
<EOL>|3526,3527
8.|3527,3529
Losartan|3531,3539
Potassium|3540,3549
50|3550,3552
mg|3553,3555
PO|3556,3558
DAILY|3559,3564
<EOL>|3566,3567
<EOL>|3567,3568
<EOL>|3569,3570
Discharge|3570,3579
Disposition|3580,3591
:|3591,3592
<EOL>|3592,3593
Extended|3593,3601
Care|3602,3606
<EOL>|3606,3607
<EOL>|3608,3609
Facility|3609,3617
:|3617,3618
<EOL>|3618,3619
_|3619,3620
_|3620,3621
_|3621,3622
<EOL>|3622,3623
<EOL>|3624,3625
Discharge|3625,3634
Diagnosis|3635,3644
:|3644,3645
<EOL>|3645,3646
Bladder|3646,3653
cancer|3654,3660
<EOL>|3660,3661
<EOL>|3661,3662
<EOL>|3663,3664
Discharge|3664,3673
Condition|3674,3683
:|3683,3684
<EOL>|3684,3685
WdWn|3685,3689
,|3689,3690
NAD|3691,3694
,|3694,3695
AVSS|3696,3700
<EOL>|3700,3701
Abdomen|3701,3708
soft|3709,3713
,|3713,3714
appropriately|3715,3728
tender|3729,3735
along|3736,3741
incision|3742,3750
<EOL>|3750,3751
Incision|3751,3759
is|3760,3762
c|3763,3764
/|3764,3765
d|3765,3766
/|3766,3767
I|3767,3768
(|3769,3770
steris|3770,3776
)|3776,3777
<EOL>|3777,3778
Stoma|3778,3783
is|3784,3786
well|3787,3791
perfused|3792,3800
;|3800,3801
Urine|3802,3807
color|3808,3813
is|3814,3816
yellow|3817,3823
<EOL>|3823,3824
Ureteral|3824,3832
stent|3833,3838
noted|3839,3844
via|3845,3848
stoma|3849,3854
<EOL>|3854,3855
JP|3855,3857
drain|3858,3863
has|3864,3867
been|3868,3872
removed|3873,3880
<EOL>|3880,3881
Bilateral|3881,3890
lower|3891,3896
extremities|3897,3908
are|3909,3912
warm|3913,3917
,|3917,3918
dry|3919,3922
,|3922,3923
well|3924,3928
perfused|3929,3937
.|3937,3938
There|3940,3945
<EOL>|3946,3947
is|3947,3949
no|3950,3952
reported|3953,3961
calf|3962,3966
pain|3967,3971
to|3972,3974
deep|3975,3979
palpation|3980,3989
.|3989,3990
No|3991,3993
edema|3994,3999
or|4000,4002
pitting|4003,4010
<EOL>|4010,4011
<EOL>|4011,4012
<EOL>|4013,4014
Discharge|4014,4023
Instructions|4024,4036
:|4036,4037
<EOL>|4037,4038
-|4038,4039
Please|4039,4045
also|4046,4050
refer|4051,4056
to|4057,4059
the|4060,4063
handout|4064,4071
of|4072,4074
instructions|4075,4087
provided|4088,4096
to|4097,4099
<EOL>|4100,4101
you|4101,4104
by|4105,4107
your|4108,4112
Urologist|4113,4122
<EOL>|4122,4123
-|4123,4124
Please|4124,4130
also|4131,4135
refer|4136,4141
to|4142,4144
the|4145,4148
instructions|4149,4161
provided|4162,4170
to|4171,4173
you|4174,4177
by|4178,4180
the|4181,4184
<EOL>|4185,4186
Ostomy|4186,4192
nurse|4193,4198
specialist|4199,4209
that|4210,4214
details|4215,4222
the|4223,4226
required|4227,4235
care|4236,4240
and|4241,4244
<EOL>|4245,4246
management|4246,4256
of|4257,4259
your|4260,4264
Urostomy|4265,4273
<EOL>|4273,4274
-|4274,4275
You|4275,4278
will|4279,4283
be|4284,4286
sent|4287,4291
home|4292,4296
with|4297,4301
Visiting|4302,4310
Nurse|4311,4316
_|4317,4318
_|4318,4319
_|4319,4320
<EOL>|4321,4322
services|4322,4330
to|4331,4333
facilitate|4334,4344
your|4345,4349
transition|4350,4360
to|4361,4363
home|4364,4368
care|4369,4373
of|4374,4376
your|4377,4381
<EOL>|4382,4383
urostomy|4383,4391
<EOL>|4391,4392
-|4392,4393
Resume|4393,4399
your|4400,4404
pre-admission|4405,4418
/|4418,4419
home|4419,4423
medications|4424,4435
except|4436,4442
as|4443,4445
noted|4446,4451
.|4451,4452
<EOL>|4453,4454
Always|4454,4460
call|4461,4465
to|4466,4468
inform|4469,4475
,|4475,4476
review|4477,4483
and|4484,4487
discuss|4488,4495
any|4496,4499
medication|4500,4510
changes|4511,4518
<EOL>|4519,4520
and|4520,4523
your|4524,4528
post-operative|4529,4543
course|4544,4550
with|4551,4555
your|4556,4560
primary|4561,4568
care|4569,4573
doctor|4574,4580
<EOL>|4580,4581
-|4581,4582
_|4582,4583
_|4583,4584
_|4584,4585
you|4586,4589
have|4590,4594
been|4595,4599
prescribed|4600,4610
IBUPROFEN|4611,4620
,|4620,4621
please|4622,4628
note|4629,4633
that|4634,4638
you|4639,4642
may|4643,4646
<EOL>|4647,4648
take|4648,4652
this|4653,4657
in|4658,4660
addition|4661,4669
to|4670,4672
the|4673,4676
prescribed|4677,4687
NARCOTIC|4688,4696
pain|4697,4701
<EOL>|4702,4703
medications|4703,4714
and|4715,4718
/|4718,4719
or|4719,4721
tylenol|4722,4729
.|4729,4730
FIRST|4731,4736
,|4736,4737
alternate|4738,4747
Tylenol|4748,4755
<EOL>|4756,4757
(|4757,4758
acetaminophen|4758,4771
)|4771,4772
and|4773,4776
Ibuprofen|4777,4786
for|4787,4790
pain|4791,4795
control|4796,4803
.|4803,4804
<EOL>|4804,4805
-|4805,4806
REPLACE|4806,4813
the|4814,4817
Tylenol|4818,4825
with|4826,4830
the|4831,4834
prescribed|4835,4845
narcotic|4846,4854
if|4855,4857
the|4858,4861
<EOL>|4862,4863
narcotic|4863,4871
is|4872,4874
combined|4875,4883
with|4884,4888
Tylenol|4889,4896
(|4897,4898
examples|4898,4906
include|4907,4914
brand|4915,4920
names|4921,4926
<EOL>|4927,4928
_|4928,4929
_|4929,4930
_|4930,4931
,|4931,4932
Tylenol|4933,4940
#|4941,4942
3|4942,4943
w|4944,4945
/|4945,4946
codeine|4947,4954
and|4955,4958
their|4959,4964
generic|4965,4972
<EOL>|4973,4974
equivalents|4974,4985
)|4985,4986
.|4986,4987
ALWAYS|4988,4994
discuss|4995,5002
your|5003,5007
medications|5008,5019
(|5020,5021
especially|5021,5031
when|5032,5036
<EOL>|5037,5038
using|5038,5043
narcotics|5044,5053
or|5054,5056
new|5057,5060
medications|5061,5072
)|5072,5073
use|5074,5077
with|5078,5082
the|5083,5086
pharmacist|5087,5097
when|5098,5102
<EOL>|5103,5104
you|5104,5107
first|5108,5113
retrieve|5114,5122
your|5123,5127
prescription|5128,5140
if|5141,5143
you|5144,5147
have|5148,5152
any|5153,5156
questions|5157,5166
.|5166,5167
<EOL>|5168,5169
Use|5169,5172
the|5173,5176
narcotic|5177,5185
pain|5186,5190
medication|5191,5201
for|5202,5205
break|5206,5211
-|5211,5212
through|5212,5219
pain|5220,5224
that|5225,5229
is|5230,5232
<EOL>|5233,5234
>|5234,5235
4|5235,5236
on|5237,5239
the|5240,5243
pain|5244,5248
scale|5249,5254
.|5254,5255
<EOL>|5255,5256
-|5256,5257
The|5257,5260
MAXIMUM|5261,5268
dose|5269,5273
of|5274,5276
Tylenol|5277,5284
(|5285,5286
ACETAMINOPHEN|5286,5299
)|5299,5300
is|5301,5303
4|5304,5305
grams|5306,5311
(|5312,5313
from|5313,5317
<EOL>|5318,5319
ALL|5319,5322
sources|5323,5330
)|5330,5331
PER|5332,5335
DAY|5336,5339
and|5340,5343
remember|5344,5352
that|5353,5357
the|5358,5361
prescribed|5362,5372
narcotic|5373,5381
<EOL>|5382,5383
pain|5383,5387
medication|5388,5398
may|5399,5402
also|5403,5407
contain|5408,5415
Tylenol|5416,5423
(|5424,5425
acetaminophen|5425,5438
)|5438,5439
so|5440,5442
this|5443,5447
<EOL>|5448,5449
needs|5449,5454
to|5455,5457
be|5458,5460
considered|5461,5471
when|5472,5476
monitoring|5477,5487
your|5488,5492
daily|5493,5498
dose|5499,5503
and|5504,5507
<EOL>|5508,5509
maximum|5509,5516
.|5516,5517
<EOL>|5517,5518
-|5518,5519
If|5519,5521
you|5522,5525
are|5526,5529
taking|5530,5536
Ibuprofen|5537,5546
(|5547,5548
Brand|5548,5553
names|5554,5559
include|5560,5567
_|5568,5569
_|5569,5570
_|5570,5571
<EOL>|5572,5573
this|5573,5577
should|5578,5584
always|5585,5591
be|5592,5594
taken|5595,5600
with|5601,5605
food|5606,5610
.|5610,5611
If|5612,5614
you|5615,5618
develop|5619,5626
stomach|5627,5634
<EOL>|5635,5636
pain|5636,5640
or|5641,5643
note|5644,5648
black|5649,5654
stool|5655,5660
,|5660,5661
stop|5662,5666
the|5667,5670
Ibuprofen|5671,5680
.|5680,5681
<EOL>|5681,5682
-|5682,5683
Please|5683,5689
do|5690,5692
NOT|5693,5696
drive|5697,5702
,|5702,5703
operate|5704,5711
dangerous|5712,5721
machinery|5722,5731
,|5731,5732
or|5733,5735
consume|5736,5743
<EOL>|5744,5745
alcohol|5745,5752
while|5753,5758
taking|5759,5765
narcotic|5766,5774
pain|5775,5779
medications|5780,5791
.|5791,5792
<EOL>|5792,5793
-|5793,5794
Do|5794,5796
NOT|5797,5800
drive|5801,5806
and|5807,5810
until|5811,5816
you|5817,5820
are|5821,5824
cleared|5825,5832
to|5833,5835
resume|5836,5842
such|5843,5847
<EOL>|5848,5849
activities|5849,5859
by|5860,5862
your|5863,5867
PCP|5868,5871
or|5872,5874
urologist|5875,5884
.|5884,5885
You|5886,5889
may|5890,5893
be|5894,5896
a|5897,5898
passenger|5899,5908
<EOL>|5908,5909
-|5909,5910
Colace|5910,5916
may|5917,5920
have|5921,5925
been|5926,5930
prescribed|5931,5941
to|5942,5944
avoid|5945,5950
post|5951,5955
surgical|5956,5964
<EOL>|5965,5966
constipation|5966,5978
and|5979,5982
constipation|5983,5995
related|5996,6003
to|6004,6006
narcotic|6007,6015
pain|6016,6020
<EOL>|6021,6022
medication|6022,6032
.|6032,6033
Discontinue|6034,6045
if|6046,6048
loose|6049,6054
stool|6055,6060
or|6061,6063
diarrhea|6064,6072
develops|6073,6081
.|6081,6082
<EOL>|6083,6084
Colace|6084,6090
is|6091,6093
a|6094,6095
stool|6096,6101
-|6101,6102
softener|6102,6110
,|6110,6111
NOT|6112,6115
a|6116,6117
laxative|6118,6126
.|6126,6127
<EOL>|6127,6128
-|6128,6129
You|6129,6132
may|6133,6136
shower|6137,6143
2|6144,6145
days|6146,6150
after|6151,6156
surgery|6157,6164
,|6164,6165
but|6166,6169
do|6170,6172
not|6173,6176
tub|6177,6180
bathe|6181,6186
,|6186,6187
<EOL>|6188,6189
swim|6189,6193
,|6193,6194
soak|6195,6199
,|6199,6200
or|6201,6203
scrub|6204,6209
incision|6210,6218
for|6219,6222
2|6223,6224
weeks|6225,6230
<EOL>|6230,6231
-|6231,6232
If|6232,6234
you|6235,6238
had|6239,6242
a|6243,6244
drain|6245,6250
or|6251,6253
skin|6254,6258
clips|6259,6264
(|6265,6266
staples|6266,6273
)|6273,6274
removed|6275,6282
from|6283,6287
your|6288,6292
<EOL>|6293,6294
abdomen|6294,6301
;|6301,6302
bandage|6303,6310
strips|6311,6317
called|6318,6324
|6325,6326
steristrips|6326,6337
|6337,6338
have|6339,6343
been|6344,6348
applied|6349,6356
<EOL>|6357,6358
to|6358,6360
close|6361,6366
the|6367,6370
wound|6371,6376
OR|6377,6379
the|6380,6383
site|6384,6388
was|6389,6392
covered|6393,6400
with|6401,6405
a|6406,6407
gauze|6408,6413
<EOL>|6414,6415
dressing|6415,6423
.|6423,6424
Allow|6425,6430
any|6431,6434
steristrips|6435,6446
/|6446,6447
bandage|6447,6454
strips|6455,6461
to|6462,6464
fall|6465,6469
off|6470,6473
on|6474,6476
<EOL>|6477,6478
their|6478,6483
own|6484,6487
_|6488,6489
_|6489,6490
_|6490,6491
days|6492,6496
)|6496,6497
.|6497,6498
PLEASE|6499,6505
REMOVE|6506,6512
any|6513,6516
"|6517,6518
gauze|6518,6523
"|6523,6524
dressings|6525,6534
within|6535,6541
<EOL>|6542,6543
two|6543,6546
days|6547,6551
of|6552,6554
discharge|6555,6564
.|6564,6565
Steristrips|6566,6577
may|6578,6581
get|6582,6585
wet|6586,6589
.|6589,6590
<EOL>|6590,6591
-|6591,6592
No|6592,6594
heavy|6595,6600
lifting|6601,6608
for|6609,6612
4|6613,6614
weeks|6615,6620
(|6621,6622
no|6622,6624
more|6625,6629
than|6630,6634
10|6635,6637
pounds|6638,6644
)|6644,6645
.|6645,6646
Do|6647,6649
"|6650,6651
not|6651,6654
"|6654,6655
<EOL>|6656,6657
be|6657,6659
sedentary|6660,6669
.|6669,6670
Walk|6671,6675
frequently|6676,6686
.|6686,6687
Light|6688,6693
household|6694,6703
chores|6704,6710
(|6711,6712
cooking|6712,6719
,|6719,6720
<EOL>|6721,6722
folding|6722,6729
laundry|6730,6737
,|6737,6738
washing|6739,6746
dishes|6747,6753
)|6753,6754
are|6755,6758
generally|6759,6768
|6769,6770
ok|6770,6772
|6772,6773
but|6774,6777
AGAIN|6778,6783
,|6783,6784
<EOL>|6785,6786
avoid|6786,6791
straining|6792,6801
,|6801,6802
pulling|6803,6810
,|6810,6811
twisting|6812,6820
(|6821,6822
do|6822,6824
NOT|6825,6828
vacuum|6829,6835
)|6835,6836
.|6836,6837
<EOL>|6837,6838
<EOL>|6838,6839
<EOL>|6840,6841
Followup|6841,6849
Instructions|6850,6862
:|6862,6863
<EOL>|6863,6864
_|6864,6865
_|6865,6866
_|6866,6867
<EOL>|6867,6868

