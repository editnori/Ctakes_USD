 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Procedure|Health Care Activity|SIMPLE_SEGMENT|43,52|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|43,57|false|false|false|C2598112||Admission Date
Finding|Body Substance|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|77,86|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|77,91|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|133,136|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|144,151|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|144,151|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|153,161|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|Allergies|185,194|false|false|false|C1717415||Allergies
Finding|Pathologic Function|Allergies|185,194|false|false|false|C0020517|Hypersensitivity|Allergies
Finding|Pathologic Function|Allergies|197,219|true|false|false|C0041755|Adverse reaction to drug|Adverse Drug Reactions
Drug|Pharmacologic Substance|Allergies|205,209|false|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|Drug
Finding|Finding|Allergies|205,209|false|false|false|C0740721|Drug problem|Drug
Finding|Pathologic Function|Allergies|205,219|true|false|false|C0041755|Adverse reaction to drug|Drug Reactions
Finding|Functional Concept|Allergies|222,231|false|false|false|C1999232|Attending (action)|Attending
Attribute|Clinical Attribute|Chief Complaint|257,276|false|false|false|C2707305||Shortness of breath
Finding|Sign or Symptom|Chief Complaint|257,276|false|false|false|C0013404|Dyspnea|Shortness of breath
Finding|Body Substance|Chief Complaint|270,276|false|false|false|C0225386|Breath|breath
Finding|Mental Process|Chief Complaint|286,292|false|false|false|C0229992|Psyche structure|mental
Attribute|Clinical Attribute|Chief Complaint|286,299|false|false|false|C0488568;C0488569||mental status
Finding|Finding|Chief Complaint|286,299|false|false|false|C0278060|Mental state|mental status
Attribute|Clinical Attribute|Chief Complaint|293,299|false|false|false|C5889824||status
Finding|Idea or Concept|Chief Complaint|293,299|false|false|false|C1546481|What subject filter - Status|status
Finding|Classification|Chief Complaint|302,307|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|308,316|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|308,316|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|320,338|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|329,338|false|false|false|C0945766||Procedure
Event|Occupational Activity|Chief Complaint|329,338|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|329,338|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|329,338|false|false|false|C0184661|Interventional procedure|Procedure
Finding|Body Substance|History of Present Illness|376,383|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|376,383|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|376,383|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|394,398|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|History of Present Illness|394,398|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Body Substance|History of Present Illness|403,410|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|403,410|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|403,410|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Conceptual Entity|History of Present Illness|416,423|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|416,423|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|History of Present Illness|416,423|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|416,426|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|History of Present Illness|427,436|false|false|false|C1527336|Sjogren's Syndrome|Sjogren's
Disorder|Disease or Syndrome|History of Present Illness|438,446|false|false|false|C0039082|Syndrome|syndrome
Finding|Finding|History of Present Illness|448,456|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|History of Present Illness|448,456|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Finding|History of Present Illness|461,483|false|false|false|C0745043|History of recent hospitalization|recent hospitalization
Procedure|Health Care Activity|History of Present Illness|468,483|false|false|false|C0019993|Hospitalization|hospitalization
Disorder|Disease or Syndrome|History of Present Illness|488,494|false|false|false|C0036690;C0243026|Sepsis;Septicemia|sepsis
Disorder|Neoplastic Process|History of Present Illness|496,505|false|false|false|C0027627|Neoplasm Metastasis|secondary
Finding|Functional Concept|History of Present Illness|496,505|false|false|false|C1522484|metastatic qualifier|secondary
Disorder|Disease or Syndrome|History of Present Illness|517,524|false|true|false|C0009319|Colitis|colitis
Attribute|Clinical Attribute|History of Present Illness|553,564|false|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|History of Present Illness|553,564|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|History of Present Illness|553,564|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|History of Present Illness|553,564|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Disorder|Disease or Syndrome|History of Present Illness|553,572|false|false|false|C1145670|Respiratory Failure|respiratory failure
Finding|Functional Concept|History of Present Illness|565,572|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|History of Present Illness|565,572|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|History of Present Illness|565,572|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|583,593|false|false|false|C0021925|Intubation (procedure)|intubation
Finding|Finding|History of Present Illness|638,645|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|History of Present Illness|638,645|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Idea or Concept|History of Present Illness|654,657|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|History of Present Illness|654,657|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Body Substance|History of Present Illness|660,667|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|660,667|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|660,667|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Procedure|Health Care Activity|History of Present Illness|719,734|false|false|false|C0019993|Hospitalization|hospitalization
Disorder|Disease or Syndrome|History of Present Illness|748,755|false|true|false|C0009319|Colitis|colitis
Finding|Body Substance|History of Present Illness|758,765|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|758,765|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|758,765|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Gene or Genome|History of Present Illness|770,773|false|false|false|C1412045|A1BG gene|ABG
Procedure|Laboratory Procedure|History of Present Illness|770,773|false|false|false|C0150411|Analysis of arterial blood gases and pH|ABG
Finding|Functional Concept|History of Present Illness|815,823|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|History of Present Illness|815,823|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|History of Present Illness|815,823|false|false|false|C4706767|Transfer (immobility management)|transfer
Finding|Finding|History of Present Illness|860,887|false|false|false|C4718286|Reports shortness of breath|reports shortness of breath
Attribute|Clinical Attribute|History of Present Illness|868,887|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|History of Present Illness|868,887|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|History of Present Illness|881,887|false|false|false|C0225386|Breath|breath
Drug|Organic Chemical|History of Present Illness|908,913|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|History of Present Illness|908,913|false|false|false|C3815497|Cough (guaifenesin)|cough
Finding|Sign or Symptom|History of Present Illness|908,913|false|false|false|C0010200|Coughing|cough
Anatomy|Body Location or Region|History of Present Illness|927,932|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|927,932|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|History of Present Illness|927,937|true|false|false|C2926613||chest pain
Finding|Sign or Symptom|History of Present Illness|927,937|true|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|History of Present Illness|933,937|true|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|933,937|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|933,937|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|History of Present Illness|950,956|true|false|false|C4255480||nausea
Finding|Sign or Symptom|History of Present Illness|950,956|true|false|false|C0027497|Nausea|nausea
Finding|Finding|History of Present Illness|950,968|true|false|false|C3843946|Nausea or vomiting|nausea or vomiting
Finding|Sign or Symptom|History of Present Illness|960,968|true|false|false|C0042963|Vomiting|vomiting
Anatomy|Body Location or Region|History of Present Illness|982,991|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|History of Present Illness|982,996|false|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|History of Present Illness|992,996|false|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|992,996|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|992,996|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Idea or Concept|History of Present Illness|1010,1017|false|false|false|C1555582|Initial (abbreviation)|initial
Finding|Functional Concept|History of Present Illness|1061,1065|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|History of Present Illness|1061,1065|false|false|false|C0582103|Medical Examination|Exam
Finding|Finding|History of Present Illness|1082,1091|false|false|false|C0231835|Tachypnea|tachypnea
Attribute|Clinical Attribute|History of Present Illness|1097,1108|false|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|History of Present Illness|1097,1108|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|History of Present Illness|1097,1108|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|History of Present Illness|1097,1108|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Attribute|Clinical Attribute|History of Present Illness|1097,1114|false|false|false|C0231832|Respiratory rate|respiratory rates
Disorder|Disease or Syndrome|History of Present Illness|1142,1147|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|History of Present Illness|1142,1147|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Finding|History of Present Illness|1142,1156|false|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|blood pressure
Finding|Organism Function|History of Present Illness|1142,1156|false|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|blood pressure
Procedure|Health Care Activity|History of Present Illness|1142,1156|false|false|false|C0005824|Blood pressure determination|blood pressure
Finding|Finding|History of Present Illness|1148,1156|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|History of Present Illness|1148,1156|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|History of Present Illness|1148,1156|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|History of Present Illness|1148,1156|false|false|false|C0033095||pressure
Finding|Finding|History of Present Illness|1176,1184|false|false|false|C0184511;C1561611;C4084203|Admission Level of Care Code - Improved;Improved;Improved - answer to question|improved
Finding|Intellectual Product|History of Present Illness|1176,1184|false|false|false|C0184511;C1561611;C4084203|Admission Level of Care Code - Improved;Improved;Improved - answer to question|improved
Finding|Finding|History of Present Illness|1194,1197|false|false|false|C5939094|Own|own
Finding|Finding|History of Present Illness|1209,1218|false|false|false|C0231835|Tachypnea|tachypnea
Drug|Organic Chemical|History of Present Illness|1220,1225|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|History of Present Illness|1220,1225|false|false|false|C3815497|Cough (guaifenesin)|cough
Finding|Sign or Symptom|History of Present Illness|1220,1225|false|false|false|C0010200|Coughing|cough
Finding|Finding|History of Present Illness|1231,1238|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|History of Present Illness|1231,1238|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Idea or Concept|History of Present Illness|1251,1258|false|false|false|C2699424|Concern|concern
Disorder|Disease or Syndrome|History of Present Illness|1263,1272|false|false|false|C0032285|Pneumonia|pneumonia
Finding|Body Substance|History of Present Illness|1275,1282|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|1275,1282|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|1275,1282|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1292,1302|false|false|false|C0042313|vancomycin|vancomycin
Drug|Antibiotic|History of Present Illness|1292,1302|false|false|false|C0042313|vancomycin|vancomycin
Procedure|Laboratory Procedure|History of Present Illness|1292,1302|false|false|false|C0489941|Vancomycin measurement|vancomycin
Drug|Antibiotic|History of Present Illness|1308,1320|false|false|false|C0282386|levofloxacin|levofloxacin
Drug|Organic Chemical|History of Present Illness|1308,1320|false|false|false|C0282386|levofloxacin|levofloxacin
Procedure|Diagnostic Procedure|History of Present Illness|1323,1326|false|false|false|C0039985|Plain chest X-ray|CXR
Procedure|Diagnostic Procedure|History of Present Illness|1362,1365|false|false|false|C0039985|Plain chest X-ray|CXR
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1392,1397|false|false|false|C1956423|Biphasic Continuous Positive Airway Pressure|BIPAP
Finding|Body Substance|History of Present Illness|1400,1407|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|1400,1407|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|1400,1407|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1418,1421|false|false|false|C3813556|Cancer/Testis Antigen|CTA
Finding|Gene or Genome|History of Present Illness|1418,1421|false|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|History of Present Illness|1418,1421|false|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Procedure|Health Care Activity|History of Present Illness|1425,1433|false|false|false|C0220825|Evaluation|evaluate
Finding|Functional Concept|History of Present Illness|1467,1475|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|History of Present Illness|1467,1475|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|History of Present Illness|1467,1475|false|false|false|C4706767|Transfer (immobility management)|transfer
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1522,1527|false|false|false|C1956423|Biphasic Continuous Positive Airway Pressure|BIPAP
Event|Activity|History of Present Illness|1536,1543|false|false|false|C1706079||arrival
Finding|Functional Concept|History of Present Illness|1536,1543|false|false|false|C1555577|arrival - ActRelationshipType|arrival
Finding|Body Substance|History of Present Illness|1557,1564|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|1557,1564|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|1557,1564|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1576,1581|false|false|false|C1956423|Biphasic Continuous Positive Airway Pressure|BiPAP
Finding|Functional Concept|History of Present Illness|1633,1645|false|false|false|C2348609|Supplement|supplemental
Finding|Finding|History of Present Illness|1633,1652|false|false|false|C4534306|Supplemental oxygen|supplemental oxygen
Drug|Biologically Active Substance|History of Present Illness|1646,1652|false|false|false|C0030054|oxygen|oxygen
Drug|Element, Ion, or Isotope|History of Present Illness|1646,1652|false|false|false|C0030054|oxygen|oxygen
Drug|Pharmacologic Substance|History of Present Illness|1646,1652|false|false|false|C0030054|oxygen|oxygen
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1646,1652|false|false|false|C0184633|Oxygen Therapy Care|oxygen
Attribute|Clinical Attribute|History of Present Illness|1667,1671|true|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|1667,1671|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1667,1671|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|History of Present Illness|1684,1689|true|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|History of Present Illness|1684,1689|true|false|false|C3815497|Cough (guaifenesin)|cough
Finding|Sign or Symptom|History of Present Illness|1684,1689|true|false|false|C0010200|Coughing|cough
Attribute|Clinical Attribute|History of Present Illness|1693,1712|true|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|History of Present Illness|1693,1712|true|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|History of Present Illness|1706,1712|false|false|false|C0225386|Breath|breath
Finding|Idea or Concept|History of Present Illness|1717,1723|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|Review
Finding|Intellectual Product|History of Present Illness|1717,1723|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|Review
Finding|Functional Concept|History of Present Illness|1717,1726|false|false|false|C0699752|Review of|Review of
Attribute|Clinical Attribute|History of Present Illness|1717,1734|false|false|false|C0488564;C0488565||Review of systems
Procedure|Health Care Activity|History of Present Illness|1717,1734|false|false|false|C0489633|Review of systems (procedure)|Review of systems
Finding|Functional Concept|History of Present Illness|1727,1734|false|false|false|C0449913|System|systems
Finding|Finding|History of Present Illness|1737,1743|false|false|false|C1299582|Unable|Unable
Finding|Body Substance|History of Present Illness|1755,1762|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|1755,1762|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|1755,1762|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1771,1776|false|false|false|C1956423|Biphasic Continuous Positive Airway Pressure|BiPAP
Disorder|Disease or Syndrome|Past Medical History|1822,1828|false|false|false|C0002871|Anemia|Anemia
Lab|Laboratory or Test Result|Past Medical History|1831,1853|false|false|false|C0694540|borderline cholesterol|Borderline cholesterol
Drug|Biologically Active Substance|Past Medical History|1842,1853|false|false|false|C0008377|cholesterol|cholesterol
Drug|Organic Chemical|Past Medical History|1842,1853|false|false|false|C0008377|cholesterol|cholesterol
Procedure|Laboratory Procedure|Past Medical History|1842,1853|false|false|false|C0201950|Cholesterol measurement|cholesterol
Finding|Sign or Symptom|Past Medical History|1866,1876|false|false|false|C0016204|Flatulence|Flatulence
Finding|Idea or Concept|Past Medical History|1879,1885|false|false|false|C0018684|Health|Health
Procedure|Health Care Activity|Past Medical History|1879,1897|false|false|false|C0262500|Health maintenance|Health Maintenance
Event|Activity|Past Medical History|1886,1897|false|false|false|C0024501|Maintenance|Maintenance
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1900,1905|false|false|false|C0018787;C4037974|Chest>Heart;Heart|Heart
Disorder|Neoplastic Process|Past Medical History|1900,1905|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|Heart
Finding|Sign or Symptom|Past Medical History|1900,1905|false|false|false|C0795691|HEART PROBLEM|Heart
Finding|Finding|Past Medical History|1900,1912|false|false|false|C0018808|Heart murmur|Heart Murmur
Finding|Finding|Past Medical History|1906,1912|false|false|false|C0018808|Heart murmur|Murmur
Disorder|Disease or Syndrome|Past Medical History|1915,1927|false|false|false|C0020538|Hypertensive disease|Hypertension
Disorder|Disease or Syndrome|Past Medical History|1930,1944|false|false|false|C0020676|Hypothyroidism|Hypothyroidism
Disorder|Disease or Syndrome|Past Medical History|1947,1967|false|false|false|C0026266|Mitral Valve Insufficiency|Mitral Regurgitation
Finding|Finding|Past Medical History|1954,1967|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|Regurgitation
Finding|Sign or Symptom|Past Medical History|1954,1967|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|Regurgitation
Phenomenon|Biologic Function|Past Medical History|1954,1967|false|false|false|C0460152|Regurgitation - mechanism|Regurgitation
Disorder|Disease or Syndrome|Past Medical History|1970,1982|false|false|false|C0029456|Osteoporosis|Osteoporosis
Finding|Finding|Past Medical History|1970,1982|false|false|false|C2911643|Encounter due to family history of osteoporosis|Osteoporosis
Disorder|Disease or Syndrome|Past Medical History|1985,1994|false|false|false|C0032285|Pneumonia|Pneumonia
Disorder|Disease or Syndrome|Past Medical History|1997,2006|false|false|false|C0037199|Sinusitis|Sinusitis
Finding|Conceptual Entity|Family Medical History|2059,2066|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|2059,2066|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Family Medical History|2059,2066|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|2059,2069|false|false|false|C0262926|Medical History|history of
Finding|Finding|Family Medical History|2059,2082|false|false|false|C0455527||history of hypertension
Disorder|Disease or Syndrome|Family Medical History|2070,2082|false|false|false|C0020538|Hypertensive disease|hypertension
Drug|Amino Acid, Peptide, or Protein|Family Medical History|2086,2096|false|false|false|C3812393|ErbB Receptors|her family
Drug|Enzyme|Family Medical History|2086,2096|false|false|false|C3812393|ErbB Receptors|her family
Finding|Receptor|Family Medical History|2086,2096|false|false|false|C3812393|ErbB Receptors|her family
Finding|Classification|Family Medical History|2090,2096|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|Family Medical History|2090,2096|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|Family Medical History|2090,2096|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|Family Medical History|2090,2096|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Attribute|Clinical Attribute|Family Medical History|2108,2114|false|false|false|C4255046||report
Finding|Intellectual Product|Family Medical History|2108,2114|false|false|false|C0684224|Report (document)|report
Procedure|Health Care Activity|Family Medical History|2108,2114|false|false|false|C0700287|Reporting|report
Finding|Conceptual Entity|Family Medical History|2125,2131|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|father
Finding|Idea or Concept|Family Medical History|2125,2131|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|father
Finding|Classification|Family Medical History|2134,2140|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|Family Medical History|2134,2140|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|Family Medical History|2134,2140|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|Family Medical History|2134,2140|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|Family Medical History|2147,2154|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|2147,2154|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Family Medical History|2147,2154|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|2147,2157|false|false|false|C0262926|Medical History|history of
Disorder|Neoplastic Process|Family Medical History|2167,2174|false|false|false|C0006826|Malignant Neoplasms|cancers
Finding|Conceptual Entity|Family Medical History|2207,2214|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|2207,2214|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Family Medical History|2207,2214|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|2207,2217|false|false|false|C0262926|Medical History|history of
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2218,2225|false|false|false|C0038351;C3714551;C4266636|Abdomen>Stomach;Stomach;Stomach structure|stomach
Disorder|Disease or Syndrome|Family Medical History|2218,2225|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Disorder|Neoplastic Process|Family Medical History|2218,2225|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Finding|Finding|Family Medical History|2218,2225|false|false|false|C0577027|Stomach problem|stomach
Procedure|Therapeutic or Preventive Procedure|Family Medical History|2218,2225|false|false|false|C0872393|Procedure on stomach|stomach
Disorder|Neoplastic Process|Family Medical History|2218,2232|false|false|false|C0024623;C0699791|Malignant neoplasm of stomach;Stomach Carcinoma|stomach cancer
Disorder|Neoplastic Process|Family Medical History|2226,2232|false|false|false|C0006826|Malignant Neoplasms|cancer
Finding|Conceptual Entity|Family Medical History|2254,2261|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|2254,2261|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Family Medical History|2254,2261|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|2254,2264|false|false|false|C0262926|Medical History|history of
Anatomy|Body Location or Region|Family Medical History|2265,2271|false|false|false|C0031354;C0230069;C3665375|Anterior portion of neck;Pharyngeal structure;Throat|throat
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2265,2271|false|false|false|C0031354;C0230069;C3665375|Anterior portion of neck;Pharyngeal structure;Throat|throat
Drug|Pharmacologic Substance|Family Medical History|2265,2271|false|false|false|C1950455|Throat Homeopathic Medication|throat
Finding|Body Substance|Family Medical History|2265,2271|false|false|false|C1547926;C1550663|Specimen Type - Throat|throat
Finding|Intellectual Product|Family Medical History|2265,2271|false|false|false|C1547926;C1550663|Specimen Type - Throat|throat
Disorder|Neoplastic Process|Family Medical History|2265,2278|false|false|false|C0740339|Throat cancer|throat cancer
Disorder|Neoplastic Process|Family Medical History|2272,2278|false|false|false|C0006826|Malignant Neoplasms|cancer
Finding|Conceptual Entity|Family Medical History|2296,2303|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|2296,2303|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Family Medical History|2296,2303|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|2296,2306|true|false|false|C0262926|Medical History|history of
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2308,2313|false|false|false|C0009368;C4071907|Abdomen+Pelvis>Colon;Colon structure (body structure)|colon
Disorder|Disease or Syndrome|Family Medical History|2308,2313|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Disorder|Neoplastic Process|Family Medical History|2308,2313|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Finding|Finding|Family Medical History|2308,2313|false|false|false|C0750873|COLON PROBLEM|colon
Disorder|Neoplastic Process|Family Medical History|2308,2321|false|false|false|C0007102|Malignant tumor of colon|colon cancers
Disorder|Neoplastic Process|Family Medical History|2314,2321|false|false|false|C0006826|Malignant Neoplasms|cancers
Finding|Conceptual Entity|Family Medical History|2323,2329|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Idea or Concept|Family Medical History|2323,2329|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Disorder|Disease or Syndrome|Family Medical History|2334,2340|false|false|false|C0038454|Cerebrovascular accident|stroke
Finding|Finding|Family Medical History|2334,2340|false|false|false|C5977286|Stroke (heart beat)|stroke
Finding|Classification|Family Medical History|2345,2351|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|Family Medical History|2345,2351|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|Family Medical History|2345,2351|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|Family Medical History|2345,2351|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|Family Medical History|2360,2366|false|false|false|C1546508|Relationship - Mother|Mother
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2374,2379|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Family Medical History|2374,2379|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Family Medical History|2374,2379|false|false|false|C0795691|HEART PROBLEM|heart
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2374,2385|false|false|false|C0018826;C1305961|Heart Valves|heart valve
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2380,2385|false|false|false|C1186983|Anatomical valve|valve
Finding|Intellectual Product|Family Medical History|2403,2407|true|false|false|C4724437|SURE Test|sure
Finding|Functional Concept|General Exam|2438,2442|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|General Exam|2438,2442|false|false|false|C0582103|Medical Examination|Exam
Procedure|Health Care Activity|General Exam|2448,2457|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Classification|General Exam|2459,2466|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|General Exam|2459,2466|false|false|false|C3812897|General medical service|General
Finding|Finding|General Exam|2468,2473|false|false|false|C0234422|Awake (finding)|Awake
Finding|Functional Concept|General Exam|2475,2486|false|false|false|C1704675|Interaction|interactive
Finding|Finding|General Exam|2507,2515|false|false|false|C1961028|Oriented to place|oriented
Event|Activity|General Exam|2520,2525|false|false|false|C1882509|put - instruction imperative|place
Finding|Functional Concept|General Exam|2520,2525|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|General Exam|2520,2525|false|false|false|C1533810||place
Finding|Finding|General Exam|2529,2533|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|General Exam|2529,2533|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|General Exam|2529,2533|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Disorder|Disease or Syndrome|General Exam|2569,2572|false|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Finding|Intellectual Product|General Exam|2569,2572|false|false|false|C2346952|Bachelor of Education|bed
Finding|Finding|General Exam|2585,2590|false|false|false|C0871754;C5702585|Frail;Frail by Myeloma Frailty Index|frail
Anatomy|Body Location or Region|General Exam|2609,2614|false|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|General Exam|2616,2622|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|General Exam|2616,2622|false|false|false|C0036412|Scleral Diseases|Sclera
Procedure|Health Care Activity|General Exam|2616,2622|false|false|false|C2228481|examination of sclera|Sclera
Finding|Finding|General Exam|2623,2632|false|false|false|C0205180|Anicteric|anicteric
Finding|Body Substance|General Exam|2638,2643|false|false|false|C0026727;C1546714;C2753459|Mucus (substance);mucus layer|mucus
Finding|Intellectual Product|General Exam|2638,2643|false|false|false|C0026727;C1546714;C2753459|Mucus (substance);mucus layer|mucus
Anatomy|Tissue|General Exam|2644,2653|false|false|false|C0025255|Membrane Tissue|membranes
Anatomy|Body Location or Region|General Exam|2657,2661|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Anatomy|Cell Component|General Exam|2657,2661|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Finding|Finding|General Exam|2657,2661|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|Neck
Finding|Functional Concept|General Exam|2663,2669|false|false|false|C0332254|Supple|supple
Finding|Finding|General Exam|2671,2674|false|false|false|C0428897|Jugular venous pressure|JVP
Anatomy|Body Part, Organ, or Organ Component|General Exam|2692,2695|true|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|General Exam|2692,2695|true|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Finding|Gene or Genome|General Exam|2692,2695|true|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Event|Activity|General Exam|2710,2714|false|false|false|C0871208|Rating (action)|rate
Finding|Idea or Concept|General Exam|2710,2714|false|false|false|C1549480|Amount type - Rate|rate
Finding|Finding|General Exam|2719,2725|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|General Exam|2719,2725|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Organ or Tissue Function|General Exam|2749,2757|false|false|false|C0039155|Systole|systolic
Finding|Finding|General Exam|2759,2765|false|false|false|C0018808|Heart murmur|murmur
Anatomy|Cell Component|General Exam|2769,2773|false|false|false|C3890171|dinoflagellate apex|apex
Drug|Amino Acid, Peptide, or Protein|General Exam|2769,2773|false|false|false|C0140145|APEX1 protein, human|apex
Drug|Enzyme|General Exam|2769,2773|false|false|false|C0140145|APEX1 protein, human|apex
Finding|Gene or Genome|General Exam|2769,2773|false|false|false|C1332102|APEX1 gene|apex
Anatomy|Body Part, Organ, or Organ Component|General Exam|2775,2780|false|false|false|C0024109|Lung|Lungs
Finding|Sign or Symptom|General Exam|2782,2786|false|false|false|C0278144|Dull pain|Dull
Drug|Chemical Viewed Functionally|General Exam|2790,2795|false|false|false|C0178499|Base|bases
Disorder|Congenital Abnormality|General Exam|2836,2852|false|false|false|C0158784|Accessory skeletal muscle|accessory muscle
Finding|Finding|General Exam|2836,2856|false|false|false|C1821466|Use of accessory muscles|accessory muscle use
Anatomy|Body Part, Organ, or Organ Component|General Exam|2846,2852|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Anatomy|Tissue|General Exam|2846,2852|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Finding|Functional Concept|General Exam|2853,2856|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|General Exam|2853,2856|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Anatomy|Body Location or Region|General Exam|2858,2865|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|General Exam|2858,2865|false|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Finding|Finding|General Exam|2858,2865|false|false|false|C0941288|Abdomen problem|Abdomen
Disorder|Disease or Syndrome|General Exam|2867,2871|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Finding|Finding|General Exam|2873,2882|false|false|false|C0700124|Dilated|distended
Finding|Finding|General Exam|2907,2915|false|false|false|C0427198|Protective muscle spasm|guarding
Anatomy|Body Part, Organ, or Organ Component|General Exam|2917,2922|false|false|false|C0021853|Intestines|bowel
Phenomenon|Natural Phenomenon or Process|General Exam|2924,2930|false|false|false|C0037709||sounds
Finding|Finding|General Exam|2931,2938|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|General Exam|2931,2938|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Sign or Symptom|General Exam|2960,2972|false|false|false|C0011991;C2129214|Diarrhea;Loose stool|watery stool
Finding|Body Substance|General Exam|2967,2972|false|false|false|C0015733|Feces|stool
Disorder|Disease or Syndrome|General Exam|2978,2983|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|General Exam|2978,2983|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Event|Activity|General Exam|3005,3010|false|false|false|C1882509|put - instruction imperative|place
Finding|Functional Concept|General Exam|3005,3010|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|General Exam|3005,3010|false|false|false|C1533810||place
Disorder|Congenital Abnormality|General Exam|3018,3021|false|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Finding|Gene or Genome|General Exam|3018,3021|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Finding|Finding|General Exam|3023,3027|false|false|false|C0582051|Feels warm|warm
Phenomenon|Natural Phenomenon or Process|General Exam|3023,3027|false|false|false|C0687712|warming process|warm
Drug|Food|General Exam|3035,3041|false|false|false|C5890763||pulses
Finding|Physiologic Function|General Exam|3035,3041|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|General Exam|3035,3041|false|false|false|C0034107|Pulse taking|pulses
Attribute|Clinical Attribute|General Exam|3051,3056|false|false|false|C1717255||edema
Finding|Pathologic Function|General Exam|3051,3056|false|false|false|C0013604|Edema|edema
Finding|Finding|General Exam|3073,3079|false|false|false|C1554187|Gender Status - Intact|intact
Disorder|Mental or Behavioral Dysfunction|General Exam|3094,3105|false|false|false|C0424101|Inattention|inattentive
Finding|Body Substance|General Exam|3107,3116|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|General Exam|3107,3116|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|General Exam|3107,3116|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|General Exam|3107,3116|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Functional Concept|General Exam|3117,3121|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|General Exam|3117,3121|false|false|false|C0582103|Medical Examination|exam
Finding|Finding|General Exam|3124,3133|false|false|false|C0442739||unchanged
Finding|Idea or Concept|General Exam|3139,3144|false|false|false|C1552828|Table Frame - above|above
Finding|Classification|General Exam|3163,3170|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|General Exam|3163,3170|false|false|false|C3812897|General medical service|General
Finding|Finding|General Exam|3172,3177|false|false|false|C0234422|Awake (finding)|Awake
Finding|Finding|General Exam|3179,3185|false|false|false|C0013144|Drowsiness|sleepy
Finding|Idea or Concept|General Exam|3203,3208|false|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Finding|Intellectual Product|General Exam|3203,3208|false|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Finding|Organism Function|General Exam|3203,3208|false|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Disorder|Disease or Syndrome|General Exam|3210,3213|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|General Exam|3210,3213|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|General Exam|3210,3213|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|3210,3213|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|General Exam|3210,3213|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Finding|Finding|General Exam|3210,3213|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Finding|Gene or Genome|General Exam|3241,3244|false|false|false|C1540289|CD200 gene|Ox2
Finding|Intellectual Product|General Exam|3246,3250|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|name
Lab|Laboratory or Test Result|General Exam|3329,3333|false|false|false|C0587081|Laboratory test finding|Labs
Procedure|Health Care Activity|General Exam|3339,3348|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Disorder|Disease or Syndrome|General Exam|3362,3367|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|3362,3367|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|3368,3371|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|3376,3379|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|3376,3379|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|3376,3379|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|3386,3389|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|3386,3389|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|3386,3389|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|3386,3389|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|3395,3398|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|3395,3398|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|3406,3409|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|General Exam|3406,3409|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|3406,3409|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|3406,3409|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|3413,3416|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|3413,3416|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|General Exam|3413,3416|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|3413,3416|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|3413,3416|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|General Exam|3422,3426|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|3442,3445|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|3462,3467|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|3462,3467|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Antibiotic|General Exam|3483,3488|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|General Exam|3483,3488|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|General Exam|3483,3488|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|General Exam|3493,3496|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|Eos
Finding|Gene or Genome|General Exam|3493,3496|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|Eos
Disorder|Disease or Syndrome|General Exam|3523,3528|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|3523,3528|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|3523,3536|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|3523,3536|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|3523,3536|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|3529,3536|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|3529,3536|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|3529,3536|false|false|false|C0017725|glucose|Glucose
Lab|Laboratory or Test Result|General Exam|3529,3536|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|3529,3536|false|false|false|C0337438|Glucose measurement|Glucose
Disorder|Disease or Syndrome|General Exam|3613,3618|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|3613,3618|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|3619,3622|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|General Exam|3619,3622|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|General Exam|3619,3622|false|false|false|C0001899|Alanine Transaminase|ALT
Finding|Gene or Genome|General Exam|3619,3622|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|General Exam|3619,3622|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|General Exam|3619,3622|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|General Exam|3619,3622|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|General Exam|3626,3629|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|General Exam|3626,3629|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|3626,3629|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|General Exam|3626,3629|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|General Exam|3626,3629|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Finding|Gene or Genome|General Exam|3626,3629|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|3633,3640|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|General Exam|3633,3640|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Disorder|Disease or Syndrome|General Exam|3670,3675|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|3670,3675|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|General Exam|3701,3706|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|3701,3706|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|3701,3714|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|General Exam|3707,3714|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|General Exam|3707,3714|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|General Exam|3707,3714|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|General Exam|3707,3714|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|General Exam|3707,3714|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Finding|Physiologic Function|General Exam|3707,3714|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|General Exam|3707,3714|false|false|false|C0201925|Calcium measurement|Calcium
Disorder|Disease or Syndrome|General Exam|3749,3754|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|3749,3754|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Attribute|Clinical Attribute|General Exam|3749,3759|false|false|false|C1383165|Blood Type|BLOOD Type
Finding|Classification|General Exam|3749,3759|false|false|false|C0005810;C2911644|Blood Group Systems;Encounter due to blood type|BLOOD Type
Finding|Finding|General Exam|3749,3759|false|false|false|C0005810;C2911644|Blood Group Systems;Encounter due to blood type|BLOOD Type
Procedure|Laboratory Procedure|General Exam|3749,3759|false|false|false|C0005844|Blood group typing (procedure)|BLOOD Type
Finding|Gene or Genome|General Exam|3755,3759|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|Type
Finding|Intellectual Product|General Exam|3755,3759|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|Type
Drug|Organic Chemical|General Exam|3760,3763|false|false|false|C0052432|artesunate|ART
Drug|Pharmacologic Substance|General Exam|3760,3763|false|false|false|C0052432|artesunate|ART
Finding|Gene or Genome|General Exam|3760,3763|false|false|false|C1412286;C3890191|AGRP gene;AGRP wt Allele|ART
Procedure|Therapeutic or Preventive Procedure|General Exam|3760,3763|false|false|false|C0872104;C1963724|Antiretroviral therapy;Assisted Reproductive Technologies|ART
Finding|Gene or Genome|General Exam|3764,3768|false|false|false|C1823816|C1orf210 gene|Temp
Procedure|Therapeutic or Preventive Procedure|General Exam|3764,3768|false|false|false|C0279848|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Temp
Finding|Finding|General Exam|3786,3790|false|false|false|C3494516|Positive end expiratory pressure (finding)|PEEP
Procedure|Therapeutic or Preventive Procedure|General Exam|3786,3790|false|false|false|C0032740|Positive End-Expiratory Pressure|PEEP
Attribute|Clinical Attribute|General Exam|3794,3798|false|false|false|C3484065||FiO2
Finding|Finding|General Exam|3794,3798|false|false|false|C0428167|Fraction of inspired oxygen|FiO2
Procedure|Diagnostic Procedure|General Exam|3794,3798|false|false|false|C1512797;C2370852|Inspired Oxygen Fraction Test;fraction of inspired oxygen (FiO2) (treatment)|FiO2
Procedure|Therapeutic or Preventive Procedure|General Exam|3794,3798|false|false|false|C1512797;C2370852|Inspired Oxygen Fraction Test;fraction of inspired oxygen (FiO2) (treatment)|FiO2
Finding|Classification|General Exam|3802,3805|false|false|false|C0391840;C4521535|Partial pressure of Oxygen;US Military enlisted E5|pO2
Finding|Molecular Function|General Exam|3802,3805|false|false|false|C0391840;C4521535|Partial pressure of Oxygen;US Military enlisted E5|pO2
Procedure|Laboratory Procedure|General Exam|3802,3805|false|false|false|C1283004|PO2 measurement|pO2
Lab|Laboratory or Test Result|General Exam|3811,3815|false|false|false|C0391839|Carbon dioxide, partial pressure|pCO2
Procedure|Laboratory Procedure|General Exam|3811,3815|false|false|false|C0201931|Carbon dioxide measurement, partial pressure|pCO2
Anatomy|Body Location or Region|General Exam|3840,3844|false|false|false|C2987514|Anatomical base|Base
Drug|Biomedical or Dental Material|General Exam|3840,3844|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|Base
Drug|Chemical Viewed Functionally|General Exam|3840,3844|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|Base
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|3840,3844|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|Base
Finding|Gene or Genome|General Exam|3840,3844|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|Base
Finding|Idea or Concept|General Exam|3840,3844|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|Base
Drug|Organic Chemical|General Exam|3845,3850|false|false|false|C5557572|Pam3Cys-GDPKHPKSF XS15|XS-15
Drug|Pharmacologic Substance|General Exam|3845,3850|false|false|false|C5557572|Pam3Cys-GDPKHPKSF XS15|XS-15
Disorder|Disease or Syndrome|General Exam|3883,3888|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|3883,3888|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|3883,3896|false|false|false|C3824990|lactate in blood (lab test)|BLOOD Lactate
Drug|Organic Chemical|General Exam|3889,3896|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Drug|Pharmacologic Substance|General Exam|3889,3896|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Procedure|Laboratory Procedure|General Exam|3889,3896|false|false|false|C0202115|Lactic acid measurement|Lactate
Finding|Body Substance|General Exam|3902,3911|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|General Exam|3902,3911|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|General Exam|3902,3911|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|General Exam|3902,3911|false|false|false|C0030685|Patient Discharge|Discharge
Lab|Laboratory or Test Result|General Exam|3912,3916|false|false|false|C0587081|Laboratory test finding|labs
Disorder|Disease or Syndrome|General Exam|3930,3935|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|3930,3935|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|3936,3939|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|3944,3947|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|3944,3947|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|3944,3947|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|3954,3957|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|3954,3957|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|3954,3957|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|3954,3957|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|3963,3966|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|3963,3966|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|3974,3977|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|General Exam|3974,3977|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|3974,3977|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|3974,3977|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|3982,3985|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|3982,3985|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|General Exam|3982,3985|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|3982,3985|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|3982,3985|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|General Exam|3991,3995|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|4010,4013|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|4030,4035|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4030,4035|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|4030,4043|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|4030,4043|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|4030,4043|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|4036,4043|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|4036,4043|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|4036,4043|false|false|false|C0017725|glucose|Glucose
Lab|Laboratory or Test Result|General Exam|4036,4043|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|4036,4043|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|General Exam|4089,4093|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|4089,4093|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|General Exam|4089,4093|false|false|false|C0202059|Bicarbonate measurement|HCO3
Finding|Conceptual Entity|General Exam|4107,4112|false|false|false|C3811161;C4049106|Micro (prefix);Microbiology - Laboratory Class|Micro
Finding|Intellectual Product|General Exam|4107,4112|false|false|false|C3811161;C4049106|Micro (prefix);Microbiology - Laboratory Class|Micro
Procedure|Laboratory Procedure|General Exam|4107,4112|false|false|false|C0085672|Microbiology procedure|Micro
Drug|Food|General Exam|4140,4145|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|Yeast
Drug|Immunologic Factor|General Exam|4140,4145|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|Yeast
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|4140,4145|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|Yeast
Drug|Pharmacologic Substance|General Exam|4140,4145|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|Yeast
Lab|Laboratory or Test Result|General Exam|4150,4166|true|false|false|C0427944|Determination of bacterial growth|bacterial growth
Finding|Finding|General Exam|4160,4166|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|growth
Finding|Organ or Tissue Function|General Exam|4160,4166|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|growth
Finding|Organism Function|General Exam|4160,4166|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|growth
Finding|Physiologic Function|General Exam|4160,4166|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|growth
Phenomenon|Phenomenon or Process|General Exam|4160,4166|true|false|false|C2911660|Growth action|growth
Anatomy|Cell Component|General Exam|4168,4175|false|false|false|C1660780|midline cell component|Midline
Finding|Gene or Genome|General Exam|4176,4179|false|false|false|C1705504;C1823282;C1825626;C1825978|ITFG1 gene;KAT5 wt Allele;METTL8 gene;TIPRL gene|tip
Procedure|Therapeutic or Preventive Procedure|General Exam|4176,4179|false|false|false|C0673828|TIP regimen|tip
Finding|Finding|General Exam|4196,4199|false|false|false|C4050242;C5202919|Pathologic Complete Response;Residual Cancer Burden Class 0|PCR
Procedure|Laboratory Procedure|General Exam|4196,4199|false|false|false|C0032520;C3853643|Polymerase Chain Reaction;Probe with target amplification technique|PCR
Procedure|Molecular Biology Research Technique|General Exam|4196,4199|false|false|false|C0032520;C3853643|Polymerase Chain Reaction;Probe with target amplification technique|PCR
Finding|Finding|General Exam|4202,4205|false|false|false|C5848551|Neg - answer|neg
Finding|Finding|General Exam|4207,4214|false|false|false|C0740845|Imaging problem|Imaging
Procedure|Diagnostic Procedure|General Exam|4207,4214|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|Imaging
Procedure|Diagnostic Procedure|General Exam|4222,4225|false|false|false|C0039985|Plain chest X-ray|CXR
Finding|Intellectual Product|General Exam|4227,4237|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|General Exam|4227,4237|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Idea or Concept|General Exam|4243,4254|true|false|false|C0750502|Significant|significant
Finding|Intellectual Product|General Exam|4255,4263|true|false|false|C1552654|Parameterized Data Type - Interval|interval
Finding|Finding|General Exam|4255,4270|true|false|false|C2041208||interval change
Finding|Functional Concept|General Exam|4264,4270|true|false|false|C0392747|Changing|change
Procedure|Therapeutic or Preventive Procedure|General Exam|4264,4270|true|false|false|C4319952|Change - procedure|change
Anatomy|Tissue|General Exam|4287,4294|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|General Exam|4287,4294|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Pathologic Function|General Exam|4287,4304|false|false|false|C0032227|Pleural effusion (disorder)|pleural effusions
Finding|Pathologic Function|General Exam|4295,4304|false|false|false|C0013687|effusion|effusions
Finding|Functional Concept|General Exam|4310,4315|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Finding|Intellectual Product|General Exam|4324,4332|false|false|false|C1546572||catheter
Anatomy|Body Location or Region|General Exam|4341,4346|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|General Exam|4341,4346|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Location or Region|General Exam|4341,4352|false|false|false|C0446470|Surface region of lower chest|lower chest
Anatomy|Body Location or Region|General Exam|4347,4352|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|General Exam|4347,4352|false|false|false|C0741025|Chest problem|chest
Finding|Finding|General Exam|4355,4363|false|false|false|C0332149|Possible|Possible
Finding|Functional Concept|General Exam|4370,4375|false|true|false|C1552823|Table Cell Horizontal Align - right|right
Disorder|Disease or Syndrome|General Exam|4383,4395|false|false|false|C0032326|Pneumothorax|pneumothorax
Finding|Intellectual Product|General Exam|4409,4419|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|General Exam|4409,4419|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Idea or Concept|General Exam|4429,4437|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|General Exam|4429,4440|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Anatomy|Body Part, Organ, or Organ Component|General Exam|4441,4450|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|General Exam|4441,4450|true|false|false|C2707265||pulmonary
Finding|Finding|General Exam|4441,4450|true|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|General Exam|4441,4459|true|false|false|C0034065|Pulmonary Embolism|pulmonary embolism
Finding|Finding|General Exam|4451,4459|true|false|false|C0013922;C1704212|Embolism;Embolus|embolism
Finding|Pathologic Function|General Exam|4451,4459|true|false|false|C0013922;C1704212|Embolism;Embolus|embolism
Anatomy|Tissue|General Exam|4476,4483|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|General Exam|4476,4483|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Pathologic Function|General Exam|4476,4493|false|false|false|C0032227|Pleural effusion (disorder)|pleural effusions
Finding|Pathologic Function|General Exam|4484,4493|false|false|false|C0013687|effusion|effusions
Finding|Finding|General Exam|4504,4512|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|General Exam|4504,4512|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Functional Concept|General Exam|4520,4524|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Event|Activity|General Exam|4566,4577|false|false|false|C4321457|Examination|examination
Procedure|Health Care Activity|General Exam|4566,4577|false|false|false|C0031809;C0582103|Medical Examination;Physical Examination|examination
Finding|Functional Concept|General Exam|4582,4587|false|false|false|C1883002|Sequence Chromatogram|trace
Finding|Functional Concept|General Exam|4595,4600|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Finding|Intellectual Product|General Exam|4652,4660|false|false|false|C1546572||catheter
Event|Activity|General Exam|4671,4676|false|false|false|C1882509|put - instruction imperative|place
Finding|Functional Concept|General Exam|4671,4676|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|General Exam|4671,4676|false|false|false|C1533810||place
Finding|Functional Concept|General Exam|4684,4689|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Disorder|Disease or Syndrome|General Exam|4698,4705|false|false|false|C0003962|Ascites|Ascites
Finding|Pathologic Function|General Exam|4698,4705|false|false|false|C5441966|Peritoneal Effusion|Ascites
Finding|Idea or Concept|Hospital Course|4738,4742|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|Hospital Course|4738,4742|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Disorder|Disease or Syndrome|Hospital Course|4793,4799|false|false|false|C0036690;C0243026|Sepsis;Septicemia|sepsis
Finding|Pathologic Function|Hospital Course|4805,4810|false|false|false|C0036974|Shock|shock
Finding|Mental Process|Hospital Course|4854,4860|false|false|false|C0229992|Psyche structure|mental
Attribute|Clinical Attribute|Hospital Course|4854,4867|false|false|false|C0488568;C0488569||mental status
Finding|Finding|Hospital Course|4854,4867|false|false|false|C0278060|Mental state|mental status
Attribute|Clinical Attribute|Hospital Course|4861,4867|false|false|false|C5889824||status
Finding|Idea or Concept|Hospital Course|4861,4867|false|false|false|C1546481|What subject filter - Status|status
Finding|Finding|Hospital Course|4869,4878|false|false|false|C0231835|Tachypnea|tachypnea
Finding|Intellectual Product|Hospital Course|4885,4889|false|false|false|C1547225|Mild Severity of Illness Code|mild
Attribute|Clinical Attribute|Hospital Course|4890,4901|false|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|Hospital Course|4890,4901|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|Hospital Course|4890,4901|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|Hospital Course|4890,4901|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Disorder|Disease or Syndrome|Hospital Course|4890,4910|false|false|false|C0001127|Acidosis, Respiratory|respiratory acidosis
Finding|Pathologic Function|Hospital Course|4902,4910|false|false|false|C0001122|Acidosis|acidosis
Finding|Finding|Hospital Course|4914,4921|false|false|false|C0242184;C1963140|Hypoxia;Hypoxia, CTCAE|Hypoxia
Finding|Pathologic Function|Hospital Course|4914,4921|false|false|false|C0242184;C1963140|Hypoxia;Hypoxia, CTCAE|Hypoxia
Finding|Finding|Hospital Course|4922,4933|false|false|false|C0020440|Hypercapnia|hypercarbia
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4958,4963|false|false|false|C1956423|Biphasic Continuous Positive Airway Pressure|BiPAP
Event|Activity|Hospital Course|4998,5008|false|false|false|C1283169||monitoring
Procedure|Health Care Activity|Hospital Course|4998,5008|false|false|false|C0150369|Preventive monitoring|monitoring
Attribute|Clinical Attribute|Hospital Course|5016,5027|false|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|Hospital Course|5016,5027|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|Hospital Course|5016,5027|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|Hospital Course|5016,5027|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Attribute|Clinical Attribute|Hospital Course|5016,5034|false|false|false|C2598168||respiratory status
Finding|Finding|Hospital Course|5016,5034|false|false|false|C1998827|Respiratory Status|respiratory status
Attribute|Clinical Attribute|Hospital Course|5028,5034|false|false|false|C5889824||status
Finding|Idea or Concept|Hospital Course|5028,5034|false|false|false|C1546481|What subject filter - Status|status
Finding|Finding|Hospital Course|5046,5050|false|false|false|C1299581|Able (qualifier value)|able
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5069,5074|false|false|false|C1956423|Biphasic Continuous Positive Airway Pressure|BiPAP
Anatomy|Body Space or Junction|Hospital Course|5078,5081|false|false|false|C0228479|Structure of intraculminate fissure|ICU
Finding|Intellectual Product|Hospital Course|5078,5081|false|false|false|C4554035|Inventory of Callous-Unemotional Traits|ICU
Finding|Idea or Concept|Hospital Course|5082,5085|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|5082,5085|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Finding|Hospital Course|5082,5087|false|false|false|C3842676|Day 2|day 2
Finding|Finding|Hospital Course|5118,5122|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Hospital Course|5118,5122|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Hospital Course|5118,5122|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Body Substance|Hospital Course|5126,5135|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|5126,5135|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|5126,5135|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|5126,5135|false|false|false|C0030685|Patient Discharge|discharge
Finding|Conceptual Entity|Hospital Course|5138,5143|false|false|false|C0015127;C1524003|Etiology aspects;Science of Etiology|Cause
Finding|Functional Concept|Hospital Course|5138,5143|false|false|false|C0015127;C1524003|Etiology aspects;Science of Etiology|Cause
Attribute|Clinical Attribute|Hospital Course|5151,5162|false|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|Hospital Course|5151,5162|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|Hospital Course|5151,5162|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|Hospital Course|5151,5162|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|Hospital Course|5164,5172|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Hospital Course|5164,5172|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Pathologic Function|Hospital Course|5203,5218|false|false|false|C3203358|Hypoventilation|hypoventilation
Disorder|Mental or Behavioral Dysfunction|Hospital Course|5225,5235|false|false|false|C2830004|Somnolence|somnolence
Finding|Finding|Hospital Course|5225,5235|false|false|false|C0013144|Drowsiness|somnolence
Drug|Organic Chemical|Hospital Course|5236,5243|false|false|false|C0163712|Relate - vinyl resin|related
Finding|Finding|Hospital Course|5236,5243|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Finding|Functional Concept|Hospital Course|5236,5243|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Finding|Finding|Hospital Course|5247,5259|false|false|false|C0542127|Oversedation|oversedation
Drug|Organic Chemical|Hospital Course|5265,5272|false|false|false|C0527258|Zyprexa|Zyprexa
Drug|Pharmacologic Substance|Hospital Course|5265,5272|false|false|false|C0527258|Zyprexa|Zyprexa
Drug|Organic Chemical|Hospital Course|5275,5282|false|false|false|C0527258|Zyprexa|Zyprexa
Drug|Pharmacologic Substance|Hospital Course|5275,5282|false|false|false|C0527258|Zyprexa|Zyprexa
Finding|Finding|Hospital Course|5300,5304|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Hospital Course|5300,5304|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Hospital Course|5300,5304|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Body Substance|Hospital Course|5308,5317|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|5308,5317|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|5308,5317|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|5308,5317|false|false|false|C0030685|Patient Discharge|discharge
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5320,5323|false|false|false|C3813556|Cancer/Testis Antigen|CTA
Finding|Gene or Genome|Hospital Course|5320,5323|false|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|Hospital Course|5320,5323|false|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Anatomy|Body Location or Region|Hospital Course|5324,5329|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|Hospital Course|5324,5329|false|false|false|C0741025|Chest problem|Chest
Finding|Classification|Hospital Course|5334,5342|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|5334,5342|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|5334,5342|false|false|false|C5237010|Expression Negative|negative
Finding|Finding|Hospital Course|5334,5346|false|false|false|C0205160|Negative|negative for
Finding|Idea or Concept|Hospital Course|5365,5370|false|false|false|C1550016|Remote control command - Clear|clear
Finding|Idea or Concept|Hospital Course|5371,5379|false|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Hospital Course|5371,5382|false|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Disorder|Disease or Syndrome|Hospital Course|5383,5392|true|false|false|C0032285|Pneumonia|pneumonia
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5425,5429|false|false|false|C0535219|SMC3 protein, human|HCAP
Drug|Biologically Active Substance|Hospital Course|5425,5429|false|false|false|C0535219|SMC3 protein, human|HCAP
Finding|Gene or Genome|Hospital Course|5425,5429|false|false|false|C1419431;C1422826;C1704469;C1822780|DCD gene;RNGTT gene;SMC3 gene;SMC3 wt Allele|HCAP
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5425,5429|false|false|false|C0056451|Cyclophosphamide/Altretamine/Doxorubicin/Cisplatin Regimen|HCAP
Drug|Antibiotic|Hospital Course|5430,5441|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Drug|Antibiotic|Hospital Course|5452,5460|false|false|false|C0055003|cefepime|cefepime
Drug|Organic Chemical|Hospital Course|5452,5460|false|false|false|C0055003|cefepime|cefepime
Finding|Body Substance|Hospital Course|5498,5507|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|5498,5507|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|5498,5507|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|5498,5507|false|false|false|C0030685|Patient Discharge|discharge
Finding|Idea or Concept|Hospital Course|5523,5531|false|true|false|C0010453|Culture (Anthropological)|cultures
Finding|Classification|Hospital Course|5538,5546|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|5538,5546|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|5538,5546|false|false|false|C5237010|Expression Negative|negative
Disorder|Disease or Syndrome|Hospital Course|5564,5577|true|false|false|C0521530|Lung consolidation|consolidation
Finding|Finding|Hospital Course|5581,5588|false|false|false|C0740845|Imaging problem|imaging
Procedure|Diagnostic Procedure|Hospital Course|5581,5588|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|imaging
Disorder|Mental or Behavioral Dysfunction|Hospital Course|5594,5602|false|false|false|C0011206|Delirium|Delirium
Finding|Finding|Hospital Course|5604,5610|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Finding|Idea or Concept|Hospital Course|5604,5610|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Finding|Finding|Hospital Course|5611,5625|false|true|false|C1837655|Multifactorial|multifactorial
Drug|Organic Chemical|Hospital Course|5645,5652|false|true|false|C0163712|Relate - vinyl resin|related
Finding|Finding|Hospital Course|5645,5652|false|true|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Finding|Functional Concept|Hospital Course|5645,5652|false|true|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Finding|Finding|Hospital Course|5657,5669|false|false|false|C0542127|Oversedation|oversedation
Drug|Organic Chemical|Hospital Course|5675,5682|false|false|false|C0527258|Zyprexa|Zyprexa
Drug|Pharmacologic Substance|Hospital Course|5675,5682|false|false|false|C0527258|Zyprexa|Zyprexa
Finding|Idea or Concept|Hospital Course|5698,5706|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Hospital Course|5698,5709|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Disorder|Disease or Syndrome|Hospital Course|5710,5719|true|false|false|C0009450|Communicable Diseases|infection
Finding|Pathologic Function|Hospital Course|5710,5719|true|false|false|C3714514|Infection|infection
Drug|Antibiotic|Hospital Course|5725,5736|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Finding|Idea or Concept|Hospital Course|5771,5776|false|false|false|C1552828|Table Frame - above|above
Finding|Classification|Hospital Course|5806,5814|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|5806,5814|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|5806,5814|false|false|false|C5237010|Expression Negative|negative
Drug|Food|Hospital Course|5829,5834|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|yeast
Drug|Immunologic Factor|Hospital Course|5829,5834|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|yeast
Drug|Indicator, Reagent, or Diagnostic Aid|Hospital Course|5829,5834|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|yeast
Drug|Pharmacologic Substance|Hospital Course|5829,5834|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|yeast
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5852,5859|false|false|false|C0042027|Urinary tract|urinary
Finding|Sign or Symptom|Hospital Course|5852,5868|false|false|false|C0426359|Urinary symptoms|urinary symptoms
Finding|Functional Concept|Hospital Course|5860,5868|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Hospital Course|5860,5868|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Mental Process|Hospital Course|5883,5889|false|false|false|C0229992|Psyche structure|mental
Attribute|Clinical Attribute|Hospital Course|5883,5896|false|false|false|C0488568;C0488569||mental status
Finding|Finding|Hospital Course|5883,5896|false|false|false|C0278060|Mental state|mental status
Finding|Finding|Hospital Course|5883,5904|false|false|false|C0856054|Mental status changes|mental status changes
Attribute|Clinical Attribute|Hospital Course|5890,5896|false|false|false|C5889824||status
Finding|Idea or Concept|Hospital Course|5890,5896|false|false|false|C1546481|What subject filter - Status|status
Finding|Functional Concept|Hospital Course|5897,5904|false|false|false|C0392747|Changing|changes
Finding|Finding|Hospital Course|5911,5919|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|probably
Finding|Idea or Concept|Hospital Course|5911,5919|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|probably
Drug|Organic Chemical|Hospital Course|5920,5927|false|false|false|C0163712|Relate - vinyl resin|related
Finding|Finding|Hospital Course|5920,5927|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Finding|Functional Concept|Hospital Course|5920,5927|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Attribute|Clinical Attribute|Hospital Course|5945,5956|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Hospital Course|5945,5956|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|Hospital Course|5945,5956|false|false|false|C4284232|Medications|medications
Finding|Finding|Hospital Course|5961,5972|false|false|false|C0020440|Hypercapnia|hypercarbia
Procedure|Health Care Activity|Hospital Course|5977,5986|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6008,6013|false|false|false|C1956423|Biphasic Continuous Positive Airway Pressure|BiPAP
Drug|Pharmacologic Substance|Hospital Course|6031,6045|false|false|false|C0040615|Antipsychotic Agents|antipsychotics
Disorder|Disease or Syndrome|Hospital Course|6057,6064|false|false|false|C0009319|Colitis|Colitis
Disorder|Disease or Syndrome|Hospital Course|6096,6103|false|false|false|C0009319|Colitis|colitis
Disorder|Disease or Syndrome|Hospital Course|6110,6116|false|false|false|C0036690;C0243026|Sepsis;Septicemia|sepsis
Finding|Functional Concept|Hospital Course|6118,6124|false|false|false|C0205341;C1705914|Repeat;Repeat Object|Repeat
Finding|Finding|Hospital Course|6132,6135|false|false|false|C4050242;C5202919|Pathologic Complete Response;Residual Cancer Burden Class 0|PCR
Procedure|Laboratory Procedure|Hospital Course|6132,6135|false|false|false|C0032520;C3853643|Polymerase Chain Reaction;Probe with target amplification technique|PCR
Procedure|Molecular Biology Research Technique|Hospital Course|6132,6135|false|false|false|C0032520;C3853643|Polymerase Chain Reaction;Probe with target amplification technique|PCR
Finding|Classification|Hospital Course|6140,6148|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|6140,6148|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|6140,6148|false|false|false|C5237010|Expression Negative|negative
Procedure|Health Care Activity|Hospital Course|6162,6177|false|false|false|C0019993|Hospitalization|hospitalization
Finding|Finding|Hospital Course|6201,6205|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|Hospital Course|6201,6205|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|Hospital Course|6201,6205|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|Hospital Course|6206,6212|false|false|false|C1705102|Volume (publication)|volume
Finding|Body Substance|Hospital Course|6213,6218|false|false|false|C0015733|Feces|stool
Finding|Conceptual Entity|Hospital Course|6219,6225|false|false|false|C1709366|system output|output
Procedure|Health Care Activity|Hospital Course|6219,6225|false|false|false|C3251815|Measurement of fluid output|output
Event|Activity|Hospital Course|6247,6252|false|false|false|C1882509|put - instruction imperative|place
Finding|Functional Concept|Hospital Course|6247,6252|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|Hospital Course|6247,6252|false|false|false|C1533810||place
Anatomy|Body System|Hospital Course|6257,6261|false|false|false|C1123023;C4520765|Skin;Skin, Human|skin
Disorder|Disease or Syndrome|Hospital Course|6257,6261|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Disorder|Neoplastic Process|Hospital Course|6257,6261|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Finding|Body Substance|Hospital Course|6257,6261|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Finding|Intellectual Product|Hospital Course|6257,6261|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Finding|Pathologic Function|Hospital Course|6257,6272|false|false|false|C0037299|Skin Ulcer|skin ulceration
Finding|Pathologic Function|Hospital Course|6262,6272|false|false|false|C0041582;C3887532|Ulcer;Ulceration|ulceration
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6303,6308|false|false|false|C0042313|vancomycin|vanco
Drug|Antibiotic|Hospital Course|6303,6308|false|false|false|C0042313|vancomycin|vanco
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6355,6359|false|false|false|C0535219|SMC3 protein, human|HCAP
Drug|Biologically Active Substance|Hospital Course|6355,6359|false|false|false|C0535219|SMC3 protein, human|HCAP
Finding|Gene or Genome|Hospital Course|6355,6359|false|false|false|C1419431;C1422826;C1704469;C1822780|DCD gene;RNGTT gene;SMC3 gene;SMC3 wt Allele|HCAP
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6355,6359|false|false|false|C0056451|Cyclophosphamide/Altretamine/Doxorubicin/Cisplatin Regimen|HCAP
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6382,6387|false|false|false|C0042313|vancomycin|vanco
Drug|Antibiotic|Hospital Course|6382,6387|false|false|false|C0042313|vancomycin|vanco
Drug|Antibiotic|Hospital Course|6448,6456|false|false|false|C0055003|cefepime|cefepime
Drug|Organic Chemical|Hospital Course|6448,6456|false|false|false|C0055003|cefepime|cefepime
Event|Activity|Hospital Course|6489,6494|false|false|false|C1882509|put - instruction imperative|place
Finding|Functional Concept|Hospital Course|6489,6494|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|Hospital Course|6489,6494|false|false|false|C1533810||place
Finding|Body Substance|Hospital Course|6498,6507|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|6498,6507|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|6498,6507|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|6498,6507|false|false|false|C0030685|Patient Discharge|discharge
Disorder|Disease or Syndrome|Hospital Course|6512,6518|false|false|false|C0002871|Anemia|Anemia
Finding|Body Substance|Hospital Course|6520,6527|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|6520,6527|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|6520,6527|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Indicator, Reagent, or Diagnostic Aid|Hospital Course|6533,6539|false|false|false|C0018302|guaiac|guaiac
Drug|Organic Chemical|Hospital Course|6533,6539|false|false|false|C0018302|guaiac|guaiac
Lab|Laboratory or Test Result|Hospital Course|6533,6548|false|false|false|C0744492|guaiac positive|guaiac positive
Finding|Finding|Hospital Course|6533,6555|false|false|false|C0266813||guaiac positive stools
Disorder|Cell or Molecular Dysfunction|Hospital Course|6540,6548|false|false|false|C4727483|BRAF Gene Rearrangement|positive
Finding|Classification|Hospital Course|6540,6548|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|Hospital Course|6540,6548|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Attribute|Clinical Attribute|Hospital Course|6549,6555|false|false|false|C0489144||stools
Finding|Body Substance|Hospital Course|6549,6555|false|false|false|C0015733|Feces|stools
Procedure|Health Care Activity|Hospital Course|6561,6570|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Finding|Hospital Course|6573,6576|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Hospital Course|6573,6576|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Procedure|Health Care Activity|Hospital Course|6587,6596|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Disorder|Neoplastic Process|Hospital Course|6610,6619|false|false|false|C0027627|Neoplasm Metastasis|secondary
Finding|Functional Concept|Hospital Course|6610,6619|false|false|false|C1522484|metastatic qualifier|secondary
Finding|Pathologic Function|Hospital Course|6623,6632|false|false|false|C0027544|Necrotic debris|sloughing
Anatomy|Tissue|Hospital Course|6638,6645|false|false|false|C0026724|Mucous Membrane|mucosal
Finding|Finding|Hospital Course|6646,6652|false|false|false|C1446325;C2089742|Oozing (Hemorrhage);oozing skin lesion|oozing
Finding|Pathologic Function|Hospital Course|6646,6652|false|false|false|C1446325;C2089742|Oozing (Hemorrhage);oozing skin lesion|oozing
Disorder|Neoplastic Process|Hospital Course|6653,6662|false|false|false|C0027627|Neoplasm Metastasis|secondary
Finding|Functional Concept|Hospital Course|6653,6662|false|false|false|C1522484|metastatic qualifier|secondary
Drug|Organic Chemical|Hospital Course|6681,6688|false|false|false|C0022924;C0376261|Lactates;lactate|lactate
Drug|Pharmacologic Substance|Hospital Course|6681,6688|false|false|false|C0022924;C0376261|Lactates;lactate|lactate
Procedure|Laboratory Procedure|Hospital Course|6681,6688|false|false|false|C0202115|Lactic acid measurement|lactate
Procedure|Health Care Activity|Hospital Course|6692,6701|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Anatomy|Body Location or Region|Hospital Course|6714,6723|false|false|false|C0000726|Abdomen|abdominal
Procedure|Diagnostic Procedure|Hospital Course|6714,6728|false|false|false|C0562238|Examination of abdomen|abdominal exam
Finding|Functional Concept|Hospital Course|6724,6728|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|Hospital Course|6724,6728|false|false|false|C0582103|Medical Examination|exam
Procedure|Laboratory Procedure|Hospital Course|6731,6734|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6731,6734|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Finding|Intellectual Product|Hospital Course|6744,6752|false|false|false|C4553760|Study Variable|variable
Finding|Intellectual Product|Hospital Course|6775,6781|false|false|false|C1547311|Patient Condition Code - Stable|stable
Disorder|Disease or Syndrome|Hospital Course|6792,6797|false|false|false|C1410088|Still|still
Drug|Biomedical or Dental Material|Hospital Course|6817,6825|false|false|false|C0168634|BaseLine dental cement|baseline
Finding|Idea or Concept|Hospital Course|6817,6825|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Finding|Finding|Hospital Course|6829,6832|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|Hospital Course|6829,6832|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Anatomy|Tissue|Hospital Course|6859,6866|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|Hospital Course|6859,6866|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Pathologic Function|Hospital Course|6859,6876|false|false|false|C0032227|Pleural effusion (disorder)|pleural effusions
Finding|Pathologic Function|Hospital Course|6867,6876|false|false|false|C0013687|effusion|effusions
Anatomy|Tissue|Hospital Course|6902,6909|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|Hospital Course|6902,6909|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Pathologic Function|Hospital Course|6911,6920|false|true|false|C0013687|effusion|effusions
Procedure|Health Care Activity|Hospital Course|6926,6941|false|true|false|C0019993|Hospitalization|hospitalization
Finding|Mental Process|Hospital Course|6945,6952|false|false|false|C0542559|contextual factors|setting
Drug|Substance|Hospital Course|6964,6969|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Hospital Course|6964,6969|false|false|false|C1546638|Fluid Specimen Code|fluid
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6971,6984|false|false|false|C0035273|Resuscitation (procedure)|resuscitation
Finding|Functional Concept|Hospital Course|6986,6991|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Tissue|Hospital Course|6992,6999|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|Hospital Course|6992,6999|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Intellectual Product|Hospital Course|7008,7016|false|false|false|C1546572||catheter
Procedure|Health Care Activity|Hospital Course|7031,7040|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Disorder|Disease or Syndrome|Hospital Course|7061,7066|false|false|false|C1410088|Still|still
Finding|Intellectual Product|Hospital Course|7067,7073|false|false|false|C1705102|Volume (publication)|volume
Finding|Functional Concept|Hospital Course|7088,7092|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|Hospital Course|7088,7092|false|false|false|C0582103|Medical Examination|exam
Drug|Organic Chemical|Hospital Course|7103,7109|false|false|false|C0074722|sodium bicarbonate|bicarb
Drug|Pharmacologic Substance|Hospital Course|7103,7109|false|false|false|C0074722|sodium bicarbonate|bicarb
Finding|Organ or Tissue Function|Hospital Course|7164,7172|false|false|false|C0012797|Diuresis|diuresis
Drug|Organic Chemical|Hospital Course|7188,7194|false|false|false|C0074722|sodium bicarbonate|bicarb
Drug|Pharmacologic Substance|Hospital Course|7188,7194|false|false|false|C0074722|sodium bicarbonate|bicarb
Finding|Functional Concept|Hospital Course|7216,7219|false|false|false|C0678226;C3146286|Due;Due to|due
Finding|Idea or Concept|Hospital Course|7216,7219|false|false|false|C0678226;C3146286|Due;Due to|due
Finding|Mental Process|Hospital Course|7224,7236|false|false|false|C0152057;C0152058|Compensation (Defense Mechanism);Compensation as a General Biological Function|compensation
Finding|Physiologic Function|Hospital Course|7224,7236|false|false|false|C0152057;C0152058|Compensation (Defense Mechanism);Compensation as a General Biological Function|compensation
Attribute|Clinical Attribute|Hospital Course|7246,7257|false|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|Hospital Course|7246,7257|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|Hospital Course|7246,7257|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|Hospital Course|7246,7257|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Disorder|Disease or Syndrome|Hospital Course|7246,7266|false|false|false|C0001127|Acidosis, Respiratory|respiratory acidosis
Finding|Pathologic Function|Hospital Course|7258,7266|false|false|false|C0001122|Acidosis|acidosis
Finding|Intellectual Product|Hospital Course|7271,7277|false|false|false|C1705102|Volume (publication)|Volume
Finding|Pathologic Function|Hospital Course|7271,7286|false|false|false|C0546817|Hypervolemia (finding)|Volume overload
Attribute|Clinical Attribute|Hospital Course|7301,7310|false|false|false|C0012000|Diastole|diastolic
Finding|Pathologic Function|Hospital Course|7301,7322|false|false|false|C0520863|Diastolic dysfunction|diastolic dysfunction
Disorder|Disease or Syndrome|Hospital Course|7311,7322|false|false|false|C3887505|DYSFUNCTION - SKIN DISORDERS|dysfunction
Finding|Conceptual Entity|Hospital Course|7311,7322|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Functional Concept|Hospital Course|7311,7322|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Pathologic Function|Hospital Course|7311,7322|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Anatomy|Fully Formed Anatomical Structure|Hospital Course|7370,7380|false|false|false|C0229960||total body
Anatomy|Anatomical Structure|Hospital Course|7376,7380|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7376,7380|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Finding|Intellectual Product|Hospital Course|7376,7380|false|false|false|C1551342|Document Body|body
Finding|Finding|Hospital Course|7393,7399|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Hospital Course|7393,7399|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Mental Process|Hospital Course|7404,7411|false|false|false|C0542559|contextual factors|setting
Finding|Intellectual Product|Hospital Course|7415,7421|false|false|false|C1705102|Volume (publication)|volume
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7422,7435|false|false|false|C0035273|Resuscitation (procedure)|resuscitation
Procedure|Health Care Activity|Hospital Course|7445,7454|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Disorder|Disease or Syndrome|Hospital Course|7460,7466|false|false|false|C0036690;C0243026|Sepsis;Septicemia|sepsis
Finding|Pathologic Function|Hospital Course|7477,7488|false|false|false|C1140999|Contraction (finding)|contraction
Finding|Pathologic Function|Hospital Course|7477,7498|false|false|false|C1737236|Contraction alkalosis|contraction alkalosis
Disorder|Disease or Syndrome|Hospital Course|7489,7498|false|false|false|C0002063|Alkalosis|alkalosis
Finding|Organ or Tissue Function|Hospital Course|7522,7530|false|false|false|C0012797|Diuresis|diuresis
Finding|Idea or Concept|Hospital Course|7543,7548|false|false|false|C1552828|Table Frame - above|above
Finding|Organ or Tissue Function|Hospital Course|7568,7576|false|false|false|C0012797|Diuresis|diuresis
Finding|Intellectual Product|Hospital Course|7577,7581|false|false|false|C1720092|Once - dosing instruction fragment|once
Finding|Finding|Hospital Course|7583,7594|false|false|false|C0020440|Hypercapnia|hypercarbia
Drug|Organic Chemical|Hospital Course|7608,7614|false|false|false|C0074722|sodium bicarbonate|bicarb
Drug|Pharmacologic Substance|Hospital Course|7608,7614|false|false|false|C0074722|sodium bicarbonate|bicarb
Disorder|Disease or Syndrome|Hospital Course|7633,7647|false|false|false|C0020676|Hypothyroidism|Hypothyroidism
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7662,7675|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Hormone|Hospital Course|7662,7675|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Organic Chemical|Hospital Course|7662,7675|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Pharmacologic Substance|Hospital Course|7662,7675|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Disorder|Disease or Syndrome|Hospital Course|7694,7706|false|false|false|C0020538|Hypertensive disease|Hypertension
Finding|Body Substance|Hospital Course|7708,7715|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|7708,7715|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|7708,7715|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7734,7744|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|Hospital Course|7734,7744|false|false|false|C0065374|lisinopril|lisinopril
Procedure|Health Care Activity|Hospital Course|7772,7781|false|true|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Mental Process|Hospital Course|7785,7792|false|false|false|C0542559|contextual factors|setting
Disorder|Disease or Syndrome|Hospital Course|7796,7802|false|false|false|C0036690;C0243026|Sepsis;Septicemia|sepsis
Attribute|Clinical Attribute|Hospital Course|7807,7815|false|false|false|C3172260||relative
Finding|Idea or Concept|Hospital Course|7807,7815|false|false|false|C1546849|Living Arrangement - Relative|relative
Finding|Finding|Hospital Course|7817,7828|false|false|false|C0020649|Hypotension|hypotension
Disorder|Disease or Syndrome|Hospital Course|7860,7864|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Finding|Body Substance|Hospital Course|7866,7873|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|7866,7873|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|7866,7873|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Organic Chemical|Hospital Course|7888,7898|false|false|false|C0028978|omeprazole|omeprazole
Drug|Pharmacologic Substance|Hospital Course|7888,7898|false|false|false|C0028978|omeprazole|omeprazole
Procedure|Health Care Activity|Hospital Course|7904,7919|false|false|false|C0019993|Hospitalization|hospitalization
Disorder|Cell or Molecular Dysfunction|Hospital Course|7964,7972|false|false|false|C4727483|BRAF Gene Rearrangement|positive
Finding|Classification|Hospital Course|7964,7972|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|Hospital Course|7964,7972|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Drug|Pharmacologic Substance|Hospital Course|8003,8013|false|false|false|C0019593|Histamine H2 Antagonists|H2 blocker
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8021,8032|false|false|false|C0199176|Prophylactic treatment|prophylaxis
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8077,8086|false|false|false|C0011206|Delirium|delirious
Procedure|Health Care Activity|Hospital Course|8092,8107|false|false|false|C0019993|Hospitalization|hospitalization
Drug|Pharmacologic Substance|Hospital Course|8127,8137|false|false|false|C0019593|Histamine H2 Antagonists|H2 blocker
Finding|Body Substance|Hospital Course|8141,8150|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|8141,8150|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|8141,8150|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|8141,8150|false|false|false|C0030685|Patient Discharge|discharge
Finding|Idea or Concept|Hospital Course|8162,8169|false|false|false|C2699424|Concern|concern
Disorder|Disease or Syndrome|Hospital Course|8206,8209|false|false|false|C1860224|ABLEPHARON-MACROSTOMIA SYNDROME|AMS
Finding|Gene or Genome|Hospital Course|8206,8209|false|false|false|C4284022|TWIST2 wt Allele|AMS
Procedure|Laboratory Procedure|Hospital Course|8206,8209|false|false|false|C4521393|Accelerator Mass Spectrometry|AMS
Event|Occupational Activity|Hospital Course|8214,8218|false|false|false|C0009219|Coding|Code
Finding|Intellectual Product|Hospital Course|8214,8218|false|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|Code
Procedure|Health Care Activity|Hospital Course|8214,8225|false|false|false|C0742531|CODE STATUS|Code status
Attribute|Clinical Attribute|Hospital Course|8219,8225|false|false|false|C5889824||status
Finding|Idea or Concept|Hospital Course|8219,8225|false|false|false|C1546481|What subject filter - Status|status
Procedure|Health Care Activity|Hospital Course|8231,8240|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Idea or Concept|Hospital Course|8250,8262|false|false|false|C1548597|Marketing basis - Transitional|Transitional
Finding|Body Substance|Hospital Course|8323,8332|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|8323,8332|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|8323,8332|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|8323,8332|false|false|false|C0030685|Patient Discharge|discharge
Finding|Finding|Hospital Course|8369,8375|false|false|false|C1299582|Unable|unable
Finding|Finding|Hospital Course|8369,8383|false|false|false|C4068785|Unable to void|unable to void
Finding|Intellectual Product|Hospital Course|8379,8383|false|false|false|C0042034;C1552835|Urination;Void - TableFrame|void
Finding|Organism Function|Hospital Course|8379,8383|false|false|false|C0042034;C1552835|Urination;Void - TableFrame|void
Finding|Organ or Tissue Function|Hospital Course|8399,8407|false|false|false|C0012797|Diuresis|diuresis
Drug|Organic Chemical|Hospital Course|8413,8419|false|false|false|C0074722|sodium bicarbonate|bicarb
Drug|Pharmacologic Substance|Hospital Course|8413,8419|false|false|false|C0074722|sodium bicarbonate|bicarb
Finding|Idea or Concept|Hospital Course|8433,8441|false|false|false|C0549178|Continuous|Continue
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8445,8450|false|false|false|C0042313|vancomycin|vanco
Drug|Antibiotic|Hospital Course|8445,8450|false|false|false|C0042313|vancomycin|vanco
Procedure|Laboratory Procedure|Hospital Course|8488,8491|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8488,8491|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Finding|Functional Concept|Hospital Course|8504,8513|false|false|false|C0333618|melanotic|melanotic
Attribute|Clinical Attribute|Hospital Course|8514,8520|false|false|false|C0489144||stools
Finding|Body Substance|Hospital Course|8514,8520|false|false|false|C0015733|Feces|stools
Anatomy|Cell Component|Hospital Course|8563,8570|false|false|false|C1660780|midline cell component|Midline
Finding|Intellectual Product|Hospital Course|8592,8600|false|false|false|C1546572||catheter
Procedure|Health Care Activity|Hospital Course|8614,8623|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Idea or Concept|Hospital Course|8629,8636|false|false|false|C1691786;C1704475|Pending - Allergy Clinical Status;Pending - referral status|pending
Finding|Intellectual Product|Hospital Course|8642,8650|false|false|false|C1546572||catheter
Drug|Substance|Hospital Course|8642,8654|false|false|false|C1292474|Catheter tip specimen|catheter tip
Finding|Intellectual Product|Hospital Course|8642,8654|false|false|false|C1546587|Catheter tip specimen code|catheter tip
Finding|Gene or Genome|Hospital Course|8651,8654|false|false|false|C1705504;C1823282;C1825626;C1825978|ITFG1 gene;KAT5 wt Allele;METTL8 gene;TIPRL gene|tip
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8651,8654|false|false|false|C0673828|TIP regimen|tip
Attribute|Clinical Attribute|Hospital Course|8660,8671|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|8660,8671|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|Hospital Course|8660,8671|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|8660,8684|false|false|false|C1627937|Medications on admission|Medications on Admission
Procedure|Health Care Activity|Hospital Course|8675,8684|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|Hospital Course|8686,8697|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|8686,8697|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|Hospital Course|8686,8697|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Hospital Course|8706,8717|false|false|false|C0082607|fluticasone|fluticasone
Drug|Pharmacologic Substance|Hospital Course|8706,8717|false|false|false|C0082607|fluticasone|fluticasone
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8725,8730|false|false|false|C0028429||nasal
Drug|Biomedical or Dental Material|Hospital Course|8725,8730|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Organic Chemical|Hospital Course|8725,8730|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Pharmacologic Substance|Hospital Course|8725,8730|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Finding|Finding|Hospital Course|8725,8730|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Functional Concept|Hospital Course|8725,8730|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Drug|Pharmacologic Substance|Hospital Course|8725,8736|false|false|false|C2608294|Nasal Spray brand of phenylephrine|nasal spray
Drug|Biomedical or Dental Material|Hospital Course|8731,8736|false|false|false|C1154182|Spray Dosage Form|spray
Event|Activity|Hospital Course|8731,8736|false|false|false|C2003858|Spray (action)|spray
Finding|Functional Concept|Hospital Course|8731,8736|false|false|false|C4521772|Spray (administration method)|spray
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8747,8750|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8747,8750|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|8747,8750|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|8747,8750|false|false|false|C1332410|BID gene|BID
Finding|Gene or Genome|Hospital Course|8751,8754|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8756,8769|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Hormone|Hospital Course|8756,8769|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Organic Chemical|Hospital Course|8756,8769|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Pharmacologic Substance|Hospital Course|8756,8769|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Organic Chemical|Hospital Course|8783,8796|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Drug|Pharmacologic Substance|Hospital Course|8783,8796|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Procedure|Laboratory Procedure|Hospital Course|8783,8796|false|false|false|C0373527|Acetaminophen measurement|acetaminophen
Finding|Gene or Genome|Hospital Course|8808,8811|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|8812,8816|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|8812,8816|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|8812,8816|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Biomedical or Dental Material|Hospital Course|8817,8826|false|false|false|C0032629|Polyvinyls|polyvinyl
Drug|Organic Chemical|Hospital Course|8817,8826|false|false|false|C0032629|Polyvinyls|polyvinyl
Drug|Biomedical or Dental Material|Hospital Course|8817,8834|false|false|false|C0032623|polyvinyl alcohol|polyvinyl alcohol
Drug|Organic Chemical|Hospital Course|8827,8834|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Drug|Pharmacologic Substance|Hospital Course|8827,8834|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Finding|Intellectual Product|Hospital Course|8827,8834|false|false|false|C1547288|Alcohol - Recreational Drug Use Code|alcohol
Drug|Biomedical or Dental Material|Hospital Course|8840,8845|false|false|false|C0991568|Drops - Drug Form|drops
Finding|Gene or Genome|Hospital Course|8855,8858|false|false|false|C1422467|CIAO3 gene|PRN
Disorder|Disease or Syndrome|Hospital Course|8859,8867|false|false|false|C0013238;C0022575|Dry Eye Syndromes;Keratoconjunctivitis Sicca|dry eyes
Drug|Pharmacologic Substance|Hospital Course|8859,8867|false|false|false|C0720056|Dry Eyes brand of ocular lubricant|dry eyes
Finding|Sign or Symptom|Hospital Course|8859,8867|false|false|false|C0314719|Dryness of eye|dry eyes
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8863,8867|false|false|false|C0015392|Eye|eyes
Attribute|Clinical Attribute|Hospital Course|8863,8867|false|false|false|C5848506||eyes
Drug|Biologically Active Substance|Hospital Course|8868,8875|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Organic Chemical|Hospital Course|8868,8875|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Pharmacologic Substance|Hospital Course|8868,8875|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Biologically Active Substance|Hospital Course|8876,8880|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Hospital Course|8876,8880|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Substance|Hospital Course|8876,8880|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Finding|Intellectual Product|Hospital Course|8876,8880|false|false|false|C1546701|line source specimen code|line
Attribute|Clinical Attribute|Hospital Course|8876,8886|false|false|false|C4036660||line flush
Finding|Functional Concept|Hospital Course|8881,8886|false|false|false|C0016382;C1696091|Flush - RouteOfAdministration;Flushing|flush
Finding|Sign or Symptom|Hospital Course|8881,8886|false|false|false|C0016382;C1696091|Flush - RouteOfAdministration;Flushing|flush
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8887,8894|false|false|false|C0528249|Humalog|Humalog
Drug|Pharmacologic Substance|Hospital Course|8887,8894|false|false|false|C0528249|Humalog|Humalog
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8895,8902|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|Hospital Course|8895,8902|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|Hospital Course|8895,8902|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Finding|Gene or Genome|Hospital Course|8895,8902|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|Hospital Course|8895,8902|false|false|false|C0202098|Insulin measurement|insulin
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8911,8916|false|false|false|C0222045|Integumentary scale|scale
Event|Activity|Hospital Course|8911,8916|false|false|false|C1947916|Scaling|scale
Finding|Conceptual Entity|Hospital Course|8911,8916|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|scale
Finding|Intellectual Product|Hospital Course|8911,8916|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|scale
Drug|Organic Chemical|Hospital Course|8917,8927|false|false|false|C0025942|miconazole|Miconazole
Drug|Pharmacologic Substance|Hospital Course|8917,8927|false|false|false|C0025942|miconazole|Miconazole
Drug|Organic Chemical|Hospital Course|8917,8935|false|false|false|C0086620|miconazole nitrate|Miconazole nitrate
Drug|Pharmacologic Substance|Hospital Course|8917,8935|false|false|false|C0086620|miconazole nitrate|Miconazole nitrate
Drug|Element, Ion, or Isotope|Hospital Course|8928,8935|false|false|false|C0028125;C0699857;C3848573|Nitrate;Nitrates;nitrate ion|nitrate
Drug|Inorganic Chemical|Hospital Course|8928,8935|false|false|false|C0028125;C0699857;C3848573|Nitrate;Nitrates;nitrate ion|nitrate
Drug|Pharmacologic Substance|Hospital Course|8928,8935|false|false|false|C0028125;C0699857;C3848573|Nitrate;Nitrates;nitrate ion|nitrate
Drug|Biomedical or Dental Material|Hospital Course|8939,8945|false|false|false|C0032861;C1382110|Powder dose form;powder physical state|powder
Drug|Substance|Hospital Course|8939,8945|false|false|false|C0032861;C1382110|Powder dose form;powder physical state|powder
Finding|Functional Concept|Hospital Course|8949,8960|false|false|false|C0870325;C1547755;C1947919;C2347934;C4048755|Application Document;Apply;Computer Application;HL7 Version 2.5 - Application;Regulatory Application|application
Finding|Idea or Concept|Hospital Course|8949,8960|false|false|false|C0870325;C1547755;C1947919;C2347934;C4048755|Application Document;Apply;Computer Application;HL7 Version 2.5 - Application;Regulatory Application|application
Finding|Intellectual Product|Hospital Course|8949,8960|false|false|false|C0870325;C1547755;C1947919;C2347934;C4048755|Application Document;Apply;Computer Application;HL7 Version 2.5 - Application;Regulatory Application|application
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8949,8960|false|false|false|C0185125|Application procedure|application
Finding|Gene or Genome|Hospital Course|8965,8968|false|false|false|C1422467|CIAO3 gene|PRN
Disorder|Disease or Syndrome|Hospital Course|8969,8973|false|false|false|C5779629|Eruption of skin (disorder)|rash
Finding|Pathologic Function|Hospital Course|8969,8973|false|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Sign or Symptom|Hospital Course|8969,8973|false|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Drug|Organic Chemical|Hospital Course|8974,8985|false|false|false|C0061851|ondansetron|ondansetron
Drug|Pharmacologic Substance|Hospital Course|8974,8985|false|false|false|C0061851|ondansetron|ondansetron
Finding|Gene or Genome|Hospital Course|8998,9001|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|9002,9008|false|false|false|C4255480||nausea
Finding|Sign or Symptom|Hospital Course|9002,9008|false|false|false|C0027497|Nausea|nausea
Drug|Organic Chemical|Hospital Course|9009,9019|false|false|false|C0171023|olanzapine|Olanzapine
Drug|Pharmacologic Substance|Hospital Course|9009,9019|false|false|false|C0171023|olanzapine|Olanzapine
Finding|Gene or Genome|Hospital Course|9044,9047|false|false|false|C1422467|CIAO3 gene|PRN
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9048,9055|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Finding|Sign or Symptom|Hospital Course|9048,9055|false|false|false|C0860603|Anxiety symptoms|anxiety
Drug|Pharmacologic Substance|Hospital Course|9056,9064|false|false|false|C1950154|Insomnia homeopathic medication|insomnia
Finding|Sign or Symptom|Hospital Course|9056,9064|false|false|false|C0917801|Sleeplessness|insomnia
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9065,9075|false|false|false|C0042313|vancomycin|Vancomycin
Drug|Antibiotic|Hospital Course|9065,9075|false|false|false|C0042313|vancomycin|Vancomycin
Procedure|Laboratory Procedure|Hospital Course|9065,9075|false|false|false|C0489941|Vancomycin measurement|Vancomycin
Finding|Body Substance|Hospital Course|9110,9119|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|9110,9119|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|9110,9119|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|9110,9119|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|9110,9131|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|9120,9131|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|9120,9131|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|Hospital Course|9120,9131|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Hospital Course|9136,9147|false|false|false|C0082607|fluticasone|fluticasone
Drug|Pharmacologic Substance|Hospital Course|9136,9147|false|false|false|C0082607|fluticasone|fluticasone
Drug|Biomedical or Dental Material|Hospital Course|9165,9170|false|false|false|C1154182|Spray Dosage Form|Spray
Event|Activity|Hospital Course|9165,9170|false|false|false|C2003858|Spray (action)|Spray
Finding|Functional Concept|Hospital Course|9165,9170|false|false|false|C4521772|Spray (administration method)|Spray
Drug|Biomedical or Dental Material|Hospital Course|9165,9182|false|false|false|C1710170|SPRAY, SUSPENSION|Spray, Suspension
Drug|Biomedical or Dental Material|Hospital Course|9172,9182|false|false|false|C0038960;C1382107|Suspension substance;Suspensions|Suspension
Drug|Substance|Hospital Course|9172,9182|false|false|false|C0038960;C1382107|Suspension substance;Suspensions|Suspension
Finding|Functional Concept|Hospital Course|9172,9182|false|false|false|C1705537|Suspension (action)|Suspension
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9199,9204|false|false|false|C0028429||Nasal
Drug|Biomedical or Dental Material|Hospital Course|9199,9204|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Organic Chemical|Hospital Course|9199,9204|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Pharmacologic Substance|Hospital Course|9199,9204|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Finding|Finding|Hospital Course|9199,9204|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Finding|Functional Concept|Hospital Course|9199,9204|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Finding|Idea or Concept|Hospital Course|9213,9216|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|9213,9216|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Attribute|Clinical Attribute|Hospital Course|9231,9240|false|false|false|C1717415||allergies
Finding|Pathologic Function|Hospital Course|9231,9240|false|false|false|C0020517|Hypersensitivity|allergies
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9247,9260|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Hormone|Hospital Course|9247,9260|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Organic Chemical|Hospital Course|9247,9260|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Pharmacologic Substance|Hospital Course|9247,9260|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Biomedical or Dental Material|Hospital Course|9268,9274|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|9288,9294|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Organic Chemical|Hospital Course|9319,9332|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Drug|Pharmacologic Substance|Hospital Course|9319,9332|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Procedure|Laboratory Procedure|Hospital Course|9319,9332|false|false|false|C0373527|Acetaminophen measurement|acetaminophen
Drug|Biomedical or Dental Material|Hospital Course|9340,9346|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|9356,9363|false|false|false|C0039225|Tablet Dosage Form|Tablets
Finding|Finding|Hospital Course|9403,9408|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|Hospital Course|9403,9408|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Attribute|Clinical Attribute|Hospital Course|9412,9416|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|9412,9416|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|9412,9416|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Biomedical or Dental Material|Hospital Course|9423,9432|false|false|false|C0032629|Polyvinyls|polyvinyl
Drug|Organic Chemical|Hospital Course|9423,9432|false|false|false|C0032629|Polyvinyls|polyvinyl
Drug|Biomedical or Dental Material|Hospital Course|9423,9440|false|false|false|C0032623|polyvinyl alcohol|polyvinyl alcohol
Drug|Organic Chemical|Hospital Course|9433,9440|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Drug|Pharmacologic Substance|Hospital Course|9433,9440|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Finding|Intellectual Product|Hospital Course|9433,9440|false|false|false|C1547288|Alcohol - Recreational Drug Use Code|alcohol
Drug|Biomedical or Dental Material|Hospital Course|9447,9452|false|false|false|C0991568|Drops - Drug Form|Drops
Drug|Biomedical or Dental Material|Hospital Course|9466,9470|false|false|false|C0991568|Drops - Drug Form|drop
Event|Activity|Hospital Course|9466,9470|false|false|false|C1705648|Dropping|drop
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9471,9481|false|false|false|C0015392|Eye|Ophthalmic
Drug|Biomedical or Dental Material|Hospital Course|9471,9481|false|false|false|C2347396|Ophthalmic Dosage Form|Ophthalmic
Finding|Functional Concept|Hospital Course|9471,9481|false|false|false|C1522230|Ophthalmic Route of Administration|Ophthalmic
Disorder|Disease or Syndrome|Hospital Course|9518,9526|false|false|false|C0013238;C0022575|Dry Eye Syndromes;Keratoconjunctivitis Sicca|dry eyes
Drug|Pharmacologic Substance|Hospital Course|9518,9526|false|false|false|C0720056|Dry Eyes brand of ocular lubricant|dry eyes
Finding|Sign or Symptom|Hospital Course|9518,9526|false|false|false|C0314719|Dryness of eye|dry eyes
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9522,9526|false|false|false|C0015392|Eye|eyes
Attribute|Clinical Attribute|Hospital Course|9522,9526|false|false|false|C5848506||eyes
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9533,9540|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|Hospital Course|9533,9540|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|Hospital Course|9533,9540|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Finding|Gene or Genome|Hospital Course|9533,9540|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|Hospital Course|9533,9540|false|false|false|C0202098|Insulin measurement|insulin
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9533,9547|false|false|false|C0293359|insulin lispro|insulin lispro
Drug|Hormone|Hospital Course|9533,9547|false|false|false|C0293359|insulin lispro|insulin lispro
Drug|Pharmacologic Substance|Hospital Course|9533,9547|false|false|false|C0293359|insulin lispro|insulin lispro
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9541,9547|false|false|false|C0293359|insulin lispro|lispro
Drug|Hormone|Hospital Course|9541,9547|false|false|false|C0293359|insulin lispro|lispro
Drug|Pharmacologic Substance|Hospital Course|9541,9547|false|false|false|C0293359|insulin lispro|lispro
Drug|Biomedical or Dental Material|Hospital Course|9560,9568|false|false|false|C0037633;C0525069;C1382100|Pharmaceutical Solutions;Solution Dosage Form;Solutions|Solution
Drug|Substance|Hospital Course|9560,9568|false|false|false|C0037633;C0525069;C1382100|Pharmaceutical Solutions;Solution Dosage Form;Solutions|Solution
Finding|Conceptual Entity|Hospital Course|9560,9568|false|false|false|C2699488|Resolution|Solution
Finding|Functional Concept|Hospital Course|9574,9581|false|false|false|C0332246|Sliding|Sliding
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9574,9587|false|false|false|C2937251|sliding scale|Sliding scale
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9582,9587|false|false|false|C0222045|Integumentary scale|scale
Event|Activity|Hospital Course|9582,9587|false|false|false|C1947916|Scaling|scale
Finding|Conceptual Entity|Hospital Course|9582,9587|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|scale
Finding|Intellectual Product|Hospital Course|9582,9587|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|scale
Finding|Functional Concept|Hospital Course|9595,9607|false|false|false|C1522438|Subcutaneous Route of Administration|Subcutaneous
Disorder|Disease or Syndrome|Hospital Course|9614,9619|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|Hospital Course|9622,9625|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|9622,9625|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Functional Concept|Hospital Course|9749,9753|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|call
Finding|Gene or Genome|Hospital Course|9749,9753|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|call
Finding|Intellectual Product|Hospital Course|9749,9753|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|call
Finding|Mental Process|Hospital Course|9749,9753|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|call
Drug|Organic Chemical|Hospital Course|9763,9773|false|false|false|C0025942|miconazole|miconazole
Drug|Pharmacologic Substance|Hospital Course|9763,9773|false|false|false|C0025942|miconazole|miconazole
Drug|Organic Chemical|Hospital Course|9763,9781|false|false|false|C0086620|miconazole nitrate|miconazole nitrate
Drug|Pharmacologic Substance|Hospital Course|9763,9781|false|false|false|C0086620|miconazole nitrate|miconazole nitrate
Drug|Element, Ion, or Isotope|Hospital Course|9774,9781|false|false|false|C0028125;C0699857;C3848573|Nitrate;Nitrates;nitrate ion|nitrate
Drug|Inorganic Chemical|Hospital Course|9774,9781|false|false|false|C0028125;C0699857;C3848573|Nitrate;Nitrates;nitrate ion|nitrate
Drug|Pharmacologic Substance|Hospital Course|9774,9781|false|false|false|C0028125;C0699857;C3848573|Nitrate;Nitrates;nitrate ion|nitrate
Drug|Biomedical or Dental Material|Hospital Course|9786,9792|false|false|false|C0032861;C1382110|Powder dose form;powder physical state|Powder
Drug|Substance|Hospital Course|9786,9792|false|false|false|C0032861;C1382110|Powder dose form;powder physical state|Powder
Finding|Functional Concept|Hospital Course|9806,9817|false|false|false|C0870325;C1547755;C1947919;C2347934;C4048755|Application Document;Apply;Computer Application;HL7 Version 2.5 - Application;Regulatory Application|application
Finding|Idea or Concept|Hospital Course|9806,9817|false|false|false|C0870325;C1547755;C1947919;C2347934;C4048755|Application Document;Apply;Computer Application;HL7 Version 2.5 - Application;Regulatory Application|application
Finding|Intellectual Product|Hospital Course|9806,9817|false|false|false|C0870325;C1547755;C1947919;C2347934;C4048755|Application Document;Apply;Computer Application;HL7 Version 2.5 - Application;Regulatory Application|application
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9806,9817|false|false|false|C0185125|Application procedure|application
Drug|Biomedical or Dental Material|Hospital Course|9819,9826|false|false|false|C1710439|Topical Dosage Form|Topical
Finding|Functional Concept|Hospital Course|9819,9826|false|false|false|C1522168|Topical Route of Administration|Topical
Disorder|Disease or Syndrome|Hospital Course|9833,9838|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|Hospital Course|9841,9844|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|9841,9844|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Disorder|Disease or Syndrome|Hospital Course|9859,9863|false|false|false|C5779629|Eruption of skin (disorder)|rash
Finding|Pathologic Function|Hospital Course|9859,9863|false|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Sign or Symptom|Hospital Course|9859,9863|false|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9870,9880|false|false|false|C0042313|vancomycin|vancomycin
Drug|Antibiotic|Hospital Course|9870,9880|false|false|false|C0042313|vancomycin|vancomycin
Procedure|Laboratory Procedure|Hospital Course|9870,9880|false|false|false|C0489941|Vancomycin measurement|vancomycin
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9888,9895|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|9888,9895|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|9888,9895|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9909,9916|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|9909,9916|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|9909,9916|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Finding|Intellectual Product|Hospital Course|9925,9930|false|false|false|C1720374|Every - dosing instruction fragment|every
Drug|Biologically Active Substance|Hospital Course|9976,9983|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Organic Chemical|Hospital Course|9976,9983|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Pharmacologic Substance|Hospital Course|9976,9983|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Biologically Active Substance|Hospital Course|9976,9993|false|false|false|C0770546|heparin, porcine|heparin (porcine)
Drug|Organic Chemical|Hospital Course|9976,9993|false|false|false|C0770546|heparin, porcine|heparin (porcine)
Drug|Pharmacologic Substance|Hospital Course|9976,9993|false|false|false|C0770546|heparin, porcine|heparin (porcine)
Finding|Finding|Hospital Course|9985,9992|false|false|false|C4554819|Porcine prosthetic valve|porcine
Drug|Biomedical or Dental Material|Hospital Course|10008,10016|false|false|false|C0037633;C0525069;C1382100|Pharmaceutical Solutions;Solution Dosage Form;Solutions|Solution
Drug|Substance|Hospital Course|10008,10016|false|false|false|C0037633;C0525069;C1382100|Pharmaceutical Solutions;Solution Dosage Form;Solutions|Solution
Finding|Conceptual Entity|Hospital Course|10008,10016|false|false|false|C2699488|Resolution|Solution
Drug|Biomedical or Dental Material|Hospital Course|10041,10050|false|false|false|C1272883|Injection|Injection
Finding|Functional Concept|Hospital Course|10041,10050|false|false|false|C1828121|Injection Route of Administration|Injection
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10041,10050|false|false|false|C0021485;C1533685|Injection of therapeutic agent;Injection procedure|Injection
Disorder|Disease or Syndrome|Hospital Course|10057,10062|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|Hospital Course|10065,10068|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|10065,10068|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|Hospital Course|10075,10084|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|Hospital Course|10075,10084|false|false|false|C0001927|albuterol|albuterol
Drug|Organic Chemical|Hospital Course|10075,10092|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Pharmacologic Substance|Hospital Course|10075,10092|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Element, Ion, or Isotope|Hospital Course|10085,10092|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Inorganic Chemical|Hospital Course|10085,10092|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Pharmacologic Substance|Hospital Course|10085,10092|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Biomedical or Dental Material|Hospital Course|10116,10124|false|false|false|C0037633;C0525069;C1382100|Pharmaceutical Solutions;Solution Dosage Form;Solutions|Solution
Drug|Substance|Hospital Course|10116,10124|false|false|false|C0037633;C0525069;C1382100|Pharmaceutical Solutions;Solution Dosage Form;Solutions|Solution
Finding|Conceptual Entity|Hospital Course|10116,10124|false|false|false|C2699488|Resolution|Solution
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10130,10142|false|false|false|C1659427|nebulization-mediated drug administration|Nebulization
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10156,10159|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|neb
Drug|Biologically Active Substance|Hospital Course|10156,10159|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|neb
Drug|Biomedical or Dental Material|Hospital Course|10156,10159|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|neb
Finding|Cell Function|Hospital Course|10156,10159|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|neb
Finding|Gene or Genome|Hospital Course|10156,10159|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|neb
Finding|Functional Concept|Hospital Course|10160,10170|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Finding|Organism Function|Hospital Course|10160,10170|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Attribute|Clinical Attribute|Hospital Course|10207,10226|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|Hospital Course|10207,10226|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|Hospital Course|10220,10226|false|false|false|C0225386|Breath|breath
Finding|Sign or Symptom|Hospital Course|10230,10238|false|false|false|C0043144|Wheezing|wheezing
Drug|Organic Chemical|Hospital Course|10246,10257|false|false|false|C0027235|ipratropium|ipratropium
Drug|Pharmacologic Substance|Hospital Course|10246,10257|false|false|false|C0027235|ipratropium|ipratropium
Drug|Organic Chemical|Hospital Course|10246,10265|false|false|false|C0700580|ipratropium bromide|ipratropium bromide
Drug|Pharmacologic Substance|Hospital Course|10246,10265|false|false|false|C0700580|ipratropium bromide|ipratropium bromide
Drug|Inorganic Chemical|Hospital Course|10258,10265|false|false|false|C0006222|Bromides|bromide
Procedure|Laboratory Procedure|Hospital Course|10258,10265|false|false|false|C0202341|Bromides measurement|bromide
Drug|Biomedical or Dental Material|Hospital Course|10273,10281|false|false|false|C0037633;C0525069;C1382100|Pharmaceutical Solutions;Solution Dosage Form;Solutions|Solution
Drug|Substance|Hospital Course|10273,10281|false|false|false|C0037633;C0525069;C1382100|Pharmaceutical Solutions;Solution Dosage Form;Solutions|Solution
Finding|Conceptual Entity|Hospital Course|10273,10281|false|false|false|C2699488|Resolution|Solution
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10295,10298|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|neb
Drug|Biologically Active Substance|Hospital Course|10295,10298|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|neb
Drug|Biomedical or Dental Material|Hospital Course|10295,10298|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|neb
Finding|Cell Function|Hospital Course|10295,10298|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|neb
Finding|Gene or Genome|Hospital Course|10295,10298|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|neb
Finding|Functional Concept|Hospital Course|10300,10310|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Finding|Organism Function|Hospital Course|10300,10310|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Attribute|Clinical Attribute|Hospital Course|10345,10364|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|Hospital Course|10345,10364|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|Hospital Course|10358,10364|false|false|false|C0225386|Breath|breath
Finding|Sign or Symptom|Hospital Course|10369,10377|false|false|false|C0043144|Wheezing|wheezing
Finding|Body Substance|Hospital Course|10384,10393|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|10384,10393|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|10384,10393|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|10384,10393|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|10384,10405|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|10384,10405|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|10394,10405|false|false|false|C2926604||Disposition
Procedure|Health Care Activity|Hospital Course|10394,10405|false|false|false|C0184758|Patient disposition|Disposition
Finding|Finding|Hospital Course|10407,10415|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|10407,10415|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Procedure|Health Care Activity|Hospital Course|10407,10420|false|false|false|C0023977|long-term care|Extended Care
Event|Activity|Hospital Course|10416,10420|false|false|false|C1947933|care activity|Care
Finding|Finding|Hospital Course|10416,10420|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|Hospital Course|10416,10420|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|Hospital Course|10423,10431|false|false|false|C4695111|ADMIN.FACILITY|Facility
Finding|Body Substance|Hospital Course|10439,10448|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|10439,10448|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|10439,10448|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|10439,10448|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|10439,10458|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|10449,10458|false|false|false|C0945731||Diagnosis
Finding|Classification|Hospital Course|10449,10458|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|10449,10458|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|10449,10458|false|false|false|C0011900|Diagnosis|Diagnosis
Finding|Mental Process|Principle Diagnosis|10487,10493|false|false|false|C0229992|Psyche structure|mental
Attribute|Clinical Attribute|Principle Diagnosis|10487,10500|false|false|false|C0488568;C0488569||mental status
Finding|Finding|Principle Diagnosis|10487,10500|false|false|false|C0278060|Mental state|mental status
Attribute|Clinical Attribute|Principle Diagnosis|10494,10500|false|false|false|C5889824||status
Finding|Idea or Concept|Principle Diagnosis|10494,10500|false|false|false|C1546481|What subject filter - Status|status
Finding|Finding|Principle Diagnosis|10501,10508|false|false|false|C0242184;C1963140|Hypoxia;Hypoxia, CTCAE|Hypoxia
Finding|Pathologic Function|Principle Diagnosis|10501,10508|false|false|false|C0242184;C1963140|Hypoxia;Hypoxia, CTCAE|Hypoxia
Disorder|Neoplastic Process|Principle Diagnosis|10510,10519|false|false|false|C0027627|Neoplasm Metastasis|Secondary
Finding|Functional Concept|Principle Diagnosis|10510,10519|false|false|false|C1522484|metastatic qualifier|Secondary
Procedure|Diagnostic Procedure|Principle Diagnosis|10520,10529|false|false|false|C0011900|Diagnosis|diagnoses
Finding|Mental Process|Discharge Condition|10577,10583|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|10577,10590|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|10577,10590|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|10584,10590|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|10584,10590|false|false|false|C1546481|What subject filter - Status|Status
Disorder|Mental or Behavioral Dysfunction|Discharge Condition|10592,10600|false|false|false|C0009676|Confusion|Confused
Finding|Finding|Discharge Condition|10592,10600|false|false|false|C0683369;C1547301|Clouded consciousness;Precaution Code - Confused|Confused
Finding|Intellectual Product|Discharge Condition|10592,10600|false|false|false|C0683369;C1547301|Clouded consciousness;Precaution Code - Confused|Confused
Attribute|Clinical Attribute|Discharge Condition|10614,10636|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|10614,10636|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Finding|Finding|Discharge Condition|10623,10636|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|10623,10636|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Sign or Symptom|Discharge Condition|10638,10647|false|false|false|C0023380|Lethargy|Lethargic
Event|Activity|Discharge Condition|10663,10671|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|10663,10671|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|10663,10671|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|10672,10678|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|10672,10678|false|false|false|C1546481|What subject filter - Status|Status
Disorder|Disease or Syndrome|Discharge Condition|10687,10690|false|false|false|C3159311|BORNHOLM EYE DISEASE|Bed
Finding|Intellectual Product|Discharge Condition|10687,10690|false|false|false|C2346952|Bachelor of Education|Bed
Finding|Social Behavior|Discharge Condition|10696,10706|false|false|false|C0018896|Helping Behavior|assistance
Finding|Finding|Discharge Condition|10720,10730|false|false|false|C2135586;C4321408|Wheelchair Usually Used;has wheelchair at home (history)|wheelchair
Finding|Gene or Genome|Discharge Instructions|10759,10763|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Finding|Intellectual Product|Discharge Instructions|10783,10791|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|Discharge Instructions|10783,10791|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|Discharge Instructions|10799,10803|false|false|false|C1947933|care activity|care
Finding|Finding|Discharge Instructions|10799,10803|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|10799,10803|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|10799,10806|false|false|false|C1555558|care of - AddressPartType|care of
Procedure|Health Care Activity|Discharge Instructions|10823,10832|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Finding|Discharge Instructions|10845,10852|false|false|false|C0242184;C1963140|Hypoxia;Hypoxia, CTCAE|hypoxia
Finding|Pathologic Function|Discharge Instructions|10845,10852|false|false|false|C0242184;C1963140|Hypoxia;Hypoxia, CTCAE|hypoxia
Finding|Finding|Discharge Instructions|10853,10864|false|false|false|C0020440|Hypercapnia|hypercarbia
Finding|Mental Process|Discharge Instructions|10877,10883|false|false|false|C0229992|Psyche structure|mental
Attribute|Clinical Attribute|Discharge Instructions|10877,10890|false|false|false|C0488568;C0488569||mental status
Finding|Finding|Discharge Instructions|10877,10890|false|false|false|C0278060|Mental state|mental status
Attribute|Clinical Attribute|Discharge Instructions|10884,10890|false|false|false|C5889824||status
Finding|Idea or Concept|Discharge Instructions|10884,10890|false|false|false|C1546481|What subject filter - Status|status
Finding|Mental Process|Discharge Instructions|10899,10905|false|false|false|C0229992|Psyche structure|mental
Attribute|Clinical Attribute|Discharge Instructions|10899,10912|false|false|false|C0488568;C0488569||mental status
Finding|Finding|Discharge Instructions|10899,10912|false|false|false|C0278060|Mental state|mental status
Attribute|Clinical Attribute|Discharge Instructions|10906,10912|false|false|false|C5889824||status
Finding|Idea or Concept|Discharge Instructions|10906,10912|false|false|false|C1546481|What subject filter - Status|status
Drug|Organic Chemical|Discharge Instructions|10943,10950|false|false|false|C0527258|Zyprexa|Zyprexa
Drug|Pharmacologic Substance|Discharge Instructions|10943,10950|false|false|false|C0527258|Zyprexa|Zyprexa
Disorder|Disease or Syndrome|Discharge Instructions|10999,11008|false|false|false|C0009450|Communicable Diseases|infection
Finding|Pathologic Function|Discharge Instructions|10999,11008|false|false|false|C3714514|Infection|infection
Finding|Finding|Discharge Instructions|11023,11027|false|false|false|C1299581|Able (qualifier value)|able
Finding|Idea or Concept|Discharge Instructions|11038,11043|false|false|false|C1550016|Remote control command - Clear|clear
Finding|Finding|Discharge Instructions|11044,11050|false|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Finding|Functional Concept|Discharge Instructions|11044,11050|false|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Finding|Intellectual Product|Discharge Instructions|11044,11050|false|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Drug|Antibiotic|Discharge Instructions|11081,11092|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Finding|Idea or Concept|Discharge Instructions|11104,11112|false|true|false|C0010453|Culture (Anthropological)|cultures
Finding|Idea or Concept|Discharge Instructions|11118,11125|false|false|false|C1691786;C1704475|Pending - Allergy Clinical Status;Pending - referral status|pending
Drug|Amino Acid, Peptide, or Protein|Discharge Instructions|11150,11155|false|false|false|C0042313|vancomycin|vanco
Drug|Antibiotic|Discharge Instructions|11150,11155|false|false|false|C0042313|vancomycin|vanco
Finding|Functional Concept|Discharge Instructions|11163,11173|false|false|false|C1524062|Additional|additional
Finding|Functional Concept|Discharge Instructions|11197,11204|false|false|false|C0392747|Changing|changes
Attribute|Clinical Attribute|Discharge Instructions|11223,11234|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|11223,11234|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|Discharge Instructions|11223,11234|false|false|false|C4284232|Medications|medications
Finding|Functional Concept|Discharge Instructions|11236,11242|false|false|false|C0392747|Changing|CHANGE
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|11236,11242|false|false|false|C4319952|Change - procedure|CHANGE
Drug|Amino Acid, Peptide, or Protein|Discharge Instructions|11243,11253|false|false|false|C0042313|vancomycin|vancomycin
Drug|Antibiotic|Discharge Instructions|11243,11253|false|false|false|C0042313|vancomycin|vancomycin
Procedure|Laboratory Procedure|Discharge Instructions|11243,11253|false|false|false|C0489941|Vancomycin measurement|vancomycin
Finding|Functional Concept|Discharge Instructions|11260,11268|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Discharge Instructions|11263,11268|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Discharge Instructions|11263,11268|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Food|Discharge Instructions|11310,11315|false|false|false|C0452588|Start brand of breakfast cereal|START
Finding|Intellectual Product|Discharge Instructions|11310,11315|false|false|false|C1552850|start - HtmlLinkType|START
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|11310,11315|false|false|false|C5447432|Collagen Tile Brachytherapy|START
Drug|Organic Chemical|Discharge Instructions|11316,11325|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|Discharge Instructions|11316,11325|false|false|false|C0001927|albuterol|albuterol
Drug|Amino Acid, Peptide, or Protein|Discharge Instructions|11326,11329|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|neb
Drug|Biologically Active Substance|Discharge Instructions|11326,11329|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|neb
Drug|Biomedical or Dental Material|Discharge Instructions|11326,11329|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|neb
Finding|Cell Function|Discharge Instructions|11326,11329|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|neb
Finding|Gene or Genome|Discharge Instructions|11326,11329|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|neb
Finding|Sign or Symptom|Discharge Instructions|11358,11361|false|false|false|C0013404|Dyspnea|SOB
Finding|Sign or Symptom|Discharge Instructions|11362,11370|false|false|false|C0043144|Wheezing|wheezing
Drug|Food|Discharge Instructions|11371,11376|false|false|false|C0452588|Start brand of breakfast cereal|START
Finding|Intellectual Product|Discharge Instructions|11371,11376|false|false|false|C1552850|start - HtmlLinkType|START
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|11371,11376|false|false|false|C5447432|Collagen Tile Brachytherapy|START
Drug|Organic Chemical|Discharge Instructions|11377,11388|false|false|false|C0027235|ipratropium|ipratropium
Drug|Pharmacologic Substance|Discharge Instructions|11377,11388|false|false|false|C0027235|ipratropium|ipratropium
Drug|Amino Acid, Peptide, or Protein|Discharge Instructions|11389,11392|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|neb
Drug|Biologically Active Substance|Discharge Instructions|11389,11392|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|neb
Drug|Biomedical or Dental Material|Discharge Instructions|11389,11392|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|neb
Finding|Cell Function|Discharge Instructions|11389,11392|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|neb
Finding|Gene or Genome|Discharge Instructions|11389,11392|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|neb
Finding|Sign or Symptom|Discharge Instructions|11421,11424|false|false|false|C0013404|Dyspnea|SOB
Finding|Sign or Symptom|Discharge Instructions|11425,11433|false|false|false|C0043144|Wheezing|wheezing
Drug|Inorganic Chemical|Discharge Instructions|11434,11438|false|false|false|C0723457|Stop brand of fluoride|STOP
Drug|Pharmacologic Substance|Discharge Instructions|11434,11438|false|false|false|C0723457|Stop brand of fluoride|STOP
Event|Activity|Discharge Instructions|11434,11438|false|false|false|C1947925|Stop (Instruction Imperative)|STOP
Finding|Gene or Genome|Discharge Instructions|11434,11438|false|false|false|C1417022|MAP6 gene|STOP
Drug|Organic Chemical|Discharge Instructions|11439,11446|false|false|false|C0527258|Zyprexa|Zyprexa
Drug|Pharmacologic Substance|Discharge Instructions|11439,11446|false|false|false|C0527258|Zyprexa|Zyprexa
Procedure|Health Care Activity|Discharge Instructions|11449,11457|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|11458,11470|false|false|false|C3263700||Instructions
Finding|Intellectual Product|Discharge Instructions|11458,11470|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

