 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|33,37
No|38,40
:|40,41
_|44,45
_|45,46
_|46,47
<EOL>|47,48
<EOL>|49,50
Admission|50,59
Date|60,64
:|64,65
_|67,68
_|68,69
_|69,70
Discharge|84,93
Date|94,98
:|98,99
_|102,103
_|103,104
_|104,105
<EOL>|105,106
<EOL>|107,108
Date|108,112
of|113,115
Birth|116,121
:|121,122
_|124,125
_|125,126
_|126,127
Sex|140,143
:|143,144
F|147,148
<EOL>|148,149
<EOL>|150,151
Service|151,158
:|158,159
MEDICINE|160,168
<EOL>|168,169
<EOL>|170,171
Allergies|171,180
:|180,181
<EOL>|182,183
Percocet|183,191
<EOL>|191,192
<EOL>|193,194
Attending|194,203
:|203,204
_|205,206
_|206,207
_|207,208
.|208,209
<EOL>|209,210
<EOL>|211,212
Chief|212,217
Complaint|218,227
:|227,228
<EOL>|228,229
abdominal|229,238
fullness|239,247
and|248,251
discomfort|252,262
<EOL>|262,263
<EOL>|264,265
Major|265,270
Surgical|271,279
or|280,282
Invasive|283,291
Procedure|292,301
:|301,302
<EOL>|302,303
_|303,304
_|304,305
_|305,306
diagnostic|307,317
paracentesis|318,330
<EOL>|330,331
_|331,332
_|332,333
_|333,334
therapeutic|335,346
paracentesis|347,359
<EOL>|359,360
<EOL>|360,361
<EOL>|362,363
History|363,370
of|371,373
Present|374,381
Illness|382,389
:|389,390
<EOL>|390,391
_|391,392
_|392,393
_|393,394
with|395,399
HIV|400,403
on|404,406
HAART|407,412
,|412,413
COPD|414,418
,|418,419
HCV|420,423
cirrhosis|424,433
complicated|434,445
by|446,448
<EOL>|449,450
ascites|450,457
and|458,461
HE|462,464
admitted|465,473
with|474,478
abdominal|479,488
distention|489,499
and|500,503
pain|504,508
.|508,509
She|510,513
<EOL>|514,515
was|515,518
admitted|519,527
to|528,530
_|531,532
_|532,533
_|533,534
for|535,538
the|539,542
same|543,547
symptoms|548,556
<EOL>|557,558
recently|558,566
and|567,570
had|571,574
3L|575,577
fluid|578,583
removed|584,591
(|592,593
no|593,595
SBP|596,599
)|599,600
three|601,606
days|607,611
ago|612,615
and|616,619
<EOL>|620,621
felt|621,625
better|626,632
.|632,633
Since|634,639
discharge|640,649
,|649,650
her|651,654
abdomen|655,662
has|663,666
become|667,673
<EOL>|674,675
increasingly|675,687
distended|688,697
with|698,702
pain|703,707
.|707,708
This|709,713
feels|714,719
similar|720,727
to|728,730
prior|731,736
<EOL>|737,738
episodes|738,746
of|747,749
ascites|750,757
.|757,758
<EOL>|760,761
Her|761,764
diuretics|765,774
were|775,779
recently|780,788
decreased|789,798
on|799,801
_|802,803
_|803,804
_|804,805
due|806,809
to|810,812
worsening|813,822
<EOL>|823,824
hyponatremia|824,836
128|837,840
and|841,844
hyperkalemia|845,857
5.1|858,861
.|861,862
Patient|863,870
states|871,877
she|878,881
has|882,885
<EOL>|886,887
been|887,891
compliant|892,901
with|902,906
her|907,910
HIV|911,914
and|915,918
diuretic|919,927
medications|928,939
but|940,943
never|944,949
<EOL>|950,951
filled|951,957
out|958,961
the|962,965
lactulose|966,975
prescription|976,988
.|988,989
She|990,993
states|994,1000
she|1001,1004
has|1005,1008
had|1009,1012
<EOL>|1013,1014
_|1014,1015
_|1015,1016
_|1016,1017
BMs|1018,1021
daily|1022,1027
at|1028,1030
home|1031,1035
.|1035,1036
She|1037,1040
has|1041,1044
had|1045,1048
some|1049,1053
visual|1054,1060
hallucinations|1061,1075
<EOL>|1076,1077
and|1077,1080
forgetfulness|1081,1094
.|1094,1095
Her|1096,1099
appetite|1100,1108
has|1109,1112
been|1113,1117
poor|1118,1122
.|1122,1123
<EOL>|1125,1126
In|1126,1128
the|1129,1132
ED|1133,1135
,|1135,1136
initial|1137,1144
vitals|1145,1151
were|1152,1156
98.9|1157,1161
88|1162,1164
116|1165,1168
/|1168,1169
88|1169,1171
18|1172,1174
97|1175,1177
%|1177,1178
RA|1179,1181
.|1181,1182
CBC|1183,1186
<EOL>|1187,1188
near|1188,1192
baseline|1193,1201
,|1201,1202
INR|1203,1206
1.4|1207,1210
,|1210,1211
Na|1212,1214
125|1215,1218
,|1218,1219
Cr|1220,1222
0.6|1223,1226
.|1226,1227
AST|1228,1231
and|1232,1235
ALT|1236,1239
mildly|1240,1246
above|1247,1252
<EOL>|1253,1254
baseline|1254,1262
182|1263,1266
and|1267,1270
126|1271,1274
and|1275,1278
albumin|1279,1286
2.8|1287,1290
.|1290,1291
Diagnostic|1292,1302
para|1303,1307
with|1308,1312
225|1313,1316
<EOL>|1317,1318
WBC|1318,1321
,|1321,1322
7|1323,1324
%|1324,1325
PMN|1326,1329
,|1329,1330
total|1331,1336
protein|1337,1344
0.3|1345,1348
.|1348,1349
UA|1350,1352
with|1353,1357
few|1358,1361
bact|1362,1366
,|1366,1367
6|1368,1369
WBC|1370,1373
,|1373,1374
mod|1375,1378
<EOL>|1379,1380
leuk|1380,1384
,|1384,1385
neg|1386,1389
nitr|1390,1394
,|1394,1395
but|1396,1399
contaminated|1400,1412
with|1413,1417
6|1418,1419
epi|1420,1423
.|1423,1424
CXR|1425,1428
clear|1429,1434
.|1434,1435
RUQ|1436,1439
US|1440,1442
<EOL>|1443,1444
with|1444,1448
no|1449,1451
PV|1452,1454
thrombus|1455,1463
,|1463,1464
moderate|1465,1473
ascites|1474,1481
.|1481,1482
She|1483,1486
was|1487,1490
given|1491,1496
ondansetron|1497,1508
<EOL>|1509,1510
4mg|1510,1513
IV|1514,1516
and|1517,1520
morphine|1521,1529
2.5|1530,1533
mg|1533,1535
IV|1536,1538
x1|1539,1541
in|1542,1544
the|1545,1548
ED|1549,1551
.|1551,1552
<EOL>|1554,1555
On|1555,1557
the|1558,1561
floor|1562,1567
,|1567,1568
she|1569,1572
is|1573,1575
feeling|1576,1583
improved|1584,1592
but|1593,1596
still|1597,1602
has|1603,1606
abdominal|1607,1616
<EOL>|1617,1618
distention|1618,1628
and|1629,1632
discomfort|1633,1643
.|1643,1644
<EOL>|1646,1647
ROS|1647,1650
:|1650,1651
+|1652,1653
Abdominal|1653,1662
distention|1663,1673
and|1674,1677
pain|1678,1682
.|1682,1683
No|1684,1686
black|1687,1692
/|1692,1693
bloody|1693,1699
stools|1700,1706
.|1706,1707
No|1708,1710
<EOL>|1711,1712
_|1712,1713
_|1713,1714
_|1714,1715
pain|1716,1720
or|1721,1723
swelling|1724,1732
.|1732,1733
No|1734,1736
fevers|1737,1743
or|1744,1746
chills|1747,1753
.|1753,1754
Denies|1755,1761
chest|1762,1767
pain|1768,1772
,|1772,1773
<EOL>|1774,1775
nausea|1775,1781
,|1781,1782
vomiting|1783,1791
.|1791,1792
No|1793,1795
dysuria|1796,1803
or|1804,1806
frequency|1807,1816
.|1816,1817
<EOL>|1818,1819
<EOL>|1820,1821
Past|1821,1825
Medical|1826,1833
History|1834,1841
:|1841,1842
<EOL>|1842,1843
1.|1843,1845
HCV|1846,1849
Cirrhosis|1850,1859
<EOL>|1861,1862
2.|1862,1864
No|1865,1867
history|1868,1875
of|1876,1878
abnormal|1879,1887
Pap|1888,1891
smears|1892,1898
.|1898,1899
<EOL>|1901,1902
3.|1902,1904
She|1905,1908
had|1909,1912
calcification|1913,1926
in|1927,1929
her|1930,1933
breast|1934,1940
,|1940,1941
which|1942,1947
was|1948,1951
removed|1952,1959
<EOL>|1961,1962
previously|1962,1972
and|1973,1976
per|1977,1980
patient|1981,1988
not|1989,1992
,|1992,1993
it|1994,1996
was|1997,2000
benign|2001,2007
.|2007,2008
<EOL>|2010,2011
4|2011,2012
.|2012,2013
For|2014,2017
HIV|2018,2021
disease|2022,2029
,|2029,2030
she|2031,2034
is|2035,2037
being|2038,2043
followed|2044,2052
by|2053,2055
Dr.|2056,2059
_|2060,2061
_|2061,2062
_|2062,2063
Dr|2064,2066
.|2066,2067
<EOL>|2069,2070
_|2070,2071
_|2071,2072
_|2072,2073
.|2073,2074
<EOL>|2076,2077
5.|2077,2079
COPD|2080,2084
<EOL>|2086,2087
6.|2087,2089
Past|2090,2094
history|2095,2102
of|2103,2105
smoking|2106,2113
.|2113,2114
<EOL>|2116,2117
7.|2117,2119
She|2120,2123
also|2124,2128
had|2129,2132
a|2133,2134
skin|2135,2139
lesion|2140,2146
,|2146,2147
which|2148,2153
was|2154,2157
biopsied|2158,2166
and|2167,2170
showed|2171,2177
<EOL>|2179,2180
skin|2180,2184
cancer|2185,2191
per|2192,2195
patient|2196,2203
report|2204,2210
and|2211,2214
is|2215,2217
scheduled|2218,2227
for|2228,2231
a|2232,2233
complete|2234,2242
<EOL>|2244,2245
removal|2245,2252
of|2253,2255
the|2256,2259
skin|2260,2264
lesion|2265,2271
in|2272,2274
_|2275,2276
_|2276,2277
_|2277,2278
of|2279,2281
this|2282,2286
year|2287,2291
.|2291,2292
<EOL>|2294,2295
8.|2295,2297
She|2298,2301
also|2302,2306
had|2307,2310
another|2311,2318
lesion|2319,2325
in|2326,2328
her|2329,2332
forehead|2333,2341
with|2342,2346
purple|2347,2353
<EOL>|2355,2356
discoloration|2356,2369
.|2369,2370
It|2371,2373
was|2374,2377
biopsied|2378,2386
to|2387,2389
exclude|2390,2397
the|2398,2401
possibility|2402,2413
of|2414,2416
<EOL>|2418,2419
_|2419,2420
_|2420,2421
_|2421,2422
'|2422,2423
s|2423,2424
sarcoma|2425,2432
,|2432,2433
the|2434,2437
results|2438,2445
is|2446,2448
pending|2449,2456
.|2456,2457
<EOL>|2459,2460
9|2460,2461
.|2461,2462
A|2463,2464
15|2465,2467
mm|2468,2470
hypoechoic|2471,2481
lesion|2482,2488
on|2489,2491
her|2492,2495
ultrasound|2496,2506
on|2507,2509
_|2510,2511
_|2511,2512
_|2512,2513
<EOL>|2515,2516
and|2516,2519
is|2520,2522
being|2523,2528
monitored|2529,2538
by|2539,2541
an|2542,2544
MRI|2545,2548
.|2548,2549
<EOL>|2551,2552
10|2552,2554
.|2554,2555
History|2556,2563
of|2564,2566
dysplasia|2567,2576
of|2577,2579
anus|2580,2584
in|2585,2587
_|2588,2589
_|2589,2590
_|2590,2591
.|2591,2592
<EOL>|2594,2595
11|2595,2597
.|2597,2598
Bipolar|2599,2606
affective|2607,2616
disorder|2617,2625
,|2625,2626
currently|2627,2636
manic|2637,2642
,|2642,2643
mild|2644,2648
,|2648,2649
and|2650,2653
PTSD|2654,2658
.|2658,2659
<EOL>|2660,2661
<EOL>|2662,2663
12.|2663,2666
History|2667,2674
of|2675,2677
cocaine|2678,2685
and|2686,2689
heroin|2690,2696
use|2697,2700
.|2700,2701
<EOL>|2703,2704
<EOL>|2704,2705
<EOL>|2706,2707
Social|2707,2713
History|2714,2721
:|2721,2722
<EOL>|2722,2723
_|2723,2724
_|2724,2725
_|2725,2726
<EOL>|2726,2727
Family|2727,2733
History|2734,2741
:|2741,2742
<EOL>|2742,2743
She|2743,2746
a|2747,2748
total|2749,2754
of|2755,2757
five|2758,2762
siblings|2763,2771
,|2771,2772
but|2773,2776
she|2777,2780
is|2781,2783
not|2784,2787
talking|2789,2796
to|2797,2799
most|2800,2804
of|2805,2807
<EOL>|2808,2809
them|2809,2813
.|2813,2814
She|2815,2818
only|2819,2823
has|2824,2827
one|2828,2831
brother|2832,2839
that|2840,2844
she|2845,2848
is|2849,2851
in|2852,2854
touch|2856,2861
with|2862,2866
and|2867,2870
<EOL>|2871,2872
lives|2872,2877
in|2878,2880
_|2881,2882
_|2882,2883
_|2883,2884
.|2884,2885
She|2886,2889
is|2890,2892
not|2893,2896
aware|2897,2902
of|2903,2905
any|2906,2909
known|2910,2915
GI|2916,2918
or|2919,2921
liver|2922,2927
<EOL>|2928,2929
disease|2929,2936
in|2937,2939
her|2940,2943
family|2944,2950
.|2950,2951
<EOL>|2953,2954
<EOL>|2955,2956
Physical|2956,2964
Exam|2965,2969
:|2969,2970
<EOL>|2970,2971
ADMISSION|2971,2980
PHYSICAL|2981,2989
EXAM|2990,2994
:|2994,2995
<EOL>|2997,2998
VS|2998,3000
:|3000,3001
T98|3002,3005
.1|3005,3007
105|3008,3011
/|3011,3012
57|3012,3014
79|3015,3017
20|3018,3020
97RA|3021,3025
44.6|3026,3030
kg|3030,3032
<EOL>|3034,3035
GENERAL|3035,3042
:|3042,3043
Thin|3044,3048
chronically|3049,3060
ill|3061,3064
appearing|3065,3074
woman|3075,3080
in|3081,3083
no|3084,3086
acute|3087,3092
<EOL>|3093,3094
distress|3094,3102
<EOL>|3104,3105
HEENT|3105,3110
:|3110,3111
Sclera|3112,3118
anicteric|3119,3128
,|3128,3129
MMM|3130,3133
,|3133,3134
no|3135,3137
oral|3138,3142
lesions|3143,3150
<EOL>|3152,3153
HEART|3153,3158
:|3158,3159
RRR|3160,3163
,|3163,3164
normal|3165,3171
S1|3172,3174
S2|3175,3177
,|3177,3178
no|3179,3181
murmurs|3182,3189
<EOL>|3191,3192
LUNGS|3192,3197
:|3197,3198
Clear|3199,3204
,|3204,3205
no|3206,3208
wheezes|3209,3216
,|3216,3217
rales|3218,3223
,|3223,3224
or|3225,3227
rhonchi|3228,3235
<EOL>|3237,3238
ABD|3238,3241
:|3241,3242
Significant|3243,3254
distention|3255,3265
with|3266,3270
visible|3271,3278
veins|3279,3284
,|3284,3285
bulging|3286,3293
flanks|3294,3300
,|3300,3301
<EOL>|3302,3303
nontender|3303,3312
to|3313,3315
palpation|3316,3325
,|3325,3326
tympanitic|3327,3337
on|3338,3340
percussion|3341,3351
,|3351,3352
normal|3353,3359
bowel|3360,3365
<EOL>|3366,3367
sounds|3367,3373
<EOL>|3375,3376
EXT|3376,3379
:|3379,3380
no|3381,3383
_|3384,3385
_|3385,3386
_|3386,3387
edema|3388,3393
,|3393,3394
2|3395,3396
+|3396,3397
DP|3398,3400
and|3401,3404
_|3405,3406
_|3406,3407
_|3407,3408
pulses|3409,3415
<EOL>|3417,3418
NEURO|3418,3423
:|3423,3424
alert|3425,3430
and|3431,3434
oriented|3435,3443
,|3443,3444
not|3445,3448
confused|3449,3457
,|3457,3458
no|3459,3461
asterixis|3462,3471
<EOL>|3471,3472
<EOL>|3472,3473
DISCHARGE|3473,3482
PE|3483,3485
:|3485,3486
<EOL>|3486,3487
VS|3487,3489
:|3489,3490
T|3491,3492
98.4|3493,3497
BP|3498,3500
95|3501,3503
/|3503,3504
55|3504,3506
(|3507,3508
SBP|3508,3511
_|3512,3513
_|3513,3514
_|3514,3515
HR|3516,3518
80|3519,3521
RR|3522,3524
18|3525,3527
O2|3528,3530
95RA|3531,3535
<EOL>|3537,3538
I|3538,3539
/|3539,3540
O|3540,3541
240|3542,3545
/|3545,3546
150|3546,3549
this|3550,3554
am|3555,3557
<EOL>|3559,3560
GENERAL|3560,3567
:|3567,3568
Thin|3569,3573
chronically|3574,3585
ill|3586,3589
appearing|3590,3599
woman|3600,3605
in|3606,3608
no|3609,3611
acute|3612,3617
<EOL>|3618,3619
distress|3619,3627
<EOL>|3629,3630
HEENT|3630,3635
:|3635,3636
Sclera|3637,3643
anicteric|3644,3653
,|3653,3654
MMM|3655,3658
,|3658,3659
no|3660,3662
oral|3663,3667
lesions|3668,3675
<EOL>|3677,3678
HEART|3678,3683
:|3683,3684
RRR|3685,3688
,|3688,3689
normal|3690,3696
S1|3697,3699
S2|3700,3702
,|3702,3703
no|3704,3706
murmurs|3707,3714
<EOL>|3716,3717
LUNGS|3717,3722
:|3722,3723
Clear|3724,3729
,|3729,3730
no|3731,3733
wheezes|3734,3741
,|3741,3742
rales|3743,3748
,|3748,3749
or|3750,3752
rhonchi|3753,3760
<EOL>|3762,3763
ABD|3763,3766
:|3766,3767
Significant|3768,3779
distention|3780,3790
with|3791,3795
visible|3796,3803
veins|3804,3809
,|3809,3810
bulging|3811,3818
flanks|3819,3825
,|3825,3826
<EOL>|3827,3828
nontender|3828,3837
to|3838,3840
palpation|3841,3850
,|3850,3851
tympanitic|3852,3862
on|3863,3865
percussion|3866,3876
,|3876,3877
normal|3878,3884
bowel|3885,3890
<EOL>|3891,3892
sounds|3892,3898
<EOL>|3900,3901
EXT|3901,3904
:|3904,3905
no|3906,3908
_|3909,3910
_|3910,3911
_|3911,3912
edema|3913,3918
,|3918,3919
2|3920,3921
+|3921,3922
DP|3923,3925
and|3926,3929
_|3930,3931
_|3931,3932
_|3932,3933
pulses|3934,3940
<EOL>|3942,3943
NEURO|3943,3948
:|3948,3949
alert|3950,3955
and|3956,3959
oriented|3960,3968
,|3968,3969
not|3970,3973
confused|3974,3982
,|3982,3983
no|3984,3986
asterixis|3987,3996
<EOL>|3996,3997
<EOL>|3998,3999
Pertinent|3999,4008
Results|4009,4016
:|4016,4017
<EOL>|4017,4018
LABS|4018,4022
ON|4023,4025
ADMISSION|4026,4035
:|4035,4036
<EOL>|4036,4037
_|4037,4038
_|4038,4039
_|4039,4040
04|4041,4043
:|4043,4044
10PM|4044,4048
BLOOD|4049,4054
_|4055,4056
_|4056,4057
_|4057,4058
<EOL>|4059,4060
_|4060,4061
_|4061,4062
_|4062,4063
Plt|4064,4067
_|4068,4069
_|4069,4070
_|4070,4071
<EOL>|4071,4072
_|4072,4073
_|4073,4074
_|4074,4075
04|4076,4078
:|4078,4079
10PM|4079,4083
BLOOD|4084,4089
_|4090,4091
_|4091,4092
_|4092,4093
<EOL>|4094,4095
_|4095,4096
_|4096,4097
_|4097,4098
<EOL>|4098,4099
_|4099,4100
_|4100,4101
_|4101,4102
04|4103,4105
:|4105,4106
10PM|4106,4110
BLOOD|4111,4116
_|4117,4118
_|4118,4119
_|4119,4120
<EOL>|4121,4122
_|4122,4123
_|4123,4124
_|4124,4125
<EOL>|4125,4126
_|4126,4127
_|4127,4128
_|4128,4129
04|4130,4132
:|4132,4133
10PM|4133,4137
BLOOD|4138,4143
_|4144,4145
_|4145,4146
_|4146,4147
<EOL>|4148,4149
_|4149,4150
_|4150,4151
_|4151,4152
<EOL>|4152,4153
_|4153,4154
_|4154,4155
_|4155,4156
04|4157,4159
:|4159,4160
10PM|4160,4164
BLOOD|4165,4170
_|4171,4172
_|4172,4173
_|4173,4174
<EOL>|4174,4175
_|4175,4176
_|4176,4177
_|4177,4178
04|4179,4181
:|4181,4182
39PM|4182,4186
BLOOD|4187,4192
_|4193,4194
_|4194,4195
_|4195,4196
<EOL>|4196,4197
<EOL>|4197,4198
LABS|4198,4202
ON|4203,4205
DISCHARGE|4206,4215
:|4215,4216
<EOL>|4216,4217
_|4217,4218
_|4218,4219
_|4219,4220
05|4221,4223
:|4223,4224
10AM|4224,4228
BLOOD|4229,4234
_|4235,4236
_|4236,4237
_|4237,4238
<EOL>|4239,4240
_|4240,4241
_|4241,4242
_|4242,4243
Plt|4244,4247
_|4248,4249
_|4249,4250
_|4250,4251
<EOL>|4251,4252
_|4252,4253
_|4253,4254
_|4254,4255
05|4256,4258
:|4258,4259
10AM|4259,4263
BLOOD|4264,4269
_|4270,4271
_|4271,4272
_|4272,4273
_|4274,4275
_|4275,4276
_|4276,4277
<EOL>|4277,4278
_|4278,4279
_|4279,4280
_|4280,4281
05|4282,4284
:|4284,4285
10AM|4285,4289
BLOOD|4290,4295
_|4296,4297
_|4297,4298
_|4298,4299
<EOL>|4300,4301
_|4301,4302
_|4302,4303
_|4303,4304
<EOL>|4304,4305
_|4305,4306
_|4306,4307
_|4307,4308
05|4309,4311
:|4311,4312
10AM|4312,4316
BLOOD|4317,4322
_|4323,4324
_|4324,4325
_|4325,4326
<EOL>|4327,4328
_|4328,4329
_|4329,4330
_|4330,4331
<EOL>|4331,4332
_|4332,4333
_|4333,4334
_|4334,4335
05|4336,4338
:|4338,4339
10AM|4339,4343
BLOOD|4344,4349
_|4350,4351
_|4351,4352
_|4352,4353
<EOL>|4353,4354
<EOL>|4354,4355
MICRO|4355,4360
:|4360,4361
<EOL>|4361,4362
_|4362,4363
_|4363,4364
_|4364,4365
10|4366,4368
:|4368,4369
39|4369,4371
pm|4372,4374
URINE|4375,4380
Source|4386,4392
:|4392,4393
_|4394,4395
_|4395,4396
_|4396,4397
.|4397,4398
<EOL>|4399,4400
<EOL>|4400,4401
*|4429,4430
*|4430,4431
FINAL|4431,4436
REPORT|4437,4443
_|4444,4445
_|4445,4446
_|4446,4447
<EOL>|4447,4448
<EOL>|4448,4449
URINE|4452,4457
CULTURE|4458,4465
(|4466,4467
Final|4467,4472
_|4473,4474
_|4474,4475
_|4475,4476
:|4476,4477
<EOL>|4478,4479
MIXED|4485,4490
BACTERIAL|4491,4500
FLORA|4501,4506
(|4507,4508
>|4509,4510
=|4510,4511
3|4512,4513
COLONY|4514,4520
TYPES|4521,4526
)|4526,4527
,|4527,4528
CONSISTENT|4529,4539
<EOL>|4540,4541
WITH|4541,4545
SKIN|4546,4550
<EOL>|4550,4551
AND|4557,4560
/|4560,4561
OR|4561,4563
GENITAL|4564,4571
CONTAMINATION|4572,4585
.|4585,4586
<EOL>|4587,4588
<EOL>|4588,4589
_|4589,4590
_|4590,4591
_|4591,4592
7|4593,4594
:|4594,4595
00|4595,4597
pm|4598,4600
PERITONEAL|4601,4611
FLUID|4612,4617
PERITONEAL|4623,4633
FLUID|4634,4639
.|4639,4640
<EOL>|4641,4642
<EOL>|4642,4643
GRAM|4646,4650
STAIN|4651,4656
(|4657,4658
Final|4658,4663
_|4664,4665
_|4665,4666
_|4666,4667
:|4667,4668
<EOL>|4669,4670
1|4676,4677
+|4677,4678
(|4682,4683
<|4683,4684
1|4684,4685
per|4686,4689
1000X|4690,4695
FIELD|4696,4701
)|4701,4702
:|4702,4703
POLYMORPHONUCLEAR|4706,4723
<EOL>|4724,4725
LEUKOCYTES|4725,4735
.|4735,4736
<EOL>|4737,4738
NO|4744,4746
MICROORGANISMS|4747,4761
SEEN|4762,4766
.|4766,4767
<EOL>|4768,4769
This|4775,4779
is|4780,4782
a|4783,4784
concentrated|4785,4797
smear|4798,4803
made|4804,4808
by|4809,4811
cytospin|4812,4820
method|4821,4827
,|4827,4828
<EOL>|4829,4830
please|4830,4836
refer|4837,4842
to|4843,4845
<EOL>|4845,4846
hematology|4852,4862
for|4863,4866
a|4867,4868
quantitative|4869,4881
white|4882,4887
blood|4888,4893
cell|4894,4898
count|4899,4904
.|4904,4905
.|4905,4906
<EOL>|4907,4908
<EOL>|4908,4909
FLUID|4912,4917
CULTURE|4918,4925
(|4926,4927
Final|4927,4932
_|4933,4934
_|4934,4935
_|4935,4936
:|4936,4937
NO|4941,4943
GROWTH|4944,4950
.|4950,4951
<EOL>|4952,4953
<EOL>|4953,4954
ANAEROBIC|4957,4966
CULTURE|4967,4974
(|4975,4976
Preliminary|4976,4987
)|4987,4988
:|4988,4989
NO|4993,4995
GROWTH|4996,5002
.|5002,5003
<EOL>|5003,5004
<EOL>|5004,5005
_|5005,5006
_|5006,5007
_|5007,5008
7|5009,5010
:|5010,5011
00|5011,5013
pm|5014,5016
PERITONEAL|5017,5027
FLUID|5028,5033
PERITONEAL|5039,5049
FLUID|5050,5055
.|5055,5056
<EOL>|5057,5058
<EOL>|5058,5059
GRAM|5062,5066
STAIN|5067,5072
(|5073,5074
Final|5074,5079
_|5080,5081
_|5081,5082
_|5082,5083
:|5083,5084
<EOL>|5085,5086
1|5092,5093
+|5093,5094
(|5098,5099
<|5099,5100
1|5100,5101
per|5102,5105
1000X|5106,5111
FIELD|5112,5117
)|5117,5118
:|5118,5119
POLYMORPHONUCLEAR|5122,5139
<EOL>|5140,5141
LEUKOCYTES|5141,5151
.|5151,5152
<EOL>|5153,5154
NO|5160,5162
MICROORGANISMS|5163,5177
SEEN|5178,5182
.|5182,5183
<EOL>|5184,5185
This|5191,5195
is|5196,5198
a|5199,5200
concentrated|5201,5213
smear|5214,5219
made|5220,5224
by|5225,5227
cytospin|5228,5236
method|5237,5243
,|5243,5244
<EOL>|5245,5246
please|5246,5252
refer|5253,5258
to|5259,5261
<EOL>|5261,5262
hematology|5268,5278
for|5279,5282
a|5283,5284
quantitative|5285,5297
white|5298,5303
blood|5304,5309
cell|5310,5314
count|5315,5320
.|5320,5321
.|5321,5322
<EOL>|5323,5324
<EOL>|5324,5325
FLUID|5328,5333
CULTURE|5334,5341
(|5342,5343
Final|5343,5348
_|5349,5350
_|5350,5351
_|5351,5352
:|5352,5353
NO|5357,5359
GROWTH|5360,5366
.|5366,5367
<EOL>|5368,5369
<EOL>|5369,5370
ANAEROBIC|5373,5382
CULTURE|5383,5390
(|5391,5392
Preliminary|5392,5403
)|5403,5404
:|5404,5405
NO|5409,5411
GROWTH|5412,5418
.|5418,5419
<EOL>|5420,5421
<EOL>|5421,5422
Diagnositc|5422,5432
Para|5433,5437
:|5437,5438
<EOL>|5438,5439
_|5439,5440
_|5440,5441
_|5441,5442
07|5443,5445
:|5445,5446
00PM|5446,5450
ASCITES|5451,5458
_|5459,5460
_|5460,5461
_|5461,5462
<EOL>|5463,5464
_|5464,5465
_|5465,5466
_|5466,5467
<EOL>|5467,5468
_|5468,5469
_|5469,5470
_|5470,5471
07|5472,5474
:|5474,5475
00PM|5475,5479
ASCITES|5480,5487
_|5488,5489
_|5489,5490
_|5490,5491
<EOL>|5491,5492
<EOL>|5492,5493
IMAGING|5493,5500
:|5500,5501
<EOL>|5501,5502
_|5502,5503
_|5503,5504
_|5504,5505
CXR|5506,5509
-|5509,5510
No|5511,5513
acute|5514,5519
cardiopulmonary|5520,5535
abnormality|5536,5547
.|5547,5548
<EOL>|5550,5551
_|5551,5552
_|5552,5553
_|5553,5554
RUQ|5555,5558
US|5559,5561
-|5561,5562
<EOL>|5564,5565
1.|5565,5567
Extremely|5568,5577
coarse|5578,5584
and|5585,5588
nodular|5589,5596
liver|5597,5602
echotexture|5603,5614
consistent|5615,5625
<EOL>|5626,5627
with|5627,5631
a|5632,5633
history|5634,5641
of|5642,5644
cirrhosis|5645,5654
.|5654,5655
<EOL>|5657,5658
2.|5658,5660
Moderate|5661,5669
ascites|5670,5677
.|5677,5678
<EOL>|5680,5681
3.|5681,5683
Patent|5684,5690
portal|5691,5697
vein|5698,5702
.|5702,5703
<EOL>|5703,5704
<EOL>|5705,5706
Brief|5706,5711
Hospital|5712,5720
Course|5721,5727
:|5727,5728
<EOL>|5728,5729
_|5729,5730
_|5730,5731
_|5731,5732
with|5733,5737
HIV|5738,5741
on|5742,5744
HAART|5745,5750
,|5750,5751
HCV|5752,5755
cirrhosis|5756,5765
with|5766,5770
ascites|5771,5778
and|5779,5782
HE|5783,5785
,|5785,5786
h|5787,5788
/|5788,5789
o|5789,5790
<EOL>|5791,5792
IVDU|5792,5796
,|5796,5797
COPD|5798,5802
,|5802,5803
bipolar|5804,5811
disorder|5812,5820
presents|5821,5829
with|5830,5834
abdominal|5835,5844
discomfort|5845,5855
<EOL>|5856,5857
due|5857,5860
to|5861,5863
_|5864,5865
_|5865,5866
_|5866,5867
ascites|5868,5875
.|5875,5876
<EOL>|5878,5879
<EOL>|5880,5881
#|5881,5882
ASCITES|5883,5890
.|5890,5891
Now|5892,5895
diuretic|5896,5904
refractory|5905,5915
given|5916,5921
last|5922,5926
tap|5927,5930
was|5931,5934
three|5935,5940
days|5941,5945
<EOL>|5946,5947
ago|5947,5950
with|5951,5955
3L|5956,5958
removed|5959,5966
and|5967,5970
she|5971,5974
has|5975,5978
already|5979,5986
built|5987,5992
up|5993,5995
moderate|5996,6004
<EOL>|6005,6006
ascites|6006,6013
.|6013,6014
Infectious|6015,6025
workup|6026,6032
negative|6033,6041
,|6041,6042
with|6043,6047
CXR|6048,6051
clear|6052,6057
,|6057,6058
UA|6059,6061
<EOL>|6062,6063
contaminated|6063,6075
but|6076,6079
not|6080,6083
grossly|6084,6091
positive|6092,6100
so|6101,6103
will|6104,6108
f|6109,6110
/|6110,6111
u|6111,6112
culture|6113,6120
,|6120,6121
<EOL>|6122,6123
diagnostic|6123,6133
para|6134,6138
with|6139,6143
only|6144,6148
225|6149,6152
WBC|6153,6156
,|6156,6157
RUQ|6158,6161
US|6162,6164
with|6165,6169
no|6170,6172
PV|6173,6175
thrombus|6176,6184
.|6184,6185
<EOL>|6186,6187
Compliant|6187,6196
with|6197,6201
diuretics|6202,6211
but|6212,6215
not|6216,6219
following|6220,6229
low|6230,6233
sodium|6234,6240
diet|6241,6245
or|6246,6248
<EOL>|6249,6250
fluid|6250,6255
restriction|6256,6267
.|6267,6268
Dr.|6269,6272
_|6273,6274
_|6274,6275
_|6275,6276
discussed|6277,6286
possible|6287,6295
TIPS|6296,6300
in|6301,6303
<EOL>|6304,6305
the|6305,6308
office|6309,6315
but|6316,6319
due|6320,6323
to|6324,6326
lung|6327,6331
disease|6332,6339
,|6339,6340
that|6341,6345
was|6346,6349
on|6350,6352
hold|6353,6357
pending|6358,6365
<EOL>|6366,6367
further|6367,6374
cardiac|6375,6382
evaluation|6383,6393
.|6393,6394
Diuretics|6395,6404
were|6405,6409
recently|6410,6418
decreased|6419,6428
<EOL>|6429,6430
due|6430,6433
to|6434,6436
hyponatremia|6437,6449
and|6450,6453
hyperkalemia|6454,6466
.|6466,6467
Held|6468,6472
spironolactone|6473,6487
for|6488,6491
<EOL>|6492,6493
now|6493,6496
due|6497,6500
to|6501,6503
K|6504,6505
5.2|6506,6509
and|6510,6513
increased|6514,6523
lasix|6524,6529
20|6530,6532
-|6533,6534
>|6534,6535
40|6536,6538
.|6538,6539
No|6540,6542
evidence|6543,6551
of|6552,6554
<EOL>|6555,6556
severe|6556,6562
hyponatremia|6563,6575
(|6576,6577
Na|6577,6579
<|6579,6580
120|6580,6583
)|6583,6584
or|6585,6587
renal|6588,6593
failure|6594,6601
Cr|6602,6604
>|6604,6605
2.0|6605,6608
to|6609,6611
stop|6612,6616
<EOL>|6617,6618
diuretics|6618,6627
at|6628,6630
present|6631,6638
.|6638,6639
Diagnostic|6640,6650
paracentesis|6651,6663
negative|6664,6672
for|6673,6676
<EOL>|6677,6678
infection|6678,6687
.|6687,6688
Ascitic|6689,6696
total|6697,6702
protein|6703,6710
0.3|6711,6714
so|6715,6717
warrants|6718,6726
SBP|6727,6730
prophylaxis|6731,6742
<EOL>|6743,6744
(|6744,6745
<|6745,6746
1.0|6746,6749
)|6749,6750
and|6751,6754
fortunately|6755,6766
already|6767,6774
on|6775,6777
Bactrim|6778,6785
for|6786,6789
PCP|6790,6793
prophylaxis|6794,6805
<EOL>|6806,6807
which|6807,6812
would|6813,6818
be|6819,6821
appropriate|6822,6833
for|6834,6837
SBP|6838,6841
ppx|6842,6845
also|6846,6850
.|6850,6851
Patient|6852,6859
did|6860,6863
admit|6864,6869
<EOL>|6870,6871
to|6871,6873
eating|6874,6880
pizza|6881,6886
and|6887,6890
some|6891,6895
_|6896,6897
_|6897,6898
_|6898,6899
food|6900,6904
prior|6905,6910
to|6911,6913
<EOL>|6914,6915
admission|6915,6924
.|6924,6925
She|6926,6929
had|6930,6933
therapeutic|6934,6945
paracentesis|6946,6958
with|6959,6963
4.3|6964,6967
L|6967,6968
removed|6969,6976
<EOL>|6977,6978
and|6978,6981
received|6982,6990
37.5|6991,6995
G|6995,6996
albumin|6997,7004
IV|7005,7007
post|7008,7012
procedure|7013,7022
.|7022,7023
She|7024,7027
felt|7028,7032
much|7033,7037
<EOL>|7038,7039
better|7039,7045
with|7046,7050
resolution|7051,7061
of|7062,7064
abdominal|7065,7074
discomfort|7075,7085
.|7085,7086
Patient|7087,7094
is|7095,7097
<EOL>|7098,7099
scheduled|7099,7108
for|7109,7112
repeat|7113,7119
paracentesis|7120,7132
as|7133,7135
outpatient|7136,7146
on|7147,7149
_|7150,7151
_|7151,7152
_|7152,7153
.|7153,7154
<EOL>|7156,7157
<EOL>|7157,7158
#|7158,7159
HEPATIC|7160,7167
ENCEPHALOPATHY|7168,7182
.|7182,7183
History|7184,7191
of|7192,7194
HE|7195,7197
from|7198,7202
Hep|7203,7206
C|7207,7208
cirrhosis|7209,7218
.|7218,7219
<EOL>|7220,7221
Now|7221,7224
with|7225,7229
mild|7230,7234
encephalopathy|7235,7249
(|7250,7251
hallucinations|7251,7265
and|7266,7269
forgetfulness|7270,7283
)|7283,7284
<EOL>|7285,7286
due|7286,7289
to|7290,7292
medication|7293,7303
noncompliance|7304,7317
,|7317,7318
but|7319,7322
not|7323,7326
acutely|7327,7334
encephalopathic|7335,7350
<EOL>|7351,7352
and|7352,7355
without|7356,7363
asterixis|7364,7373
on|7374,7376
exam|7377,7381
.|7381,7382
Infectious|7383,7393
workup|7394,7400
negative|7401,7409
thus|7410,7414
<EOL>|7415,7416
far|7416,7419
.|7419,7420
Continue|7421,7429
lactulose|7430,7439
30mL|7440,7444
TID|7445,7448
and|7449,7452
titrate|7453,7460
to|7461,7463
3|7464,7465
BMs|7466,7469
daily|7470,7475
and|7476,7479
<EOL>|7480,7481
continue|7481,7489
rifaximin|7490,7499
550mg|7500,7505
BID|7506,7509
.|7509,7510
<EOL>|7511,7512
<EOL>|7513,7514
#|7514,7515
HYPONATREMIA|7516,7528
.|7528,7529
Na|7530,7532
125|7533,7536
on|7537,7539
admission|7540,7549
,|7549,7550
128|7551,7554
four|7555,7559
days|7560,7564
ago|7565,7568
,|7568,7569
and|7570,7573
135|7574,7577
<EOL>|7578,7579
one|7579,7582
month|7583,7588
ago|7589,7592
.|7592,7593
Likely|7594,7600
due|7601,7604
to|7605,7607
third|7608,7613
spacing|7614,7621
from|7622,7626
worsening|7627,7636
<EOL>|7637,7638
ascites|7638,7645
and|7646,7649
fluid|7650,7655
overload|7656,7664
.|7664,7665
1.5|7666,7669
L|7669,7670
fluid|7671,7676
restriction|7677,7688
,|7688,7689
low|7690,7693
salt|7694,7698
<EOL>|7699,7700
diet|7700,7704
.|7704,7705
S|7706,7707
/|7707,7708
p|7708,7709
therapeutic|7710,7721
paracentesis|7722,7734
with|7735,7739
albumin|7740,7747
replacement|7748,7759
.|7759,7760
<EOL>|7760,7761
<EOL>|7761,7762
#|7762,7763
CIRRHOSIS|7764,7773
,|7773,7774
HEPATITIS|7775,7784
C.|7785,7787
MELD|7788,7792
score|7793,7798
of|7799,7801
10|7802,7804
and|7805,7808
Child|7809,7814
's|7814,7816
_|7817,7818
_|7818,7819
_|7819,7820
<EOL>|7821,7822
class|7822,7827
B|7828,7829
on|7830,7832
this|7833,7837
admission|7838,7847
.|7847,7848
Now|7849,7852
decompensated|7853,7866
due|7867,7870
to|7871,7873
ascites|7874,7881
.|7881,7882
<EOL>|7883,7884
Hepatitis|7884,7893
C|7894,7895
genotype|7896,7904
IIIB|7905,7909
.|7909,7910
Dr.|7911,7914
_|7915,7916
_|7916,7917
_|7917,7918
starting|7919,7927
<EOL>|7928,7929
_|7929,7930
_|7930,7931
_|7931,7932
and|7933,7936
_|7937,7938
_|7938,7939
_|7939,7940
with|7941,7945
patient|7946,7953
in|7954,7956
clinic|7957,7963
and|7964,7967
the|7968,7971
<EOL>|7972,7973
insurance|7973,7982
process|7983,7990
was|7991,7994
started|7995,8002
by|8003,8005
her|8006,8009
office|8010,8016
.|8016,8017
No|8018,8020
history|8021,8028
of|8029,8031
EGD|8032,8035
,|8035,8036
<EOL>|8037,8038
needs|8038,8043
this|8044,8048
as|8049,8051
outpatient|8052,8062
for|8063,8066
varices|8067,8074
screening|8075,8084
.|8084,8085
<EOL>|8087,8088
<EOL>|8089,8090
#|8090,8091
NUTRITION|8092,8101
.|8101,8102
Unclear|8103,8110
if|8111,8113
truly|8114,8119
compliant|8120,8129
with|8130,8134
low|8135,8138
salt|8139,8143
diet|8144,8148
.|8148,8149
Poor|8150,8154
<EOL>|8155,8156
oral|8156,8160
intake|8161,8167
.|8167,8168
Low|8169,8172
albumin|8173,8180
2.8|8181,8184
on|8185,8187
admission|8188,8197
.|8197,8198
Met|8199,8202
with|8203,8207
nutrition|8208,8217
.|8217,8218
<EOL>|8219,8220
<EOL>|8221,8222
#|8222,8223
COAGULOPATHY|8224,8236
.|8236,8237
INR|8238,8241
1.4|8242,8245
four|8246,8250
days|8251,8255
ago|8256,8259
.|8259,8260
No|8261,8263
evidence|8264,8272
of|8273,8275
active|8276,8282
<EOL>|8283,8284
bleeding|8284,8292
.|8292,8293
Very|8294,8298
mild|8299,8303
thrombocytopenia|8304,8320
with|8321,8325
plts|8326,8330
143|8331,8334
.|8334,8335
<EOL>|8337,8338
<EOL>|8339,8340
#|8340,8341
HIV|8342,8345
.|8345,8346
Most|8347,8351
recent|8352,8358
CD4|8359,8362
173|8363,8366
.|8366,8367
On|8368,8370
HAART|8371,8376
.|8376,8377
No|8378,8380
established|8381,8392
ID|8393,8395
<EOL>|8396,8397
provider|8397,8405
.|8405,8406
Continue|8407,8415
Truvada|8416,8423
and|8424,8427
Isentress|8428,8437
,|8437,8438
Bactrim|8439,8446
DS|8447,8449
daily|8450,8455
for|8456,8459
<EOL>|8460,8461
PCP|8461,8464
_|8465,8466
_|8466,8467
_|8467,8468
.|8468,8469
Needs|8470,8475
outpatient|8476,8486
ID|8487,8489
appointment|8490,8501
<EOL>|8503,8504
<EOL>|8504,8505
#|8505,8506
COPD|8507,8511
.|8511,8512
Stable|8513,8519
.|8519,8520
States|8521,8527
she|8528,8531
is|8532,8534
on|8535,8537
intermittent|8538,8550
home|8551,8555
O2|8556,8558
for|8559,8562
<EOL>|8563,8564
comfort|8564,8571
at|8572,8574
night|8575,8580
and|8581,8584
with|8585,8589
abdominal|8590,8599
distentiom|8600,8610
.|8610,8611
Continued|8612,8621
home|8622,8626
<EOL>|8627,8628
COPD|8628,8632
meds|8633,8637
and|8638,8641
home|8642,8646
O2|8647,8649
as|8650,8652
needed|8653,8659
<EOL>|8660,8661
<EOL>|8661,8662
*|8662,8663
*|8663,8664
Transitional|8664,8676
Issues|8677,8683
*|8683,8684
*|8684,8685
<EOL>|8685,8686
-|8686,8687
Discontinued|8688,8700
spironolactone|8701,8715
_|8716,8717
_|8717,8718
_|8718,8719
elevated|8720,8728
potassium|8729,8738
<EOL>|8738,8739
-|8739,8740
Increased|8741,8750
furosemide|8751,8761
to|8762,8764
40mg|8765,8769
daily|8770,8775
<EOL>|8775,8776
-|8776,8777
Please|8778,8784
recheck|8785,8792
electrolytes|8793,8805
at|8806,8808
next|8809,8813
visit|8814,8819
<EOL>|8819,8820
-|8820,8821
Had|8822,8825
paracentesis|8826,8838
_|8839,8840
_|8840,8841
_|8841,8842
with|8843,8847
4.3|8848,8851
L|8852,8853
removed|8854,8861
,|8861,8862
received|8863,8871
37.5|8872,8876
G|8876,8877
<EOL>|8878,8879
albumin|8879,8886
<EOL>|8886,8887
-|8887,8888
Needs|8889,8894
outpatient|8895,8905
ID|8906,8908
provider|8909,8917
<EOL>|8917,8918
-|8918,8919
_|8920,8921
_|8921,8922
_|8922,8923
needs|8924,8929
more|8930,8934
frequent|8935,8943
paracentesis|8944,8956
<EOL>|8956,8957
<EOL>|8958,8959
Medications|8959,8970
on|8971,8973
Admission|8974,8983
:|8983,8984
<EOL>|8984,8985
The|8985,8988
Preadmission|8989,9001
Medication|9002,9012
list|9013,9017
is|9018,9020
accurate|9021,9029
and|9030,9033
complete|9034,9042
.|9042,9043
<EOL>|9043,9044
1.|9044,9046
Albuterol|9047,9056
Inhaler|9057,9064
2|9065,9066
PUFF|9067,9071
IH|9072,9074
Q6H|9075,9078
:|9078,9079
PRN|9079,9082
wheezing|9083,9091
,|9091,9092
SOB|9093,9096
<EOL>|9097,9098
2.|9098,9100
_|9101,9102
_|9102,9103
_|9103,9104
(|9105,9106
Truvada|9106,9113
)|9113,9114
1|9115,9116
TAB|9117,9120
PO|9121,9123
DAILY|9124,9129
<EOL>|9130,9131
3.|9131,9133
Furosemide|9134,9144
20|9145,9147
mg|9148,9150
PO|9151,9153
DAILY|9154,9159
<EOL>|9160,9161
4.|9161,9163
Raltegravir|9164,9175
400|9176,9179
mg|9180,9182
PO|9183,9185
BID|9186,9189
<EOL>|9190,9191
5.|9191,9193
Spironolactone|9194,9208
50|9209,9211
mg|9212,9214
PO|9215,9217
DAILY|9218,9223
<EOL>|9224,9225
6.|9225,9227
Acetaminophen|9228,9241
500|9242,9245
mg|9246,9248
PO|9249,9251
Q6H|9252,9255
:|9255,9256
PRN|9256,9259
pain|9260,9264
,|9264,9265
fever|9265,9270
<EOL>|9271,9272
7.|9272,9274
Tiotropium|9275,9285
Bromide|9286,9293
1|9294,9295
CAP|9296,9299
IH|9300,9302
DAILY|9303,9308
<EOL>|9309,9310
8.|9310,9312
Rifaximin|9313,9322
550|9323,9326
mg|9327,9329
PO|9330,9332
BID|9333,9336
<EOL>|9337,9338
9.|9338,9340
Calcium|9341,9348
Carbonate|9349,9358
1250|9359,9363
mg|9364,9366
PO|9367,9369
BID|9370,9373
<EOL>|9374,9375
10.|9375,9378
Lactulose|9379,9388
15|9389,9391
mL|9392,9394
PO|9395,9397
TID|9398,9401
<EOL>|9402,9403
11.|9403,9406
Sulfameth|9407,9416
/|9416,9417
Trimethoprim|9417,9429
DS|9430,9432
1|9433,9434
TAB|9435,9438
PO|9439,9441
DAILY|9442,9447
<EOL>|9448,9449
<EOL>|9449,9450
<EOL>|9451,9452
Discharge|9452,9461
Medications|9462,9473
:|9473,9474
<EOL>|9474,9475
1.|9475,9477
Acetaminophen|9478,9491
500|9492,9495
mg|9496,9498
PO|9499,9501
Q6H|9502,9505
:|9505,9506
PRN|9506,9509
pain|9510,9514
,|9514,9515
fever|9515,9520
<EOL>|9521,9522
2.|9522,9524
Albuterol|9525,9534
Inhaler|9535,9542
2|9543,9544
PUFF|9545,9549
IH|9550,9552
Q6H|9553,9556
:|9556,9557
PRN|9557,9560
wheezing|9561,9569
,|9569,9570
SOB|9571,9574
<EOL>|9575,9576
3|9576,9577
.|9577,9578
Calcium|9579,9586
Carbonate|9587,9596
1250|9597,9601
mg|9602,9604
PO|9605,9607
BID|9608,9611
<EOL>|9612,9613
4.|9613,9615
_|9616,9617
_|9617,9618
_|9618,9619
(|9620,9621
Truvada|9621,9628
)|9628,9629
1|9630,9631
TAB|9632,9635
PO|9636,9638
DAILY|9639,9644
<EOL>|9645,9646
5.|9646,9648
Furosemide|9649,9659
40|9660,9662
mg|9663,9665
PO|9666,9668
DAILY|9669,9674
<EOL>|9675,9676
6.|9676,9678
Lactulose|9679,9688
15|9689,9691
mL|9692,9694
PO|9695,9697
TID|9698,9701
<EOL>|9702,9703
7.|9703,9705
Raltegravir|9706,9717
400|9718,9721
mg|9722,9724
PO|9725,9727
BID|9728,9731
<EOL>|9732,9733
8.|9733,9735
Rifaximin|9736,9745
550|9746,9749
mg|9750,9752
PO|9753,9755
BID|9756,9759
<EOL>|9760,9761
9.|9761,9763
Sulfameth|9764,9773
/|9773,9774
Trimethoprim|9774,9786
DS|9787,9789
1|9790,9791
TAB|9792,9795
PO|9796,9798
DAILY|9799,9804
<EOL>|9805,9806
10.|9806,9809
Tiotropium|9810,9820
Bromide|9821,9828
1|9829,9830
CAP|9831,9834
IH|9835,9837
DAILY|9838,9843
<EOL>|9844,9845
<EOL>|9845,9846
<EOL>|9847,9848
Discharge|9848,9857
Disposition|9858,9869
:|9869,9870
<EOL>|9870,9871
Home|9871,9875
<EOL>|9875,9876
<EOL>|9877,9878
Discharge|9878,9887
Diagnosis|9888,9897
:|9897,9898
<EOL>|9898,9899
Primary|9899,9906
:|9906,9907
diuretic|9909,9917
refractory|9918,9928
ascites|9929,9936
<EOL>|9936,9937
Secondary|9937,9946
:|9946,9947
HCV|9948,9951
cirrhosis|9952,9961
,|9961,9962
HIV|9963,9966
,|9966,9967
hyponatremia|9968,9980
,|9980,9981
COPD|9982,9986
<EOL>|9986,9987
<EOL>|9987,9988
<EOL>|9989,9990
Discharge|9990,9999
Condition|10000,10009
:|10009,10010
<EOL>|10010,10011
Mental|10011,10017
Status|10018,10024
:|10024,10025
Clear|10026,10031
and|10032,10035
coherent|10036,10044
.|10044,10045
<EOL>|10045,10046
Level|10046,10051
of|10052,10054
Consciousness|10055,10068
:|10068,10069
Alert|10070,10075
and|10076,10079
interactive|10080,10091
.|10091,10092
<EOL>|10092,10093
Activity|10093,10101
Status|10102,10108
:|10108,10109
Ambulatory|10110,10120
-|10121,10122
Independent|10123,10134
.|10134,10135
<EOL>|10135,10136
<EOL>|10136,10137
<EOL>|10138,10139
Discharge|10139,10148
Instructions|10149,10161
:|10161,10162
<EOL>|10162,10163
Dear|10163,10167
_|10168,10169
_|10169,10170
_|10170,10171
,|10171,10172
<EOL>|10172,10173
<EOL>|10173,10174
_|10174,10175
_|10175,10176
_|10176,10177
was|10178,10181
a|10182,10183
pleasure|10184,10192
to|10193,10195
take|10196,10200
care|10201,10205
of|10206,10208
you|10209,10212
at|10213,10215
_|10216,10217
_|10217,10218
_|10218,10219
<EOL>|10220,10221
_|10221,10222
_|10222,10223
_|10223,10224
.|10224,10225
You|10226,10229
were|10230,10234
admitted|10235,10243
with|10244,10248
abdominal|10249,10258
fullness|10259,10267
and|10268,10271
<EOL>|10272,10273
pain|10273,10277
from|10278,10282
your|10283,10287
ascites|10288,10295
.|10295,10296
You|10297,10300
had|10301,10304
a|10305,10306
diagnostic|10307,10317
and|10318,10321
therapeutic|10322,10333
<EOL>|10334,10335
paracentesis|10335,10347
with|10348,10352
4.3|10353,10356
L|10357,10358
removed|10359,10366
.|10366,10367
Your|10368,10372
spironolactone|10373,10387
was|10388,10391
<EOL>|10392,10393
discontinued|10393,10405
because|10406,10413
your|10414,10418
potassium|10419,10428
was|10429,10432
high|10433,10437
.|10437,10438
Your|10439,10443
lasix|10444,10449
was|10450,10453
<EOL>|10454,10455
increased|10455,10464
to|10465,10467
40mg|10468,10472
daily|10473,10478
.|10478,10479
You|10480,10483
are|10484,10487
scheduled|10488,10497
for|10498,10501
another|10502,10509
<EOL>|10510,10511
paracentesis|10511,10523
on|10524,10526
_|10527,10528
_|10528,10529
_|10529,10530
prior|10531,10536
to|10537,10539
your|10540,10544
other|10545,10550
appointments|10551,10563
that|10564,10568
day|10569,10572
.|10572,10573
<EOL>|10574,10575
Please|10575,10581
call|10582,10586
tomorrow|10587,10595
to|10596,10598
find|10599,10603
out|10604,10607
the|10608,10611
time|10612,10616
of|10617,10619
the|10620,10623
paracentesis|10624,10636
.|10636,10637
<EOL>|10638,10639
Please|10639,10645
continue|10646,10654
to|10655,10657
follow|10658,10664
a|10665,10666
low|10667,10670
sodium|10671,10677
diet|10678,10682
and|10683,10686
fluid|10687,10692
<EOL>|10693,10694
restriction|10694,10705
.|10705,10706
You|10707,10710
should|10711,10717
call|10718,10722
your|10723,10727
liver|10728,10733
doctor|10734,10740
or|10741,10743
return|10744,10750
to|10751,10753
the|10754,10757
<EOL>|10758,10759
emergency|10759,10768
room|10769,10773
if|10774,10776
you|10777,10780
have|10781,10785
abdominal|10786,10795
pain|10796,10800
,|10800,10801
fever|10802,10807
,|10807,10808
chills|10809,10815
,|10815,10816
<EOL>|10817,10818
confusion|10818,10827
,|10827,10828
or|10829,10831
other|10832,10837
concerning|10838,10848
symptoms|10849,10857
.|10857,10858
<EOL>|10858,10859
<EOL>|10859,10860
Sincerely|10860,10869
,|10869,10870
<EOL>|10870,10871
Your|10871,10875
_|10876,10877
_|10877,10878
_|10878,10879
medical|10880,10887
team|10888,10892
<EOL>|10892,10893
<EOL>|10894,10895
Followup|10895,10903
Instructions|10904,10916
:|10916,10917
<EOL>|10917,10918
_|10918,10919
_|10919,10920
_|10920,10921
<EOL>|10921,10922

