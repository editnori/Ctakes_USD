 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Procedure|Health Care Activity|SIMPLE_SEGMENT|43,52|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|43,57|false|false|false|C2598112||Admission Date
Finding|Body Substance|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|77,86|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|77,91|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|133,136|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|144,151|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|144,151|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|153,161|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|SIMPLE_SEGMENT|164,173|false|false|false|C1717415||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|164,173|false|false|false|C0020517|Hypersensitivity|Allergies
Drug|Antibiotic|SIMPLE_SEGMENT|176,185|false|false|false|C0066005;C1314417|INJECTION, MEROPENEM, 100 MG ADMINISTERED;meropenem|meropenem
Drug|Clinical Drug|SIMPLE_SEGMENT|176,185|false|false|false|C0066005;C1314417|INJECTION, MEROPENEM, 100 MG ADMINISTERED;meropenem|meropenem
Drug|Organic Chemical|SIMPLE_SEGMENT|176,185|false|false|false|C0066005;C1314417|INJECTION, MEROPENEM, 100 MG ADMINISTERED;meropenem|meropenem
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|188,199|false|false|false|C0161486;C2876539|Poisoning by penicillin;Poisoning by, adverse effect of and underdosing of penicillins|Penicillins
Drug|Antibiotic|SIMPLE_SEGMENT|188,199|false|false|false|C0030842|penicillins|Penicillins
Drug|Organic Chemical|SIMPLE_SEGMENT|188,199|false|false|false|C0030842|penicillins|Penicillins
Finding|Pathologic Function|SIMPLE_SEGMENT|188,199|false|false|false|C0413443|Adverse reaction to penicillins|Penicillins
Finding|Functional Concept|SIMPLE_SEGMENT|202,211|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|SIMPLE_SEGMENT|220,235|false|false|false|C0277786|Chief complaint (finding)|Chief Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|226,235|false|false|false|C3864418||Complaint
Finding|Finding|SIMPLE_SEGMENT|226,235|false|false|false|C5441521|Complaint (finding)|Complaint
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|237,242|false|false|false|C0018932|Hematochezia|BRBPR
Finding|Classification|SIMPLE_SEGMENT|245,250|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|SIMPLE_SEGMENT|251,259|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|251,259|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|263,281|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|272,281|false|false|false|C0945766||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|272,281|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|272,281|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|272,281|false|false|false|C0184661|Interventional procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|283,290|false|false|false|C1550015;C1609614;C4318470|Order aborted;aborted - ActStatus;aborted - QueryStatusCode|aborted
Finding|Intellectual Product|SIMPLE_SEGMENT|283,290|false|false|false|C1550015;C1609614;C4318470|Order aborted;aborted - ActStatus;aborted - QueryStatusCode|aborted
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|291,313|false|false|false|C0016234|Flexible fiberoptic sigmoidoscopy|flexible sigmoidoscopy
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|300,313|false|false|false|C0037075;C1548917|Consent Type - Sigmoidoscopy;Sigmoidoscopy (procedure)|sigmoidoscopy
Procedure|Health Care Activity|SIMPLE_SEGMENT|300,313|false|false|false|C0037075;C1548917|Consent Type - Sigmoidoscopy;Sigmoidoscopy (procedure)|sigmoidoscopy
Event|Event|SIMPLE_SEGMENT|314,321|false|false|false|C1516084|Attempt|attempt
Finding|Body Substance|SIMPLE_SEGMENT|330,335|false|false|false|C0015733|Feces|stool
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|339,344|false|false|false|C1550319|Vault|vault
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|351,373|false|false|false|C0016234|Flexible fiberoptic sigmoidoscopy|Flexible sigmoidoscopy
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|360,373|false|false|false|C0037075;C1548917|Consent Type - Sigmoidoscopy;Sigmoidoscopy (procedure)|sigmoidoscopy
Procedure|Health Care Activity|SIMPLE_SEGMENT|360,373|false|false|false|C0037075;C1548917|Consent Type - Sigmoidoscopy;Sigmoidoscopy (procedure)|sigmoidoscopy
Finding|Conceptual Entity|SIMPLE_SEGMENT|381,388|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|381,388|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|381,388|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|381,391|false|false|false|C0262926|Medical History|History of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|381,407|false|false|false|C0488508||History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|381,407|false|false|false|C0262512|History of present illness (finding)|History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|392,399|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Idea or Concept|SIMPLE_SEGMENT|392,399|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Finding|SIMPLE_SEGMENT|392,407|false|false|false|C4264312|Present illness|Present Illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|400,407|false|false|false|C0221423|Illness (finding)|Illness
Finding|Idea or Concept|SIMPLE_SEGMENT|424,428|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|SIMPLE_SEGMENT|424,428|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Finding|SIMPLE_SEGMENT|445,465|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|past medical history
Finding|Functional Concept|SIMPLE_SEGMENT|450,457|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Idea or Concept|SIMPLE_SEGMENT|450,457|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Intellectual Product|SIMPLE_SEGMENT|450,457|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|450,457|false|false|false|C0199168|Medical service|medical
Finding|Finding|SIMPLE_SEGMENT|450,465|false|false|false|C0262926|Medical History|medical history
Finding|Finding|SIMPLE_SEGMENT|450,468|false|false|false|C0262926|Medical History|medical history of
Finding|Conceptual Entity|SIMPLE_SEGMENT|458,465|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|458,465|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|458,465|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|458,468|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|479,493|false|false|false|C0020676|Hypothyroidism|hypothyroidism
Attribute|Clinical Attribute|SIMPLE_SEGMENT|502,511|false|false|false|C0945731||diagnosis
Finding|Classification|SIMPLE_SEGMENT|502,511|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|502,511|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|502,511|false|false|false|C0011900|Diagnosis|diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|518,529|false|false|false|C0332459;C4551657|Compressed structure|compression
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|518,529|false|false|false|C0728907|Compression|compression
Procedure|Machine Activity|SIMPLE_SEGMENT|518,529|false|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|518,529|false|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|530,538|false|false|false|C0016658|Fracture|fracture
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|552,561|false|false|false|C0009450|Communicable Diseases|infection
Finding|Pathologic Function|SIMPLE_SEGMENT|552,561|false|false|false|C3714514|Infection|infection
Finding|Finding|SIMPLE_SEGMENT|579,585|false|false|false|C0423899;C1414153;C3539536|ARID1B wt Allele;ARID3A gene;Above average intellect|bright
Finding|Gene or Genome|SIMPLE_SEGMENT|579,585|false|false|false|C0423899;C1414153;C3539536|ARID1B wt Allele;ARID3A gene;Above average intellect|bright
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|579,589|false|false|false|C1096868|DC Red No. 8|bright red
Drug|Organic Chemical|SIMPLE_SEGMENT|579,589|false|false|false|C1096868|DC Red No. 8|bright red
Finding|Finding|SIMPLE_SEGMENT|579,589|false|false|false|C1272329|Bright red color (finding)|bright red
Finding|Finding|SIMPLE_SEGMENT|586,589|false|false|false|C0332575;C1414207;C1416378|DYRK3 gene;IK gene;Redness|red
Finding|Gene or Genome|SIMPLE_SEGMENT|586,589|false|false|false|C0332575;C1414207;C1416378|DYRK3 gene;IK gene;Redness|red
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|591,596|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|SIMPLE_SEGMENT|591,596|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Functional Concept|SIMPLE_SEGMENT|597,607|false|false|false|C1527425;C4048189|Per rectum;Rectal Route of Administration|per rectum
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|601,607|false|false|false|C0034896;C4482211|Pelvis>Rectum;Rectum|rectum
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|601,607|false|false|false|C0034882;C0154062;C0496867;C0496908|Benign neoplasm of rectum;Carcinoma in situ of rectum;Neoplasm of uncertain or unknown behavior of rectum;Rectal Diseases|rectum
Disorder|Neoplastic Process|SIMPLE_SEGMENT|601,607|false|false|false|C0034882;C0154062;C0496867;C0496908|Benign neoplasm of rectum;Carcinoma in situ of rectum;Neoplasm of uncertain or unknown behavior of rectum;Rectal Diseases|rectum
Procedure|Health Care Activity|SIMPLE_SEGMENT|601,607|false|false|false|C0869814|Procedure on rectum|rectum
Finding|Body Substance|SIMPLE_SEGMENT|610,617|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|610,617|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|610,617|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|645,657|false|false|false|C0449450|Presentation|presentation
Finding|Functional Concept|SIMPLE_SEGMENT|684,689|false|false|false|C1442792|State|state
Finding|Finding|SIMPLE_SEGMENT|684,699|false|false|false|C0683314|personal health|state of health
Finding|Idea or Concept|SIMPLE_SEGMENT|693,699|false|false|false|C0018684|Health|health
Finding|Idea or Concept|SIMPLE_SEGMENT|706,710|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|706,710|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|706,710|false|false|false|C1553498|home health encounter|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|706,717|false|false|false|C1553498|home health encounter|home health
Finding|Idea or Concept|SIMPLE_SEGMENT|711,717|false|false|false|C0018684|Health|health
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|718,721|false|false|false|C1454018|AICDA protein, human|aid
Drug|Enzyme|SIMPLE_SEGMENT|718,721|false|false|false|C1454018|AICDA protein, human|aid
Finding|Gene or Genome|SIMPLE_SEGMENT|718,721|false|false|false|C1421876;C3540469|AICDA gene;AICDA wt Allele|aid
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|718,721|false|false|false|C0021588;C0280108|AID - Artificial insemination by donor;dacarbazine/doxorubicin/ifosfamide protocol|aid
Finding|Finding|SIMPLE_SEGMENT|722,728|false|false|false|C5452990|Helped|helped
Finding|Gene or Genome|SIMPLE_SEGMENT|771,776|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Finding|Intellectual Product|SIMPLE_SEGMENT|777,783|false|false|false|C1705102|Volume (publication)|volume
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|790,795|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|SIMPLE_SEGMENT|790,795|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Functional Concept|SIMPLE_SEGMENT|796,806|false|false|false|C1527425;C4048189|Per rectum;Rectal Route of Administration|per rectum
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|800,806|false|false|false|C0034896;C4482211|Pelvis>Rectum;Rectum|rectum
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|800,806|false|false|false|C0034882;C0154062;C0496867;C0496908|Benign neoplasm of rectum;Carcinoma in situ of rectum;Neoplasm of uncertain or unknown behavior of rectum;Rectal Diseases|rectum
Disorder|Neoplastic Process|SIMPLE_SEGMENT|800,806|false|false|false|C0034882;C0154062;C0496867;C0496908|Benign neoplasm of rectum;Carcinoma in situ of rectum;Neoplasm of uncertain or unknown behavior of rectum;Rectal Diseases|rectum
Procedure|Health Care Activity|SIMPLE_SEGMENT|800,806|false|false|false|C0869814|Procedure on rectum|rectum
Finding|Idea or Concept|SIMPLE_SEGMENT|818,822|false|false|false|C1552851|next - HtmlLinkType|next
Finding|Intellectual Product|SIMPLE_SEGMENT|839,843|false|false|false|C1720594|Then - dosing instruction fragment|then
Finding|Idea or Concept|SIMPLE_SEGMENT|872,876|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|SIMPLE_SEGMENT|872,876|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|SIMPLE_SEGMENT|872,876|false|false|false|C1553498|home health encounter|Home
Procedure|Health Care Activity|SIMPLE_SEGMENT|872,883|false|false|false|C1553498|home health encounter|Home health
Finding|Idea or Concept|SIMPLE_SEGMENT|877,883|false|false|false|C0018684|Health|health
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|884,887|false|false|false|C1454018|AICDA protein, human|aid
Drug|Enzyme|SIMPLE_SEGMENT|884,887|false|false|false|C1454018|AICDA protein, human|aid
Finding|Gene or Genome|SIMPLE_SEGMENT|884,887|false|false|false|C1421876;C3540469|AICDA gene;AICDA wt Allele|aid
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|884,887|false|false|false|C0021588;C0280108|AID - Artificial insemination by donor;dacarbazine/doxorubicin/ifosfamide protocol|aid
Finding|Classification|SIMPLE_SEGMENT|903,909|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|903,909|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|903,909|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|903,909|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|914,918|false|false|false|C1720594|Then - dosing instruction fragment|then
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|985,989|false|false|false|C0587081|Laboratory test finding|Labs
Anatomy|Cell|SIMPLE_SEGMENT|1007,1010|false|false|false|C0023516|Leukocytes|WBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1017,1020|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1017,1020|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|1017,1020|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1017,1020|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1026,1029|false|false|false|C0201617|Primed lymphocyte test|Plt
Drug|Organic Chemical|SIMPLE_SEGMENT|1050,1057|false|false|false|C0022924;C0376261|Lactates;lactate|lactate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1050,1057|false|false|false|C0022924;C0376261|Lactates;lactate|lactate
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1050,1057|false|false|false|C0202115|Lactic acid measurement|lactate
Finding|Finding|SIMPLE_SEGMENT|1066,1069|false|false|false|C5848551|Neg - answer|neg
Finding|Functional Concept|SIMPLE_SEGMENT|1083,1087|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|1083,1087|false|false|false|C0582103|Medical Examination|Exam
Finding|Finding|SIMPLE_SEGMENT|1100,1111|false|false|false|C0039231;C3827868|Tachycardia;Tachycardia by ECG Finding|tachycardia
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1121,1126|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|SIMPLE_SEGMENT|1121,1126|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1127,1133|false|false|false|C0034896;C4482211|Pelvis>Rectum;Rectum|rectum
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1127,1133|false|false|false|C0034882;C0154062;C0496867;C0496908|Benign neoplasm of rectum;Carcinoma in situ of rectum;Neoplasm of uncertain or unknown behavior of rectum;Rectal Diseases|rectum
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1127,1133|false|false|false|C0034882;C0154062;C0496867;C0496908|Benign neoplasm of rectum;Carcinoma in situ of rectum;Neoplasm of uncertain or unknown behavior of rectum;Rectal Diseases|rectum
Procedure|Health Care Activity|SIMPLE_SEGMENT|1127,1133|false|false|false|C0869814|Procedure on rectum|rectum
Finding|Gene or Genome|SIMPLE_SEGMENT|1142,1147|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1148,1159|true|false|false|C0019112|Hemorrhoids|hemorrhoids
Drug|Organic Chemical|SIMPLE_SEGMENT|1161,1164|false|false|false|C0032478;C0032483|polyethylene glycol 400;polyethylene glycols|PEG
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1161,1164|false|false|false|C0032478;C0032483|polyethylene glycol 400;polyethylene glycols|PEG
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1161,1164|false|false|false|C0176751;C4300182|PEG Study;Percutaneous endoscopic gastrostomy|PEG
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1161,1164|false|false|false|C0176751;C4300182|PEG Study;Percutaneous endoscopic gastrostomy|PEG
Finding|Intellectual Product|SIMPLE_SEGMENT|1165,1171|false|false|false|C1546689||lavage
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1165,1171|false|false|false|C0022100|Irrigation|lavage
Finding|Classification|SIMPLE_SEGMENT|1184,1192|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|1184,1192|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1184,1192|false|false|false|C5237010|Expression Negative|negative
Finding|Finding|SIMPLE_SEGMENT|1184,1196|false|false|false|C0205160|Negative|negative for
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1197,1202|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|SIMPLE_SEGMENT|1197,1202|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Drug|Organic Chemical|SIMPLE_SEGMENT|1259,1265|false|false|false|C0699678|Flagyl|flagyl
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1259,1265|false|false|false|C0699678|Flagyl|flagyl
Finding|Gene or Genome|SIMPLE_SEGMENT|1303,1306|false|false|false|C1427027|DHDDS gene|HDS
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1308,1311|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1308,1311|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1329,1333|false|false|false|C0005790|Blood coagulation tests|Coag
Finding|Conceptual Entity|SIMPLE_SEGMENT|1356,1366|false|false|false|C1521721|Supportive assistance|supportive
Procedure|Health Care Activity|SIMPLE_SEGMENT|1356,1371|false|false|false|C0030231;C0344211|Palliative Care;Supportive care|supportive care
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1356,1371|false|false|false|C0030231;C0344211|Palliative Care;Supportive care|supportive care
Event|Activity|SIMPLE_SEGMENT|1367,1371|false|false|false|C1947933|care activity|care
Finding|Finding|SIMPLE_SEGMENT|1367,1371|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|1367,1371|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Drug|Substance|SIMPLE_SEGMENT|1377,1383|false|false|false|C0302908|Liquid substance|fluids
Finding|Body Substance|SIMPLE_SEGMENT|1377,1383|false|false|false|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1377,1383|false|false|false|C0016286|Fluid Therapy|fluids
Finding|Functional Concept|SIMPLE_SEGMENT|1388,1399|false|false|false|C0199960||transfusion
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1388,1399|false|false|false|C0005841;C1879316|Blood Transfusion;Transfusion (procedure)|transfusion
Finding|Pathologic Function|SIMPLE_SEGMENT|1423,1431|false|false|false|C0019080|Hemorrhage|bleeding
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|1435,1446|false|false|false|C0019010|Hemodynamics|hemodynamic
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1435,1446|false|false|false|C4281788|hemodynamics (procedure)|hemodynamic
Finding|Functional Concept|SIMPLE_SEGMENT|1447,1454|false|false|false|C0392747|Changing|changes
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1467,1470|false|false|false|C3813556|Cancer/Testis Antigen|CTA
Finding|Gene or Genome|SIMPLE_SEGMENT|1467,1470|false|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1467,1470|false|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Finding|Idea or Concept|SIMPLE_SEGMENT|1475,1482|false|false|false|C2699424|Concern|concern
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1486,1494|false|false|false|C0203057|Upper gastrointestinal tract series|upper GI
Finding|Pathologic Function|SIMPLE_SEGMENT|1486,1503|false|true|true|C0041909|Upper gastrointestinal hemorrhage|upper GI bleeding
Finding|Pathologic Function|SIMPLE_SEGMENT|1492,1503|false|false|false|C0017181|Gastrointestinal Hemorrhage|GI bleeding
Finding|Pathologic Function|SIMPLE_SEGMENT|1495,1503|false|false|false|C0019080|Hemorrhage|bleeding
Finding|Intellectual Product|SIMPLE_SEGMENT|1509,1515|false|false|false|C1546689||lavage
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1509,1515|false|false|false|C0022100|Irrigation|lavage
Drug|Organic Chemical|SIMPLE_SEGMENT|1520,1523|false|false|false|C0032478;C0032483|polyethylene glycol 400;polyethylene glycols|PEG
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1520,1523|false|false|false|C0032478;C0032483|polyethylene glycol 400;polyethylene glycols|PEG
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1520,1523|false|false|false|C0176751;C4300182|PEG Study;Percutaneous endoscopic gastrostomy|PEG
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1520,1523|false|false|false|C0176751;C4300182|PEG Study;Percutaneous endoscopic gastrostomy|PEG
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1537,1540|false|false|false|C0358591|Proton Pump Inhibitors|PPI
Finding|Physiologic Function|SIMPLE_SEGMENT|1537,1540|false|false|false|C0871125|Prepulse Inhibition|PPI
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|1544,1552|false|false|false|C4727483|BRAF Gene Rearrangement|positive
Finding|Classification|SIMPLE_SEGMENT|1544,1552|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|SIMPLE_SEGMENT|1544,1552|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Body Substance|SIMPLE_SEGMENT|1556,1563|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1556,1563|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1556,1563|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Inorganic Chemical|SIMPLE_SEGMENT|1584,1590|false|false|false|C0036082|Saline Solution|saline
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1584,1590|false|false|false|C0036082|Saline Solution|saline
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1584,1590|false|false|false|C0450082|Saline method|saline
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1611,1619|false|false|false|C0013227|Pharmaceutical Preparations|medicine
Event|Activity|SIMPLE_SEGMENT|1624,1631|false|false|false|C1706079||arrival
Finding|Functional Concept|SIMPLE_SEGMENT|1624,1631|false|false|false|C1555577|arrival - ActRelationshipType|arrival
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|1639,1644|false|false|false|C3714591|Floor (anatomic)|floor
Finding|Body Substance|SIMPLE_SEGMENT|1645,1652|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1645,1652|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1645,1652|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1662,1667|false|false|false|C1552828|Table Frame - above|above
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1686,1695|false|false|false|C0945731||diagnosis
Finding|Classification|SIMPLE_SEGMENT|1686,1695|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|1686,1695|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1686,1695|false|false|false|C0011900|Diagnosis|diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|1702,1713|false|false|false|C0332459;C4551657|Compressed structure|compression
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|1702,1713|false|false|false|C0728907|Compression|compression
Procedure|Machine Activity|SIMPLE_SEGMENT|1702,1713|false|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1702,1713|false|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Finding|Pathologic Function|SIMPLE_SEGMENT|1702,1722|false|false|false|C0521169|Compression fracture|compression fracture
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|1714,1722|false|false|false|C0016658|Fracture|fracture
Finding|Finding|SIMPLE_SEGMENT|1740,1750|false|false|false|C1299586|Has difficulty doing (qualifier value)|difficulty
Drug|Organic Chemical|SIMPLE_SEGMENT|1769,1772|false|false|false|C0032478;C0032483|polyethylene glycol 400;polyethylene glycols|PEG
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1769,1772|false|false|false|C0032478;C0032483|polyethylene glycol 400;polyethylene glycols|PEG
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1769,1772|false|false|false|C0176751;C4300182|PEG Study;Percutaneous endoscopic gastrostomy|PEG
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1769,1772|false|false|false|C0176751;C4300182|PEG Study;Percutaneous endoscopic gastrostomy|PEG
Finding|Functional Concept|SIMPLE_SEGMENT|1773,1777|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|tube
Finding|Gene or Genome|SIMPLE_SEGMENT|1773,1777|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|tube
Finding|Finding|SIMPLE_SEGMENT|1778,1785|false|false|false|C4534363|At home|at home
Finding|Idea or Concept|SIMPLE_SEGMENT|1781,1785|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|1781,1785|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|1781,1785|false|false|false|C1553498|home health encounter|home
Finding|Idea or Concept|SIMPLE_SEGMENT|1802,1808|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Finding|Intellectual Product|SIMPLE_SEGMENT|1802,1808|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Finding|Functional Concept|SIMPLE_SEGMENT|1802,1811|false|false|false|C0699752|Review of|review of
Finding|Functional Concept|SIMPLE_SEGMENT|1812,1819|false|false|false|C0449913|System|systems
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|1820,1828|false|false|false|C4727483|BRAF Gene Rearrangement|positive
Finding|Classification|SIMPLE_SEGMENT|1820,1828|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|SIMPLE_SEGMENT|1820,1828|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Classification|SIMPLE_SEGMENT|1852,1860|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|1852,1860|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1852,1860|false|false|false|C5237010|Expression Negative|negative
Finding|Finding|SIMPLE_SEGMENT|1866,1886|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Finding|Functional Concept|SIMPLE_SEGMENT|1871,1878|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|1871,1878|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|1871,1878|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|1871,1878|false|false|false|C0199168|Medical service|Medical
Finding|Finding|SIMPLE_SEGMENT|1871,1886|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1879,1886|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1879,1886|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|1879,1886|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1897,1911|false|false|false|C0020676|Hypothyroidism|Hypothyroidism
Finding|Finding|SIMPLE_SEGMENT|1916,1922|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|SIMPLE_SEGMENT|1916,1922|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1929,1936|false|false|false|C0033684|Proteins|Protein
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1929,1936|false|false|false|C0033684|Proteins|Protein
Finding|Conceptual Entity|SIMPLE_SEGMENT|1929,1936|false|false|false|C1521746|Protein Info|Protein
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1929,1936|false|false|false|C0202202|Protein measurement|Protein
Finding|Pathologic Function|SIMPLE_SEGMENT|1929,1957|false|false|false|C0033677|Protein-Energy Malnutrition|Protein calorie malnutrition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1945,1957|false|false|false|C0162429|Malnutrition|malnutrition
Drug|Organic Chemical|SIMPLE_SEGMENT|1962,1965|false|false|false|C0032478;C0032483|polyethylene glycol 400;polyethylene glycols|PEG
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1962,1965|false|false|false|C0032478;C0032483|polyethylene glycol 400;polyethylene glycols|PEG
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1962,1965|false|false|false|C0176751;C4300182|PEG Study;Percutaneous endoscopic gastrostomy|PEG
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1962,1965|false|false|false|C0176751;C4300182|PEG Study;Percutaneous endoscopic gastrostomy|PEG
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1966,1978|false|false|false|C0029456|Osteoporosis|Osteoporosis
Finding|Finding|SIMPLE_SEGMENT|1966,1978|false|false|false|C2911643|Encounter due to family history of osteoporosis|Osteoporosis
Finding|Functional Concept|SIMPLE_SEGMENT|1986,1997|false|false|false|C0332459;C4551657|Compressed structure|compression
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|1986,1997|false|false|false|C0728907|Compression|compression
Procedure|Machine Activity|SIMPLE_SEGMENT|1986,1997|false|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1986,1997|false|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Finding|Pathologic Function|SIMPLE_SEGMENT|1986,2006|false|false|false|C0521169|Compression fracture|compression fracture
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|1998,2006|false|false|false|C0016658|Fracture|fracture
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|2007,2017|false|false|false|C0011570;C0011581;C0344315;C0812393|Cancer patients and suicide and depression;Depressed mood;Depressive disorder;Mental Depression|Depression
Finding|Functional Concept|SIMPLE_SEGMENT|2007,2017|false|false|false|C0460137;C1579931|Depression - motion|Depression
Finding|Sign or Symptom|SIMPLE_SEGMENT|2007,2017|false|false|false|C0460137;C1579931|Depression - motion|Depression
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2018,2029|false|false|false|C0019112|Hemorrhoids|Hemorrhoids
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2041,2047|false|false|false|C0002871|Anemia|anemia
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2049,2063|false|false|false|C0006267|Bronchiectasis|Bronchiectasis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2069,2077|false|false|false|C0019360|Herpes zoster (disorder)|Shingles
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|2079,2087|false|false|false|C0011265;C0497327|Dementia;Presenile dementia|Dementia
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2098,2118|false|false|false|C0026266|Mitral Valve Insufficiency|Mitral regurgitation
Finding|Finding|SIMPLE_SEGMENT|2105,2118|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|SIMPLE_SEGMENT|2105,2118|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|SIMPLE_SEGMENT|2105,2118|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Finding|Functional Concept|SIMPLE_SEGMENT|2123,2129|false|false|false|C0728831|Social|Social
Finding|Finding|SIMPLE_SEGMENT|2123,2137|false|false|false|C0424945;C3714536|Social History;Social and personal history|Social History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2130,2137|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2130,2137|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2130,2137|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Classification|SIMPLE_SEGMENT|2143,2149|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|SIMPLE_SEGMENT|2143,2149|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|SIMPLE_SEGMENT|2143,2149|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|SIMPLE_SEGMENT|2143,2149|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Finding|SIMPLE_SEGMENT|2143,2157|false|false|false|C0241889|Family Medical History|Family History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2150,2157|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2150,2157|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2150,2157|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2176,2182|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Idea or Concept|SIMPLE_SEGMENT|2176,2182|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2187,2198|false|false|false|C0019112|Hemorrhoids|hemorrhoids
Finding|Conceptual Entity|SIMPLE_SEGMENT|2204,2211|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|2204,2211|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|2204,2211|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|2204,2214|false|false|false|C0262926|Medical History|history of
Finding|Finding|SIMPLE_SEGMENT|2204,2221|true|false|false|C0455471|History of malignant neoplasm|history of cancer
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2215,2221|true|false|false|C0006826|Malignant Neoplasms|cancer
Finding|Pathologic Function|SIMPLE_SEGMENT|2223,2234|false|false|false|C0017181|Gastrointestinal Hemorrhage|GI bleeding
Finding|Pathologic Function|SIMPLE_SEGMENT|2226,2234|false|false|false|C0019080|Hemorrhage|bleeding
Finding|Finding|SIMPLE_SEGMENT|2240,2248|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|2240,2248|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|2240,2248|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|2240,2253|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2240,2253|false|false|false|C0031809|Physical Examination|Physical Exam
Finding|Functional Concept|SIMPLE_SEGMENT|2249,2253|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2249,2253|false|false|false|C0582103|Medical Examination|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2255,2264|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Finding|Classification|SIMPLE_SEGMENT|2310,2313|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Finding|Gene or Genome|SIMPLE_SEGMENT|2310,2313|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2326,2329|false|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Finding|Intellectual Product|SIMPLE_SEGMENT|2326,2329|false|false|false|C2346952|Bachelor of Education|bed
Finding|Finding|SIMPLE_SEGMENT|2331,2342|false|false|false|C5546696|Feeling comfortable|comfortable
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2344,2348|false|false|false|C4750744|Acute limbic encephalitis following transplant|pale
Finding|Finding|SIMPLE_SEGMENT|2344,2348|false|false|false|C0241137;C0678215|Body pale (finding);Pallor of skin|pale
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2349,2353|false|false|false|C0015392|Eye|Eyes
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2349,2353|false|false|false|C5848506||Eyes
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2361,2364|false|false|false|C0150934;C0175196|Ear, nose and throat;Structure of entorhinal cortex|ENT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2361,2364|false|false|false|C0150934;C0175196|Ear, nose and throat;Structure of entorhinal cortex|ENT
Finding|Gene or Genome|SIMPLE_SEGMENT|2361,2364|false|false|false|C0262471;C1417861;C3889152|ENT problem;NT5E gene;NT5E wt Allele|ENT
Finding|Sign or Symptom|SIMPLE_SEGMENT|2361,2364|false|false|false|C0262471;C1417861;C3889152|ENT problem;NT5E gene;NT5E wt Allele|ENT
Finding|Idea or Concept|SIMPLE_SEGMENT|2370,2375|false|false|false|C1550016|Remote control command - Clear|clear
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2377,2380|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2377,2380|false|false|false|C0026987|Myelofibrosis|MMM
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2381,2386|false|false|false|C0018787;C4037974|Chest>Heart;Heart|Heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2381,2386|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|Heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|2381,2386|false|false|false|C0795691|HEART PROBLEM|Heart
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|2418,2426|false|false|false|C0039155|Systole|systolic
Finding|Finding|SIMPLE_SEGMENT|2418,2433|false|false|false|C0232257|Systolic Murmurs|systolic murmur
Finding|Finding|SIMPLE_SEGMENT|2427,2433|false|false|false|C0018808|Heart murmur|murmur
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2445,2451|false|false|false|C0004454|Axilla|axilla
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2454,2459|false|false|false|C0024109|Lung|Lungs
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2462,2465|false|false|false|C3813556|Cancer/Testis Antigen|CTA
Finding|Gene or Genome|SIMPLE_SEGMENT|2462,2465|false|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2462,2465|false|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2478,2481|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|Abd
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|2478,2481|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|Abd
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2484,2488|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2512,2517|false|false|false|C0021853|Intestines|bowel
Finding|Finding|SIMPLE_SEGMENT|2512,2524|false|false|false|C0232693|Bowel sounds|bowel sounds
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|2518,2524|false|false|false|C0037709||sounds
Drug|Organic Chemical|SIMPLE_SEGMENT|2526,2529|false|false|false|C0032478;C0032483|polyethylene glycol 400;polyethylene glycols|PEG
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2526,2529|false|false|false|C0032478;C0032483|polyethylene glycol 400;polyethylene glycols|PEG
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2526,2529|false|false|false|C0176751;C4300182|PEG Study;Percutaneous endoscopic gastrostomy|PEG
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2526,2529|false|false|false|C0176751;C4300182|PEG Study;Percutaneous endoscopic gastrostomy|PEG
Event|Activity|SIMPLE_SEGMENT|2533,2538|false|false|false|C1882509|put - instruction imperative|place
Finding|Functional Concept|SIMPLE_SEGMENT|2533,2538|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|SIMPLE_SEGMENT|2533,2538|false|false|false|C1533810||place
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2539,2545|false|false|false|C0034896;C4482211|Pelvis>Rectum;Rectum|Rectum
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2539,2545|false|false|false|C0034882;C0154062;C0496867;C0496908|Benign neoplasm of rectum;Carcinoma in situ of rectum;Neoplasm of uncertain or unknown behavior of rectum;Rectal Diseases|Rectum
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2539,2545|false|false|false|C0034882;C0154062;C0496867;C0496908|Benign neoplasm of rectum;Carcinoma in situ of rectum;Neoplasm of uncertain or unknown behavior of rectum;Rectal Diseases|Rectum
Procedure|Health Care Activity|SIMPLE_SEGMENT|2539,2545|false|false|false|C0869814|Procedure on rectum|Rectum
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2560,2565|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|SIMPLE_SEGMENT|2560,2565|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2569,2574|false|false|false|C1550319|Vault|vault
Finding|Gene or Genome|SIMPLE_SEGMENT|2579,2584|true|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2585,2596|true|false|false|C0019112|Hemorrhoids|hemorrhoids
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|2606,2609|false|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Finding|Gene or Genome|SIMPLE_SEGMENT|2606,2609|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Finding|Functional Concept|SIMPLE_SEGMENT|2612,2617|false|false|false|C1883002|Sequence Chromatogram|trace
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2618,2623|false|false|false|C1717255||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|2618,2623|false|false|false|C0013604|Edema|edema
Anatomy|Body System|SIMPLE_SEGMENT|2636,2640|false|false|false|C1123023;C4520765|Skin;Skin, Human|Skin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2636,2640|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|Skin
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2636,2640|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|Skin
Finding|Body Substance|SIMPLE_SEGMENT|2636,2640|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|Skin
Finding|Intellectual Product|SIMPLE_SEGMENT|2636,2640|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|Skin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2644,2648|false|false|false|C4750744|Acute limbic encephalitis following transplant|pale
Finding|Finding|SIMPLE_SEGMENT|2644,2648|false|false|false|C0241137;C0678215|Body pale (finding);Pallor of skin|pale
Finding|Sign or Symptom|SIMPLE_SEGMENT|2653,2659|true|false|false|C0015230;C5779628|Exanthema;Skin rash|rashes
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2660,2664|false|false|false|C0042373|Vascular Diseases|Vasc
Finding|Conceptual Entity|SIMPLE_SEGMENT|2673,2679|false|false|false|C0442038;C0920847|Circumpennate;Radial|radial
Drug|Food|SIMPLE_SEGMENT|2680,2686|false|false|false|C5890763||pulses
Finding|Physiologic Function|SIMPLE_SEGMENT|2680,2686|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|SIMPLE_SEGMENT|2680,2686|false|false|false|C0034107|Pulse taking|pulses
Finding|Gene or Genome|SIMPLE_SEGMENT|2695,2699|false|false|false|C1425523|AOX2P gene|AOx2
Finding|Intellectual Product|SIMPLE_SEGMENT|2708,2712|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|name
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2732,2747|false|false|false|C0278454|All extremities|all extremities
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2736,2747|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|2748,2753|false|false|false|C0004936;C1306597|Mental disorders;Psychiatric problem|Psych
Finding|Body Substance|SIMPLE_SEGMENT|2769,2778|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|2769,2778|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|2769,2778|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|2769,2778|false|false|false|C0030685|Patient Discharge|DISCHARGE
Finding|Classification|SIMPLE_SEGMENT|2808,2811|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Finding|Gene or Genome|SIMPLE_SEGMENT|2808,2811|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2824,2827|false|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Finding|Intellectual Product|SIMPLE_SEGMENT|2824,2827|false|false|false|C2346952|Bachelor of Education|bed
Finding|Finding|SIMPLE_SEGMENT|2829,2840|false|false|false|C5546696|Feeling comfortable|comfortable
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2851,2855|false|false|false|C0015392|Eye|Eyes
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2851,2855|false|false|false|C5848506||Eyes
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2863,2866|false|false|false|C0150934;C0175196|Ear, nose and throat;Structure of entorhinal cortex|ENT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2863,2866|false|false|false|C0150934;C0175196|Ear, nose and throat;Structure of entorhinal cortex|ENT
Finding|Gene or Genome|SIMPLE_SEGMENT|2863,2866|false|false|false|C0262471;C1417861;C3889152|ENT problem;NT5E gene;NT5E wt Allele|ENT
Finding|Sign or Symptom|SIMPLE_SEGMENT|2863,2866|false|false|false|C0262471;C1417861;C3889152|ENT problem;NT5E gene;NT5E wt Allele|ENT
Finding|Idea or Concept|SIMPLE_SEGMENT|2872,2877|false|false|false|C1550016|Remote control command - Clear|clear
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2879,2882|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2879,2882|false|false|false|C0026987|Myelofibrosis|MMM
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2883,2888|false|false|false|C0018787;C4037974|Chest>Heart;Heart|Heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2883,2888|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|Heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|2883,2888|false|false|false|C0795691|HEART PROBLEM|Heart
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|2902,2910|false|false|false|C0039155|Systole|systolic
Finding|Finding|SIMPLE_SEGMENT|2902,2917|false|false|false|C0232257|Systolic Murmurs|systolic murmur
Finding|Finding|SIMPLE_SEGMENT|2911,2917|false|false|false|C0018808|Heart murmur|murmur
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2929,2935|false|false|false|C0004454|Axilla|axilla
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2938,2943|false|false|false|C0024109|Lung|Lungs
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2946,2949|false|false|false|C3813556|Cancer/Testis Antigen|CTA
Finding|Gene or Genome|SIMPLE_SEGMENT|2946,2949|false|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2946,2949|false|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Finding|Finding|SIMPLE_SEGMENT|2963,2972|false|false|false|C0442739||unchanged
Finding|Idea or Concept|SIMPLE_SEGMENT|2978,2981|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|2978,2981|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2988,2991|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|Abd
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|2988,2991|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|Abd
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2994,2998|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3022,3027|false|false|false|C0021853|Intestines|bowel
Finding|Finding|SIMPLE_SEGMENT|3022,3034|false|false|false|C0232693|Bowel sounds|bowel sounds
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3028,3034|false|false|false|C0037709||sounds
Drug|Organic Chemical|SIMPLE_SEGMENT|3036,3039|false|false|false|C0032478;C0032483|polyethylene glycol 400;polyethylene glycols|PEG
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3036,3039|false|false|false|C0032478;C0032483|polyethylene glycol 400;polyethylene glycols|PEG
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3036,3039|false|false|false|C0176751;C4300182|PEG Study;Percutaneous endoscopic gastrostomy|PEG
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3036,3039|false|false|false|C0176751;C4300182|PEG Study;Percutaneous endoscopic gastrostomy|PEG
Event|Activity|SIMPLE_SEGMENT|3043,3048|false|false|false|C1882509|put - instruction imperative|place
Finding|Functional Concept|SIMPLE_SEGMENT|3043,3048|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|SIMPLE_SEGMENT|3043,3048|false|false|false|C1533810||place
Finding|Finding|SIMPLE_SEGMENT|3051,3060|false|false|false|C0442739||unchanged
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|3077,3080|false|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Finding|Gene or Genome|SIMPLE_SEGMENT|3077,3080|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3086,3091|true|false|false|C1717255||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|3086,3091|true|false|false|C0013604|Edema|edema
Anatomy|Body System|SIMPLE_SEGMENT|3093,3097|false|false|false|C1123023;C4520765|Skin;Skin, Human|Skin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3093,3097|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|Skin
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3093,3097|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|Skin
Finding|Body Substance|SIMPLE_SEGMENT|3093,3097|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|Skin
Finding|Intellectual Product|SIMPLE_SEGMENT|3093,3097|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|Skin
Finding|Sign or Symptom|SIMPLE_SEGMENT|3103,3109|true|false|false|C0015230;C5779628|Exanthema;Skin rash|rashes
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3110,3114|false|false|false|C0042373|Vascular Diseases|Vasc
Finding|Conceptual Entity|SIMPLE_SEGMENT|3123,3129|false|false|false|C0442038;C0920847|Circumpennate;Radial|radial
Drug|Food|SIMPLE_SEGMENT|3130,3136|false|false|false|C5890763||pulses
Finding|Physiologic Function|SIMPLE_SEGMENT|3130,3136|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|SIMPLE_SEGMENT|3130,3136|false|false|false|C0034107|Pulse taking|pulses
Finding|Intellectual Product|SIMPLE_SEGMENT|3156,3160|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|name
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3180,3195|false|false|false|C0278454|All extremities|all extremities
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3184,3195|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|3196,3201|false|false|false|C0004936;C1306597|Mental disorders;Psychiatric problem|Psych
Procedure|Health Care Activity|SIMPLE_SEGMENT|3237,3246|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3259,3264|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3259,3264|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|3265,3268|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|3275,3278|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3275,3278|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3275,3278|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3285,3288|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3285,3288|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|3285,3288|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3285,3288|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3294,3297|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3294,3297|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|3305,3308|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3305,3308|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3305,3308|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3305,3308|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|3312,3315|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3312,3315|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|3312,3315|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|3312,3315|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3312,3315|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3321,3325|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3353,3356|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3373,3378|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3373,3378|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|3373,3386|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3373,3386|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3373,3386|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3379,3386|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|3379,3386|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3379,3386|false|false|false|C0017725|glucose|Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3379,3386|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3379,3386|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|SIMPLE_SEGMENT|3430,3434|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3430,3434|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3430,3434|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3459,3464|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3459,3464|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3465,3468|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3465,3468|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|SIMPLE_SEGMENT|3465,3468|false|false|false|C0001899|Alanine Transaminase|ALT
Finding|Gene or Genome|SIMPLE_SEGMENT|3465,3468|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|SIMPLE_SEGMENT|3465,3468|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|SIMPLE_SEGMENT|3465,3468|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3465,3468|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|3472,3475|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3472,3475|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3472,3475|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3472,3475|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|SIMPLE_SEGMENT|3472,3475|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Finding|Gene or Genome|SIMPLE_SEGMENT|3472,3475|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3479,3486|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|SIMPLE_SEGMENT|3479,3486|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Finding|Body Substance|SIMPLE_SEGMENT|3503,3512|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|3503,3512|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|3503,3512|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|3503,3512|false|false|false|C0030685|Patient Discharge|DISCHARGE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3525,3530|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3525,3530|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|3531,3534|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|3539,3542|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3539,3542|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3539,3542|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3549,3552|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3549,3552|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|3549,3552|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3549,3552|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3559,3562|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3559,3562|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|3570,3573|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3570,3573|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3570,3573|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3570,3573|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|3577,3580|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3577,3580|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|3577,3580|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|3577,3580|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3577,3580|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3586,3590|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3617,3620|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3637,3642|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3637,3642|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|3637,3650|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3637,3650|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3637,3650|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3643,3650|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|3643,3650|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3643,3650|false|false|false|C0017725|glucose|Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3643,3650|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3643,3650|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|SIMPLE_SEGMENT|3696,3700|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3696,3700|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3696,3700|false|false|false|C0202059|Bicarbonate measurement|HCO3
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3714,3736|false|false|false|C0016234|Flexible fiberoptic sigmoidoscopy|Flexible Sigmoidoscopy
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3723,3736|false|false|false|C0037075;C1548917|Consent Type - Sigmoidoscopy;Sigmoidoscopy (procedure)|Sigmoidoscopy
Procedure|Health Care Activity|SIMPLE_SEGMENT|3723,3736|false|false|false|C0037075;C1548917|Consent Type - Sigmoidoscopy;Sigmoidoscopy (procedure)|Sigmoidoscopy
Anatomy|Tissue|SIMPLE_SEGMENT|3743,3749|false|false|false|C0026724|Mucous Membrane|Mucosa
Finding|Intellectual Product|SIMPLE_SEGMENT|3743,3749|false|false|false|C1561514||Mucosa
Anatomy|Tissue|SIMPLE_SEGMENT|3758,3764|false|false|false|C0026724|Mucous Membrane|mucosa
Finding|Intellectual Product|SIMPLE_SEGMENT|3758,3764|false|false|false|C1561514||mucosa
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3782,3788|false|false|false|C0034896;C4482211|Pelvis>Rectum;Rectum|rectum
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3782,3788|false|false|false|C0034882;C0154062;C0496867;C0496908|Benign neoplasm of rectum;Carcinoma in situ of rectum;Neoplasm of uncertain or unknown behavior of rectum;Rectal Diseases|rectum
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3782,3788|false|false|false|C0034882;C0154062;C0496867;C0496908|Benign neoplasm of rectum;Carcinoma in situ of rectum;Neoplasm of uncertain or unknown behavior of rectum;Rectal Diseases|rectum
Procedure|Health Care Activity|SIMPLE_SEGMENT|3782,3788|false|false|false|C0869814|Procedure on rectum|rectum
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3782,3806|false|false|false|C0521377|Rectum and sigmoid colon|rectum and sigmoid colon
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3793,3800|false|false|false|C0227391|Sigmoid colon|sigmoid
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3793,3806|false|false|false|C0227391|Sigmoid colon|sigmoid colon
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3793,3806|false|false|false|C0153436;C0496864|Benign neoplasm of sigmoid colon;Malignant neoplasm of sigmoid colon|sigmoid colon
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3801,3806|false|false|false|C0009368;C4071907|Abdomen+Pelvis>Colon;Colon structure (body structure)|colon
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3801,3806|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3801,3806|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Finding|Finding|SIMPLE_SEGMENT|3801,3806|false|false|false|C0750873|COLON PROBLEM|colon
Finding|Pathologic Function|SIMPLE_SEGMENT|3820,3828|true|false|false|C0019080|Hemorrhage|bleeding
Finding|Finding|SIMPLE_SEGMENT|3829,3836|true|false|false|C0449416|Source|sources
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3840,3845|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|SIMPLE_SEGMENT|3840,3845|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3876,3883|false|false|false|C0227391|Sigmoid colon|sigmoid
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3876,3889|false|false|false|C0227391|Sigmoid colon|sigmoid colon
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3876,3889|false|false|false|C0153436;C0496864|Benign neoplasm of sigmoid colon;Malignant neoplasm of sigmoid colon|sigmoid colon
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3884,3889|false|false|false|C0009368;C4071907|Abdomen+Pelvis>Colon;Colon structure (body structure)|colon
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3884,3889|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3884,3889|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Finding|Finding|SIMPLE_SEGMENT|3884,3889|false|false|false|C0750873|COLON PROBLEM|colon
Finding|Intellectual Product|SIMPLE_SEGMENT|3915,3919|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|poor
Event|Activity|SIMPLE_SEGMENT|3920,3924|false|false|false|C1521827|Preparation|prep
Finding|Gene or Genome|SIMPLE_SEGMENT|3920,3924|false|false|false|C1418885;C1425030;C4319962|PITRM1 gene;PITRM1 wt Allele;PREP gene|prep
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3920,3924|false|false|false|C5400798||prep
Finding|Intellectual Product|SIMPLE_SEGMENT|3928,3938|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|Impression
Finding|Mental Process|SIMPLE_SEGMENT|3928,3938|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|Impression
Anatomy|Tissue|SIMPLE_SEGMENT|3947,3953|false|false|false|C0026724|Mucous Membrane|mucosa
Finding|Intellectual Product|SIMPLE_SEGMENT|3947,3953|false|false|false|C1561514||mucosa
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3961,3967|false|false|false|C0034896;C4482211|Pelvis>Rectum;Rectum|rectum
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3961,3967|false|false|false|C0034882;C0154062;C0496867;C0496908|Benign neoplasm of rectum;Carcinoma in situ of rectum;Neoplasm of uncertain or unknown behavior of rectum;Rectal Diseases|rectum
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3961,3967|false|false|false|C0034882;C0154062;C0496867;C0496908|Benign neoplasm of rectum;Carcinoma in situ of rectum;Neoplasm of uncertain or unknown behavior of rectum;Rectal Diseases|rectum
Procedure|Health Care Activity|SIMPLE_SEGMENT|3961,3967|false|false|false|C0869814|Procedure on rectum|rectum
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3961,3985|false|false|false|C0521377|Rectum and sigmoid colon|rectum and sigmoid colon
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3972,3979|false|false|false|C0227391|Sigmoid colon|sigmoid
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3972,3985|false|false|false|C0227391|Sigmoid colon|sigmoid colon
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3972,3985|false|false|false|C0153436;C0496864|Benign neoplasm of sigmoid colon;Malignant neoplasm of sigmoid colon|sigmoid colon
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3980,3985|false|false|false|C0009368;C4071907|Abdomen+Pelvis>Colon;Colon structure (body structure)|colon
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3980,3985|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3980,3985|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Finding|Finding|SIMPLE_SEGMENT|3980,3985|false|false|false|C0750873|COLON PROBLEM|colon
Finding|Pathologic Function|SIMPLE_SEGMENT|3989,3997|true|false|false|C0019080|Hemorrhage|bleeding
Finding|Finding|SIMPLE_SEGMENT|3998,4005|true|false|false|C0449416|Source|sources
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4009,4014|true|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|SIMPLE_SEGMENT|4009,4014|true|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4045,4052|false|false|false|C0227391|Sigmoid colon|sigmoid
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4045,4058|false|false|false|C0227391|Sigmoid colon|sigmoid colon
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4045,4058|false|false|false|C0153436;C0496864|Benign neoplasm of sigmoid colon;Malignant neoplasm of sigmoid colon|sigmoid colon
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4053,4058|false|false|false|C0009368;C4071907|Abdomen+Pelvis>Colon;Colon structure (body structure)|colon
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4053,4058|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4053,4058|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Finding|Finding|SIMPLE_SEGMENT|4053,4058|false|false|false|C0750873|COLON PROBLEM|colon
Finding|Intellectual Product|SIMPLE_SEGMENT|4084,4088|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|poor
Event|Activity|SIMPLE_SEGMENT|4089,4093|false|false|false|C1521827|Preparation|prep
Finding|Gene or Genome|SIMPLE_SEGMENT|4089,4093|false|false|false|C1418885;C1425030;C4319962|PITRM1 gene;PITRM1 wt Allele;PREP gene|prep
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4089,4093|false|false|false|C5400798||prep
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4112,4125|false|false|false|C0037075;C1548917|Consent Type - Sigmoidoscopy;Sigmoidoscopy (procedure)|sigmoidoscopy
Procedure|Health Care Activity|SIMPLE_SEGMENT|4112,4125|false|false|false|C0037075;C1548917|Consent Type - Sigmoidoscopy;Sigmoidoscopy (procedure)|sigmoidoscopy
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4129,4136|false|false|false|C0227391|Sigmoid colon|sigmoid
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4129,4142|false|false|false|C0227391|Sigmoid colon|sigmoid colon
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4129,4142|false|false|false|C0153436;C0496864|Benign neoplasm of sigmoid colon;Malignant neoplasm of sigmoid colon|sigmoid colon
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4137,4142|false|false|false|C0009368;C4071907|Abdomen+Pelvis>Colon;Colon structure (body structure)|colon
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4137,4142|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4137,4142|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Finding|Finding|SIMPLE_SEGMENT|4137,4142|false|false|false|C0750873|COLON PROBLEM|colon
Finding|Idea or Concept|SIMPLE_SEGMENT|4153,4168|false|false|false|C0034866|Recommendation|Recommendations
Finding|Pathologic Function|SIMPLE_SEGMENT|4173,4181|false|false|false|C0019080|Hemorrhage|bleeding
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4212,4223|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Procedure|Health Care Activity|SIMPLE_SEGMENT|4212,4223|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Event|Activity|SIMPLE_SEGMENT|4229,4233|false|false|false|C1521827|Preparation|prep
Finding|Gene or Genome|SIMPLE_SEGMENT|4229,4233|false|false|false|C1418885;C1425030;C4319962|PITRM1 gene;PITRM1 wt Allele;PREP gene|prep
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4229,4233|false|false|false|C5400798||prep
Finding|Intellectual Product|SIMPLE_SEGMENT|4239,4244|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|Brief
Finding|Idea or Concept|SIMPLE_SEGMENT|4245,4253|false|false|false|C1547192|Organization unit type - Hospital|Hospital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4245,4260|false|false|false|C0488549||Hospital Course
Finding|Finding|SIMPLE_SEGMENT|4245,4260|false|false|false|C0489547|Hospital course|Hospital Course
Finding|Idea or Concept|SIMPLE_SEGMENT|4277,4281|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|SIMPLE_SEGMENT|4277,4281|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Finding|SIMPLE_SEGMENT|4298,4318|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|past medical history
Finding|Functional Concept|SIMPLE_SEGMENT|4303,4310|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Idea or Concept|SIMPLE_SEGMENT|4303,4310|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Intellectual Product|SIMPLE_SEGMENT|4303,4310|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|4303,4310|false|false|false|C0199168|Medical service|medical
Finding|Finding|SIMPLE_SEGMENT|4303,4318|false|false|false|C0262926|Medical History|medical history
Finding|Finding|SIMPLE_SEGMENT|4303,4321|false|false|false|C0262926|Medical History|medical history of
Finding|Conceptual Entity|SIMPLE_SEGMENT|4311,4318|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|4311,4318|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|4311,4318|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|4311,4321|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4333,4344|false|false|false|C0019112|Hemorrhoids|hemorrhoids
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4358,4367|false|false|false|C0009450|Communicable Diseases|infection
Finding|Pathologic Function|SIMPLE_SEGMENT|4358,4367|false|false|false|C3714514|Infection|infection
Finding|Finding|SIMPLE_SEGMENT|4388,4394|false|false|false|C0423899;C1414153;C3539536|ARID1B wt Allele;ARID3A gene;Above average intellect|bright
Finding|Gene or Genome|SIMPLE_SEGMENT|4388,4394|false|false|false|C0423899;C1414153;C3539536|ARID1B wt Allele;ARID3A gene;Above average intellect|bright
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|4388,4398|false|false|false|C1096868|DC Red No. 8|bright red
Drug|Organic Chemical|SIMPLE_SEGMENT|4388,4398|false|false|false|C1096868|DC Red No. 8|bright red
Finding|Finding|SIMPLE_SEGMENT|4388,4398|false|false|false|C1272329|Bright red color (finding)|bright red
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4388,4415|false|false|false|C0018932|Hematochezia|bright red blood per rectum
Finding|Finding|SIMPLE_SEGMENT|4395,4398|false|false|false|C0332575;C1414207;C1416378|DYRK3 gene;IK gene;Redness|red
Finding|Gene or Genome|SIMPLE_SEGMENT|4395,4398|false|false|false|C0332575;C1414207;C1416378|DYRK3 gene;IK gene;Redness|red
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4399,4404|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|SIMPLE_SEGMENT|4399,4404|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Pathologic Function|SIMPLE_SEGMENT|4399,4415|false|false|false|C0267596|Rectal hemorrhage|blood per rectum
Finding|Functional Concept|SIMPLE_SEGMENT|4405,4415|false|false|false|C1527425;C4048189|Per rectum;Rectal Route of Administration|per rectum
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4409,4415|false|false|false|C0034896;C4482211|Pelvis>Rectum;Rectum|rectum
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4409,4415|false|false|false|C0034882;C0154062;C0496867;C0496908|Benign neoplasm of rectum;Carcinoma in situ of rectum;Neoplasm of uncertain or unknown behavior of rectum;Rectal Diseases|rectum
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4409,4415|false|false|false|C0034882;C0154062;C0496867;C0496908|Benign neoplasm of rectum;Carcinoma in situ of rectum;Neoplasm of uncertain or unknown behavior of rectum;Rectal Diseases|rectum
Procedure|Health Care Activity|SIMPLE_SEGMENT|4409,4415|false|false|false|C0869814|Procedure on rectum|rectum
Finding|Idea or Concept|SIMPLE_SEGMENT|4416,4423|false|false|false|C0039869;C4319827|Thought|thought
Finding|Mental Process|SIMPLE_SEGMENT|4416,4423|false|false|false|C0039869;C4319827|Thought|thought
Finding|Intellectual Product|SIMPLE_SEGMENT|4430,4435|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4436,4441|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|4436,4441|false|false|false|C2003888|Lower (action)|lower
Finding|Pathologic Function|SIMPLE_SEGMENT|4446,4451|false|false|false|C0019080|Hemorrhage|bleed
Procedure|Health Care Activity|SIMPLE_SEGMENT|4486,4498|true|false|false|C0184661;C0886296;C1273869|Intervention regimes;Interventional procedure;Nursing interventions|intervention
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4486,4498|true|false|false|C0184661;C0886296;C1273869|Intervention regimes;Interventional procedure;Nursing interventions|intervention
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4500,4506|false|false|false|C5889824||status
Finding|Idea or Concept|SIMPLE_SEGMENT|4500,4506|false|false|false|C1546481|What subject filter - Status|status
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4513,4535|false|false|false|C0016234|Flexible fiberoptic sigmoidoscopy|flexible sigmoidoscopy
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4522,4535|false|false|false|C0037075;C1548917|Consent Type - Sigmoidoscopy;Sigmoidoscopy (procedure)|sigmoidoscopy
Procedure|Health Care Activity|SIMPLE_SEGMENT|4522,4535|false|false|false|C0037075;C1548917|Consent Type - Sigmoidoscopy;Sigmoidoscopy (procedure)|sigmoidoscopy
Finding|Conceptual Entity|SIMPLE_SEGMENT|4544,4556|false|false|false|C1705683|Identifiable Class|identifiable
Finding|Finding|SIMPLE_SEGMENT|4557,4563|true|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Finding|Functional Concept|SIMPLE_SEGMENT|4557,4563|true|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Finding|Intellectual Product|SIMPLE_SEGMENT|4557,4563|true|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Finding|Intellectual Product|SIMPLE_SEGMENT|4576,4582|false|false|false|C1547311|Patient Condition Code - Stable|stable
Finding|Finding|SIMPLE_SEGMENT|4606,4610|false|false|false|C1299581|Able (qualifier value)|able
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4632,4637|false|false|false|C0034991|Rehabilitation therapy|rehab
Finding|Intellectual Product|SIMPLE_SEGMENT|4638,4646|false|false|false|C4695111|ADMIN.FACILITY|facility
Finding|Intellectual Product|SIMPLE_SEGMENT|4651,4656|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|Acute
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4651,4665|false|false|false|C0266807|Acute gastrointestinal hemorrhage|Acute GI Bleed
Finding|Pathologic Function|SIMPLE_SEGMENT|4657,4665|false|false|false|C0017181|Gastrointestinal Hemorrhage|GI Bleed
Finding|Pathologic Function|SIMPLE_SEGMENT|4660,4665|false|false|false|C0019080|Hemorrhage|Bleed
Finding|Body Substance|SIMPLE_SEGMENT|4672,4679|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|4672,4679|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|4672,4679|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|4695,4700|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4713,4718|false|false|false|C0018932|Hematochezia|BRBPR
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4734,4739|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|4734,4739|false|false|false|C2003888|Lower (action)|lower
Finding|Finding|SIMPLE_SEGMENT|4743,4749|false|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Finding|Functional Concept|SIMPLE_SEGMENT|4743,4749|false|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Finding|Intellectual Product|SIMPLE_SEGMENT|4743,4749|false|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Finding|Body Substance|SIMPLE_SEGMENT|4752,4759|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|4752,4759|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|4752,4759|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Finding|SIMPLE_SEGMENT|4792,4795|true|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|4792,4795|true|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4809,4815|true|false|false|C0002871|Anemia|anemia
Finding|Social Behavior|SIMPLE_SEGMENT|4824,4834|false|false|false|C2584313|Discussion (communication)|discussion
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4824,4834|false|false|false|C0557061|Discussion (procedure)|discussion
Finding|Classification|SIMPLE_SEGMENT|4841,4847|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|4841,4847|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|4841,4847|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|4841,4847|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Body Substance|SIMPLE_SEGMENT|4852,4859|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|4852,4859|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|4852,4859|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4920,4942|false|false|false|C0016234|Flexible fiberoptic sigmoidoscopy|flexible sigmoidoscopy
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4929,4942|false|false|false|C0037075;C1548917|Consent Type - Sigmoidoscopy;Sigmoidoscopy (procedure)|sigmoidoscopy
Procedure|Health Care Activity|SIMPLE_SEGMENT|4929,4942|false|false|false|C0037075;C1548917|Consent Type - Sigmoidoscopy;Sigmoidoscopy (procedure)|sigmoidoscopy
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4949,4960|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Procedure|Health Care Activity|SIMPLE_SEGMENT|4949,4960|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Finding|Body Substance|SIMPLE_SEGMENT|4987,4994|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|4987,4994|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|4987,4994|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Functional Concept|SIMPLE_SEGMENT|5005,5012|false|false|false|C1550015;C1609614;C4318470|Order aborted;aborted - ActStatus;aborted - QueryStatusCode|aborted
Finding|Intellectual Product|SIMPLE_SEGMENT|5005,5012|false|false|false|C1550015;C1609614;C4318470|Order aborted;aborted - ActStatus;aborted - QueryStatusCode|aborted
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5023,5036|false|false|false|C0037075;C1548917|Consent Type - Sigmoidoscopy;Sigmoidoscopy (procedure)|sigmoidoscopy
Procedure|Health Care Activity|SIMPLE_SEGMENT|5023,5036|false|false|false|C0037075;C1548917|Consent Type - Sigmoidoscopy;Sigmoidoscopy (procedure)|sigmoidoscopy
Finding|Finding|SIMPLE_SEGMENT|5064,5071|false|false|false|C3845930|Copious|copious
Finding|Body Substance|SIMPLE_SEGMENT|5072,5077|false|false|false|C0015733|Feces|stool
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5082,5088|false|false|false|C1272938|Rectal Dosage Form|rectal
Finding|Finding|SIMPLE_SEGMENT|5082,5088|false|false|false|C1527425;C4521903|Rectal (intended site);Rectal Route of Administration|rectal
Finding|Functional Concept|SIMPLE_SEGMENT|5082,5088|false|false|false|C1527425;C4521903|Rectal (intended site);Rectal Route of Administration|rectal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5089,5094|false|false|false|C1550319|Vault|vault
Finding|Intellectual Product|SIMPLE_SEGMENT|5100,5104|false|false|false|C1720594|Then - dosing instruction fragment|then
Finding|Social Behavior|SIMPLE_SEGMENT|5115,5125|false|false|false|C0597535|Success|successful
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5136,5149|false|false|false|C0037075;C1548917|Consent Type - Sigmoidoscopy;Sigmoidoscopy (procedure)|sigmoidoscopy
Procedure|Health Care Activity|SIMPLE_SEGMENT|5136,5149|false|false|false|C0037075;C1548917|Consent Type - Sigmoidoscopy;Sigmoidoscopy (procedure)|sigmoidoscopy
Finding|Conceptual Entity|SIMPLE_SEGMENT|5165,5177|false|false|false|C1705683|Identifiable Class|identifiable
Finding|Finding|SIMPLE_SEGMENT|5178,5184|false|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Finding|Functional Concept|SIMPLE_SEGMENT|5178,5184|false|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Finding|Intellectual Product|SIMPLE_SEGMENT|5178,5184|false|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Finding|Pathologic Function|SIMPLE_SEGMENT|5194,5202|false|false|false|C0019080|Hemorrhage|bleeding
Procedure|Health Care Activity|SIMPLE_SEGMENT|5210,5219|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5220,5223|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5220,5223|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|5220,5223|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5220,5223|false|false|false|C0019029|Hemoglobin concentration|Hgb
Finding|Body Substance|SIMPLE_SEGMENT|5229,5238|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|5229,5238|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|5229,5238|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|5229,5238|false|false|false|C0030685|Patient Discharge|discharge
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5239,5249|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5239,5249|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Organic Chemical|SIMPLE_SEGMENT|5239,5249|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5239,5249|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Finding|Finding|SIMPLE_SEGMENT|5239,5249|false|false|false|C1561562|Hemoglobin finding|hemoglobin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5239,5249|false|false|false|C0518015|Hemoglobin measurement|hemoglobin
Finding|Classification|SIMPLE_SEGMENT|5285,5295|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|5285,5295|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5296,5307|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Procedure|Health Care Activity|SIMPLE_SEGMENT|5296,5307|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Finding|Idea or Concept|SIMPLE_SEGMENT|5312,5322|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|5312,5327|false|false|false|C0332290|Consistent with|consistent with
Finding|Body Substance|SIMPLE_SEGMENT|5328,5335|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|5328,5335|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|5328,5335|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5351,5363|false|false|false|C0029456|Osteoporosis|Osteoporosis
Finding|Finding|SIMPLE_SEGMENT|5351,5363|false|false|false|C2911643|Encounter due to family history of osteoporosis|Osteoporosis
Finding|Intellectual Product|SIMPLE_SEGMENT|5366,5373|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|5366,5373|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Finding|Functional Concept|SIMPLE_SEGMENT|5377,5388|false|false|false|C0332459;C4551657|Compressed structure|compression
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|5377,5388|false|false|false|C0728907|Compression|compression
Procedure|Machine Activity|SIMPLE_SEGMENT|5377,5388|false|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5377,5388|false|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Finding|Pathologic Function|SIMPLE_SEGMENT|5377,5397|false|false|false|C0521169|Compression fracture|compression fracture
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|5389,5397|false|false|false|C0016658|Fracture|fracture
Finding|Body Substance|SIMPLE_SEGMENT|5418,5425|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|5418,5425|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|5418,5425|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|SIMPLE_SEGMENT|5441,5452|false|false|false|C0332459;C4551657|Compressed structure|compression
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|5441,5452|false|false|false|C0728907|Compression|compression
Procedure|Machine Activity|SIMPLE_SEGMENT|5441,5452|false|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5441,5452|false|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Finding|Pathologic Function|SIMPLE_SEGMENT|5441,5461|false|false|false|C0521169|Compression fracture|compression fracture
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|5453,5461|false|false|false|C0016658|Fracture|fracture
Finding|Classification|SIMPLE_SEGMENT|5466,5476|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|5466,5476|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Procedure|Health Care Activity|SIMPLE_SEGMENT|5486,5495|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Body Substance|SIMPLE_SEGMENT|5497,5504|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|5497,5504|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|5497,5504|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Procedure|Health Care Activity|SIMPLE_SEGMENT|5551,5560|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Social Behavior|SIMPLE_SEGMENT|5572,5582|false|false|false|C0018896|Helping Behavior|assistance
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|5588,5592|false|false|false|C0001288|Activity of daily living (function)|ADLs
Finding|Body Substance|SIMPLE_SEGMENT|5595,5602|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|5595,5602|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|5595,5602|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5635,5640|false|false|false|C0034991|Rehabilitation therapy|rehab
Finding|Idea or Concept|SIMPLE_SEGMENT|5653,5657|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|5653,5657|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|5653,5657|false|false|false|C1553498|home health encounter|home
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5659,5666|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|5659,5666|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5659,5666|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5659,5666|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|5659,5666|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|5659,5666|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5659,5666|false|false|false|C0201925|Calcium measurement|Calcium
Drug|Organic Chemical|SIMPLE_SEGMENT|5673,5680|false|false|false|C0042890|Vitamins|vitamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5673,5680|false|false|false|C0042890|Vitamins|vitamin
Drug|Vitamin|SIMPLE_SEGMENT|5673,5680|false|false|false|C0042890|Vitamins|vitamin
Drug|Hormone|SIMPLE_SEGMENT|5673,5682|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|vitamin D
Drug|Organic Chemical|SIMPLE_SEGMENT|5673,5682|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|vitamin D
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5673,5682|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|vitamin D
Drug|Vitamin|SIMPLE_SEGMENT|5673,5682|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|vitamin D
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5673,5682|false|false|false|C0919758|Vitamin D measurement|vitamin D
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5684,5694|false|false|false|C0006668;C0770558;C1704385;C2825090;C4520796|Calcitonin Precursor, human;Calcitonin [EPC];Recombinant Calcitonin;calcitonin;human calcitonin|calcitonin
Drug|Hormone|SIMPLE_SEGMENT|5684,5694|false|false|false|C0006668;C0770558;C1704385;C2825090;C4520796|Calcitonin Precursor, human;Calcitonin [EPC];Recombinant Calcitonin;calcitonin;human calcitonin|calcitonin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5684,5694|false|false|false|C0006668;C0770558;C1704385;C2825090;C4520796|Calcitonin Precursor, human;Calcitonin [EPC];Recombinant Calcitonin;calcitonin;human calcitonin|calcitonin
Finding|Gene or Genome|SIMPLE_SEGMENT|5684,5694|false|false|false|C1367551|CALCA gene|calcitonin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5684,5694|false|false|false|C0201924|Calcitonin measurement|calcitonin
Drug|Organic Chemical|SIMPLE_SEGMENT|5707,5714|false|false|false|C0699142|Tylenol|Tylenol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5707,5714|false|false|false|C0699142|Tylenol|Tylenol
Drug|Organic Chemical|SIMPLE_SEGMENT|5720,5728|false|false|false|C0040610|tramadol|tramadol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5720,5728|false|false|false|C0040610|tramadol|tramadol
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5720,5728|false|false|false|C1266765|Tramadol measurement (procedure)|tramadol
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5733,5737|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|5733,5737|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|5733,5737|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|SIMPLE_SEGMENT|5733,5745|false|false|false|C5548091|Demonstrates adequate pain control|pain control
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5733,5745|false|false|false|C0002766;C1304888|Pain control;Pain management (procedure)|pain control
Drug|Organic Chemical|SIMPLE_SEGMENT|5738,5745|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5738,5745|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Substance|SIMPLE_SEGMENT|5738,5745|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Finding|Conceptual Entity|SIMPLE_SEGMENT|5738,5745|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Functional Concept|SIMPLE_SEGMENT|5738,5745|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Idea or Concept|SIMPLE_SEGMENT|5738,5745|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Idea or Concept|SIMPLE_SEGMENT|5751,5755|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Finding|Finding|SIMPLE_SEGMENT|5751,5762|false|false|false|C0541990|good effect|good effect
Finding|Intellectual Product|SIMPLE_SEGMENT|5767,5774|false|false|false|C1547296|Chronic - Admission Level of Care Code|Chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|5767,5774|false|false|false|C1555457|Provision of recurring care for chronic illness|Chronic
Finding|Finding|SIMPLE_SEGMENT|5775,5781|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|Severe
Finding|Intellectual Product|SIMPLE_SEGMENT|5775,5781|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|Severe
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5775,5810|false|false|false|C1283368||Severe Protein Calorie Malnutrition
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5782,5789|false|false|false|C0033684|Proteins|Protein
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5782,5789|false|false|false|C0033684|Proteins|Protein
Finding|Conceptual Entity|SIMPLE_SEGMENT|5782,5789|false|false|false|C1521746|Protein Info|Protein
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5782,5789|false|false|false|C0202202|Protein measurement|Protein
Finding|Pathologic Function|SIMPLE_SEGMENT|5782,5810|false|false|false|C0033677|Protein-Energy Malnutrition|Protein Calorie Malnutrition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5798,5810|false|false|false|C0162429|Malnutrition|Malnutrition
Finding|Social Behavior|SIMPLE_SEGMENT|5817,5827|false|false|false|C2584313|Discussion (communication)|discussion
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5817,5827|false|false|false|C0557061|Discussion (procedure)|discussion
Finding|Classification|SIMPLE_SEGMENT|5834,5840|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|5834,5840|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|5834,5840|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|5834,5840|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|5845,5851|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Finding|Intellectual Product|SIMPLE_SEGMENT|5845,5851|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Finding|Functional Concept|SIMPLE_SEGMENT|5845,5854|false|false|false|C0699752|Review of|review of
Finding|Intellectual Product|SIMPLE_SEGMENT|5855,5860|false|false|false|C0684240|Charts (publication)|chart
Finding|Body Substance|SIMPLE_SEGMENT|5862,5869|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|5862,5869|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|5862,5869|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|SIMPLE_SEGMENT|5862,5873|false|false|false|C0332310|Has patient|patient has
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5879,5885|false|false|false|C0944911||weight
Finding|Finding|SIMPLE_SEGMENT|5879,5885|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|SIMPLE_SEGMENT|5879,5885|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|SIMPLE_SEGMENT|5879,5885|false|false|false|C1305866|Weighing patient|weight
Drug|Organic Chemical|SIMPLE_SEGMENT|5895,5898|false|false|false|C0032478;C0032483|polyethylene glycol 400;polyethylene glycols|PEG
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5895,5898|false|false|false|C0032478;C0032483|polyethylene glycol 400;polyethylene glycols|PEG
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5895,5898|false|false|false|C0176751;C4300182|PEG Study;Percutaneous endoscopic gastrostomy|PEG
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5895,5898|false|false|false|C0176751;C4300182|PEG Study;Percutaneous endoscopic gastrostomy|PEG
Procedure|Health Care Activity|SIMPLE_SEGMENT|5899,5908|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5899,5908|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Finding|Body Substance|SIMPLE_SEGMENT|5913,5918|false|false|false|C1186706;C1550436|Bolus of ingested food;Response Modality - Bolus|bolus
Finding|Intellectual Product|SIMPLE_SEGMENT|5913,5918|false|false|false|C1186706;C1550436|Bolus of ingested food;Response Modality - Bolus|bolus
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5913,5918|false|false|false|C1511237|bolus infusion|bolus
Finding|Functional Concept|SIMPLE_SEGMENT|5919,5923|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|tube
Finding|Gene or Genome|SIMPLE_SEGMENT|5919,5923|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|tube
Finding|Functional Concept|SIMPLE_SEGMENT|5924,5929|false|false|false|C1510670|Feeds|feeds
Finding|Finding|SIMPLE_SEGMENT|5939,5949|false|false|false|C1299586|Has difficulty doing (qualifier value)|difficulty
Finding|Functional Concept|SIMPLE_SEGMENT|5966,5972|false|false|false|C1512806|Intake|intake
Procedure|Health Care Activity|SIMPLE_SEGMENT|5966,5972|false|false|false|C3251814;C4521161|Intake (treatment);Measurement of fluid intake|intake
Finding|Finding|SIMPLE_SEGMENT|5996,6003|false|false|false|C4534363|At home|At home
Finding|Idea or Concept|SIMPLE_SEGMENT|5999,6003|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|5999,6003|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|5999,6003|false|false|false|C1553498|home health encounter|home
Finding|Body Substance|SIMPLE_SEGMENT|6004,6011|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|6004,6011|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|6004,6011|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|SIMPLE_SEGMENT|6004,6015|false|false|false|C0332310|Has patient|patient has
Drug|Food|SIMPLE_SEGMENT|6057,6063|false|false|false|C1875551|NUTREN|Nutren
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6074,6077|false|false|false|C0228225|Structure of calcar avis|Cal
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6074,6077|false|false|false|C1135160|monoclonal antibody CAL|Cal
Drug|Immunologic Factor|SIMPLE_SEGMENT|6074,6077|false|false|false|C1135160|monoclonal antibody CAL|Cal
Finding|Gene or Genome|SIMPLE_SEGMENT|6074,6077|false|false|false|C1425021;C1825283;C3273482;C5890925|FBLIM1 wt Allele;FBLP1 gene;GOPC gene;GOPC wt Allele|Cal
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|6084,6087|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6084,6087|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6084,6087|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|SIMPLE_SEGMENT|6084,6087|false|false|false|C1332410|BID gene|BID
Finding|Body Substance|SIMPLE_SEGMENT|6095,6102|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|6095,6102|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|6095,6102|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Finding|SIMPLE_SEGMENT|6111,6120|false|false|false|C0392209;C0518896;C1442959|Nutrition (function);Nutrition outcomes;Nutritional status|nutrition
Finding|Intellectual Product|SIMPLE_SEGMENT|6111,6120|false|false|false|C0392209;C0518896;C1442959|Nutrition (function);Nutrition outcomes;Nutritional status|nutrition
Finding|Organism Function|SIMPLE_SEGMENT|6111,6120|false|false|false|C0392209;C0518896;C1442959|Nutrition (function);Nutrition outcomes;Nutritional status|nutrition
Procedure|Research Activity|SIMPLE_SEGMENT|6111,6120|false|false|false|C0600072;C1521729|Feeding and dietary regimes;Nutritional Study|nutrition
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6111,6120|false|false|false|C0600072;C1521729|Feeding and dietary regimes;Nutritional Study|nutrition
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|6164,6168|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6164,6168|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|6164,6168|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|6164,6168|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6169,6184|false|false|false|C0242297|Dietary Supplementation|supplementation
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|6198,6203|false|false|false|C1998602|Meal (occasion for eating)|meals
Finding|Finding|SIMPLE_SEGMENT|6207,6211|false|false|false|C5575035|Well (answer to question)|well
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|6219,6229|false|false|false|C0011570;C0011581;C0344315;C0812393|Cancer patients and suicide and depression;Depressed mood;Depressive disorder;Mental Depression|Depression
Finding|Functional Concept|SIMPLE_SEGMENT|6219,6229|false|false|false|C0460137;C1579931|Depression - motion|Depression
Finding|Sign or Symptom|SIMPLE_SEGMENT|6219,6229|false|false|false|C0460137;C1579931|Depression - motion|Depression
Finding|Idea or Concept|SIMPLE_SEGMENT|6242,6246|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|6242,6246|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|6242,6246|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|6247,6256|false|false|false|C0085208|bupropion|BuPROPion
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6247,6256|false|false|false|C0085208|bupropion|BuPROPion
Drug|Organic Chemical|SIMPLE_SEGMENT|6261,6272|false|false|false|C0049506|mirtazapine|mirtazapine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6261,6272|false|false|false|C0049506|mirtazapine|mirtazapine
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6304,6317|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Hormone|SIMPLE_SEGMENT|6304,6317|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Organic Chemical|SIMPLE_SEGMENT|6304,6317|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6304,6317|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Finding|Idea or Concept|SIMPLE_SEGMENT|6320,6332|false|false|false|C1548597|Marketing basis - Transitional|Transitional
Event|Occupational Activity|SIMPLE_SEGMENT|6342,6346|false|false|false|C0009219|Coding|Code
Finding|Intellectual Product|SIMPLE_SEGMENT|6342,6346|false|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|Code
Procedure|Health Care Activity|SIMPLE_SEGMENT|6342,6353|false|false|false|C0742531|CODE STATUS|Code status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6347,6353|false|false|false|C5889824||status
Finding|Idea or Concept|SIMPLE_SEGMENT|6347,6353|false|false|false|C1546481|What subject filter - Status|status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6356,6359|false|false|false|C4285234||DNR
Drug|Antibiotic|SIMPLE_SEGMENT|6356,6359|false|false|false|C0011015|daunorubicin|DNR
Drug|Organic Chemical|SIMPLE_SEGMENT|6356,6359|false|false|false|C0011015|daunorubicin|DNR
Finding|Finding|SIMPLE_SEGMENT|6356,6359|false|false|false|C0079252;C0582114|Do not resuscitate status;Do-Not-Resuscitate Orders|DNR
Finding|Intellectual Product|SIMPLE_SEGMENT|6356,6359|false|false|false|C0079252;C0582114|Do not resuscitate status;Do-Not-Resuscitate Orders|DNR
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6380,6385|false|false|false|C0034991|Rehabilitation therapy|rehab
Finding|Finding|SIMPLE_SEGMENT|6391,6397|true|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Finding|Functional Concept|SIMPLE_SEGMENT|6391,6397|true|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Finding|Intellectual Product|SIMPLE_SEGMENT|6391,6397|true|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Finding|Pathologic Function|SIMPLE_SEGMENT|6402,6410|true|false|false|C0019080|Hemorrhage|bleeding
Procedure|Health Care Activity|SIMPLE_SEGMENT|6427,6436|false|true|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Idea or Concept|SIMPLE_SEGMENT|6442,6450|false|false|false|C0750591|consider|consider
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6459,6470|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Procedure|Health Care Activity|SIMPLE_SEGMENT|6459,6470|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Finding|Finding|SIMPLE_SEGMENT|6483,6489|false|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Finding|Functional Concept|SIMPLE_SEGMENT|6483,6489|false|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Finding|Intellectual Product|SIMPLE_SEGMENT|6483,6489|false|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Finding|Pathologic Function|SIMPLE_SEGMENT|6493,6501|false|false|false|C0019080|Hemorrhage|bleeding
Finding|Idea or Concept|SIMPLE_SEGMENT|6531,6541|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|6531,6546|false|false|false|C0332290|Consistent with|consistent with
Finding|Body Substance|SIMPLE_SEGMENT|6547,6554|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|6547,6554|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|6547,6554|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6557,6562|false|false|false|C2979882||goals
Finding|Idea or Concept|SIMPLE_SEGMENT|6557,6562|false|false|false|C0018017;C0679840;C1546459|What subject filter - Goals;objective (goal);treatment goals|goals
Finding|Intellectual Product|SIMPLE_SEGMENT|6557,6562|false|false|false|C0018017;C0679840;C1546459|What subject filter - Goals;objective (goal);treatment goals|goals
Procedure|Health Care Activity|SIMPLE_SEGMENT|6557,6570|false|false|false|C2930505|Goals of Care|goals of care
Event|Activity|SIMPLE_SEGMENT|6566,6570|false|false|false|C1947933|care activity|care
Finding|Finding|SIMPLE_SEGMENT|6566,6570|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|6566,6570|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Social Behavior|SIMPLE_SEGMENT|6588,6601|false|false|false|C0870494|encouragement|encouragement
Finding|Functional Concept|SIMPLE_SEGMENT|6608,6614|false|false|false|C1512806|Intake|intake
Procedure|Health Care Activity|SIMPLE_SEGMENT|6608,6614|false|false|false|C3251814;C4521161|Intake (treatment);Measurement of fluid intake|intake
Drug|Organic Chemical|SIMPLE_SEGMENT|6619,6622|false|false|false|C0032478;C0032483|polyethylene glycol 400;polyethylene glycols|PEG
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6619,6622|false|false|false|C0032478;C0032483|polyethylene glycol 400;polyethylene glycols|PEG
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6619,6622|false|false|false|C0176751;C4300182|PEG Study;Percutaneous endoscopic gastrostomy|PEG
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6619,6622|false|false|false|C0176751;C4300182|PEG Study;Percutaneous endoscopic gastrostomy|PEG
Finding|Functional Concept|SIMPLE_SEGMENT|6623,6627|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|tube
Finding|Gene or Genome|SIMPLE_SEGMENT|6623,6627|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|tube
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6629,6644|false|false|false|C0242297|Dietary Supplementation|supplementation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6655,6667|false|false|false|C0162429|Malnutrition|malnutrition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6671,6682|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6671,6682|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|6671,6682|false|false|false|C4284232|Medications|Medications
Finding|Finding|SIMPLE_SEGMENT|6671,6695|false|false|false|C1627937|Medications on admission|Medications on Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|6686,6695|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6714,6724|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|6714,6724|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|6714,6729|false|false|false|C0746470|MEDICATION LIST|Medication list
Finding|Intellectual Product|SIMPLE_SEGMENT|6725,6729|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Drug|Organic Chemical|SIMPLE_SEGMENT|6746,6754|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6746,6754|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|SIMPLE_SEGMENT|6746,6754|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Finding|Functional Concept|SIMPLE_SEGMENT|6746,6754|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|SIMPLE_SEGMENT|6746,6754|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Organic Chemical|SIMPLE_SEGMENT|6759,6768|false|false|false|C0085208|bupropion|BuPROPion
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6759,6768|false|false|false|C0085208|bupropion|BuPROPion
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6805,6812|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|6805,6812|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|6805,6812|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6805,6812|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|6805,6812|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|6805,6812|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6805,6812|false|false|false|C0201925|Calcium measurement|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6805,6820|false|false|false|C3864384|Calcium 500+D|Calcium 500 + D
Drug|Vitamin|SIMPLE_SEGMENT|6805,6820|false|false|false|C3864384|Calcium 500+D|Calcium 500 + D
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6822,6829|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|6822,6829|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|6822,6829|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6822,6829|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Vitamin|SIMPLE_SEGMENT|6822,6829|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|6822,6829|false|false|false|C4553026|Calcium metabolic function|calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6822,6829|false|false|false|C0201925|Calcium measurement|calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|6822,6839|false|false|false|C0006681|calcium carbonate|calcium carbonate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6822,6839|false|false|false|C0006681|calcium carbonate|calcium carbonate
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|6830,6839|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|carbonate
Drug|Organic Chemical|SIMPLE_SEGMENT|6830,6839|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|carbonate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6830,6839|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|carbonate
Drug|Organic Chemical|SIMPLE_SEGMENT|6840,6847|false|false|false|C0042890|Vitamins|vitamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6840,6847|false|false|false|C0042890|Vitamins|vitamin
Drug|Vitamin|SIMPLE_SEGMENT|6840,6847|false|false|false|C0042890|Vitamins|vitamin
Drug|Organic Chemical|SIMPLE_SEGMENT|6840,6850|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6840,6850|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Drug|Vitamin|SIMPLE_SEGMENT|6840,6850|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|6879,6883|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6879,6883|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|6879,6883|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|6879,6883|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6894,6907|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Hormone|SIMPLE_SEGMENT|6894,6907|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Organic Chemical|SIMPLE_SEGMENT|6894,6907|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6894,6907|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6894,6914|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Hormone|SIMPLE_SEGMENT|6894,6914|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6894,6914|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6908,6914|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|6908,6914|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6908,6914|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|6908,6914|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6908,6914|false|false|false|C0337443|Sodium measurement|Sodium
Drug|Organic Chemical|SIMPLE_SEGMENT|6935,6946|false|false|false|C0049506|mirtazapine|Mirtazapine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6935,6946|false|false|false|C0049506|mirtazapine|Mirtazapine
Drug|Organic Chemical|SIMPLE_SEGMENT|6964,6972|false|false|false|C0040610|tramadol|TraMADol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6964,6972|false|false|false|C0040610|tramadol|TraMADol
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6964,6972|false|false|false|C1266765|Tramadol measurement (procedure)|TraMADol
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|6982,6985|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6982,6985|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6982,6985|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|SIMPLE_SEGMENT|6982,6985|false|false|false|C1332410|BID gene|BID
Finding|Gene or Genome|SIMPLE_SEGMENT|6986,6989|false|false|false|C1422467|CIAO3 gene|PRN
Finding|Sign or Symptom|SIMPLE_SEGMENT|6990,6999|false|true|false|C0004604|Back Pain|back pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6995,6999|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|6995,6999|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|6995,6999|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|SIMPLE_SEGMENT|7004,7017|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7004,7017|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7004,7017|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|SIMPLE_SEGMENT|7032,7035|false|false|false|C1422467|CIAO3 gene|PRN
Finding|Sign or Symptom|SIMPLE_SEGMENT|7036,7045|false|true|false|C0004604|Back Pain|back pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7041,7045|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|7041,7045|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|7041,7045|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|SIMPLE_SEGMENT|7050,7061|false|false|false|C0102118|alendronate|Alendronate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7050,7061|false|false|false|C0102118|alendronate|Alendronate
Drug|Organic Chemical|SIMPLE_SEGMENT|7050,7068|false|false|false|C0700482|alendronate sodium|Alendronate Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7050,7068|false|false|false|C0700482|alendronate sodium|Alendronate Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7062,7068|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|7062,7068|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7062,7068|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|7062,7068|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7062,7068|false|false|false|C0337443|Sodium measurement|Sodium
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7087,7097|false|false|false|C0006668;C0770558;C1704385;C2825090;C4520796|Calcitonin Precursor, human;Calcitonin [EPC];Recombinant Calcitonin;calcitonin;human calcitonin|Calcitonin
Drug|Hormone|SIMPLE_SEGMENT|7087,7097|false|false|false|C0006668;C0770558;C1704385;C2825090;C4520796|Calcitonin Precursor, human;Calcitonin [EPC];Recombinant Calcitonin;calcitonin;human calcitonin|Calcitonin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7087,7097|false|false|false|C0006668;C0770558;C1704385;C2825090;C4520796|Calcitonin Precursor, human;Calcitonin [EPC];Recombinant Calcitonin;calcitonin;human calcitonin|Calcitonin
Finding|Gene or Genome|SIMPLE_SEGMENT|7087,7097|false|false|false|C1367551|CALCA gene|Calcitonin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7087,7097|false|false|false|C0201924|Calcitonin measurement|Calcitonin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7087,7104|false|false|false|C0073994|salmon calcitonin|Calcitonin Salmon
Drug|Hormone|SIMPLE_SEGMENT|7087,7104|false|false|false|C0073994|salmon calcitonin|Calcitonin Salmon
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7087,7104|false|false|false|C0073994|salmon calcitonin|Calcitonin Salmon
Drug|Food|SIMPLE_SEGMENT|7098,7104|false|false|false|C0459210;C2702377;C4521768|Salmon (substance);salmon allergenic extract|Salmon
Drug|Immunologic Factor|SIMPLE_SEGMENT|7098,7104|false|false|false|C0459210;C2702377;C4521768|Salmon (substance);salmon allergenic extract|Salmon
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7098,7104|false|false|false|C0459210;C2702377;C4521768|Salmon (substance);salmon allergenic extract|Salmon
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7114,7117|false|false|false|C0027609|Neonatal Abstinence Syndrome|NAS
Drug|Organic Chemical|SIMPLE_SEGMENT|7114,7117|false|false|false|C0067783;C0068453|N-acetylserotonin;Tobacco containing mixture|NAS
Drug|Substance|SIMPLE_SEGMENT|7114,7117|false|false|false|C0067783;C0068453|N-acetylserotonin;Tobacco containing mixture|NAS
Finding|Finding|SIMPLE_SEGMENT|7114,7117|false|false|false|C5552704||NAS
Drug|Organic Chemical|SIMPLE_SEGMENT|7128,7141|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7128,7141|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|SIMPLE_SEGMENT|7128,7141|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7144,7147|false|false|false|C0039225|Tablet Dosage Form|TAB
Drug|Organic Chemical|SIMPLE_SEGMENT|7162,7170|false|false|false|C0040610|tramadol|TraMADol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7162,7170|false|false|false|C0040610|tramadol|TraMADol
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7162,7170|false|false|false|C1266765|Tramadol measurement (procedure)|TraMADol
Finding|Gene or Genome|SIMPLE_SEGMENT|7185,7188|false|false|false|C1422467|CIAO3 gene|PRN
Finding|Sign or Symptom|SIMPLE_SEGMENT|7189,7198|false|true|false|C0004604|Back Pain|back pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7194,7198|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|7194,7198|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|7194,7198|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7204,7220|false|false|false|C0003921;C2608262;C3853661|Artificial Tears;Lubricant Eye Drops;artificial tears (medication)|Artificial Tears
Finding|Body Substance|SIMPLE_SEGMENT|7215,7220|false|false|false|C0039409;C1547924;C1611838|Tears (substance);Tears specimen|Tears
Finding|Intellectual Product|SIMPLE_SEGMENT|7215,7220|false|false|false|C0039409;C1547924;C1611838|Tears (substance);Tears specimen|Tears
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7225,7229|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|SIMPLE_SEGMENT|7225,7229|false|false|false|C1705648|Dropping|DROP
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7230,7239|false|false|false|C0229118|Structure of both eyes|BOTH EYES
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7235,7239|false|false|false|C0015392|Eye|EYES
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7235,7239|false|false|false|C5848506||EYES
Finding|Body Substance|SIMPLE_SEGMENT|7248,7257|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|7248,7257|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|7248,7257|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|7248,7257|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|7248,7269|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7258,7269|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7258,7269|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|7258,7269|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|SIMPLE_SEGMENT|7274,7287|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7274,7287|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7274,7287|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|SIMPLE_SEGMENT|7303,7306|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7307,7311|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|7307,7311|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|7307,7311|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|SIMPLE_SEGMENT|7316,7325|false|false|false|C0085208|bupropion|BuPROPion
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7316,7325|false|false|false|C0085208|bupropion|BuPROPion
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7362,7372|false|false|false|C0006668;C0770558;C1704385;C2825090;C4520796|Calcitonin Precursor, human;Calcitonin [EPC];Recombinant Calcitonin;calcitonin;human calcitonin|Calcitonin
Drug|Hormone|SIMPLE_SEGMENT|7362,7372|false|false|false|C0006668;C0770558;C1704385;C2825090;C4520796|Calcitonin Precursor, human;Calcitonin [EPC];Recombinant Calcitonin;calcitonin;human calcitonin|Calcitonin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7362,7372|false|false|false|C0006668;C0770558;C1704385;C2825090;C4520796|Calcitonin Precursor, human;Calcitonin [EPC];Recombinant Calcitonin;calcitonin;human calcitonin|Calcitonin
Finding|Gene or Genome|SIMPLE_SEGMENT|7362,7372|false|false|false|C1367551|CALCA gene|Calcitonin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7362,7372|false|false|false|C0201924|Calcitonin measurement|Calcitonin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7362,7379|false|false|false|C0073994|salmon calcitonin|Calcitonin Salmon
Drug|Hormone|SIMPLE_SEGMENT|7362,7379|false|false|false|C0073994|salmon calcitonin|Calcitonin Salmon
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7362,7379|false|false|false|C0073994|salmon calcitonin|Calcitonin Salmon
Drug|Food|SIMPLE_SEGMENT|7373,7379|false|false|false|C0459210;C2702377;C4521768|Salmon (substance);salmon allergenic extract|Salmon
Drug|Immunologic Factor|SIMPLE_SEGMENT|7373,7379|false|false|false|C0459210;C2702377;C4521768|Salmon (substance);salmon allergenic extract|Salmon
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7373,7379|false|false|false|C0459210;C2702377;C4521768|Salmon (substance);salmon allergenic extract|Salmon
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7389,7392|false|false|false|C0027609|Neonatal Abstinence Syndrome|NAS
Drug|Organic Chemical|SIMPLE_SEGMENT|7389,7392|false|false|false|C0067783;C0068453|N-acetylserotonin;Tobacco containing mixture|NAS
Drug|Substance|SIMPLE_SEGMENT|7389,7392|false|false|false|C0067783;C0068453|N-acetylserotonin;Tobacco containing mixture|NAS
Finding|Finding|SIMPLE_SEGMENT|7389,7392|false|false|false|C5552704||NAS
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7403,7416|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Hormone|SIMPLE_SEGMENT|7403,7416|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Organic Chemical|SIMPLE_SEGMENT|7403,7416|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7403,7416|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7403,7423|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Hormone|SIMPLE_SEGMENT|7403,7423|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7403,7423|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7417,7423|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|7417,7423|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7417,7423|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|7417,7423|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7417,7423|false|false|false|C0337443|Sodium measurement|Sodium
Drug|Organic Chemical|SIMPLE_SEGMENT|7444,7455|false|false|false|C0049506|mirtazapine|Mirtazapine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7444,7455|false|false|false|C0049506|mirtazapine|Mirtazapine
Drug|Organic Chemical|SIMPLE_SEGMENT|7473,7486|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7473,7486|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|SIMPLE_SEGMENT|7473,7486|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7489,7492|false|false|false|C0039225|Tablet Dosage Form|TAB
Drug|Organic Chemical|SIMPLE_SEGMENT|7506,7514|false|false|false|C0040610|tramadol|TraMADol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7506,7514|false|false|false|C0040610|tramadol|TraMADol
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7506,7514|false|false|false|C1266765|Tramadol measurement (procedure)|TraMADol
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|7524,7527|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7524,7527|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7524,7527|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|SIMPLE_SEGMENT|7524,7527|false|false|false|C1332410|BID gene|BID
Finding|Gene or Genome|SIMPLE_SEGMENT|7528,7531|false|false|false|C1422467|CIAO3 gene|PRN
Finding|Sign or Symptom|SIMPLE_SEGMENT|7532,7541|false|true|false|C0004604|Back Pain|back pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7537,7541|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|7537,7541|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|7537,7541|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|SIMPLE_SEGMENT|7546,7557|false|false|false|C0102118|alendronate|Alendronate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7546,7557|false|false|false|C0102118|alendronate|Alendronate
Drug|Organic Chemical|SIMPLE_SEGMENT|7546,7564|false|false|false|C0700482|alendronate sodium|Alendronate Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7546,7564|false|false|false|C0700482|alendronate sodium|Alendronate Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7558,7564|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|7558,7564|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7558,7564|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|7558,7564|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7558,7564|false|false|false|C0337443|Sodium measurement|Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7583,7590|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|7583,7590|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|7583,7590|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7583,7590|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|7583,7590|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|7583,7590|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7583,7590|false|false|false|C0201925|Calcium measurement|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7583,7598|false|false|false|C3864384|Calcium 500+D|Calcium 500 + D
Drug|Vitamin|SIMPLE_SEGMENT|7583,7598|false|false|false|C3864384|Calcium 500+D|Calcium 500 + D
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7600,7607|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|7600,7607|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|7600,7607|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7600,7607|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Vitamin|SIMPLE_SEGMENT|7600,7607|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|7600,7607|false|false|false|C4553026|Calcium metabolic function|calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7600,7607|false|false|false|C0201925|Calcium measurement|calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|7600,7617|false|false|false|C0006681|calcium carbonate|calcium carbonate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7600,7617|false|false|false|C0006681|calcium carbonate|calcium carbonate
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|7608,7617|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|carbonate
Drug|Organic Chemical|SIMPLE_SEGMENT|7608,7617|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|carbonate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7608,7617|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|carbonate
Drug|Organic Chemical|SIMPLE_SEGMENT|7618,7625|false|false|false|C0042890|Vitamins|vitamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7618,7625|false|false|false|C0042890|Vitamins|vitamin
Drug|Vitamin|SIMPLE_SEGMENT|7618,7625|false|false|false|C0042890|Vitamins|vitamin
Drug|Organic Chemical|SIMPLE_SEGMENT|7618,7628|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7618,7628|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Drug|Vitamin|SIMPLE_SEGMENT|7618,7628|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|7657,7661|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7657,7661|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|7657,7661|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|7657,7661|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Drug|Organic Chemical|SIMPLE_SEGMENT|7673,7681|false|false|false|C0040610|tramadol|TraMADol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7673,7681|false|false|false|C0040610|tramadol|TraMADol
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7673,7681|false|false|false|C1266765|Tramadol measurement (procedure)|TraMADol
Finding|Gene or Genome|SIMPLE_SEGMENT|7696,7699|false|false|false|C1422467|CIAO3 gene|PRN
Finding|Sign or Symptom|SIMPLE_SEGMENT|7700,7709|false|true|false|C0004604|Back Pain|back pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7705,7709|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|7705,7709|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|7705,7709|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7715,7731|false|false|false|C0003921;C2608262;C3853661|Artificial Tears;Lubricant Eye Drops;artificial tears (medication)|Artificial Tears
Finding|Body Substance|SIMPLE_SEGMENT|7726,7731|false|false|false|C0039409;C1547924;C1611838|Tears (substance);Tears specimen|Tears
Finding|Intellectual Product|SIMPLE_SEGMENT|7726,7731|false|false|false|C0039409;C1547924;C1611838|Tears (substance);Tears specimen|Tears
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7736,7740|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|SIMPLE_SEGMENT|7736,7740|false|false|false|C1705648|Dropping|DROP
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7741,7750|false|false|false|C0229118|Structure of both eyes|BOTH EYES
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7746,7750|false|false|false|C0015392|Eye|EYES
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7746,7750|false|false|false|C5848506||EYES
Finding|Body Substance|SIMPLE_SEGMENT|7759,7768|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|7759,7768|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|7759,7768|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|7759,7768|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7759,7780|false|false|false|C4019243||Discharge Disposition
Finding|Finding|SIMPLE_SEGMENT|7759,7780|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7769,7780|false|false|false|C2926604||Disposition
Procedure|Health Care Activity|SIMPLE_SEGMENT|7769,7780|false|false|false|C0184758|Patient disposition|Disposition
Finding|Finding|SIMPLE_SEGMENT|7782,7790|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|SIMPLE_SEGMENT|7782,7790|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Procedure|Health Care Activity|SIMPLE_SEGMENT|7782,7795|false|false|false|C0023977|long-term care|Extended Care
Event|Activity|SIMPLE_SEGMENT|7791,7795|false|false|false|C1947933|care activity|Care
Finding|Finding|SIMPLE_SEGMENT|7791,7795|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|SIMPLE_SEGMENT|7791,7795|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|SIMPLE_SEGMENT|7798,7806|false|false|false|C4695111|ADMIN.FACILITY|Facility
Finding|Body Substance|SIMPLE_SEGMENT|7814,7823|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|7814,7823|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|7814,7823|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|7814,7823|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|7814,7833|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7824,7833|false|false|false|C0945731||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|7824,7833|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|7824,7833|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7824,7833|false|false|false|C0011900|Diagnosis|Diagnosis
Finding|Intellectual Product|SIMPLE_SEGMENT|7837,7842|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|Acute
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7837,7851|false|false|false|C0266807|Acute gastrointestinal hemorrhage|Acute GI Bleed
Finding|Pathologic Function|SIMPLE_SEGMENT|7843,7851|false|false|false|C0017181|Gastrointestinal Hemorrhage|GI Bleed
Finding|Pathologic Function|SIMPLE_SEGMENT|7846,7851|false|false|false|C0019080|Hemorrhage|Bleed
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|7859,7869|false|false|false|C0011570;C0011581;C0344315;C0812393|Cancer patients and suicide and depression;Depressed mood;Depressive disorder;Mental Depression|Depression
Finding|Functional Concept|SIMPLE_SEGMENT|7859,7869|false|false|false|C0460137;C1579931|Depression - motion|Depression
Finding|Sign or Symptom|SIMPLE_SEGMENT|7859,7869|false|false|false|C0460137;C1579931|Depression - motion|Depression
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7872,7884|false|false|false|C0029456|Osteoporosis|Osteoporosis
Finding|Finding|SIMPLE_SEGMENT|7872,7884|false|false|false|C2911643|Encounter due to family history of osteoporosis|Osteoporosis
Finding|Intellectual Product|SIMPLE_SEGMENT|7887,7894|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|7887,7894|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Finding|Functional Concept|SIMPLE_SEGMENT|7898,7909|false|false|false|C0332459;C4551657|Compressed structure|compression
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|7898,7909|false|false|false|C0728907|Compression|compression
Procedure|Machine Activity|SIMPLE_SEGMENT|7898,7909|false|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7898,7909|false|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Finding|Pathologic Function|SIMPLE_SEGMENT|7898,7918|false|false|false|C0521169|Compression fracture|compression fracture
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|7910,7918|false|false|false|C0016658|Fracture|fracture
Finding|Intellectual Product|SIMPLE_SEGMENT|7938,7945|false|false|false|C1547296|Chronic - Admission Level of Care Code|Chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|7938,7945|false|false|false|C1555457|Provision of recurring care for chronic illness|Chronic
Finding|Finding|SIMPLE_SEGMENT|7946,7952|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|Severe
Finding|Intellectual Product|SIMPLE_SEGMENT|7946,7952|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|Severe
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7946,7981|false|false|false|C1283368||Severe Protein Calorie Malnutrition
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7953,7960|false|false|false|C0033684|Proteins|Protein
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7953,7960|false|false|false|C0033684|Proteins|Protein
Finding|Conceptual Entity|SIMPLE_SEGMENT|7953,7960|false|false|false|C1521746|Protein Info|Protein
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7953,7960|false|false|false|C0202202|Protein measurement|Protein
Finding|Pathologic Function|SIMPLE_SEGMENT|7953,7981|false|false|false|C0033677|Protein-Energy Malnutrition|Protein Calorie Malnutrition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7969,7981|false|false|false|C0162429|Malnutrition|Malnutrition
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|7984,7992|false|false|false|C0011265;C0497327|Dementia;Presenile dementia|Dementia
Finding|Body Substance|SIMPLE_SEGMENT|7996,8005|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|7996,8005|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|7996,8005|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|7996,8005|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8006,8015|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8006,8015|false|false|false|C0012634|Disease|Condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|8006,8015|false|false|false|C1705253|Logical Condition|Condition
Finding|Mental Process|SIMPLE_SEGMENT|8017,8023|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8017,8030|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|SIMPLE_SEGMENT|8017,8030|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8024,8030|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|8024,8030|false|false|false|C1546481|What subject filter - Status|Status
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|8032,8040|false|false|false|C0009676|Confusion|Confused
Finding|Finding|SIMPLE_SEGMENT|8032,8040|false|false|false|C0683369;C1547301|Clouded consciousness;Precaution Code - Confused|Confused
Finding|Intellectual Product|SIMPLE_SEGMENT|8032,8040|false|false|false|C0683369;C1547301|Clouded consciousness;Precaution Code - Confused|Confused
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8054,8076|false|false|false|C4050479||Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|8054,8076|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|8063,8076|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|SIMPLE_SEGMENT|8063,8076|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8078,8083|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|8078,8083|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8078,8083|false|false|false|C0718338|Alert brand of caffeine|Alert
Finding|Finding|SIMPLE_SEGMENT|8078,8083|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|8078,8083|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|8078,8083|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|8088,8099|false|false|false|C1704675|Interaction|interactive
Event|Activity|SIMPLE_SEGMENT|8101,8109|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|8101,8109|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|SIMPLE_SEGMENT|8101,8109|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8110,8116|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|8110,8116|false|false|false|C1546481|What subject filter - Status|Status
Finding|Functional Concept|SIMPLE_SEGMENT|8118,8128|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|SIMPLE_SEGMENT|8118,8128|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|SIMPLE_SEGMENT|8118,8128|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|SIMPLE_SEGMENT|8118,8128|false|false|false|C1561560|ambulatory encounter|Ambulatory
Finding|Social Behavior|SIMPLE_SEGMENT|8140,8150|false|false|false|C0018896|Helping Behavior|assistance
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8154,8157|false|false|false|C1454018|AICDA protein, human|aid
Drug|Enzyme|SIMPLE_SEGMENT|8154,8157|false|false|false|C1454018|AICDA protein, human|aid
Finding|Gene or Genome|SIMPLE_SEGMENT|8154,8157|false|false|false|C1421876;C3540469|AICDA gene;AICDA wt Allele|aid
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8154,8157|false|false|false|C0021588;C0280108|AID - Artificial insemination by donor;dacarbazine/doxorubicin/ifosfamide protocol|aid
Finding|Body Substance|SIMPLE_SEGMENT|8180,8189|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|8180,8189|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|8180,8189|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|8180,8189|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8180,8202|false|false|false|C3669312||Discharge Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|8180,8202|false|false|false|C4282220|Discharge instructions|Discharge Instructions
Procedure|Health Care Activity|SIMPLE_SEGMENT|8180,8202|false|false|false|C2266673|hospital discharge instructions (treatment)|Discharge Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8190,8202|false|false|false|C3263700||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|8190,8202|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|8224,8232|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|SIMPLE_SEGMENT|8224,8232|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Intellectual Product|SIMPLE_SEGMENT|8281,8297|false|false|false|C1314977|Gastrointestinal attachment|gastrointestinal
Finding|Pathologic Function|SIMPLE_SEGMENT|8281,8306|false|false|false|C0017181|Gastrointestinal Hemorrhage|gastrointestinal bleeding
Finding|Pathologic Function|SIMPLE_SEGMENT|8298,8306|false|false|false|C0019080|Hemorrhage|bleeding
Finding|Finding|SIMPLE_SEGMENT|8389,8394|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|SIMPLE_SEGMENT|8389,8394|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Finding|SIMPLE_SEGMENT|8400,8406|false|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Finding|Functional Concept|SIMPLE_SEGMENT|8400,8406|false|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Finding|Intellectual Product|SIMPLE_SEGMENT|8400,8406|false|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Finding|Pathologic Function|SIMPLE_SEGMENT|8416,8424|false|false|false|C0019080|Hemorrhage|bleeding
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8455,8460|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|SIMPLE_SEGMENT|8455,8460|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Intellectual Product|SIMPLE_SEGMENT|8474,8480|false|false|false|C1547311|Patient Condition Code - Stable|stable
Finding|Finding|SIMPLE_SEGMENT|8495,8514|false|false|false|C2314972|Ready for discharge|ready for discharge
Finding|Body Substance|SIMPLE_SEGMENT|8505,8514|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|8505,8514|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|8505,8514|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|8505,8514|false|false|false|C0030685|Patient Discharge|discharge
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8505,8519|false|false|false|C0184713|Discharge to home|discharge home
Finding|Idea or Concept|SIMPLE_SEGMENT|8515,8519|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|8515,8519|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|8515,8519|false|false|false|C1553498|home health encounter|home
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8563,8574|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Procedure|Health Care Activity|SIMPLE_SEGMENT|8563,8574|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Finding|Finding|SIMPLE_SEGMENT|8592,8598|false|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Finding|Functional Concept|SIMPLE_SEGMENT|8592,8598|false|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Finding|Intellectual Product|SIMPLE_SEGMENT|8592,8598|false|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Finding|Pathologic Function|SIMPLE_SEGMENT|8607,8615|false|false|false|C0019080|Hemorrhage|bleeding
Finding|Classification|SIMPLE_SEGMENT|8679,8685|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|8679,8685|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|8679,8685|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|8679,8685|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|8690,8702|false|false|false|C1547426|Location Service Code - Primary Care|primary care
Procedure|Health Care Activity|SIMPLE_SEGMENT|8690,8702|false|false|false|C0033137|Primary Health Care|primary care
Event|Activity|SIMPLE_SEGMENT|8698,8702|false|false|false|C1947933|care activity|care
Finding|Finding|SIMPLE_SEGMENT|8698,8702|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|8698,8702|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|8703,8709|false|false|false|C2348314|Doctor - Title|doctor
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8744,8749|false|false|false|C2979882||goals
Finding|Idea or Concept|SIMPLE_SEGMENT|8744,8749|false|false|false|C0018017;C0679840;C1546459|What subject filter - Goals;objective (goal);treatment goals|goals
Finding|Intellectual Product|SIMPLE_SEGMENT|8744,8749|false|false|false|C0018017;C0679840;C1546459|What subject filter - Goals;objective (goal);treatment goals|goals
Procedure|Health Care Activity|SIMPLE_SEGMENT|8744,8757|false|false|false|C2930505|Goals of Care|goals of care
Event|Activity|SIMPLE_SEGMENT|8753,8757|false|false|false|C1947933|care activity|care
Finding|Finding|SIMPLE_SEGMENT|8753,8757|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|8753,8757|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Procedure|Health Care Activity|SIMPLE_SEGMENT|8761,8769|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8770,8782|false|false|false|C3263700||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|8770,8782|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

