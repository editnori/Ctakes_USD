 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|26,30
No|31,33
:|33,34
_|37,38
_|38,39
_|39,40
<EOL>|40,41
<EOL>|42,43
Admission|43,52
Date|53,57
:|57,58
_|60,61
_|61,62
_|62,63
Discharge|77,86
Date|87,91
:|91,92
_|95,96
_|96,97
_|97,98
<EOL>|98,99
<EOL>|100,101
Date|101,105
of|106,108
Birth|109,114
:|114,115
_|117,118
_|118,119
_|119,120
Sex|133,136
:|136,137
F|140,141
<EOL>|141,142
<EOL>|143,144
Service|144,151
:|151,152
MEDICINE|153,161
<EOL>|161,162
<EOL>|163,164
Allergies|164,173
:|173,174
<EOL>|175,176
No|176,178
Known|179,184
Allergies|185,194
/|195,196
Adverse|197,204
Drug|205,209
Reactions|210,219
<EOL>|219,220
<EOL>|221,222
Attending|222,231
:|231,232
_|233,234
_|234,235
_|235,236
.|236,237
<EOL>|237,238
<EOL>|239,240
Chief|240,245
Complaint|246,255
:|255,256
<EOL>|256,257
Fevers|257,263
and|264,267
chills|268,274
<EOL>|274,275
<EOL>|276,277
Major|277,282
Surgical|283,291
or|292,294
Invasive|295,303
Procedure|304,313
:|313,314
<EOL>|314,315
_|315,316
_|316,317
_|317,318
-|319,320
-|320,321
stent|322,327
exchange|328,336
<EOL>|336,337
<EOL>|337,338
<EOL>|339,340
History|340,347
of|348,350
Present|351,358
Illness|359,366
:|366,367
<EOL>|367,368
Ms.|368,371
_|372,373
_|373,374
_|374,375
is|376,378
a|379,380
_|381,382
_|382,383
_|383,384
female|385,391
with|392,396
the|397,400
past|401,405
<EOL>|405,406
medical|406,413
history|414,421
notable|422,429
for|430,433
history|434,441
of|442,444
bladder|445,452
cancer|453,459
status|460,466
<EOL>|467,468
post|468,472
<EOL>|472,473
robotic|473,480
TAH|481,484
-|484,485
BSO|485,488
,|488,489
lap|490,493
radical|494,501
cystectomy|502,512
with|513,517
ileal|518,523
loop|524,528
<EOL>|529,530
diversion|530,539
<EOL>|539,540
and|540,543
anterior|544,552
vaginectomy|553,564
in|565,567
_|568,569
_|569,570
_|570,571
complicated|572,583
by|584,586
abdominal|587,596
<EOL>|596,597
fluid|597,602
requiring|603,612
placement|613,622
of|623,625
drainage|626,634
catheters|635,644
,|644,645
further|646,653
<EOL>|653,654
complicated|654,665
by|666,668
a|669,670
severe|671,677
bilateral|678,687
hydronephrosis|688,702
requiring|703,712
<EOL>|712,713
bilateral|713,722
urostomy|723,731
tube|732,736
placement|737,746
and|747,750
then|751,755
ultimately|756,766
ureteral|767,775
<EOL>|775,776
stent|776,781
placements|782,792
with|793,797
improvement|798,809
who|810,813
presented|814,823
to|824,826
the|827,830
hospital|831,839
<EOL>|839,840
for|840,843
routine|844,851
stent|852,857
exchange|858,866
and|867,870
cystoscopy|871,881
.|881,882
The|884,887
patient|888,895
<EOL>|896,897
underwent|897,906
<EOL>|906,907
an|907,909
uncomplicated|910,923
procedure|924,933
but|934,937
then|938,942
postoperatively|943,958
in|959,961
the|962,965
PACU|966,970
<EOL>|970,971
she|971,974
developed|975,984
a|985,986
fever|987,992
to|993,995
102.4|996,1001
and|1002,1005
was|1006,1009
tachycardic|1010,1021
105|1022,1025
and|1026,1029
as|1030,1032
<EOL>|1032,1033
such|1033,1037
was|1038,1041
felt|1042,1046
to|1047,1049
need|1050,1054
admission|1055,1064
for|1065,1068
treatment|1069,1078
of|1079,1081
sepsis|1082,1088
.|1088,1089
At|1091,1093
<EOL>|1094,1095
that|1095,1099
<EOL>|1099,1100
time|1100,1104
she|1105,1108
was|1109,1112
given|1113,1118
ampicillin|1119,1129
and|1130,1133
gentamicin|1134,1144
given|1145,1150
her|1151,1154
history|1155,1162
<EOL>|1163,1164
of|1164,1166
<EOL>|1166,1167
drug|1167,1171
resistant|1172,1181
organisms|1182,1191
.|1191,1192
She|1194,1197
reported|1198,1206
at|1207,1209
that|1210,1214
time|1215,1219
she|1220,1223
was|1224,1227
<EOL>|1227,1228
feeling|1228,1235
feverish|1236,1244
and|1245,1248
chills|1249,1255
with|1256,1260
nausea|1261,1267
and|1268,1271
vomiting|1272,1280
x1|1281,1283
.|1283,1284
She|1286,1289
<EOL>|1289,1290
received|1290,1298
IV|1299,1301
fluids|1302,1308
and|1309,1312
her|1313,1316
IV|1317,1319
antibiotics|1320,1331
and|1332,1335
her|1336,1339
symptoms|1340,1348
<EOL>|1348,1349
improved|1349,1357
.|1357,1358
She|1360,1363
was|1364,1367
admitted|1368,1376
to|1377,1379
the|1380,1383
medical|1384,1391
service|1392,1399
for|1400,1403
further|1404,1411
<EOL>|1411,1412
evaluation|1412,1422
and|1423,1426
management|1427,1437
<EOL>|1437,1438
<EOL>|1438,1439
On|1439,1441
the|1442,1445
floor|1446,1451
the|1452,1455
patient|1456,1463
reports|1464,1471
that|1472,1476
she|1477,1480
continues|1481,1490
to|1491,1493
have|1494,1498
<EOL>|1498,1499
persistent|1499,1509
chills|1510,1516
.|1516,1517
She|1519,1522
feels|1523,1528
slightly|1529,1537
nauseous|1538,1546
.|1546,1547
She|1549,1552
denies|1553,1559
any|1560,1563
<EOL>|1563,1564
abdominal|1564,1573
pain|1574,1578
.|1578,1579
She|1581,1584
otherwise|1585,1594
reports|1595,1602
that|1603,1607
she|1608,1611
is|1612,1614
feeling|1615,1622
<EOL>|1623,1624
better|1624,1630
<EOL>|1630,1631
than|1631,1635
she|1636,1639
did|1640,1643
immediately|1644,1655
postprocedural|1656,1670
but|1671,1674
is|1675,1677
still|1678,1683
<EOL>|1683,1684
significantly|1684,1697
off|1698,1701
of|1702,1704
her|1705,1708
baseline|1709,1717
.|1717,1718
She|1720,1723
reports|1724,1731
that|1732,1736
she|1737,1740
has|1741,1744
a|1745,1746
<EOL>|1746,1747
history|1747,1754
of|1755,1757
urinary|1758,1765
tract|1766,1771
infections|1772,1782
and|1783,1786
was|1787,1790
most|1791,1795
recently|1796,1804
on|1805,1807
<EOL>|1807,1808
ciprofloxacin|1808,1821
and|1822,1825
_|1826,1827
_|1827,1828
_|1828,1829
.|1829,1830
She|1832,1835
reports|1836,1843
that|1844,1848
she|1849,1852
was|1853,1856
on|1857,1859
<EOL>|1859,1860
this|1860,1864
medication|1865,1875
for|1876,1879
7|1880,1881
-|1881,1882
day|1882,1885
course|1886,1892
.|1892,1893
No|1895,1897
_|1898,1899
_|1899,1900
_|1900,1901
acute|1902,1907
complaints|1908,1918
.|1918,1919
<EOL>|1919,1920
<EOL>|1920,1921
<EOL>|1922,1923
Past|1923,1927
Medical|1928,1935
History|1936,1943
:|1943,1944
<EOL>|1944,1945
-|1945,1946
Hypertension|1947,1959
<EOL>|1961,1962
-|1963,1964
s|1965,1966
/|1966,1967
p|1967,1968
lap|1969,1972
chole|1973,1978
<EOL>|1980,1981
-|1982,1983
s|1984,1985
/|1985,1986
p|1986,1987
left|1988,1992
knee|1993,1997
replacement|1998,2009
<EOL>|2011,2012
-|2013,2014
s|2015,2016
/|2016,2017
p|2017,2018
laminectomy|2019,2030
of|2031,2033
L5|2034,2036
-|2036,2037
S1|2037,2039
at|2040,2042
age|2043,2046
_|2047,2048
_|2048,2049
_|2049,2050
<EOL>|2052,2053
-|2054,2055
Bladder|2056,2063
Cancer|2064,2070
high|2071,2075
grade|2076,2081
TCC|2082,2085
,|2085,2086
T1|2087,2089
diagnosed|2090,2099
in|2100,2102
_|2103,2104
_|2104,2105
_|2105,2106
,|2106,2107
then|2108,2112
<EOL>|2113,2114
_|2114,2115
_|2115,2116
_|2116,2117
pelvic|2118,2124
MRI|2125,2128
w|2129,2130
/|2130,2131
invasion|2131,2139
into|2140,2144
bladder|2145,2152
wall|2153,2157
,|2157,2158
perivesical|2159,2170
<EOL>|2171,2172
soft|2172,2176
tissue|2177,2183
and|2184,2187
anterior|2188,2196
vaginal|2197,2204
wall|2205,2209
c|2210,2211
/|2211,2212
w|2212,2213
T4|2214,2216
staging|2217,2224
<EOL>|2226,2227
-|2228,2229
s|2230,2231
/|2231,2232
p|2232,2233
hysterectomy|2234,2246
and|2247,2250
bilateral|2251,2260
oophorectomy|2261,2273
for|2274,2277
large|2278,2283
uterus|2284,2290
<EOL>|2291,2292
w|2292,2293
/|2293,2294
fibroid|2294,2301
,|2301,2302
s|2303,2304
/|2304,2305
p|2305,2306
laparascopic|2307,2319
b|2320,2321
/|2321,2322
l|2322,2323
pelvic|2324,2330
lymph|2331,2336
node|2337,2341
resection|2342,2351
,|2351,2352
s|2353,2354
/|2354,2355
p|2355,2356
<EOL>|2357,2358
<EOL>|2358,2359
radical|2359,2366
cystectomy|2367,2377
and|2378,2381
anterior|2382,2390
vaginectomy|2391,2402
with|2403,2407
vaginal|2408,2415
<EOL>|2416,2417
reconstruction|2417,2431
with|2432,2436
ileal|2437,2442
conduit|2443,2450
creation|2451,2459
_|2460,2461
_|2461,2462
_|2462,2463
,|2463,2464
course|2465,2471
<EOL>|2472,2473
complicated|2473,2484
by|2485,2487
bacteremia|2488,2498
and|2499,2502
development|2503,2514
of|2515,2517
intra-abdominal|2518,2533
<EOL>|2534,2535
fluid|2535,2540
collection|2541,2551
,|2551,2552
no|2553,2555
s|2556,2557
/|2557,2558
p|2558,2559
drain|2560,2565
placement|2566,2575
by|2576,2578
_|2579,2580
_|2580,2581
_|2581,2582
_|2583,2584
_|2584,2585
_|2585,2586
<EOL>|2588,2589
-|2590,2591
h|2592,2593
/|2593,2594
o|2594,2595
LLE|2596,2599
DVT|2600,2603
and|2604,2607
PE|2608,2610
no|2611,2613
longer|2614,2620
on|2621,2623
anticoagulation|2624,2639
.|2639,2640
<EOL>|2641,2642
<EOL>|2643,2644
Social|2644,2650
History|2651,2658
:|2658,2659
<EOL>|2659,2660
_|2660,2661
_|2661,2662
_|2662,2663
<EOL>|2663,2664
Family|2664,2670
History|2671,2678
:|2678,2679
<EOL>|2679,2680
Negative|2680,2688
for|2689,2692
bladder|2693,2700
CA|2701,2703
.|2703,2704
<EOL>|2704,2705
<EOL>|2705,2706
<EOL>|2707,2708
Physical|2708,2716
Exam|2717,2721
:|2721,2722
<EOL>|2722,2723
ADMISSION|2723,2732
EXAM|2733,2737
:|2737,2738
<EOL>|2738,2739
<EOL>|2739,2740
VITALS|2740,2746
:|2746,2747
_|2748,2749
_|2749,2750
_|2750,2751
2227|2752,2756
Temp|2757,2761
:|2761,2762
99.3|2763,2767
PO|2768,2770
BP|2771,2773
:|2773,2774
119|2775,2778
/|2778,2779
54|2779,2781
HR|2782,2784
:|2784,2785
80|2786,2788
RR|2789,2791
:|2791,2792
16|2793,2795
O2|2796,2798
<EOL>|2798,2799
sat|2799,2802
:|2802,2803
98|2804,2806
%|2806,2807
O2|2808,2810
delivery|2811,2819
:|2819,2820
RA|2821,2823
Dyspnea|2824,2831
:|2831,2832
0|2833,2834
RASS|2835,2839
:|2839,2840
0|2841,2842
Pain|2843,2847
Score|2848,2853
:|2853,2854
_|2855,2856
_|2856,2857
_|2857,2858
<EOL>|2859,2860
GENERAL|2860,2867
:|2867,2868
Alert|2869,2874
and|2875,2878
in|2879,2881
no|2882,2884
apparent|2885,2893
distress|2894,2902
,|2902,2903
facial|2904,2910
twitches|2911,2919
<EOL>|2919,2920
EYES|2920,2924
:|2924,2925
Anicteric|2926,2935
,|2935,2936
pupils|2937,2943
equally|2944,2951
round|2952,2957
<EOL>|2957,2958
ENT|2958,2961
:|2961,2962
Ears|2963,2967
and|2968,2971
nose|2972,2976
without|2977,2984
visible|2985,2992
erythema|2993,3001
,|3001,3002
masses|3003,3009
,|3009,3010
or|3011,3013
trauma|3014,3020
.|3020,3021
<EOL>|3022,3023
Oropharynx|3023,3033
without|3034,3041
visible|3042,3049
lesion|3050,3056
,|3056,3057
erythema|3058,3066
or|3067,3069
exudate|3070,3077
<EOL>|3077,3078
CV|3078,3080
:|3080,3081
Heart|3082,3087
regular|3088,3095
,|3095,3096
no|3097,3099
murmur|3100,3106
,|3106,3107
no|3108,3110
S3|3111,3113
,|3113,3114
no|3115,3117
S4|3118,3120
.|3120,3121
No|3123,3125
JVD|3126,3129
.|3129,3130
<EOL>|3130,3131
RESP|3131,3135
:|3135,3136
Lungs|3137,3142
clear|3143,3148
to|3149,3151
auscultation|3152,3164
with|3165,3169
good|3170,3174
air|3175,3178
movement|3179,3187
<EOL>|3187,3188
bilaterally|3188,3199
.|3199,3200
Breathing|3202,3211
is|3212,3214
non-labored|3215,3226
<EOL>|3226,3227
GI|3227,3229
:|3229,3230
Abdomen|3231,3238
soft|3239,3243
,|3243,3244
non-distended|3245,3258
,|3258,3259
non-tender|3260,3270
to|3271,3273
palpation|3274,3283
.|3283,3284
Bowel|3286,3291
<EOL>|3291,3292
sounds|3292,3298
present|3299,3306
.|3306,3307
No|3309,3311
HSM|3312,3315
<EOL>|3315,3316
GU|3316,3318
:|3318,3319
No|3320,3322
suprapubic|3323,3333
fullness|3334,3342
or|3343,3345
tenderness|3346,3356
to|3357,3359
palpation|3360,3369
,|3369,3370
foley|3371,3376
<EOL>|3376,3377
catheter|3377,3385
in|3386,3388
place|3389,3394
<EOL>|3394,3395
MSK|3395,3398
:|3398,3399
Neck|3400,3404
supple|3405,3411
,|3411,3412
moves|3413,3418
all|3419,3422
extremities|3423,3434
,|3434,3435
strength|3436,3444
grossly|3445,3452
full|3453,3457
<EOL>|3457,3458
and|3458,3461
symmetric|3462,3471
bilaterally|3472,3483
in|3484,3486
all|3487,3490
limbs|3491,3496
<EOL>|3496,3497
SKIN|3497,3501
:|3501,3502
No|3503,3505
rashes|3506,3512
or|3513,3515
ulcerations|3516,3527
noted|3528,3533
<EOL>|3533,3534
NEURO|3534,3539
:|3539,3540
Alert|3541,3546
,|3546,3547
oriented|3548,3556
,|3556,3557
face|3558,3562
symmetric|3563,3572
,|3572,3573
gaze|3574,3578
conjugate|3579,3588
with|3589,3593
<EOL>|3594,3595
EOMI|3595,3599
,|3599,3600
<EOL>|3600,3601
speech|3601,3607
fluent|3608,3614
,|3614,3615
moves|3616,3621
all|3622,3625
limbs|3626,3631
,|3631,3632
sensation|3633,3642
to|3643,3645
light|3646,3651
touch|3652,3657
grossly|3658,3665
<EOL>|3665,3666
intact|3666,3672
throughout|3673,3683
<EOL>|3683,3684
PSYCH|3684,3689
:|3689,3690
pleasant|3691,3699
,|3699,3700
appropriate|3701,3712
affect|3713,3719
<EOL>|3719,3720
<EOL>|3720,3721
DISCHARGE|3721,3730
EXAM|3731,3735
:|3735,3736
<EOL>|3736,3737
<EOL>|3737,3738
AVSS|3738,3742
,|3742,3743
ambulating|3744,3754
comfortably|3755,3766
at|3767,3769
baseline|3770,3778
.|3778,3779
Urostomy|3780,3788
bag|3789,3792
in|3793,3795
place|3796,3801
<EOL>|3802,3803
with|3803,3807
no|3808,3810
surround|3811,3819
erythema|3820,3828
or|3829,3831
pain|3832,3836
.|3836,3837
<EOL>|3837,3838
<EOL>|3839,3840
Pertinent|3840,3849
Results|3850,3857
:|3857,3858
<EOL>|3858,3859
LABORATORY|3859,3869
RESULTS|3870,3877
:|3877,3878
<EOL>|3878,3879
<EOL>|3879,3880
_|3880,3881
_|3881,3882
_|3882,3883
05|3884,3886
:|3886,3887
30AM|3887,3891
BLOOD|3892,3897
WBC|3898,3901
-|3901,3902
16|3902,3904
.|3904,3905
5|3905,3906
*|3906,3907
RBC|3908,3911
-|3911,3912
3|3912,3913
.|3913,3914
23|3914,3916
*|3916,3917
Hgb|3918,3921
-|3921,3922
9|3922,3923
.|3923,3924
8|3924,3925
*|3925,3926
Hct|3927,3930
-|3930,3931
31|3931,3933
.|3933,3934
8|3934,3935
*|3935,3936
<EOL>|3937,3938
MCV|3938,3941
-|3941,3942
99|3942,3944
*|3944,3945
MCH|3946,3949
-|3949,3950
30.3|3950,3954
MCHC|3955,3959
-|3959,3960
30|3960,3962
.|3962,3963
8|3963,3964
*|3964,3965
RDW|3966,3969
-|3969,3970
14.5|3970,3974
RDWSD|3975,3980
-|3980,3981
52|3981,3983
.|3983,3984
3|3984,3985
*|3985,3986
Plt|3987,3990
_|3991,3992
_|3992,3993
_|3993,3994
<EOL>|3994,3995
_|3995,3996
_|3996,3997
_|3997,3998
06|3999,4001
:|4001,4002
09AM|4002,4006
BLOOD|4007,4012
WBC|4013,4016
-|4016,4017
14|4017,4019
.|4019,4020
1|4020,4021
*|4021,4022
RBC|4023,4026
-|4026,4027
3|4027,4028
.|4028,4029
39|4029,4031
*|4031,4032
Hgb|4033,4036
-|4036,4037
10|4037,4039
.|4039,4040
2|4040,4041
*|4041,4042
Hct|4043,4046
-|4046,4047
33|4047,4049
.|4049,4050
2|4050,4051
*|4051,4052
<EOL>|4053,4054
MCV|4054,4057
-|4057,4058
98|4058,4060
MCH|4061,4064
-|4064,4065
30.1|4065,4069
MCHC|4070,4074
-|4074,4075
30|4075,4077
.|4077,4078
7|4078,4079
*|4079,4080
RDW|4081,4084
-|4084,4085
14.6|4085,4089
RDWSD|4090,4095
-|4095,4096
52|4096,4098
.|4098,4099
7|4099,4100
*|4100,4101
Plt|4102,4105
_|4106,4107
_|4107,4108
_|4108,4109
<EOL>|4109,4110
_|4110,4111
_|4111,4112
_|4112,4113
06|4114,4116
:|4116,4117
10AM|4117,4121
BLOOD|4122,4127
WBC|4128,4131
-|4131,4132
10.0|4132,4136
RBC|4137,4140
-|4140,4141
3|4141,4142
.|4142,4143
55|4143,4145
*|4145,4146
Hgb|4147,4150
-|4150,4151
10|4151,4153
.|4153,4154
5|4154,4155
*|4155,4156
Hct|4157,4160
-|4160,4161
33|4161,4163
.|4163,4164
6|4164,4165
*|4165,4166
<EOL>|4167,4168
MCV|4168,4171
-|4171,4172
95|4172,4174
MCH|4175,4178
-|4178,4179
29.6|4179,4183
MCHC|4184,4188
-|4188,4189
31|4189,4191
.|4191,4192
3|4192,4193
*|4193,4194
RDW|4195,4198
-|4198,4199
14.1|4199,4203
RDWSD|4204,4209
-|4209,4210
49|4210,4212
.|4212,4213
9|4213,4214
*|4214,4215
Plt|4216,4219
_|4220,4221
_|4221,4222
_|4222,4223
<EOL>|4223,4224
_|4224,4225
_|4225,4226
_|4226,4227
05|4228,4230
:|4230,4231
30AM|4231,4235
BLOOD|4236,4241
Glucose|4242,4249
-|4249,4250
115|4250,4253
*|4253,4254
UreaN|4255,4260
-|4260,4261
34|4261,4263
*|4263,4264
Creat|4265,4270
-|4270,4271
1|4271,4272
.|4272,4273
6|4273,4274
*|4274,4275
Na|4276,4278
-|4278,4279
142|4279,4282
<EOL>|4283,4284
K|4284,4285
-|4285,4286
4.2|4286,4289
Cl|4290,4292
-|4292,4293
106|4293,4296
HCO3|4297,4301
-|4301,4302
22|4302,4304
AnGap|4305,4310
-|4310,4311
14|4311,4313
<EOL>|4313,4314
_|4314,4315
_|4315,4316
_|4316,4317
06|4318,4320
:|4320,4321
10AM|4321,4325
BLOOD|4326,4331
Glucose|4332,4339
-|4339,4340
99|4340,4342
UreaN|4343,4348
-|4348,4349
29|4349,4351
*|4351,4352
Creat|4353,4358
-|4358,4359
1|4359,4360
.|4360,4361
3|4361,4362
*|4362,4363
Na|4364,4366
-|4366,4367
141|4367,4370
<EOL>|4371,4372
K|4372,4373
-|4373,4374
3.8|4374,4377
Cl|4378,4380
-|4380,4381
104|4381,4384
HCO3|4385,4389
-|4389,4390
23|4390,4392
AnGap|4393,4398
-|4398,4399
14|4399,4401
<EOL>|4401,4402
_|4402,4403
_|4403,4404
_|4404,4405
05|4406,4408
:|4408,4409
30AM|4409,4413
BLOOD|4414,4419
Calcium|4420,4427
-|4427,4428
8|4428,4429
.|4429,4430
1|4430,4431
*|4431,4432
Phos|4433,4437
-|4437,4438
3.4|4438,4441
Mg|4442,4444
-|4444,4445
1.8|4445,4448
<EOL>|4448,4449
<EOL>|4449,4450
MICROBIOLOGY|4450,4462
:|4462,4463
<EOL>|4463,4464
<EOL>|4464,4465
_|4465,4466
_|4466,4467
_|4467,4468
3|4469,4470
:|4470,4471
00|4471,4473
pm|4474,4476
URINE|4477,4482
Site|4487,4491
:|4491,4492
CYSTOSCOPY|4493,4503
RIGHT|4509,4514
KIDNEY|4515,4521
<EOL>|4522,4523
WASH|4523,4527
.|4527,4528
<EOL>|4529,4530
<EOL>|4530,4531
*|4559,4560
*|4560,4561
FINAL|4561,4566
REPORT|4567,4573
_|4574,4575
_|4575,4576
_|4576,4577
<EOL>|4577,4578
<EOL>|4578,4579
URINE|4582,4587
CULTURE|4588,4595
(|4596,4597
Final|4597,4602
_|4603,4604
_|4604,4605
_|4605,4606
:|4606,4607
<EOL>|4608,4609
ENTEROCOCCUS|4615,4627
FAECIUM|4628,4635
.|4635,4636
>|4640,4641
10,000|4641,4647
CFU|4648,4651
/|4651,4652
ML|4652,4654
.|4654,4655
<EOL>|4656,4657
_|4666,4667
_|4667,4668
_|4668,4669
(|4670,4671
_|4671,4672
_|4672,4673
_|4673,4674
)|4674,4675
REQUESTS|4676,4684
SUSCEPTIBILITY|4685,4699
TESTING|4700,4707
<EOL>|4708,4709
_|4709,4710
_|4710,4711
_|4711,4712
.|4712,4713
<EOL>|4714,4715
STAPHYLOCOCCUS|4721,4735
,|4735,4736
COAGULASE|4737,4746
NEGATIVE|4747,4755
.|4755,4756
1,000|4760,4765
-|4766,4767
10,000|4768,4774
<EOL>|4775,4776
CFU|4776,4779
/|4779,4780
ML|4780,4782
.|4782,4783
<EOL>|4784,4785
CORYNEBACTERIUM|4791,4806
SPECIES|4807,4814
(|4815,4816
DIPHTHEROIDS|4816,4828
)|4828,4829
.|4829,4830
1,000|4834,4839
-|4840,4841
10,000|4842,4848
<EOL>|4849,4850
CFU|4850,4853
/|4853,4854
ML|4854,4856
.|4856,4857
<EOL>|4858,4859
<EOL>|4859,4860
SENSITIVITIES|4890,4903
:|4903,4904
MIC|4905,4908
expressed|4909,4918
in|4919,4921
<EOL>|4922,4923
MCG|4923,4926
/|4926,4927
ML|4927,4929
<EOL>|4929,4930
<EOL>|4952,4953
_|4953,4954
_|4954,4955
_|4955,4956
_|4956,4957
_|4957,4958
_|4958,4959
_|4959,4960
_|4960,4961
_|4961,4962
_|4962,4963
_|4963,4964
_|4964,4965
_|4965,4966
_|4966,4967
_|4967,4968
_|4968,4969
_|4969,4970
_|4970,4971
_|4971,4972
_|4972,4973
_|4973,4974
_|4974,4975
_|4975,4976
_|4976,4977
_|4977,4978
_|4978,4979
_|4979,4980
_|4980,4981
_|4981,4982
_|4982,4983
_|4983,4984
_|4984,4985
_|4985,4986
_|4986,4987
_|4987,4988
_|4988,4989
_|4989,4990
_|4990,4991
_|4991,4992
_|4992,4993
_|4993,4994
_|4994,4995
_|4995,4996
_|4996,4997
_|4997,4998
_|4998,4999
_|4999,5000
_|5000,5001
_|5001,5002
_|5002,5003
_|5003,5004
_|5004,5005
_|5005,5006
_|5006,5007
_|5007,5008
_|5008,5009
_|5009,5010
<EOL>|5010,5011
ENTEROCOCCUS|5040,5052
FAECIUM|5053,5060
<EOL>|5060,5061
||5090,5091
<EOL>|5094,5095
AMPICILLIN|5095,5105
-|5105,5106
-|5106,5107
-|5107,5108
-|5108,5109
-|5109,5110
-|5110,5111
-|5111,5112
-|5112,5113
-|5113,5114
-|5114,5115
-|5115,5116
-|5116,5117
8|5122,5123
S|5124,5125
<EOL>|5125,5126
NITROFURANTOIN|5126,5140
-|5140,5141
-|5141,5142
-|5142,5143
-|5143,5144
-|5144,5145
-|5145,5146
-|5146,5147
-|5147,5148
<|5150,5151
=|5151,5152
16|5152,5154
S|5155,5156
<EOL>|5156,5157
TETRACYCLINE|5157,5169
-|5169,5170
-|5170,5171
-|5171,5172
-|5172,5173
-|5173,5174
-|5174,5175
-|5175,5176
-|5176,5177
-|5177,5178
-|5178,5179
=|5181,5182
>|5182,5183
16|5183,5185
R|5186,5187
<EOL>|5187,5188
VANCOMYCIN|5188,5198
-|5198,5199
-|5199,5200
-|5200,5201
-|5201,5202
-|5202,5203
-|5203,5204
-|5204,5205
-|5205,5206
-|5206,5207
-|5207,5208
-|5208,5209
-|5209,5210
2|5215,5216
S|5217,5218
<EOL>|5218,5219
<EOL>|5219,5220
Blood|5220,5225
cultures|5226,5234
NGTD|5235,5239
<EOL>|5239,5240
<EOL>|5241,5242
Brief|5242,5247
Hospital|5248,5256
Course|5257,5263
:|5263,5264
<EOL>|5264,5265
Ms.|5265,5268
_|5269,5270
_|5270,5271
_|5271,5272
was|5273,5276
admitted|5277,5285
with|5286,5290
sepsis|5291,5297
from|5298,5302
a|5303,5304
urinary|5305,5312
tract|5313,5318
<EOL>|5319,5320
infection|5320,5329
after|5330,5335
her|5336,5339
stent|5340,5345
exchange|5346,5354
.|5354,5355
She|5356,5359
was|5360,5363
placed|5364,5370
empirically|5371,5382
<EOL>|5383,5384
on|5384,5386
vancomycin|5387,5397
and|5398,5401
cefepime|5402,5410
(|5411,5412
narrowed|5412,5420
to|5421,5423
vanc|5424,5428
/|5428,5429
ceftriaxone|5429,5440
on|5441,5443
<EOL>|5444,5445
HD|5445,5447
#|5447,5448
1|5448,5449
)|5449,5450
,|5450,5451
because|5452,5459
of|5460,5462
her|5463,5466
history|5467,5474
of|5475,5477
resistant|5478,5487
organisms|5488,5497
.|5497,5498
She|5499,5502
<EOL>|5503,5504
rapidly|5504,5511
improved|5512,5520
.|5520,5521
Her|5522,5525
urine|5526,5531
grew|5532,5536
E.|5537,5539
faecium|5540,5547
,|5547,5548
sensitive|5549,5558
to|5559,5561
<EOL>|5562,5563
ampicillin|5563,5573
.|5573,5574
Therefore|5575,5584
,|5584,5585
a|5586,5587
PICC|5588,5592
line|5593,5597
was|5598,5601
placed|5602,5608
,|5608,5609
and|5610,5613
she|5614,5617
will|5618,5622
<EOL>|5623,5624
complete|5624,5632
two|5633,5636
weeks|5637,5642
total|5643,5648
of|5649,5651
ampicillin|5652,5662
for|5663,5666
a|5667,5668
complicated|5669,5680
urinary|5681,5688
<EOL>|5689,5690
tract|5690,5695
infection|5696,5705
(|5706,5707
additional|5707,5717
day|5718,5721
days|5722,5726
)|5726,5727
.|5727,5728
She|5729,5732
will|5733,5737
follow|5738,5744
up|5745,5747
with|5748,5752
<EOL>|5753,5754
Dr.|5754,5757
_|5758,5759
_|5759,5760
_|5760,5761
as|5762,5764
an|5765,5767
outpatient|5768,5778
.|5778,5779
She|5780,5783
will|5784,5788
stop|5789,5793
her|5794,5797
prophylactic|5798,5810
TMP|5811,5814
<EOL>|5815,5816
while|5816,5821
on|5822,5824
ampicillin|5825,5835
,|5835,5836
but|5837,5840
then|5841,5845
resume|5846,5852
after|5853,5858
finishing|5859,5868
her|5869,5872
course|5873,5879
.|5879,5880
<EOL>|5880,5881
-|5881,5882
ampicillin|5883,5893
500|5894,5897
mg|5898,5900
TID|5901,5904
x|5905,5906
9|5907,5908
additional|5909,5919
days|5920,5924
<EOL>|5924,5925
-|5925,5926
restart|5927,5934
TMP|5935,5938
100|5939,5942
mg|5943,5945
daily|5946,5951
for|5952,5955
ppx|5956,5959
after|5960,5965
antibiotic|5966,5976
course|5977,5983
<EOL>|5983,5984
-|5984,5985
follow|5986,5992
up|5993,5995
with|5996,6000
Dr.|6001,6004
_|6005,6006
_|6006,6007
_|6007,6008
<EOL>|6008,6009
<EOL>|6009,6010
_|6010,6011
_|6011,6012
_|6012,6013
problems|6014,6022
addressed|6023,6032
this|6033,6037
hospitalization|6038,6053
:|6053,6054
<EOL>|6054,6055
<EOL>|6055,6056
1.|6056,6058
_|6059,6060
_|6060,6061
_|6061,6062
.|6062,6063
Ms.|6064,6067
_|6068,6069
_|6069,6070
_|6070,6071
initially|6072,6081
had|6082,6085
an|6086,6088
_|6089,6090
_|6090,6091
_|6091,6092
,|6092,6093
likely|6094,6100
prerenal|6101,6109
from|6110,6114
<EOL>|6115,6116
her|6116,6119
sepsis|6120,6126
.|6126,6127
She|6128,6131
received|6132,6140
IV|6141,6143
fluids|6144,6150
and|6151,6154
antibiotics|6155,6166
as|6167,6169
above|6170,6175
,|6175,6176
and|6177,6180
<EOL>|6181,6182
her|6182,6185
creatinine|6186,6196
down|6197,6201
-|6201,6202
trended|6202,6209
.|6209,6210
Losartan|6211,6219
was|6220,6223
initially|6224,6233
held|6234,6238
,|6238,6239
but|6240,6243
<EOL>|6244,6245
restarted|6245,6254
on|6255,6257
discharge|6258,6267
.|6267,6268
<EOL>|6268,6269
<EOL>|6269,6270
2.|6270,6272
Hyperlipidemia|6273,6287
:|6287,6288
continued|6289,6298
atorvastatin|6299,6311
10|6312,6314
mg|6315,6317
daily|6318,6323
<EOL>|6323,6324
<EOL>|6324,6325
3.|6325,6327
Hypothyroidism|6328,6342
:|6342,6343
continue|6344,6352
levothyroxine|6353,6366
175|6367,6370
mcg|6371,6374
daily|6375,6380
<EOL>|6380,6381
<EOL>|6381,6382
>|6382,6383
30|6384,6386
minutes|6387,6394
spent|6395,6400
on|6401,6403
discharge|6404,6413
activities|6414,6424
.|6424,6425
<EOL>|6425,6426
<EOL>|6426,6427
<EOL>|6428,6429
Medications|6429,6440
on|6441,6443
Admission|6444,6453
:|6453,6454
<EOL>|6454,6455
The|6455,6458
Preadmission|6459,6471
Medication|6472,6482
list|6483,6487
is|6488,6490
accurate|6491,6499
and|6500,6503
complete|6504,6512
.|6512,6513
<EOL>|6513,6514
1.|6514,6516
Acetaminophen|6517,6530
650|6531,6534
mg|6535,6537
PO|6538,6540
Q6H|6541,6544
:|6544,6545
PRN|6545,6548
Pain|6549,6553
-|6554,6555
Mild|6556,6560
/|6560,6561
Fever|6561,6566
<EOL>|6567,6568
2.|6568,6570
Atorvastatin|6571,6583
10|6584,6586
mg|6587,6589
PO|6590,6592
QPM|6593,6596
<EOL>|6597,6598
3.|6598,6600
Cyanocobalamin|6601,6615
1000|6616,6620
mcg|6621,6624
PO|6625,6627
DAILY|6628,6633
<EOL>|6634,6635
4.|6635,6637
Docusate|6638,6646
Sodium|6647,6653
100|6654,6657
mg|6658,6660
PO|6661,6663
BID|6664,6667
<EOL>|6668,6669
5.|6669,6671
Levothyroxine|6672,6685
Sodium|6686,6692
175|6693,6696
mcg|6697,6700
PO|6701,6703
DAILY|6704,6709
<EOL>|6710,6711
6.|6711,6713
LORazepam|6714,6723
0.5|6724,6727
mg|6728,6730
PO|6731,6733
Q12H|6734,6738
:|6738,6739
PRN|6739,6742
anxiety|6743,6750
<EOL>|6751,6752
7.|6752,6754
Losartan|6755,6763
Potassium|6764,6773
50|6774,6776
mg|6777,6779
PO|6780,6782
BID|6783,6786
<EOL>|6787,6788
8.|6788,6790
Multivitamins|6791,6804
1|6805,6806
TAB|6807,6810
PO|6811,6813
DAILY|6814,6819
<EOL>|6820,6821
9.|6821,6823
Polyethylene|6824,6836
Glycol|6837,6843
17|6844,6846
g|6847,6848
PO|6849,6851
DAILY|6852,6857
:|6857,6858
PRN|6858,6861
Constipation|6862,6874
-|6875,6876
First|6877,6882
<EOL>|6883,6884
Line|6884,6888
<EOL>|6889,6890
10.|6890,6893
Trimethoprim|6894,6906
100|6907,6910
mg|6911,6913
PO|6914,6916
Q24H|6917,6921
<EOL>|6922,6923
<EOL>|6923,6924
<EOL>|6925,6926
Discharge|6926,6935
Medications|6936,6947
:|6947,6948
<EOL>|6948,6949
1.|6949,6951
Ampicillin|6953,6963
500|6964,6967
mg|6968,6970
IV|6971,6973
Q8H|6974,6977
<EOL>|6978,6979
RX|6979,6981
*|6982,6983
ampicillin|6983,6993
sodium|6994,7000
500|7001,7004
mg|7005,7007
500|7008,7011
mg|7012,7014
IV|7015,7017
Every|7018,7023
eight|7024,7029
hours|7030,7035
Disp|7036,7040
<EOL>|7041,7042
#|7042,7043
*|7043,7044
15|7044,7046
Vial|7047,7051
Refills|7052,7059
:|7059,7060
*|7060,7061
0|7061,7062
<EOL>|7062,7063
RX|7063,7065
*|7066,7067
ampicillin|7067,7077
sodium|7078,7084
500|7085,7088
mg|7089,7091
500|7092,7095
mg|7096,7098
IV|7099,7101
Every|7102,7107
eight|7108,7113
hours|7114,7119
Disp|7120,7124
<EOL>|7125,7126
#|7126,7127
*|7127,7128
27|7128,7130
Vial|7131,7135
Refills|7136,7143
:|7143,7144
*|7144,7145
0|7145,7146
<EOL>|7147,7148
2.|7148,7150
Acetaminophen|7152,7165
650|7166,7169
mg|7170,7172
PO|7173,7175
Q6H|7176,7179
:|7179,7180
PRN|7180,7183
Pain|7184,7188
-|7189,7190
Mild|7191,7195
/|7195,7196
Fever|7196,7201
<EOL>|7203,7204
3.|7204,7206
Atorvastatin|7208,7220
10|7221,7223
mg|7224,7226
PO|7227,7229
QPM|7230,7233
<EOL>|7235,7236
4.|7236,7238
Cyanocobalamin|7240,7254
1000|7255,7259
mcg|7260,7263
PO|7264,7266
DAILY|7267,7272
<EOL>|7274,7275
5.|7275,7277
Docusate|7279,7287
Sodium|7288,7294
100|7295,7298
mg|7299,7301
PO|7302,7304
BID|7305,7308
<EOL>|7310,7311
6.|7311,7313
Levothyroxine|7315,7328
Sodium|7329,7335
175|7336,7339
mcg|7340,7343
PO|7344,7346
DAILY|7347,7352
<EOL>|7354,7355
7.|7355,7357
LORazepam|7359,7368
0.5|7369,7372
mg|7373,7375
PO|7376,7378
Q12H|7379,7383
:|7383,7384
PRN|7384,7387
anxiety|7388,7395
<EOL>|7397,7398
8.|7398,7400
Losartan|7402,7410
Potassium|7411,7420
50|7421,7423
mg|7424,7426
PO|7427,7429
BID|7430,7433
<EOL>|7435,7436
9.|7436,7438
Multivitamins|7440,7453
1|7454,7455
TAB|7456,7459
PO|7460,7462
DAILY|7463,7468
<EOL>|7470,7471
10.|7471,7474
Polyethylene|7476,7488
Glycol|7489,7495
17|7496,7498
g|7499,7500
PO|7501,7503
DAILY|7504,7509
:|7509,7510
PRN|7510,7513
Constipation|7514,7526
-|7527,7528
First|7529,7534
<EOL>|7535,7536
Line|7536,7540
<EOL>|7542,7543
11.|7543,7546
HELD|7547,7551
-|7551,7552
Trimethoprim|7553,7565
100|7566,7569
mg|7570,7572
PO|7573,7575
Q24H|7576,7580
This|7582,7586
medication|7587,7597
was|7598,7601
held|7602,7606
.|7606,7607
<EOL>|7608,7609
Do|7609,7611
not|7612,7615
restart|7616,7623
Trimethoprim|7624,7636
until|7637,7642
after|7643,7648
you|7649,7652
finish|7653,7659
your|7660,7664
<EOL>|7665,7666
ampicillin|7666,7676
.|7676,7677
<EOL>|7677,7678
<EOL>|7678,7679
<EOL>|7680,7681
Discharge|7681,7690
Disposition|7691,7702
:|7702,7703
<EOL>|7703,7704
Extended|7704,7712
Care|7713,7717
<EOL>|7717,7718
<EOL>|7719,7720
Facility|7720,7728
:|7728,7729
<EOL>|7729,7730
_|7730,7731
_|7731,7732
_|7732,7733
<EOL>|7733,7734
<EOL>|7735,7736
Discharge|7736,7745
Diagnosis|7746,7755
:|7755,7756
<EOL>|7756,7757
Complicated|7757,7768
E.|7769,7771
faecium|7772,7779
UTI|7780,7783
<EOL>|7783,7784
<EOL>|7784,7785
<EOL>|7786,7787
Discharge|7787,7796
Condition|7797,7806
:|7806,7807
<EOL>|7807,7808
Mental|7808,7814
Status|7815,7821
:|7821,7822
Clear|7823,7828
and|7829,7832
coherent|7833,7841
.|7841,7842
<EOL>|7842,7843
Level|7843,7848
of|7849,7851
Consciousness|7852,7865
:|7865,7866
Alert|7867,7872
and|7873,7876
interactive|7877,7888
.|7888,7889
<EOL>|7889,7890
Activity|7890,7898
Status|7899,7905
:|7905,7906
Ambulatory|7907,7917
-|7918,7919
Independent|7920,7931
.|7931,7932
<EOL>|7932,7933
<EOL>|7934,7935
Discharge|7935,7944
Instructions|7945,7957
:|7957,7958
<EOL>|7958,7959
You|7959,7962
were|7963,7967
admitted|7968,7976
to|7977,7979
the|7980,7983
hospital|7984,7992
after|7993,7998
you|7999,8002
developed|8003,8012
fevers|8013,8019
and|8020,8023
<EOL>|8024,8025
chills|8025,8031
after|8032,8037
you|8038,8041
developed|8042,8051
fevers|8052,8058
and|8059,8062
chills|8063,8069
from|8070,8074
your|8075,8079
stent|8080,8085
<EOL>|8086,8087
exchange|8087,8095
.|8095,8096
Your|8097,8101
urine|8102,8107
grew|8108,8112
the|8113,8116
enterococcus|8117,8129
species|8130,8137
-|8138,8139
-|8139,8140
the|8141,8144
source|8145,8151
<EOL>|8152,8153
of|8153,8155
your|8156,8160
infection|8161,8170
.|8170,8171
Because|8172,8179
it|8180,8182
was|8183,8186
enterococcus|8187,8199
,|8199,8200
a|8201,8202
PICC|8203,8207
line|8208,8212
was|8213,8216
<EOL>|8217,8218
placed|8218,8224
and|8225,8228
you|8229,8232
will|8233,8237
finish|8238,8244
a|8245,8246
total|8247,8252
14|8253,8255
-|8255,8256
day|8256,8259
course|8260,8266
of|8267,8269
IV|8270,8272
<EOL>|8273,8274
ampicillin|8274,8284
.|8284,8285
<EOL>|8285,8286
<EOL>|8286,8287
You|8287,8290
also|8291,8295
had|8296,8299
kidney|8300,8306
injury|8307,8313
,|8313,8314
likely|8315,8321
from|8322,8326
infection|8327,8336
,|8336,8337
that|8338,8342
resolved|8343,8351
<EOL>|8352,8353
with|8353,8357
antibiotics|8358,8369
and|8370,8373
fluids|8374,8380
.|8380,8381
It|8382,8384
was|8385,8388
a|8389,8390
pleasure|8391,8399
taking|8400,8406
care|8407,8411
of|8412,8414
<EOL>|8415,8416
you|8416,8419
!|8419,8420
<EOL>|8420,8421
<EOL>|8422,8423
Followup|8423,8431
Instructions|8432,8444
:|8444,8445
<EOL>|8445,8446
_|8446,8447
_|8447,8448
_|8448,8449
<EOL>|8449,8450

