 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|46,55|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|46,55|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|46,60|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|80,89|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|80,89|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|80,94|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|136,139|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|147,154|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|147,154|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|156,164|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|SIMPLE_SEGMENT|167,176|false|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|167,176|false|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|167,176|false|false|false|C0020517|Hypersensitivity|Allergies
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|179,189|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|179,189|false|false|false|C0065374|lisinopril|lisinopril
Event|Event|SIMPLE_SEGMENT|179,189|false|false|false|||lisinopril
Event|Event|SIMPLE_SEGMENT|192,201|false|false|false|||Attending
Finding|Functional Concept|SIMPLE_SEGMENT|192,201|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|SIMPLE_SEGMENT|209,224|false|false|false|C0277786|Chief complaint (finding)|Chief Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|215,224|false|false|false|C3864418||Complaint
Event|Event|SIMPLE_SEGMENT|215,224|false|false|false|||Complaint
Finding|Finding|SIMPLE_SEGMENT|215,224|false|false|false|C5441521|Complaint (finding)|Complaint
Anatomy|Body Location or Region|SIMPLE_SEGMENT|226,231|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|SIMPLE_SEGMENT|226,231|false|false|false|C0741025|Chest problem|Chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|226,236|false|false|false|C2926613||Chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|226,236|false|false|false|C0008031|Chest Pain|Chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|232,236|false|true|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|232,236|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|232,236|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|232,236|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Classification|SIMPLE_SEGMENT|239,244|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|SIMPLE_SEGMENT|245,253|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|245,253|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|257,275|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|266,275|false|false|false|C0945766||Procedure
Event|Event|SIMPLE_SEGMENT|266,275|false|false|false|||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|266,275|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|266,275|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|266,275|false|false|false|C0184661|Interventional procedure|Procedure
Event|Event|SIMPLE_SEGMENT|284,291|true|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|284,291|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|284,291|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|284,291|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|284,294|true|false|false|C0262926|Medical History|History of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|284,310|true|false|false|C0488508||History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|284,310|true|false|false|C0262512|History of present illness (finding)|History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|295,302|true|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Idea or Concept|SIMPLE_SEGMENT|295,302|true|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Finding|SIMPLE_SEGMENT|295,310|true|false|false|C4264312|Present illness|Present Illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|303,310|true|false|false|C0221423|Illness (finding)|Illness
Finding|Idea or Concept|SIMPLE_SEGMENT|329,333|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|SIMPLE_SEGMENT|329,333|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Event|Event|SIMPLE_SEGMENT|334,337|false|false|false|||old
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|359,366|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|359,366|false|false|false|C1314974|Cardiac attachment|cardiac
Event|Event|SIMPLE_SEGMENT|367,374|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|367,374|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|367,374|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|367,374|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Anatomy|Body Location or Region|SIMPLE_SEGMENT|398,404|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|398,404|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|405,408|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|405,408|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|405,408|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|405,408|false|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|405,408|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|405,408|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|405,408|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|405,408|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Event|Event|SIMPLE_SEGMENT|413,421|false|false|false|||stenting
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|413,421|false|false|false|C2348535|Stenting|stenting
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|429,432|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|429,432|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|SIMPLE_SEGMENT|429,432|false|false|false|||LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|429,432|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Finding|Pathologic Function|SIMPLE_SEGMENT|442,458|false|false|false|C3272317|Stent restenosis|stent restenosis
Event|Event|SIMPLE_SEGMENT|448,458|false|false|false|||restenosis
Finding|Pathologic Function|SIMPLE_SEGMENT|448,458|false|false|false|C0333186|Restenosis|restenosis
Event|Event|SIMPLE_SEGMENT|463,471|false|false|false|||stenting
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|463,471|false|false|false|C2348535|Stenting|stenting
Event|Event|SIMPLE_SEGMENT|487,491|false|false|false|||CABG
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|487,491|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Finding|Finding|SIMPLE_SEGMENT|510,518|false|false|false|C0028778;C1947917|Obstruction;Occluded|occluded
Finding|Functional Concept|SIMPLE_SEGMENT|510,518|false|false|false|C0028778;C1947917|Obstruction;Occluded|occluded
Finding|Intellectual Product|SIMPLE_SEGMENT|531,537|false|false|false|C0030650|Legal patent|patent
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|543,546|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|543,546|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|SIMPLE_SEGMENT|543,546|false|false|false|||LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|543,546|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Finding|Functional Concept|SIMPLE_SEGMENT|567,584|false|false|false|C3853134|Poorly controlled|poorly controlled
Event|Event|SIMPLE_SEGMENT|574,584|false|false|false|||controlled
Finding|Gene or Genome|SIMPLE_SEGMENT|585,589|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Finding|Intellectual Product|SIMPLE_SEGMENT|585,589|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Finding|Classification|SIMPLE_SEGMENT|585,591|false|false|false|C0441730|Type 2|type 2
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|585,600|false|false|false|C0011860|Diabetes Mellitus, Non-Insulin-Dependent|type 2 diabetes
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|585,609|false|false|false|C0011860|Diabetes Mellitus, Non-Insulin-Dependent|type 2 diabetes mellitus
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|592,600|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|diabetes
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|592,609|false|false|false|C0011849|Diabetes Mellitus|diabetes mellitus
Event|Event|SIMPLE_SEGMENT|601,609|false|false|false|||mellitus
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|612,624|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|SIMPLE_SEGMENT|612,624|false|false|false|||hypertension
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|626,630|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|626,630|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|SIMPLE_SEGMENT|626,630|false|false|false|||COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|626,630|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|632,636|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Event|Event|SIMPLE_SEGMENT|632,636|false|false|false|||GERD
Event|Event|SIMPLE_SEGMENT|642,652|false|false|false|||presenting
Finding|Finding|SIMPLE_SEGMENT|658,661|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|658,661|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Anatomy|Body Location or Region|SIMPLE_SEGMENT|662,667|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|662,667|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|662,672|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|662,672|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|668,672|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|668,672|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|668,672|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|668,672|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Idea or Concept|SIMPLE_SEGMENT|691,694|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|691,694|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|698,710|false|false|false|||presentation
Finding|Idea or Concept|SIMPLE_SEGMENT|698,710|false|false|false|C0449450|Presentation|presentation
Event|Event|SIMPLE_SEGMENT|720,727|false|false|false|||resting
Finding|Finding|SIMPLE_SEGMENT|728,735|false|false|false|C4534363|At home|at home
Event|Event|SIMPLE_SEGMENT|731,735|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|731,735|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|731,735|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|731,735|false|false|false|C1553498|home health encounter|home
Event|Event|SIMPLE_SEGMENT|750,755|false|false|false|||onset
Finding|Finding|SIMPLE_SEGMENT|759,765|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|SIMPLE_SEGMENT|759,765|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Finding|SIMPLE_SEGMENT|766,779|false|false|false|C0278145;C1444775|Sharp sensation quality;Stabbing pain|stabbing pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|766,779|false|false|false|C0278145;C1444775|Sharp sensation quality;Stabbing pain|stabbing pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|775,779|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|775,779|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|775,779|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|775,779|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Functional Concept|SIMPLE_SEGMENT|780,784|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|792,799|false|false|false|C0038293|Sternum|sternum
Attribute|Clinical Attribute|SIMPLE_SEGMENT|807,811|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|807,811|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|807,811|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|807,811|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|812,820|false|false|false|||radiated
Anatomy|Body Location or Region|SIMPLE_SEGMENT|832,837|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|832,837|false|false|false|C0741025|Chest problem|chest
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|853,856|true|false|false|C0446516;C1140618;C1269078|Upper Extremity;Upper arm|arm
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|853,856|true|true|false|C3495676|Anorectal Malformations|arm
Event|Event|SIMPLE_SEGMENT|853,856|true|false|false|||arm
Finding|Gene or Genome|SIMPLE_SEGMENT|853,856|true|true|false|C1824218;C3715044|AKR1A1 wt Allele;ARMC9 gene|arm
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|853,856|true|true|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Research Activity|SIMPLE_SEGMENT|853,856|true|true|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|853,856|true|true|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|860,863|true|false|false|C0022359|Jaw|jaw
Event|Event|SIMPLE_SEGMENT|870,874|false|false|false|||took
Drug|Organic Chemical|SIMPLE_SEGMENT|877,890|false|false|false|C0017887|nitroglycerin|nitroglycerin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|877,890|false|false|false|C0017887|nitroglycerin|nitroglycerin
Event|Event|SIMPLE_SEGMENT|877,890|false|false|false|||nitroglycerin
Event|Event|SIMPLE_SEGMENT|898,906|false|false|false|||improved
Attribute|Clinical Attribute|SIMPLE_SEGMENT|911,915|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|911,915|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|911,915|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|911,915|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|931,938|false|false|false|||reports
Attribute|Clinical Attribute|SIMPLE_SEGMENT|948,952|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|948,952|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|948,952|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|948,952|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|953,957|false|false|false|||came
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|961,966|false|false|false|C0678544||waves
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|975,984|false|false|false|C0886384|5 minutes Office visit|5 minutes
Event|Event|SIMPLE_SEGMENT|977,984|false|false|false|||minutes
Finding|Functional Concept|SIMPLE_SEGMENT|1005,1009|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1010,1015|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|1010,1015|false|false|false|C0741025|Chest problem|chest
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1010,1020|false|false|false|C0205076;C4266615|Chest wall structure;Chest>Chest wall|chest wall
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1010,1020|false|false|false|C0205076;C4266615|Chest wall structure;Chest>Chest wall|chest wall
Finding|Finding|SIMPLE_SEGMENT|1010,1031|false|false|false|C0239008|Chest wall tenderness|chest wall tenderness
Event|Event|SIMPLE_SEGMENT|1021,1031|false|false|false|||tenderness
Finding|Mental Process|SIMPLE_SEGMENT|1021,1031|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|SIMPLE_SEGMENT|1021,1031|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Event|Event|SIMPLE_SEGMENT|1045,1053|true|false|false|||remember
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1073,1078|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|1073,1078|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1073,1083|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1073,1083|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1079,1083|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|1079,1083|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|1079,1083|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1079,1083|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1103,1107|true|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|1103,1107|true|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|1103,1107|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1103,1107|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|1125,1135|true|false|false|||exertional
Finding|Sign or Symptom|SIMPLE_SEGMENT|1125,1135|true|false|false|C0239313|exercise induced|exertional
Finding|Finding|SIMPLE_SEGMENT|1141,1146|false|false|false|C1444775;C1539835;C3890003|SPEN gene;SPEN wt Allele;Sharp sensation quality|sharp
Finding|Gene or Genome|SIMPLE_SEGMENT|1141,1146|false|false|false|C1444775;C1539835;C3890003|SPEN gene;SPEN wt Allele;Sharp sensation quality|sharp
Event|Event|SIMPLE_SEGMENT|1147,1152|false|false|false|||pains
Finding|Sign or Symptom|SIMPLE_SEGMENT|1147,1152|false|false|false|C0030193|Pain|pains
Event|Event|SIMPLE_SEGMENT|1153,1161|false|false|false|||occurred
Event|Event|SIMPLE_SEGMENT|1175,1180|false|false|false|||lying
Event|Event|SIMPLE_SEGMENT|1192,1196|false|false|false|||says
Event|Governmental or Regulatory Activity|SIMPLE_SEGMENT|1201,1205|false|false|false|C1510751|Academic Research Enhancement Awards|area
Event|Event|SIMPLE_SEGMENT|1214,1220|false|false|false|||tender
Event|Event|SIMPLE_SEGMENT|1222,1227|false|false|false|||Lying
Finding|Individual Behavior|SIMPLE_SEGMENT|1222,1227|false|false|false|C0600261|Telling untruths|Lying
Finding|Functional Concept|SIMPLE_SEGMENT|1235,1239|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Event|Event|SIMPLE_SEGMENT|1245,1251|false|false|false|||causes
Finding|Functional Concept|SIMPLE_SEGMENT|1245,1251|false|false|false|C0015127;C1314792|Etiology;Etiology aspects|causes
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1253,1257|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|1253,1257|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|1253,1257|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1253,1257|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Intellectual Product|SIMPLE_SEGMENT|1267,1278|false|false|false|C2984057|Have Nausea|have nausea
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1272,1278|false|false|false|C4255480||nausea
Event|Event|SIMPLE_SEGMENT|1272,1278|false|false|false|||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|1272,1278|false|false|false|C0027497|Nausea|nausea
Event|Event|SIMPLE_SEGMENT|1290,1298|false|false|false|||mornings
Event|Event|SIMPLE_SEGMENT|1305,1313|false|false|false|||resolved
Event|Event|SIMPLE_SEGMENT|1327,1335|true|false|false|||vomiting
Finding|Sign or Symptom|SIMPLE_SEGMENT|1327,1335|true|false|false|C0042963|Vomiting|vomiting
Event|Event|SIMPLE_SEGMENT|1337,1348|true|false|false|||diaphoresis
Finding|Finding|SIMPLE_SEGMENT|1337,1348|true|false|false|C0700590|Increased sweating|diaphoresis
Event|Event|SIMPLE_SEGMENT|1350,1356|true|false|false|||fevers
Finding|Sign or Symptom|SIMPLE_SEGMENT|1350,1356|true|false|false|C0015967|Fever|fevers
Event|Event|SIMPLE_SEGMENT|1360,1366|true|false|false|||chills
Finding|Sign or Symptom|SIMPLE_SEGMENT|1360,1366|true|false|false|C0085593|Chills|chills
Event|Event|SIMPLE_SEGMENT|1376,1378|false|false|false|||an
Event|Event|SIMPLE_SEGMENT|1380,1387|false|false|false|||episode
Event|Event|SIMPLE_SEGMENT|1391,1399|false|false|false|||diarrhea
Finding|Finding|SIMPLE_SEGMENT|1391,1399|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|SIMPLE_SEGMENT|1391,1399|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1418,1427|true|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|SIMPLE_SEGMENT|1418,1432|true|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1428,1432|true|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|1428,1432|true|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|1428,1432|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1428,1432|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|SIMPLE_SEGMENT|1464,1471|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1464,1471|false|false|false|C0004057|aspirin|aspirin
Event|Event|SIMPLE_SEGMENT|1464,1471|false|false|false|||aspirin
Finding|Idea or Concept|SIMPLE_SEGMENT|1479,1482|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|1479,1482|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|1486,1498|false|false|false|||presentation
Finding|Idea or Concept|SIMPLE_SEGMENT|1486,1498|false|false|false|C0449450|Presentation|presentation
Finding|Idea or Concept|SIMPLE_SEGMENT|1515,1522|false|false|false|C1555582|Initial (abbreviation)|initial
Event|Event|SIMPLE_SEGMENT|1523,1529|false|false|false|||vitals
Event|Event|SIMPLE_SEGMENT|1544,1546|false|false|false|||HR
Event|Event|SIMPLE_SEGMENT|1587,1591|false|false|false|||FSBG
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1601,1605|false|false|false|C0587081|Laboratory test finding|Labs
Event|Event|SIMPLE_SEGMENT|1606,1613|false|false|false|||notable
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1618,1626|false|false|false|C0041199|Troponin|Troponin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1618,1626|false|false|false|C0041199|Troponin|Troponin
Event|Event|SIMPLE_SEGMENT|1618,1626|false|false|false|||Troponin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1618,1626|false|false|false|C0523952|Troponin measurement|Troponin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1618,1628|false|false|false|C0077404|Troponin T|Troponin-T
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1618,1628|false|false|false|C0077404|Troponin T|Troponin-T
Event|Event|SIMPLE_SEGMENT|1627,1628|false|false|false|||T
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1638,1643|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|SIMPLE_SEGMENT|1638,1643|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|SIMPLE_SEGMENT|1638,1643|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1638,1643|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Event|Event|SIMPLE_SEGMENT|1641,1643|false|false|false|||MB
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1649,1656|false|false|false|C0060323|Fibrin fragment D|D-Dimer
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1649,1656|false|false|false|C0060323|Fibrin fragment D|D-Dimer
Drug|Chemical Viewed Structurally|SIMPLE_SEGMENT|1651,1656|false|false|false|C0596448|dimer|Dimer
Event|Event|SIMPLE_SEGMENT|1651,1656|false|false|false|||Dimer
Event|Event|SIMPLE_SEGMENT|1670,1672|false|false|false|||Mg
Event|Event|SIMPLE_SEGMENT|1685,1689|false|false|false|||LFTs
Anatomy|Cell Component|SIMPLE_SEGMENT|1691,1694|false|false|false|C2263086|Nuclear cap binding complex location|CBC
Event|Event|SIMPLE_SEGMENT|1691,1694|false|false|false|||CBC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1691,1694|false|false|false|C0009555|Complete Blood Count|CBC
Event|Event|SIMPLE_SEGMENT|1697,1701|false|false|false|||Chem
Finding|Functional Concept|SIMPLE_SEGMENT|1697,1701|false|false|false|C0079107|chemical aspects|Chem
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1697,1701|false|false|false|C0201682|Chemical procedure|Chem
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1697,1703|false|false|false|C2237045|Basic metabolic panel|Chem 7
Event|Event|SIMPLE_SEGMENT|1711,1714|false|false|false|||WNL
Event|Event|SIMPLE_SEGMENT|1716,1719|true|false|false|||CXR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1716,1719|true|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|SIMPLE_SEGMENT|1720,1726|true|false|false|||showed
Finding|Intellectual Product|SIMPLE_SEGMENT|1730,1735|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1736,1751|true|false|false|C0553534|Cardiopulmonary|cardiopulmonary
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1736,1751|true|false|false|C4072686|Cardiovascular disease+Pulmonary disease|cardiopulmonary
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|1753,1764|true|false|false|C0000768|Congenital Abnormality|abnormality
Event|Event|SIMPLE_SEGMENT|1753,1764|true|false|false|||abnormality
Finding|Finding|SIMPLE_SEGMENT|1753,1764|true|false|false|C1704258|Abnormality|abnormality
Event|Event|SIMPLE_SEGMENT|1774,1788|true|false|false|||echocardiogram
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1774,1788|true|false|false|C0013516|Echocardiography|echocardiogram
Event|Event|SIMPLE_SEGMENT|1789,1795|true|false|false|||showed
Event|Event|SIMPLE_SEGMENT|1799,1810|true|false|false|||substantial
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1812,1823|true|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1812,1823|true|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1812,1832|true|false|false|C0031039|Pericardial effusion|pericardial effusion
Finding|Body Substance|SIMPLE_SEGMENT|1812,1832|true|false|false|C1253937|Pericardial effusion body substance|pericardial effusion
Event|Event|SIMPLE_SEGMENT|1824,1832|true|false|false|||effusion
Finding|Body Substance|SIMPLE_SEGMENT|1824,1832|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|SIMPLE_SEGMENT|1824,1832|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|1824,1832|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Event|Event|SIMPLE_SEGMENT|1836,1845|true|false|false|||tamponade
Finding|Functional Concept|SIMPLE_SEGMENT|1836,1845|true|false|false|C0332459|Compressed structure|tamponade
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1836,1845|true|false|false|C0579016||tamponade
Finding|Body Substance|SIMPLE_SEGMENT|1847,1854|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1847,1854|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1847,1854|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Organic Chemical|SIMPLE_SEGMENT|1865,1876|false|false|false|C0082607|fluticasone|fluticasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1865,1876|false|false|false|C0082607|fluticasone|fluticasone
Event|Event|SIMPLE_SEGMENT|1865,1876|false|false|false|||fluticasone
Drug|Organic Chemical|SIMPLE_SEGMENT|1878,1888|false|false|false|C0033474;C0392214|Propionates;propionate|propionate
Event|Event|SIMPLE_SEGMENT|1889,1896|false|false|false|||inhaled
Drug|Organic Chemical|SIMPLE_SEGMENT|1898,1907|false|false|false|C0030049|oxycodone|OxyCODONE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1898,1907|false|false|false|C0030049|oxycodone|OxyCODONE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1898,1907|false|false|false|C0524222|Oxycodone measurement|OxyCODONE
Drug|Organic Chemical|SIMPLE_SEGMENT|1909,1922|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1909,1922|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|SIMPLE_SEGMENT|1909,1922|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1909,1922|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1937,1946|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|Magnesium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|1937,1946|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|Magnesium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|1937,1946|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|Magnesium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1937,1946|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|Magnesium
Event|Event|SIMPLE_SEGMENT|1937,1946|false|false|false|||Magnesium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1937,1946|false|false|false|C0373675|Magnesium measurement|Magnesium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|1937,1954|false|false|false|C0024480|magnesium sulfate|Magnesium Sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1937,1954|false|false|false|C0024480|magnesium sulfate|Magnesium Sulfate
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|1947,1954|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Inorganic Chemical|SIMPLE_SEGMENT|1947,1954|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1947,1954|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Event|Activity|SIMPLE_SEGMENT|1969,1976|false|false|false|C1706079||arrival
Event|Event|SIMPLE_SEGMENT|1969,1976|false|false|false|||arrival
Finding|Functional Concept|SIMPLE_SEGMENT|1969,1976|false|false|false|C1555577|arrival - ActRelationshipType|arrival
Anatomy|Body System|SIMPLE_SEGMENT|1984,1994|false|false|false|C0007226|Cardiovascular system|cardiology
Finding|Body Substance|SIMPLE_SEGMENT|2005,2012|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|2005,2012|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|2005,2012|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|2013,2021|false|false|false|||reported
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2032,2036|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|2032,2036|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|2032,2036|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|2032,2036|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2041,2046|false|false|false|C1410088|Still|still
Event|Event|SIMPLE_SEGMENT|2060,2064|false|false|false|||felt
Event|Event|SIMPLE_SEGMENT|2088,2093|false|false|false|||worse
Finding|Finding|SIMPLE_SEGMENT|2088,2093|false|false|false|C1457868;C1550463|Observation Interpretation - worse;Worse|worse
Finding|Idea or Concept|SIMPLE_SEGMENT|2088,2093|false|false|false|C1457868;C1550463|Observation Interpretation - worse;Worse|worse
Event|Governmental or Regulatory Activity|SIMPLE_SEGMENT|2108,2112|false|false|false|C1510751|Academic Research Enhancement Awards|area
Event|Event|SIMPLE_SEGMENT|2117,2123|false|false|false|||tender
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2136,2145|true|false|false|C5885990||breathing
Finding|Finding|SIMPLE_SEGMENT|2136,2145|true|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|SIMPLE_SEGMENT|2136,2145|true|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|SIMPLE_SEGMENT|2136,2145|true|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|SIMPLE_SEGMENT|2136,2145|true|false|false|C1160636|respiratory system process|breathing
Event|Event|SIMPLE_SEGMENT|2146,2156|true|false|false|||complaints
Finding|Finding|SIMPLE_SEGMENT|2146,2156|true|false|false|C5441521|Complaint (finding)|complaints
Event|Event|SIMPLE_SEGMENT|2163,2167|false|false|false|||felt
Finding|Finding|SIMPLE_SEGMENT|2168,2176|false|false|false|C2984078;C3889124|A little bit;Only a Little|a little
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2170,2176|false|false|false|C0023882|Little's Disease|little
Event|Event|SIMPLE_SEGMENT|2170,2176|false|false|false|||little
Finding|Finding|SIMPLE_SEGMENT|2170,2176|false|false|false|C3889124|Only a Little|little
Finding|Functional Concept|SIMPLE_SEGMENT|2177,2186|false|false|false|C1533708|Congested|congested
Event|Event|SIMPLE_SEGMENT|2192,2199|false|false|false|||evening
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2209,2213|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|2209,2213|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|2209,2213|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|2209,2213|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|2214,2221|false|false|false|||started
Finding|Finding|SIMPLE_SEGMENT|2225,2245|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Event|Event|SIMPLE_SEGMENT|2230,2237|false|false|false|||Medical
Finding|Functional Concept|SIMPLE_SEGMENT|2230,2237|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|2230,2237|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|2230,2237|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|2230,2237|false|false|false|C0199168|Medical service|Medical
Finding|Finding|SIMPLE_SEGMENT|2230,2245|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2238,2245|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2238,2245|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2238,2245|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2248,2252|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2248,2252|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|SIMPLE_SEGMENT|2248,2252|false|false|false|||COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|2248,2252|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2254,2257|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2254,2257|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|2254,2257|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|2254,2257|false|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|2254,2257|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2254,2257|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|2254,2257|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2254,2257|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Event|Event|SIMPLE_SEGMENT|2262,2266|false|false|false|||CABG
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2262,2266|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Event|Event|SIMPLE_SEGMENT|2271,2279|false|false|false|||stenting
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2271,2279|false|false|false|C2348535|Stenting|stenting
Finding|Idea or Concept|SIMPLE_SEGMENT|2284,2289|false|false|false|C1552828|Table Frame - above|above
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|2291,2301|false|false|false|C0011570;C0011581;C0344315;C0812393|Cancer patients and suicide and depression;Depressed mood;Depressive disorder;Mental Depression|Depression
Event|Event|SIMPLE_SEGMENT|2291,2301|false|false|false|||Depression
Finding|Functional Concept|SIMPLE_SEGMENT|2291,2301|false|false|false|C0460137;C1579931|Depression - motion|Depression
Finding|Sign or Symptom|SIMPLE_SEGMENT|2291,2301|false|false|false|C0460137;C1579931|Depression - motion|Depression
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2311,2315|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Event|Event|SIMPLE_SEGMENT|2311,2315|false|false|false|||GERD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2319,2331|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|SIMPLE_SEGMENT|2319,2331|false|false|false|||Hypertension
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2333,2342|false|false|false|C0149931|Migraine Disorders|Migraines
Event|Event|SIMPLE_SEGMENT|2333,2342|false|false|false|||Migraines
Finding|Intellectual Product|SIMPLE_SEGMENT|2344,2351|false|false|false|C1547296|Chronic - Admission Level of Care Code|Chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|2344,2351|false|false|false|C1555457|Provision of recurring care for chronic illness|Chronic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2344,2365|false|false|false|C0748678|shoulder pain chronic|Chronic shoulder pain
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2352,2360|false|false|false|C0037004;C4299050|Shoulder;Upper extremity>Shoulder|shoulder
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2352,2360|false|false|false|C0221590;C0869975|Examination of shoulder(s);Procedures on Shoulder|shoulder
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2352,2360|false|false|false|C0221590;C0869975|Examination of shoulder(s);Procedures on Shoulder|shoulder
Finding|Sign or Symptom|SIMPLE_SEGMENT|2352,2365|false|false|false|C0037011|Shoulder Pain|shoulder pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2361,2365|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|2361,2365|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|2361,2365|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|2361,2365|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|2369,2378|false|false|false|C0027415|Narcotics|narcotics
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2369,2378|false|false|false|C0027415|Narcotics|narcotics
Event|Event|SIMPLE_SEGMENT|2369,2378|false|false|false|||narcotics
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2380,2383|false|false|false|C0520679|Sleep Apnea, Obstructive|OSA
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2380,2383|false|false|false|C0764906|OSA protein, Drosophila|OSA
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2380,2383|false|false|false|C0764906|OSA protein, Drosophila|OSA
Event|Event|SIMPLE_SEGMENT|2380,2383|false|false|false|||OSA
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2385,2406|false|false|false|C0031117;C4721453|Peripheral Nervous System Diseases;Peripheral Neuropathy|Peripheral neuropathy
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2396,2406|false|false|false|C0442874|Neuropathy|neuropathy
Event|Event|SIMPLE_SEGMENT|2396,2406|false|false|false|||neuropathy
Finding|Sign or Symptom|SIMPLE_SEGMENT|2408,2416|false|false|false|C0085631;C3887611|Agitation;Restlessness|Restless
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2408,2420|false|false|false|C0035258|Restless Legs Syndrome|Restless leg
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2417,2420|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Finding|Functional Concept|SIMPLE_SEGMENT|2423,2429|false|false|false|C0728831|Social|Social
Finding|Finding|SIMPLE_SEGMENT|2423,2437|false|false|false|C0424945;C3714536|Social History;Social and personal history|Social History
Event|Event|SIMPLE_SEGMENT|2430,2437|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2430,2437|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2430,2437|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2430,2437|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Classification|SIMPLE_SEGMENT|2443,2449|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|SIMPLE_SEGMENT|2443,2449|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|SIMPLE_SEGMENT|2443,2449|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|SIMPLE_SEGMENT|2443,2449|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Finding|SIMPLE_SEGMENT|2443,2457|false|false|false|C0241889|Family Medical History|Family History
Event|Event|SIMPLE_SEGMENT|2450,2457|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2450,2457|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2450,2457|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2450,2457|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Body Substance|SIMPLE_SEGMENT|2459,2466|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|2459,2466|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|2459,2466|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|2471,2475|false|false|false|||ward
Event|Event|SIMPLE_SEGMENT|2496,2500|true|false|false|||know
Event|Event|SIMPLE_SEGMENT|2506,2513|true|false|false|||details
Finding|Classification|SIMPLE_SEGMENT|2518,2524|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|2518,2524|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|2518,2524|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|2518,2524|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Finding|SIMPLE_SEGMENT|2518,2532|true|false|false|C0241889|Family Medical History|family history
Event|Event|SIMPLE_SEGMENT|2525,2532|true|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|2525,2532|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|2525,2532|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|2525,2532|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Event|Event|SIMPLE_SEGMENT|2534,2540|false|false|false|||Mother
Finding|Idea or Concept|SIMPLE_SEGMENT|2534,2540|false|false|false|C1546508|Relationship - Mother|Mother
Finding|Finding|SIMPLE_SEGMENT|2546,2554|false|false|false|C0332149|Possible|possible
Drug|Organic Chemical|SIMPLE_SEGMENT|2555,2562|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2555,2562|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Event|Event|SIMPLE_SEGMENT|2555,2562|false|false|false|||alcohol
Finding|Intellectual Product|SIMPLE_SEGMENT|2555,2562|false|false|false|C1547288|Alcohol - Recreational Drug Use Code|alcohol
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|2555,2568|false|true|false|C0085762|Alcohol abuse|alcohol abuse
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|2563,2568|false|false|false|C0013146|Drug abuse|abuse
Event|Event|SIMPLE_SEGMENT|2563,2568|false|false|false|||abuse
Event|Event|SIMPLE_SEGMENT|2563,2568|false|false|false|C1546935|Abuse|abuse
Finding|Finding|SIMPLE_SEGMENT|2563,2568|false|false|false|C0562381|Victim of abuse (finding)|abuse
Finding|Conceptual Entity|SIMPLE_SEGMENT|2570,2576|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Idea or Concept|SIMPLE_SEGMENT|2570,2576|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Event|Event|SIMPLE_SEGMENT|2578,2586|false|false|false|||deceased
Finding|Finding|SIMPLE_SEGMENT|2578,2586|false|false|false|C0011065;C1549464;C1704456|Cessation of life;Deceased - ActIneligibilityReason;Deceased - Military Status|deceased
Finding|Organism Function|SIMPLE_SEGMENT|2578,2586|false|false|false|C0011065;C1549464;C1704456|Cessation of life;Deceased - ActIneligibilityReason;Deceased - Military Status|deceased
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2599,2606|false|false|false|C0019829|Hodgkin Disease|Hodgkin
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2599,2616|false|false|false|C0019829|Hodgkin Disease|Hodgkin's Disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2609,2616|false|false|false|C0012634|Disease|Disease
Event|Event|SIMPLE_SEGMENT|2609,2616|false|false|false|||Disease
Event|Event|SIMPLE_SEGMENT|2625,2632|false|false|false|||records
Finding|Idea or Concept|SIMPLE_SEGMENT|2625,2632|false|false|false|C0034869;C1548330|Quantity limited request - Records;Records|records
Finding|Intellectual Product|SIMPLE_SEGMENT|2625,2632|false|false|false|C0034869;C1548330|Quantity limited request - Records;Records|records
Event|Event|SIMPLE_SEGMENT|2636,2644|false|false|false|||Physical
Finding|Finding|SIMPLE_SEGMENT|2636,2644|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|2636,2644|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|2636,2644|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|2636,2649|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2636,2649|false|false|false|C0031809|Physical Examination|Physical Exam
Event|Event|SIMPLE_SEGMENT|2645,2649|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|2645,2649|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2645,2649|false|false|false|C0582103|Medical Examination|Exam
Event|Event|SIMPLE_SEGMENT|2654,2663|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|2654,2663|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|SIMPLE_SEGMENT|2664,2671|false|false|false|||General
Finding|Classification|SIMPLE_SEGMENT|2664,2671|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|SIMPLE_SEGMENT|2664,2671|false|false|false|C3812897|General medical service|General
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2673,2678|false|false|false|C0028754|Obesity|Obese
Event|Event|SIMPLE_SEGMENT|2673,2678|false|false|false|||Obese
Finding|Intellectual Product|SIMPLE_SEGMENT|2679,2685|false|false|false|C1552826|Table Cell Vertical Align - middle|middle
Event|Event|SIMPLE_SEGMENT|2686,2690|false|false|false|||aged
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2702,2707|true|false|false|C5890168||alert
Drug|Organic Chemical|SIMPLE_SEGMENT|2702,2707|true|false|false|C0718338|Alert brand of caffeine|alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2702,2707|true|false|false|C0718338|Alert brand of caffeine|alert
Event|Event|SIMPLE_SEGMENT|2702,2707|true|false|false|||alert
Finding|Finding|SIMPLE_SEGMENT|2702,2707|true|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Functional Concept|SIMPLE_SEGMENT|2702,2707|true|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Intellectual Product|SIMPLE_SEGMENT|2702,2707|true|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Event|Event|SIMPLE_SEGMENT|2709,2717|true|false|false|||oriented
Finding|Finding|SIMPLE_SEGMENT|2709,2717|true|false|false|C1961028|Oriented to place|oriented
Finding|Intellectual Product|SIMPLE_SEGMENT|2726,2731|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|SIMPLE_SEGMENT|2732,2740|true|false|false|||distress
Finding|Finding|SIMPLE_SEGMENT|2732,2740|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|SIMPLE_SEGMENT|2732,2740|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Drug|Food|SIMPLE_SEGMENT|2741,2746|true|false|false|C1875856|Vital High Nitrogen Enteral Nutrition|Vital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2741,2752|true|false|false|C0488614;C0518766|Vital signs|Vital Signs
Procedure|Health Care Activity|SIMPLE_SEGMENT|2741,2752|true|false|false|C0150404|Taking vital signs|Vital Signs
Event|Event|SIMPLE_SEGMENT|2747,2752|true|false|false|||Signs
Finding|Finding|SIMPLE_SEGMENT|2747,2752|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|Signs
Finding|Functional Concept|SIMPLE_SEGMENT|2747,2752|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|Signs
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2801,2807|false|false|false|C0944911||Weight
Event|Event|SIMPLE_SEGMENT|2801,2807|false|false|false|||Weight
Finding|Finding|SIMPLE_SEGMENT|2801,2807|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|Weight
Finding|Sign or Symptom|SIMPLE_SEGMENT|2801,2807|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|Weight
Procedure|Health Care Activity|SIMPLE_SEGMENT|2801,2807|false|false|false|C1305866|Weighing patient|Weight
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2815,2820|false|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2822,2828|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2822,2828|false|false|false|C0036412|Scleral Diseases|Sclera
Event|Event|SIMPLE_SEGMENT|2822,2828|false|false|false|||Sclera
Procedure|Health Care Activity|SIMPLE_SEGMENT|2822,2828|false|false|false|C2228481|examination of sclera|Sclera
Event|Event|SIMPLE_SEGMENT|2829,2838|false|false|false|||anicteric
Finding|Finding|SIMPLE_SEGMENT|2829,2838|false|false|false|C0205180|Anicteric|anicteric
Finding|Body Substance|SIMPLE_SEGMENT|2840,2846|false|false|false|C0026727;C2753459|Mucus (substance);mucus layer|mucous
Anatomy|Tissue|SIMPLE_SEGMENT|2840,2856|false|false|false|C0026724|Mucous Membrane|mucous membranes
Finding|Finding|SIMPLE_SEGMENT|2840,2856|false|false|false|C2230150|moisture of mucous membranes (physical finding)|mucous membranes
Anatomy|Tissue|SIMPLE_SEGMENT|2847,2856|false|false|false|C0025255|Membrane Tissue|membranes
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2864,2874|false|false|false|C0521367|Oropharyngeal|oropharynx
Event|Event|SIMPLE_SEGMENT|2876,2881|false|false|false|||clear
Finding|Idea or Concept|SIMPLE_SEGMENT|2876,2881|false|false|false|C1550016|Remote control command - Clear|clear
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2882,2886|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|SIMPLE_SEGMENT|2882,2886|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Event|Event|SIMPLE_SEGMENT|2882,2886|false|false|false|||NECK
Finding|Finding|SIMPLE_SEGMENT|2882,2886|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Event|Event|SIMPLE_SEGMENT|2888,2897|false|false|false|||difficult
Finding|Finding|SIMPLE_SEGMENT|2888,2897|false|false|false|C0332218|Difficult (qualifier value)|difficult
Event|Event|SIMPLE_SEGMENT|2901,2911|false|false|false|||appreciate
Event|Event|SIMPLE_SEGMENT|2912,2915|false|false|false|||JVP
Finding|Finding|SIMPLE_SEGMENT|2912,2915|false|false|false|C0428897|Jugular venous pressure|JVP
Event|Activity|SIMPLE_SEGMENT|2928,2932|false|false|false|C0871208|Rating (action)|rate
Event|Event|SIMPLE_SEGMENT|2928,2932|false|false|false|||rate
Finding|Idea or Concept|SIMPLE_SEGMENT|2928,2932|false|false|false|C1549480|Amount type - Rate|rate
Event|Event|SIMPLE_SEGMENT|2937,2943|false|false|false|||rhythm
Finding|Finding|SIMPLE_SEGMENT|2937,2943|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|SIMPLE_SEGMENT|2937,2943|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Event|Event|SIMPLE_SEGMENT|2964,2971|true|false|false|||murmurs
Finding|Finding|SIMPLE_SEGMENT|2964,2971|true|false|false|C0018808|Heart murmur|murmurs
Event|Event|SIMPLE_SEGMENT|2973,2977|true|false|false|||rubs
Finding|Finding|SIMPLE_SEGMENT|2973,2977|true|false|false|C0232267|Pericardial friction rub|rubs
Event|Event|SIMPLE_SEGMENT|2980,2987|true|false|false|||gallops
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2988,2993|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|SIMPLE_SEGMENT|2988,2993|false|false|false|C0741025|Chest problem|Chest
Event|Event|SIMPLE_SEGMENT|2995,3005|false|false|false|||Tenderness
Finding|Mental Process|SIMPLE_SEGMENT|2995,3005|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|Tenderness
Finding|Sign or Symptom|SIMPLE_SEGMENT|2995,3005|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|Tenderness
Event|Event|SIMPLE_SEGMENT|3009,3018|false|false|false|||palpation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3009,3018|false|false|false|C0030247|Palpation|palpation
Finding|Functional Concept|SIMPLE_SEGMENT|3026,3030|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3026,3045|false|false|false|C0694647|left anterior chest|left anterior chest
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3031,3039|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3031,3045|false|false|false|C0230132|Anterior chest wall structure|anterior chest
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3031,3050|false|false|false|C0230132;C1305714|Anterior chest wall structure|anterior chest wall
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3031,3050|false|false|false|C0230132;C1305714|Anterior chest wall structure|anterior chest wall
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3040,3045|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|3040,3045|false|false|false|C0741025|Chest problem|chest
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3040,3050|false|false|false|C0205076;C4266615|Chest wall structure;Chest>Chest wall|chest wall
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3040,3050|false|false|false|C0205076;C4266615|Chest wall structure;Chest>Chest wall|chest wall
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3051,3056|false|false|false|C0024109|Lung|Lungs
Event|Event|SIMPLE_SEGMENT|3058,3063|true|false|false|||Clear
Finding|Idea or Concept|SIMPLE_SEGMENT|3058,3063|true|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|SIMPLE_SEGMENT|3067,3079|true|false|false|||auscultation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3067,3079|true|false|false|C0004339|Auscultation|auscultation
Event|Event|SIMPLE_SEGMENT|3096,3103|true|false|false|||wheezes
Finding|Sign or Symptom|SIMPLE_SEGMENT|3096,3103|true|false|false|C0043144|Wheezing|wheezes
Event|Event|SIMPLE_SEGMENT|3105,3110|true|false|false|||rales
Finding|Finding|SIMPLE_SEGMENT|3105,3110|true|false|false|C0034642;C0240859|Basilar Rales;Rales|rales
Event|Event|SIMPLE_SEGMENT|3113,3120|true|false|false|||rhonchi
Finding|Finding|SIMPLE_SEGMENT|3113,3120|true|false|false|C0035508|Rhonchi|rhonchi
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3121,3128|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3121,3128|false|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Event|Event|SIMPLE_SEGMENT|3121,3128|false|false|false|||Abdomen
Finding|Finding|SIMPLE_SEGMENT|3121,3128|false|false|false|C0941288|Abdomen problem|Abdomen
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3130,3134|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Event|Event|SIMPLE_SEGMENT|3130,3134|false|false|false|||Soft
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3163,3168|false|false|false|C0028754|Obesity|obese
Event|Event|SIMPLE_SEGMENT|3163,3168|false|false|false|||obese
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|3182,3185|true|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Event|Event|SIMPLE_SEGMENT|3182,3185|true|false|false|||Ext
Finding|Gene or Genome|SIMPLE_SEGMENT|3182,3185|true|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Event|Event|SIMPLE_SEGMENT|3187,3191|false|false|false|||Warm
Finding|Finding|SIMPLE_SEGMENT|3187,3191|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3187,3191|false|false|false|C0687712|warming process|Warm
Finding|Finding|SIMPLE_SEGMENT|3193,3197|false|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|3198,3206|false|false|false|||perfused
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|3211,3219|true|false|false|C0149651|Clubbing|clubbing
Event|Event|SIMPLE_SEGMENT|3211,3219|true|false|false|||clubbing
Event|Event|SIMPLE_SEGMENT|3221,3229|true|false|false|||cyanosis
Finding|Sign or Symptom|SIMPLE_SEGMENT|3221,3229|true|false|false|C0010520|Cyanosis|cyanosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3233,3238|true|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|3233,3238|true|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|3233,3238|true|false|false|C0013604|Edema|edema
Event|Event|SIMPLE_SEGMENT|3240,3244|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|3240,3244|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|3240,3244|false|false|false|C0582103|Medical Examination|Exam
Event|Event|SIMPLE_SEGMENT|3245,3254|false|false|false|||unchanged
Finding|Finding|SIMPLE_SEGMENT|3245,3254|false|false|false|C0442739||unchanged
Event|Event|SIMPLE_SEGMENT|3258,3267|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|3258,3267|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|3258,3267|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|3258,3267|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|3258,3267|false|false|false|C0030685|Patient Discharge|discharge
Finding|Functional Concept|SIMPLE_SEGMENT|3269,3273|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3274,3279|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|3274,3279|false|false|false|C0741025|Chest problem|chest
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3274,3284|false|false|false|C0205076;C4266615|Chest wall structure;Chest>Chest wall|chest wall
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3274,3284|false|false|false|C0205076;C4266615|Chest wall structure;Chest>Chest wall|chest wall
Event|Event|SIMPLE_SEGMENT|3285,3291|false|false|false|||tender
Event|Event|SIMPLE_SEGMENT|3298,3307|false|false|false|||palpation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3298,3307|false|false|false|C0030247|Palpation|palpation
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3313,3317|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|3313,3317|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|3313,3317|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|3313,3317|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|3324,3330|false|false|false|||change
Finding|Functional Concept|SIMPLE_SEGMENT|3324,3330|false|false|false|C0392747|Changing|change
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3324,3330|false|false|false|C4319952|Change - procedure|change
Finding|Functional Concept|SIMPLE_SEGMENT|3324,3333|false|false|false|C0392747|Changing|change in
Event|Event|SIMPLE_SEGMENT|3334,3342|false|false|false|||position
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3376,3381|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3376,3381|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3376,3381|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|3382,3385|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|3390,3393|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3390,3393|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3390,3393|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3400,3403|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3400,3403|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|3400,3403|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3400,3403|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3409,3412|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3409,3412|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|3419,3422|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|3419,3422|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3419,3422|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3419,3422|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3419,3422|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|3426,3429|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3426,3429|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|3426,3429|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|3426,3429|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|3426,3429|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3426,3429|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3436,3440|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3466,3469|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3487,3492|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3487,3492|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3487,3492|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|3487,3500|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3487,3500|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3487,3500|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3493,3500|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|3493,3500|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3493,3500|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|3493,3500|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3493,3500|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3493,3500|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|SIMPLE_SEGMENT|3547,3551|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3547,3551|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3547,3551|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3576,3581|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3576,3581|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3576,3581|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3582,3585|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3582,3585|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|SIMPLE_SEGMENT|3582,3585|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|SIMPLE_SEGMENT|3582,3585|false|false|false|||ALT
Finding|Gene or Genome|SIMPLE_SEGMENT|3582,3585|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|SIMPLE_SEGMENT|3582,3585|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|SIMPLE_SEGMENT|3582,3585|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3582,3585|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|3589,3592|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3589,3592|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3589,3592|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3589,3592|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|SIMPLE_SEGMENT|3589,3592|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|SIMPLE_SEGMENT|3589,3592|false|false|false|||AST
Finding|Gene or Genome|SIMPLE_SEGMENT|3589,3592|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3599,3602|false|false|false|C0010287|Creatine Kinase|CPK
Drug|Enzyme|SIMPLE_SEGMENT|3599,3602|false|false|false|C0010287|Creatine Kinase|CPK
Event|Event|SIMPLE_SEGMENT|3599,3602|false|false|false|||CPK
Finding|Gene or Genome|SIMPLE_SEGMENT|3599,3602|false|false|false|C1418571|PIK3C2A gene|CPK
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3599,3602|false|false|false|C0201973|Creatine kinase measurement|CPK
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3607,3614|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|SIMPLE_SEGMENT|3607,3614|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3643,3648|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3643,3648|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3643,3648|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3643,3656|false|false|false|C0853248|Blood albumin|BLOOD Albumin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3649,3656|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3649,3656|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3649,3656|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Event|Event|SIMPLE_SEGMENT|3649,3656|false|false|false|||Albumin
Finding|Gene or Genome|SIMPLE_SEGMENT|3649,3656|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Finding|Physiologic Function|SIMPLE_SEGMENT|3649,3656|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3649,3656|false|false|false|C0201838|Albumin measurement|Albumin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3661,3668|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|3661,3668|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|3661,3668|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3661,3668|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|3661,3668|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|SIMPLE_SEGMENT|3661,3668|false|false|false|||Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|3661,3668|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3661,3668|false|false|false|C0201925|Calcium measurement|Calcium
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3703,3708|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3703,3708|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3703,3708|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3709,3716|false|false|false|C0060323|Fibrin fragment D|D-Dimer
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3709,3716|false|false|false|C0060323|Fibrin fragment D|D-Dimer
Drug|Chemical Viewed Structurally|SIMPLE_SEGMENT|3711,3716|false|false|false|C0596448|dimer|Dimer
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3733,3738|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3733,3738|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3733,3738|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3739,3744|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|SIMPLE_SEGMENT|3739,3744|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|SIMPLE_SEGMENT|3739,3744|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3739,3744|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Event|Event|SIMPLE_SEGMENT|3742,3744|false|false|false|||MB
Finding|Gene or Genome|SIMPLE_SEGMENT|3742,3746|false|false|false|C1413238;C3273407|CD79A gene;CD79A wt Allele|MB-1
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3774,3779|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3774,3779|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3774,3779|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3780,3785|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|SIMPLE_SEGMENT|3780,3785|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|SIMPLE_SEGMENT|3780,3785|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3780,3785|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3816,3821|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3816,3821|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3816,3821|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|3822,3825|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|3830,3833|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3830,3833|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3830,3833|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3840,3843|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3840,3843|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|3840,3843|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3840,3843|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3849,3852|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3849,3852|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|3860,3863|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|3860,3863|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3860,3863|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3860,3863|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3860,3863|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|3867,3870|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3867,3870|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|3867,3870|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|3867,3870|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|3867,3870|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3867,3870|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3877,3881|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3907,3910|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3927,3932|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3927,3932|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3927,3932|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|3927,3940|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3927,3940|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3927,3940|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3933,3940|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|3933,3940|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3933,3940|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|3933,3940|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3933,3940|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3933,3940|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|SIMPLE_SEGMENT|3988,3992|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3988,3992|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3988,3992|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4017,4022|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4017,4022|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4017,4022|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4017,4030|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4023,4030|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4023,4030|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4023,4030|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4023,4030|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|4023,4030|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|SIMPLE_SEGMENT|4023,4030|false|false|false|||Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|4023,4030|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4023,4030|false|false|false|C0201925|Calcium measurement|Calcium
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4052,4055|false|false|false|C0018064|Equine Gonadotropins|ECG
Drug|Hormone|SIMPLE_SEGMENT|4052,4055|false|false|false|C0018064|Equine Gonadotropins|ECG
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4052,4055|false|false|false|C0018064|Equine Gonadotropins|ECG
Event|Event|SIMPLE_SEGMENT|4052,4055|false|false|false|||ECG
Finding|Intellectual Product|SIMPLE_SEGMENT|4052,4055|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|ECG
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4052,4055|false|false|false|C1623258|Electrocardiography|ECG
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4072,4080|false|false|false|C0168634|BaseLine dental cement|Baseline
Event|Event|SIMPLE_SEGMENT|4072,4080|false|false|false|||Baseline
Finding|Idea or Concept|SIMPLE_SEGMENT|4072,4080|false|false|false|C1552824|baseline - TableCellVerticalAlign|Baseline
Event|Event|SIMPLE_SEGMENT|4081,4089|false|false|false|||artifact
Phenomenon|Human-caused Phenomenon or Process|SIMPLE_SEGMENT|4081,4089|false|false|false|C0085089|Morphologic artifact|artifact
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4091,4096|false|false|false|C0030471;C1305231|Nasal sinus;Sinus - general anatomical term|Sinus
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|4091,4096|false|false|false|C0016169|pathologic fistula|Sinus
Drug|Organic Chemical|SIMPLE_SEGMENT|4091,4096|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|Sinus
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4091,4096|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|Sinus
Finding|Finding|SIMPLE_SEGMENT|4091,4103|false|false|false|C0232201;C2041122|Sinus rhythm|Sinus rhythm
Event|Event|SIMPLE_SEGMENT|4097,4103|false|false|false|||rhythm
Finding|Finding|SIMPLE_SEGMENT|4097,4103|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|SIMPLE_SEGMENT|4097,4103|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4116,4128|false|false|false|C0488345;C0520877|PR interval feature|P-R interval
Event|Event|SIMPLE_SEGMENT|4120,4128|false|false|false|||interval
Finding|Intellectual Product|SIMPLE_SEGMENT|4120,4128|false|false|false|C1552654|Parameterized Data Type - Interval|interval
Event|Event|SIMPLE_SEGMENT|4130,4142|false|false|false|||prolongation
Event|Event|SIMPLE_SEGMENT|4154,4161|false|false|false|||voltage
Event|Event|SIMPLE_SEGMENT|4177,4180|false|false|false|||aVL
Finding|Pathologic Function|SIMPLE_SEGMENT|4177,4180|false|false|false|C5237386|Atypical Vascular Proliferation|aVL
Event|Event|SIMPLE_SEGMENT|4200,4208|true|false|false|||criteria
Finding|Idea or Concept|SIMPLE_SEGMENT|4200,4208|true|false|false|C0243161|criteria|criteria
Finding|Functional Concept|SIMPLE_SEGMENT|4213,4217|true|false|false|C1552822|Table Cell Horizontal Align - left|left
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4213,4241|true|false|false|C3484363||left ventricular hypertrophy
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4213,4241|true|false|false|C0149721|Left Ventricular Hypertrophy|left ventricular hypertrophy
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4218,4229|true|false|false|C0018827|Heart Ventricle|ventricular
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4218,4241|true|false|false|C0340279|Ventricular hypertrophy|ventricular hypertrophy
Event|Event|SIMPLE_SEGMENT|4230,4241|true|false|false|||hypertrophy
Finding|Pathologic Function|SIMPLE_SEGMENT|4230,4241|true|false|false|C0020564|Hypertrophy|hypertrophy
Finding|Finding|SIMPLE_SEGMENT|4261,4271|false|false|false|C0429029|ST segment|ST segment
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|4272,4283|false|false|false|C0011570|Mental Depression|depressions
Event|Event|SIMPLE_SEGMENT|4272,4283|false|false|false|||depressions
Finding|Finding|SIMPLE_SEGMENT|4288,4294|false|false|false|C0429103|T wave feature|T wave
Finding|Gene or Genome|SIMPLE_SEGMENT|4290,4294|false|false|false|C1421479|WASF1 gene|wave
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|4290,4294|false|false|false|C0678544||wave
Event|Event|SIMPLE_SEGMENT|4295,4305|false|false|false|||inversions
Finding|Intellectual Product|SIMPLE_SEGMENT|4295,4305|false|false|false|C3481518|Inversions|inversions
Event|Event|SIMPLE_SEGMENT|4322,4325|false|false|false|||aVL
Finding|Pathologic Function|SIMPLE_SEGMENT|4322,4325|false|false|false|C5237386|Atypical Vascular Proliferation|aVL
Event|Event|SIMPLE_SEGMENT|4346,4351|false|false|false|||leads
Event|Event|SIMPLE_SEGMENT|4353,4361|false|false|false|||Compared
Event|Activity|SIMPLE_SEGMENT|4398,4402|false|false|false|C0871208|Rating (action)|rate
Event|Event|SIMPLE_SEGMENT|4398,4402|false|false|false|||rate
Finding|Idea or Concept|SIMPLE_SEGMENT|4398,4402|false|false|false|C1549480|Amount type - Rate|rate
Finding|Intellectual Product|SIMPLE_SEGMENT|4403,4407|false|false|false|C1720594|Then - dosing instruction fragment|then
Finding|Finding|SIMPLE_SEGMENT|4423,4429|false|false|false|C0429103|T wave feature|T wave
Finding|Gene or Genome|SIMPLE_SEGMENT|4425,4429|false|false|false|C1421479|WASF1 gene|wave
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|4425,4429|false|false|false|C0678544||wave
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|4430,4443|false|false|false|C0000768|Congenital Abnormality|abnormalities
Event|Event|SIMPLE_SEGMENT|4430,4443|false|false|false|||abnormalities
Finding|Functional Concept|SIMPLE_SEGMENT|4430,4443|false|false|false|C0000769|teratologic|abnormalities
Event|Event|SIMPLE_SEGMENT|4450,4457|false|false|false|||similar
Finding|Functional Concept|SIMPLE_SEGMENT|4468,4472|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4468,4496|false|false|false|C3484363||left ventricular hypertrophy
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4468,4496|false|false|false|C0149721|Left Ventricular Hypertrophy|left ventricular hypertrophy
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4473,4484|false|false|false|C0018827|Heart Ventricle|ventricular
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4473,4496|false|false|false|C0340279|Ventricular hypertrophy|ventricular hypertrophy
Event|Event|SIMPLE_SEGMENT|4485,4496|false|false|false|||hypertrophy
Finding|Pathologic Function|SIMPLE_SEGMENT|4485,4496|false|false|false|C0020564|Hypertrophy|hypertrophy
Finding|Intellectual Product|SIMPLE_SEGMENT|4509,4517|false|false|false|C1315013|Clinical NEC (not elsewhere classified in LNC)|Clinical
Event|Event|SIMPLE_SEGMENT|4518,4529|false|false|false|||correlation
Event|Event|SIMPLE_SEGMENT|4533,4542|false|false|false|||suggested
Event|Event|SIMPLE_SEGMENT|4545,4548|false|false|false|||CXR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4545,4548|false|false|false|C0039985|Plain chest X-ray|CXR
Finding|Body Substance|SIMPLE_SEGMENT|4553,4560|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|4553,4560|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|4553,4560|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4564,4570|false|false|false|C5889824||status
Event|Event|SIMPLE_SEGMENT|4564,4570|false|false|false|||status
Finding|Idea or Concept|SIMPLE_SEGMENT|4564,4570|false|false|false|C1546481|What subject filter - Status|status
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4576,4593|false|false|false|C1282959|Median Sternotomy|median sternotomy
Event|Event|SIMPLE_SEGMENT|4583,4593|false|false|false|||sternotomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4583,4593|false|false|false|C0185792|Sternotomy (procedure)|sternotomy
Event|Event|SIMPLE_SEGMENT|4598,4602|false|false|false|||CABG
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4598,4602|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4604,4609|false|false|false|C0018787;C4037974|Chest>Heart;Heart|Heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4604,4609|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|Heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|4604,4609|false|false|false|C0795691|HEART PROBLEM|Heart
Finding|Finding|SIMPLE_SEGMENT|4604,4614|false|false|false|C0744689|heart size|Heart size
Event|Event|SIMPLE_SEGMENT|4619,4625|false|false|false|||normal
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4627,4638|false|false|false|C0025066|Mediastinum|Mediastinal
Event|Event|SIMPLE_SEGMENT|4649,4657|false|false|false|||contours
Event|Event|SIMPLE_SEGMENT|4662,4671|false|false|false|||unchanged
Finding|Finding|SIMPLE_SEGMENT|4662,4671|false|false|false|C0442739||unchanged
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4673,4682|false|false|false|C0024109|Lung|Pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4673,4682|false|false|false|C2707265||Pulmonary
Finding|Finding|SIMPLE_SEGMENT|4673,4682|false|false|false|C4522268|Pulmonary (intended site)|Pulmonary
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|4684,4695|false|false|false|C3714653|Vasculature|vasculature
Event|Event|SIMPLE_SEGMENT|4699,4705|false|false|false|||normal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4716,4729|true|false|false|C0521530|Lung consolidation|consolidation
Event|Event|SIMPLE_SEGMENT|4716,4729|true|false|false|||consolidation
Anatomy|Tissue|SIMPLE_SEGMENT|4731,4738|true|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4731,4738|true|false|false|C0032226|Pleural Diseases|pleural
Finding|Body Substance|SIMPLE_SEGMENT|4731,4747|true|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Finding|Finding|SIMPLE_SEGMENT|4731,4747|true|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|4731,4747|true|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Event|Event|SIMPLE_SEGMENT|4739,4747|true|false|false|||effusion
Finding|Body Substance|SIMPLE_SEGMENT|4739,4747|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|SIMPLE_SEGMENT|4739,4747|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|4739,4747|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4752,4764|false|false|false|C0032326|Pneumothorax|pneumothorax
Event|Event|SIMPLE_SEGMENT|4752,4764|false|false|false|||pneumothorax
Event|Event|SIMPLE_SEGMENT|4768,4772|false|false|false|||seen
Finding|Intellectual Product|SIMPLE_SEGMENT|4777,4782|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4783,4790|true|false|false|C0262950;C4520924|Bone Tissue, Human;Skeletal bone|osseous
Anatomy|Tissue|SIMPLE_SEGMENT|4783,4790|true|false|false|C0262950;C4520924|Bone Tissue, Human;Skeletal bone|osseous
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|4791,4802|true|false|false|C0000768|Congenital Abnormality|abnormality
Event|Event|SIMPLE_SEGMENT|4791,4802|true|false|false|||abnormality
Finding|Finding|SIMPLE_SEGMENT|4791,4802|true|false|false|C1704258|Abnormality|abnormality
Event|Event|SIMPLE_SEGMENT|4807,4815|true|false|false|||detected
Event|Event|SIMPLE_SEGMENT|4817,4827|false|false|false|||IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|4817,4827|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|4817,4827|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|4832,4837|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4838,4853|true|false|false|C0553534|Cardiopulmonary|cardiopulmonary
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4838,4853|true|false|false|C4072686|Cardiovascular disease+Pulmonary disease|cardiopulmonary
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|4854,4865|true|false|false|C0000768|Congenital Abnormality|abnormality
Event|Event|SIMPLE_SEGMENT|4854,4865|true|false|false|||abnormality
Finding|Finding|SIMPLE_SEGMENT|4854,4865|true|false|false|C1704258|Abnormality|abnormality
Drug|Organic Chemical|SIMPLE_SEGMENT|4868,4880|false|false|false|C0012582|dipyridamole|Dipyridamole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4868,4880|false|false|false|C0012582|dipyridamole|Dipyridamole
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4881,4885|false|false|false|C5557372|Multiplexed Ion Beam Imaging|MIBI
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4886,4892|false|false|false|C1718621|W stress|Stress
Drug|Organic Chemical|SIMPLE_SEGMENT|4886,4892|false|false|false|C0723460|Stress bismuth subsalicylate|Stress
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4886,4892|false|false|false|C0723460|Stress bismuth subsalicylate|Stress
Finding|Finding|SIMPLE_SEGMENT|4886,4892|false|false|false|C0038435|Stress|Stress
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4886,4897|false|false|false|C0015260;C3494508|Exercise stress test;Stress Test|Stress test
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4893,4897|false|false|false|C4318744|Test - temporal region|test
Event|Event|SIMPLE_SEGMENT|4893,4897|false|false|false|||test
Finding|Functional Concept|SIMPLE_SEGMENT|4893,4897|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Finding|Intellectual Product|SIMPLE_SEGMENT|4893,4897|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4893,4897|false|false|false|C0456984|Test Result|test
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4893,4897|false|false|false|C0022885|Laboratory Procedures|test
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4924,4927|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|SIMPLE_SEGMENT|4924,4927|false|false|false|||HTN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4933,4936|false|false|false|C0085096|Peripheral Vascular Diseases|PVD
Event|Event|SIMPLE_SEGMENT|4933,4936|false|false|false|||PVD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4933,4936|false|false|false|C4521226|Pomalidomide/Bortezomib/Dexamethasone Regimen|PVD
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4941,4950|false|false|false|C0012000|Diastole|diastolic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4941,4954|false|false|false|C2183328|diastolic congestive heart failure|diastolic CHF
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4951,4954|false|false|false|C0262212|Choroidal fissure|CHF
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4951,4954|false|false|false|C0018802|Congestive heart failure|CHF
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4977,4981|false|false|false|C0228147|Structure of cisterna pontis|PCIs
Event|Event|SIMPLE_SEGMENT|4986,4990|false|false|false|||CABG
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4986,4990|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|5020,5029|false|false|false|C0001168|Complete obstruction|occlusion
Event|Event|SIMPLE_SEGMENT|5020,5029|false|false|false|||occlusion
Finding|Finding|SIMPLE_SEGMENT|5020,5029|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Functional Concept|SIMPLE_SEGMENT|5020,5029|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|5020,5029|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Pathologic Function|SIMPLE_SEGMENT|5020,5029|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Event|Event|SIMPLE_SEGMENT|5035,5043|false|false|false|||referred
Event|Event|SIMPLE_SEGMENT|5047,5055|false|false|false|||evaluate
Finding|Finding|SIMPLE_SEGMENT|5059,5067|false|false|false|C0741302|atypia morphology|atypical
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5068,5073|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|5068,5073|false|false|false|C0741025|Chest problem|chest
Finding|Sign or Symptom|SIMPLE_SEGMENT|5068,5084|false|false|false|C0235710|Chest discomfort|chest discomfort
Event|Event|SIMPLE_SEGMENT|5074,5084|false|false|false|||discomfort
Finding|Sign or Symptom|SIMPLE_SEGMENT|5074,5084|false|false|false|C2364135|Discomfort|discomfort
Finding|Body Substance|SIMPLE_SEGMENT|5091,5098|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|5091,5098|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|5091,5098|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|5103,5115|false|false|false|||administered
Finding|Conceptual Entity|SIMPLE_SEGMENT|5125,5131|false|false|false|C1532757|kg/min|kg/min
Drug|Organic Chemical|SIMPLE_SEGMENT|5135,5145|false|false|false|C0700020|Persantine|Persantine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5135,5145|false|false|false|C0700020|Persantine|Persantine
Event|Event|SIMPLE_SEGMENT|5135,5145|false|false|false|||Persantine
Event|Event|SIMPLE_SEGMENT|5154,5161|false|false|false|||minutes
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5176,5185|false|false|false|C0945766||procedure
Event|Event|SIMPLE_SEGMENT|5176,5185|false|false|false|||procedure
Event|Occupational Activity|SIMPLE_SEGMENT|5176,5185|false|false|false|C1546467|Act Class - procedure|procedure
Finding|Functional Concept|SIMPLE_SEGMENT|5176,5185|false|false|false|C2700391|Procedure (set of actions)|procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5176,5185|false|false|false|C0184661|Interventional procedure|procedure
Finding|Body Substance|SIMPLE_SEGMENT|5190,5197|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|5190,5197|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|5190,5197|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|5198,5206|false|false|false|||reported
Event|Event|SIMPLE_SEGMENT|5210,5218|false|false|false|||isolated
Finding|Functional Concept|SIMPLE_SEGMENT|5210,5218|false|false|false|C0205409;C1548221|Bed Status - Isolated;Isolated|isolated
Finding|Idea or Concept|SIMPLE_SEGMENT|5210,5218|false|false|false|C0205409;C1548221|Bed Status - Isolated;Isolated|isolated
Finding|Functional Concept|SIMPLE_SEGMENT|5220,5224|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5231,5236|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|5231,5236|false|false|false|C0741025|Chest problem|chest
Finding|Sign or Symptom|SIMPLE_SEGMENT|5231,5247|false|false|false|C0235710|Chest discomfort|chest discomfort
Event|Event|SIMPLE_SEGMENT|5237,5247|false|false|false|||discomfort
Finding|Sign or Symptom|SIMPLE_SEGMENT|5237,5247|false|false|false|C2364135|Discomfort|discomfort
Event|Event|SIMPLE_SEGMENT|5262,5269|false|false|false|||present
Finding|Finding|SIMPLE_SEGMENT|5262,5269|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|SIMPLE_SEGMENT|5262,5269|false|false|false|C0150312;C0449450|Present;Presentation|present
Event|Event|SIMPLE_SEGMENT|5277,5286|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|5277,5286|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|SIMPLE_SEGMENT|5295,5301|false|false|false|||tender
Finding|Intellectual Product|SIMPLE_SEGMENT|5305,5309|false|false|false|C1547225|Mild Severity of Illness Code|mild
Event|Event|SIMPLE_SEGMENT|5310,5319|false|false|false|||palpation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5310,5319|false|false|false|C0030247|Palpation|palpation
Event|Event|SIMPLE_SEGMENT|5332,5342|true|false|false|||discomfort
Finding|Sign or Symptom|SIMPLE_SEGMENT|5332,5342|true|false|false|C2364135|Discomfort|discomfort
Event|Event|SIMPLE_SEGMENT|5351,5357|true|false|false|||change
Event|Event|SIMPLE_SEGMENT|5361,5370|true|false|false|||intensity
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5382,5391|true|false|false|C0945766||procedure
Event|Event|SIMPLE_SEGMENT|5382,5391|true|false|false|||procedure
Event|Occupational Activity|SIMPLE_SEGMENT|5382,5391|true|false|false|C1546467|Act Class - procedure|procedure
Finding|Functional Concept|SIMPLE_SEGMENT|5382,5391|true|false|false|C2700391|Procedure (set of actions)|procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5382,5391|true|false|false|C0184661|Interventional procedure|procedure
Event|Event|SIMPLE_SEGMENT|5401,5409|false|false|false|||presence
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5401,5409|false|false|false|C0392148|Providing presence (regime/therapy)|presence
Finding|Finding|SIMPLE_SEGMENT|5401,5412|false|false|false|C0150312|Present|presence of
Finding|Finding|SIMPLE_SEGMENT|5424,5430|true|false|false|C0429103|T wave feature|T wave
Finding|Finding|SIMPLE_SEGMENT|5424,5438|true|false|false|C5780423|T wave changes|T wave changes
Finding|Gene or Genome|SIMPLE_SEGMENT|5426,5430|true|false|false|C1421479|WASF1 gene|wave
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|5426,5430|true|false|false|C0678544||wave
Event|Event|SIMPLE_SEGMENT|5431,5438|true|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|5431,5438|true|false|false|C0392747|Changing|changes
Finding|Functional Concept|SIMPLE_SEGMENT|5443,5453|true|false|false|C1524062|Additional|additional
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5454,5457|true|false|false|C0018064|Equine Gonadotropins|ECG
Drug|Hormone|SIMPLE_SEGMENT|5454,5457|true|false|false|C0018064|Equine Gonadotropins|ECG
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5454,5457|true|false|false|C0018064|Equine Gonadotropins|ECG
Event|Event|SIMPLE_SEGMENT|5454,5457|true|false|false|||ECG
Finding|Intellectual Product|SIMPLE_SEGMENT|5454,5457|true|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|ECG
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5454,5457|true|false|false|C1623258|Electrocardiography|ECG
Event|Event|SIMPLE_SEGMENT|5459,5466|true|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|5459,5466|true|false|false|C0392747|Changing|changes
Event|Event|SIMPLE_SEGMENT|5472,5477|true|false|false|||noted
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5489,5498|false|false|false|C0945766||procedure
Event|Event|SIMPLE_SEGMENT|5489,5498|false|false|false|||procedure
Event|Occupational Activity|SIMPLE_SEGMENT|5489,5498|false|false|false|C1546467|Act Class - procedure|procedure
Finding|Functional Concept|SIMPLE_SEGMENT|5489,5498|false|false|false|C2700391|Procedure (set of actions)|procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5489,5498|false|false|false|C0184661|Interventional procedure|procedure
Event|Event|SIMPLE_SEGMENT|5504,5515|false|false|false|||hemodynamic
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|5504,5515|false|false|false|C0019010|Hemodynamics|hemodynamic
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5504,5515|false|false|false|C4281788|hemodynamics (procedure)|hemodynamic
Event|Event|SIMPLE_SEGMENT|5517,5525|false|false|false|||response
Finding|Finding|SIMPLE_SEGMENT|5517,5525|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Intellectual Product|SIMPLE_SEGMENT|5517,5525|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Mental Process|SIMPLE_SEGMENT|5517,5525|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Drug|Organic Chemical|SIMPLE_SEGMENT|5533,5543|false|false|false|C0700020|Persantine|Persantine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5533,5543|false|false|false|C0700020|Persantine|Persantine
Event|Event|SIMPLE_SEGMENT|5544,5552|false|false|false|||infusion
Finding|Functional Concept|SIMPLE_SEGMENT|5544,5552|false|false|false|C1827465|Infusion route|infusion
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5544,5552|false|false|false|C0574032|Infusion procedures|infusion
Event|Event|SIMPLE_SEGMENT|5557,5568|false|false|false|||appropriate
Finding|Body Substance|SIMPLE_SEGMENT|5590,5597|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|5590,5597|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|5590,5597|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|5602,5614|false|false|false|||administered
Drug|Organic Chemical|SIMPLE_SEGMENT|5622,5635|false|false|false|C0002575|aminophylline|Aminophylline
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5622,5635|false|false|false|C0002575|aminophylline|Aminophylline
Event|Event|SIMPLE_SEGMENT|5622,5635|false|false|false|||Aminophylline
Event|Event|SIMPLE_SEGMENT|5641,5651|false|false|false|||IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|5641,5651|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|5641,5651|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Gene or Genome|SIMPLE_SEGMENT|5665,5669|true|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Finding|Intellectual Product|SIMPLE_SEGMENT|5665,5669|true|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Event|Event|SIMPLE_SEGMENT|5670,5678|true|false|false|||symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|5670,5678|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|5670,5678|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|5687,5697|true|false|false|C1524062|Additional|additional
Event|Event|SIMPLE_SEGMENT|5710,5717|true|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|5710,5717|true|false|false|C0392747|Changing|changes
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5723,5731|true|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|SIMPLE_SEGMENT|5723,5731|true|false|false|||baseline
Finding|Idea or Concept|SIMPLE_SEGMENT|5723,5731|true|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Event|Event|SIMPLE_SEGMENT|5733,5740|false|false|false|||Imaging
Finding|Finding|SIMPLE_SEGMENT|5733,5740|false|false|false|C0740845|Imaging problem|Imaging
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5733,5740|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|Imaging
Finding|Functional Concept|SIMPLE_SEGMENT|5744,5748|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5744,5767|false|false|false|C0503990|Cavity of left ventricle|Left ventricular cavity
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5744,5772|false|false|false|C0455830|Left ventricular cavity size|Left ventricular cavity size
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5749,5760|false|false|false|C0018827|Heart Ventricle|ventricular
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5749,5767|false|false|false|C0507083|Cavity of ventricle|ventricular cavity
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5761,5767|false|false|false|C0333343|Body cavities|cavity
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|5761,5767|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5761,5767|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Event|Event|SIMPLE_SEGMENT|5776,5782|false|false|false|||normal
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5786,5790|false|false|false|C1742913|REST protein, human|Rest
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5786,5790|false|false|false|C1742913|REST protein, human|Rest
Event|Event|SIMPLE_SEGMENT|5786,5790|false|false|false|||Rest
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|5786,5790|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|Rest
Finding|Gene or Genome|SIMPLE_SEGMENT|5786,5790|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|Rest
Finding|Molecular Function|SIMPLE_SEGMENT|5786,5790|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|Rest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5795,5801|false|false|false|C1718621|W stress|stress
Drug|Organic Chemical|SIMPLE_SEGMENT|5795,5801|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5795,5801|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Event|Event|SIMPLE_SEGMENT|5795,5801|false|false|false|||stress
Finding|Finding|SIMPLE_SEGMENT|5795,5801|false|false|false|C0038435|Stress|stress
Finding|Functional Concept|SIMPLE_SEGMENT|5802,5811|false|false|false|C4281794;C4723760|Perfusion (biological);Perfusion route|perfusion
Finding|Organism Function|SIMPLE_SEGMENT|5802,5811|false|false|false|C4281794;C4723760|Perfusion (biological);Perfusion route|perfusion
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5802,5811|false|false|false|C0031001;C4721534|Chemotherapeutic Perfusion;Perfusion (procedure)|perfusion
Event|Event|SIMPLE_SEGMENT|5812,5818|false|false|false|||images
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|5834,5840|false|false|false|C1522485|Tracer|tracer
Event|Event|SIMPLE_SEGMENT|5841,5847|false|false|false|||uptake
Finding|Cell Function|SIMPLE_SEGMENT|5841,5847|false|false|false|C0243144;C3888108;C3893696|Import into cell;Uptake;import across plasma membrane|uptake
Finding|Physiologic Function|SIMPLE_SEGMENT|5841,5847|false|false|false|C0243144;C3888108;C3893696|Import into cell;Uptake;import across plasma membrane|uptake
Finding|Functional Concept|SIMPLE_SEGMENT|5864,5868|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5864,5891|false|false|false|C0225899|Myocardium of left ventricle|left ventricular myocardium
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5869,5880|false|false|false|C0018827|Heart Ventricle|ventricular
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5869,5891|false|false|false|C0225880|Structure of myocardium of ventricle|ventricular myocardium
Anatomy|Tissue|SIMPLE_SEGMENT|5881,5891|false|false|false|C0027061|Myocardium|myocardium
Event|Event|SIMPLE_SEGMENT|5910,5915|false|false|false|||noted
Event|Event|SIMPLE_SEGMENT|5916,5925|false|false|false|||perfusion
Finding|Functional Concept|SIMPLE_SEGMENT|5916,5925|false|false|false|C4281794;C4723760|Perfusion (biological);Perfusion route|perfusion
Finding|Organism Function|SIMPLE_SEGMENT|5916,5925|false|false|false|C4281794;C4723760|Perfusion (biological);Perfusion route|perfusion
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5916,5925|false|false|false|C0031001;C4721534|Chemotherapeutic Perfusion;Perfusion (procedure)|perfusion
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5926,5932|false|false|false|C1861101|THYROID HORMONE PLASMA MEMBRANE TRANSPORT DEFECT|defect
Event|Event|SIMPLE_SEGMENT|5926,5932|false|false|false|||defect
Finding|Functional Concept|SIMPLE_SEGMENT|5926,5932|false|false|false|C1457869|Defect|defect
Event|Event|SIMPLE_SEGMENT|5933,5942|false|false|false|||involving
Event|Event|SIMPLE_SEGMENT|5971,5979|false|false|false|||resolved
Finding|Finding|SIMPLE_SEGMENT|5983,5988|false|false|false|C4266464|Gated|Gated
Event|Event|SIMPLE_SEGMENT|5989,5995|false|false|false|||images
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6010,6021|false|false|false|C1980023|Wall motion|wall motion
Event|Event|SIMPLE_SEGMENT|6015,6021|false|false|false|||motion
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|6015,6021|false|false|false|C0026597|Motion|motion
Event|Event|SIMPLE_SEGMENT|6038,6042|false|false|false|||left
Finding|Functional Concept|SIMPLE_SEGMENT|6038,6042|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6044,6055|false|false|false|C0018827|Heart Ventricle|ventricular
Finding|Physiologic Function|SIMPLE_SEGMENT|6044,6064|false|false|false|C2733340|Ventricular ejection|ventricular ejection
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6044,6073|false|false|false|C0042508|Ventricular Ejection Fraction|ventricular ejection fraction
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6056,6064|false|false|false|C0812388|Ejection time|ejection
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|6056,6064|false|false|false|C0336969|Ejection as a Sports activity|ejection
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|6056,6064|false|false|false|C0302131|Ejection as a Circumstance of Injury|ejection
Finding|Finding|SIMPLE_SEGMENT|6056,6073|false|false|false|C2020641;C2700378|Ejection fraction;stress echo measurements ejection fraction|ejection fraction
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6056,6073|false|false|false|C0489482|Ejection fraction (procedure)|ejection fraction
Event|Event|SIMPLE_SEGMENT|6065,6073|false|false|false|||fraction
Finding|Intellectual Product|SIMPLE_SEGMENT|6065,6073|false|false|false|C1554103|MDFAttributeType - Fraction|fraction
Event|Event|SIMPLE_SEGMENT|6082,6092|false|false|false|||IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|6082,6092|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|6082,6092|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Anatomy|Tissue|SIMPLE_SEGMENT|6101,6111|false|false|false|C0027061|Myocardium|myocardial
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6101,6127|false|false|false|C0841688|myocardial perfusion study|myocardial perfusion study
Event|Event|SIMPLE_SEGMENT|6112,6121|false|false|false|||perfusion
Finding|Functional Concept|SIMPLE_SEGMENT|6112,6121|false|false|false|C4281794;C4723760|Perfusion (biological);Perfusion route|perfusion
Finding|Organism Function|SIMPLE_SEGMENT|6112,6121|false|false|false|C4281794;C4723760|Perfusion (biological);Perfusion route|perfusion
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6112,6121|false|false|false|C0031001;C4721534|Chemotherapeutic Perfusion;Perfusion (procedure)|perfusion
Event|Event|SIMPLE_SEGMENT|6122,6127|false|false|false|||study
Finding|Intellectual Product|SIMPLE_SEGMENT|6122,6127|false|false|false|C1705923|Study Object|study
Procedure|Research Activity|SIMPLE_SEGMENT|6122,6127|false|false|false|C0008972;C0947630;C2603343|Clinical Research;Scientific Study;Study|study
Finding|Intellectual Product|SIMPLE_SEGMENT|6129,6137|false|false|false|C1552654|Parameterized Data Type - Interval|Interval
Event|Event|SIMPLE_SEGMENT|6139,6152|false|false|false|||normalization
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6162,6165|false|false|false|C2987138|Methylcytosine Dioxygenase TET1|LCx
Drug|Enzyme|SIMPLE_SEGMENT|6162,6165|false|false|false|C2987138|Methylcytosine Dioxygenase TET1|LCx
Finding|Gene or Genome|SIMPLE_SEGMENT|6162,6165|false|false|false|C1428863;C2987137|TET1 gene;TET1 wt Allele|LCx
Event|Event|SIMPLE_SEGMENT|6176,6185|false|false|false|||perfusion
Finding|Functional Concept|SIMPLE_SEGMENT|6176,6185|false|false|false|C4281794;C4723760|Perfusion (biological);Perfusion route|perfusion
Finding|Organism Function|SIMPLE_SEGMENT|6176,6185|false|false|false|C4281794;C4723760|Perfusion (biological);Perfusion route|perfusion
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6176,6185|false|false|false|C0031001;C4721534|Chemotherapeutic Perfusion;Perfusion (procedure)|perfusion
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6186,6192|false|false|false|C1861101|THYROID HORMONE PLASMA MEMBRANE TRANSPORT DEFECT|defect
Event|Event|SIMPLE_SEGMENT|6186,6192|false|false|false|||defect
Finding|Functional Concept|SIMPLE_SEGMENT|6186,6192|false|false|false|C1457869|Defect|defect
Finding|Intellectual Product|SIMPLE_SEGMENT|6196,6201|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|Brief
Finding|Idea or Concept|SIMPLE_SEGMENT|6202,6210|false|false|false|C1547192|Organization unit type - Hospital|Hospital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6202,6217|false|false|false|C0488549||Hospital Course
Finding|Finding|SIMPLE_SEGMENT|6202,6217|false|false|false|C0489547|Hospital course|Hospital Course
Finding|Gene or Genome|SIMPLE_SEGMENT|6238,6242|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Finding|Intellectual Product|SIMPLE_SEGMENT|6238,6242|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Finding|Classification|SIMPLE_SEGMENT|6238,6244|false|false|false|C0441730|Type 2|type 2
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6238,6253|false|false|false|C0011860|Diabetes Mellitus, Non-Insulin-Dependent|type 2 diabetes
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6238,6262|false|false|false|C0011860|Diabetes Mellitus, Non-Insulin-Dependent|type 2 diabetes mellitus
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6245,6253|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|diabetes
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6245,6262|false|false|false|C0011849|Diabetes Mellitus|diabetes mellitus
Event|Event|SIMPLE_SEGMENT|6254,6262|false|false|false|||mellitus
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6266,6273|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|SIMPLE_SEGMENT|6266,6273|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6266,6273|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|SIMPLE_SEGMENT|6266,6273|false|false|false|||insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|6266,6273|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6266,6273|false|false|false|C0202098|Insulin measurement|insulin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6275,6278|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6275,6278|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|6275,6278|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|6275,6278|false|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|6275,6278|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6275,6278|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|6275,6278|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6275,6278|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Event|Event|SIMPLE_SEGMENT|6284,6286|false|false|false|||MI
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|6301,6305|false|false|false|C0228147|Structure of cisterna pontis|PCIs
Event|Event|SIMPLE_SEGMENT|6310,6314|false|false|false|||CABG
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6310,6314|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6325,6328|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6325,6328|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|SIMPLE_SEGMENT|6325,6328|false|false|false|||LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|6325,6328|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Event|Event|SIMPLE_SEGMENT|6352,6357|false|false|false|||known
Finding|Finding|SIMPLE_SEGMENT|6358,6366|false|false|false|C0028778;C1947917|Obstruction;Occluded|occluded
Finding|Functional Concept|SIMPLE_SEGMENT|6358,6366|false|false|false|C0028778;C1947917|Obstruction;Occluded|occluded
Finding|Intellectual Product|SIMPLE_SEGMENT|6376,6383|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|6376,6383|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6376,6397|false|false|false|C0340288|Stable angina|chronic stable angina
Finding|Intellectual Product|SIMPLE_SEGMENT|6384,6390|false|false|false|C1547311|Patient Condition Code - Stable|stable
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6384,6397|false|false|false|C0340288|Stable angina|stable angina
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6391,6397|false|false|false|C2926611||angina
Event|Event|SIMPLE_SEGMENT|6391,6397|false|false|false|||angina
Finding|Finding|SIMPLE_SEGMENT|6391,6397|false|false|false|C0002962;C2024883|Angina Pectoris|angina
Finding|Sign or Symptom|SIMPLE_SEGMENT|6391,6397|false|false|false|C0002962;C2024883|Angina Pectoris|angina
Event|Event|SIMPLE_SEGMENT|6399,6407|false|false|false|||admitted
Event|Event|SIMPLE_SEGMENT|6413,6421|false|false|false|||atypical
Finding|Finding|SIMPLE_SEGMENT|6413,6421|false|false|false|C0741302|atypia morphology|atypical
Event|Event|SIMPLE_SEGMENT|6423,6431|false|false|false|||stabbing
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6439,6444|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|6439,6444|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6439,6449|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|6439,6449|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6445,6449|false|true|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|6445,6449|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|6445,6449|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|6445,6449|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6454,6459|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|SIMPLE_SEGMENT|6454,6459|false|false|false|C0741025|Chest problem|Chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6454,6464|false|false|false|C2926613||Chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|6454,6464|false|false|false|C0008031|Chest Pain|Chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6460,6464|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|6460,6464|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|6460,6464|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|6460,6464|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Body Substance|SIMPLE_SEGMENT|6480,6487|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|6480,6487|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|6480,6487|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|6492,6499|false|false|false|||started
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6505,6512|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Organic Chemical|SIMPLE_SEGMENT|6505,6512|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6505,6512|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Event|Event|SIMPLE_SEGMENT|6505,6512|false|false|false|||heparin
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|6529,6532|false|false|false|C0262187|anterior calcarine sulcus (human only)|ACS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6529,6532|false|false|false|C0742343;C0796147|Acrocallosal Syndrome;Acute Chest Syndrome|ACS
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6529,6532|false|false|false|C4042561|ACSS2 protein, human|ACS
Drug|Enzyme|SIMPLE_SEGMENT|6529,6532|false|false|false|C4042561|ACSS2 protein, human|ACS
Event|Event|SIMPLE_SEGMENT|6529,6532|false|false|false|||ACS
Finding|Gene or Genome|SIMPLE_SEGMENT|6529,6532|false|false|false|C1150760;C1424787;C1825842;C1842089;C2266615;C4318612;C5400867;C5551036|ACCS gene;ACS - Activity Card Sort;ACSS2 gene;ACSS2 wt Allele;American Community Survey;CO-methylating acetyl-CoA synthase activity;PLA2G15 gene;acetate-CoA ligase activity|ACS
Finding|Intellectual Product|SIMPLE_SEGMENT|6529,6532|false|false|false|C1150760;C1424787;C1825842;C1842089;C2266615;C4318612;C5400867;C5551036|ACCS gene;ACS - Activity Card Sort;ACSS2 gene;ACSS2 wt Allele;American Community Survey;CO-methylating acetyl-CoA synthase activity;PLA2G15 gene;acetate-CoA ligase activity|ACS
Finding|Molecular Function|SIMPLE_SEGMENT|6529,6532|false|false|false|C1150760;C1424787;C1825842;C1842089;C2266615;C4318612;C5400867;C5551036|ACCS gene;ACS - Activity Card Sort;ACSS2 gene;ACSS2 wt Allele;American Community Survey;CO-methylating acetyl-CoA synthase activity;PLA2G15 gene;acetate-CoA ligase activity|ACS
Finding|Finding|SIMPLE_SEGMENT|6533,6541|false|false|false|C0442711;C1507394;C1522729;C2348563;C3715209|Clinical trial protocol document;Library Protocol;Protocol - answer to question;Protocols documentation;Study Protocol|protocol
Finding|Intellectual Product|SIMPLE_SEGMENT|6533,6541|false|false|false|C0442711;C1507394;C1522729;C2348563;C3715209|Clinical trial protocol document;Library Protocol;Protocol - answer to question;Protocols documentation;Study Protocol|protocol
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6542,6553|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6542,6553|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|6542,6553|false|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|6542,6553|false|false|false|C4284232|Medications|medications
Finding|Idea or Concept|SIMPLE_SEGMENT|6559,6563|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|6559,6563|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|6559,6563|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|6564,6572|false|false|false|C0126174|losartan|losartan
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6564,6572|false|false|false|C0126174|losartan|losartan
Event|Event|SIMPLE_SEGMENT|6564,6572|false|false|false|||losartan
Drug|Organic Chemical|SIMPLE_SEGMENT|6578,6588|false|false|false|C0016860|furosemide|furosemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6578,6588|false|false|false|C0016860|furosemide|furosemide
Event|Event|SIMPLE_SEGMENT|6578,6588|false|false|false|||furosemide
Event|Event|SIMPLE_SEGMENT|6594,6598|false|false|false|||held
Finding|Finding|SIMPLE_SEGMENT|6606,6609|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|SIMPLE_SEGMENT|6606,6609|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Finding|SIMPLE_SEGMENT|6606,6625|false|false|false|C0020649|Hypotension|low blood pressures
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6610,6615|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|6610,6615|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|6610,6615|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Finding|SIMPLE_SEGMENT|6610,6625|false|false|false|C1272641|Systemic arterial pressure|blood pressures
Event|Event|SIMPLE_SEGMENT|6616,6625|false|false|false|||pressures
Finding|Finding|SIMPLE_SEGMENT|6616,6625|false|false|false|C0460139|Pressure (finding)|pressures
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|6616,6625|false|false|false|C0033095||pressures
Event|Event|SIMPLE_SEGMENT|6627,6636|false|false|false|||Suspicion
Finding|Mental Process|SIMPLE_SEGMENT|6627,6636|false|false|false|C0242114|Suspicion|Suspicion
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6642,6649|true|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|6642,6649|true|false|false|C1314974|Cardiac attachment|cardiac
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6642,6658|true|false|false|C0741922|CARDIAC ETIOLOGY|cardiac etiology
Event|Event|SIMPLE_SEGMENT|6650,6658|true|false|false|||etiology
Finding|Conceptual Entity|SIMPLE_SEGMENT|6650,6658|true|false|false|C0015127;C1314792;C1524003|Etiology;Etiology aspects;Science of Etiology|etiology
Finding|Functional Concept|SIMPLE_SEGMENT|6650,6658|true|false|false|C0015127;C1314792;C1524003|Etiology;Etiology aspects;Science of Etiology|etiology
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6662,6667|true|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|6662,6667|true|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6662,6672|true|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|6662,6672|true|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6668,6672|true|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|6668,6672|true|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|6668,6672|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|6668,6672|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|6692,6696|true|false|false|||high
Finding|Finding|SIMPLE_SEGMENT|6692,6696|true|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|SIMPLE_SEGMENT|6692,6696|true|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|SIMPLE_SEGMENT|6692,6696|true|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Event|Event|SIMPLE_SEGMENT|6719,6726|false|false|false|||ongoing
Finding|Idea or Concept|SIMPLE_SEGMENT|6719,6726|false|false|false|C0549178|Continuous|ongoing
Finding|Functional Concept|SIMPLE_SEGMENT|6731,6735|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6742,6747|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|6742,6747|false|false|false|C0741025|Chest problem|chest
Finding|Sign or Symptom|SIMPLE_SEGMENT|6742,6758|false|false|false|C0235710|Chest discomfort|chest discomfort
Event|Event|SIMPLE_SEGMENT|6748,6758|false|false|false|||discomfort
Finding|Sign or Symptom|SIMPLE_SEGMENT|6748,6758|false|false|false|C2364135|Discomfort|discomfort
Event|Event|SIMPLE_SEGMENT|6759,6770|false|false|false|||exacerbated
Event|Event|SIMPLE_SEGMENT|6775,6782|false|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|6775,6782|false|false|false|C0392747|Changing|changes
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6804,6809|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|6804,6809|false|false|false|C0741025|Chest problem|chest
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6804,6814|false|false|false|C0205076;C4266615|Chest wall structure;Chest>Chest wall|chest wall
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6804,6814|false|false|false|C0205076;C4266615|Chest wall structure;Chest>Chest wall|chest wall
Finding|Finding|SIMPLE_SEGMENT|6804,6825|false|false|false|C0239008|Chest wall tenderness|chest wall tenderness
Event|Event|SIMPLE_SEGMENT|6815,6825|false|false|false|||tenderness
Finding|Mental Process|SIMPLE_SEGMENT|6815,6825|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|SIMPLE_SEGMENT|6815,6825|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6829,6834|false|false|false|C1570446|TNFSF14 protein, human|light
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6829,6834|false|false|false|C1570446|TNFSF14 protein, human|light
Event|Event|SIMPLE_SEGMENT|6829,6834|false|false|false|||light
Finding|Finding|SIMPLE_SEGMENT|6829,6834|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Functional Concept|SIMPLE_SEGMENT|6829,6834|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Gene or Genome|SIMPLE_SEGMENT|6829,6834|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|6829,6834|false|false|false|C0023693|Light|light
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6829,6834|false|false|false|C0031765|Phototherapy|light
Event|Event|SIMPLE_SEGMENT|6836,6845|false|false|false|||palpation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6836,6845|false|false|false|C0030247|Palpation|palpation
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6865,6870|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|6865,6870|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6865,6875|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|6865,6875|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6871,6875|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|6871,6875|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|6871,6875|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|6871,6875|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6877,6885|false|false|false|C0041199|Troponin|troponin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6877,6885|false|false|false|C0041199|Troponin|troponin
Event|Event|SIMPLE_SEGMENT|6877,6885|false|false|false|||troponin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6877,6885|false|false|false|C0523952|Troponin measurement|troponin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6877,6887|false|false|false|C0077404|Troponin T|troponin-T
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6877,6887|false|false|false|C0077404|Troponin T|troponin-T
Event|Event|SIMPLE_SEGMENT|6886,6887|false|false|false|||T
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6892,6897|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|SIMPLE_SEGMENT|6892,6897|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|SIMPLE_SEGMENT|6892,6897|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6892,6897|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Event|Event|SIMPLE_SEGMENT|6895,6897|false|false|false|||MB
Event|Event|SIMPLE_SEGMENT|6899,6907|false|false|false|||negative
Finding|Classification|SIMPLE_SEGMENT|6899,6907|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|6899,6907|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6899,6907|false|false|false|C5237010|Expression Negative|negative
Event|Event|SIMPLE_SEGMENT|6915,6919|false|false|false|||EKGs
Finding|Intellectual Product|SIMPLE_SEGMENT|6915,6919|false|false|false|C0013798|Electrocardiogram|EKGs
Finding|Idea or Concept|SIMPLE_SEGMENT|6920,6926|false|false|false|C0750554|MOSTLY|mostly
Event|Event|SIMPLE_SEGMENT|6927,6936|false|false|false|||unchanged
Finding|Finding|SIMPLE_SEGMENT|6927,6936|false|false|false|C0442739||unchanged
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6966,6969|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6966,6969|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|6966,6969|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|6966,6969|false|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|6966,6969|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6966,6969|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|6966,6969|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6966,6969|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6973,6984|false|false|false|C0042402;C3537240|Vasodilator Agents;Vasodilator [EPC]|vasodilator
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6985,7004|false|false|false|C2825165|Nuclear stress test|nuclear stress test
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6993,6999|false|false|false|C1718621|W stress|stress
Drug|Organic Chemical|SIMPLE_SEGMENT|6993,6999|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6993,6999|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Finding|Finding|SIMPLE_SEGMENT|6993,6999|false|false|false|C0038435|Stress|stress
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6993,7004|false|false|false|C0015260;C3494508|Exercise stress test;Stress Test|stress test
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7000,7004|false|false|false|C4318744|Test - temporal region|test
Event|Event|SIMPLE_SEGMENT|7000,7004|false|false|false|||test
Finding|Functional Concept|SIMPLE_SEGMENT|7000,7004|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Finding|Intellectual Product|SIMPLE_SEGMENT|7000,7004|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|7000,7004|false|false|false|C0456984|Test Result|test
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7000,7004|false|false|false|C0022885|Laboratory Procedures|test
Event|Event|SIMPLE_SEGMENT|7028,7038|false|false|false|||reassuring
Procedure|Health Care Activity|SIMPLE_SEGMENT|7028,7038|false|false|false|C0557055|Reassuring (procedure)|reassuring
Event|Event|SIMPLE_SEGMENT|7044,7054|true|false|false|||discomfort
Finding|Sign or Symptom|SIMPLE_SEGMENT|7044,7054|true|false|false|C2364135|Discomfort|discomfort
Event|Event|SIMPLE_SEGMENT|7063,7069|true|false|false|||change
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7095,7101|true|false|false|C1718621|W stress|stress
Drug|Organic Chemical|SIMPLE_SEGMENT|7095,7101|true|false|false|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7095,7101|true|false|false|C0723460|Stress bismuth subsalicylate|stress
Finding|Finding|SIMPLE_SEGMENT|7095,7101|true|false|false|C0038435|Stress|stress
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7095,7106|true|false|false|C0015260;C3494508|Exercise stress test;Stress Test|stress test
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7102,7106|false|false|false|C4318744|Test - temporal region|test
Finding|Functional Concept|SIMPLE_SEGMENT|7102,7106|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Finding|Intellectual Product|SIMPLE_SEGMENT|7102,7106|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|7102,7106|false|false|false|C0456984|Test Result|test
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7102,7106|false|false|false|C0022885|Laboratory Procedures|test
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7102,7111|false|false|false|C0038577|Substance Abuse Detection|test drug
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7107,7111|false|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|drug
Event|Event|SIMPLE_SEGMENT|7107,7111|false|false|false|||drug
Finding|Finding|SIMPLE_SEGMENT|7107,7111|false|false|false|C0740721|Drug problem|drug
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7107,7120|false|false|false|C0392877|infusion of drug|drug infusion
Event|Event|SIMPLE_SEGMENT|7112,7120|false|false|false|||infusion
Finding|Functional Concept|SIMPLE_SEGMENT|7112,7120|false|false|false|C1827465|Infusion route|infusion
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7112,7120|false|false|false|C0574032|Infusion procedures|infusion
Event|Event|SIMPLE_SEGMENT|7129,7137|false|false|false|||presence
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7129,7137|false|false|false|C0392148|Providing presence (regime/therapy)|presence
Finding|Finding|SIMPLE_SEGMENT|7129,7140|false|false|false|C0150312|Present|presence of
Finding|Gene or Genome|SIMPLE_SEGMENT|7155,7159|true|false|false|C1421479|WASF1 gene|wave
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|7155,7159|true|false|false|C0678544||wave
Event|Event|SIMPLE_SEGMENT|7160,7167|true|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|7160,7167|true|false|false|C0392747|Changing|changes
Finding|Functional Concept|SIMPLE_SEGMENT|7172,7182|true|false|false|C1524062|Additional|additional
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7183,7186|true|false|false|C0018064|Equine Gonadotropins|ECG
Drug|Hormone|SIMPLE_SEGMENT|7183,7186|true|false|false|C0018064|Equine Gonadotropins|ECG
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7183,7186|true|false|false|C0018064|Equine Gonadotropins|ECG
Event|Event|SIMPLE_SEGMENT|7183,7186|true|false|false|||ECG
Finding|Intellectual Product|SIMPLE_SEGMENT|7183,7186|true|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|ECG
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7183,7186|true|false|false|C1623258|Electrocardiography|ECG
Event|Event|SIMPLE_SEGMENT|7187,7194|true|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|7187,7194|true|false|false|C0392747|Changing|changes
Event|Event|SIMPLE_SEGMENT|7200,7205|true|false|false|||noted
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7218,7227|false|false|false|C0945766||procedure
Event|Event|SIMPLE_SEGMENT|7218,7227|false|false|false|||procedure
Event|Occupational Activity|SIMPLE_SEGMENT|7218,7227|false|false|false|C1546467|Act Class - procedure|procedure
Finding|Functional Concept|SIMPLE_SEGMENT|7218,7227|false|false|false|C2700391|Procedure (set of actions)|procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7218,7227|false|false|false|C0184661|Interventional procedure|procedure
Event|Event|SIMPLE_SEGMENT|7233,7244|false|false|false|||hemodynamic
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|7233,7244|false|false|false|C0019010|Hemodynamics|hemodynamic
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7233,7244|false|false|false|C4281788|hemodynamics (procedure)|hemodynamic
Event|Event|SIMPLE_SEGMENT|7245,7253|false|false|false|||response
Finding|Finding|SIMPLE_SEGMENT|7245,7253|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Intellectual Product|SIMPLE_SEGMENT|7245,7253|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Mental Process|SIMPLE_SEGMENT|7245,7253|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Drug|Organic Chemical|SIMPLE_SEGMENT|7261,7271|false|false|false|C0700020|Persantine|Persantine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7261,7271|false|false|false|C0700020|Persantine|Persantine
Event|Event|SIMPLE_SEGMENT|7272,7280|false|false|false|||infusion
Finding|Functional Concept|SIMPLE_SEGMENT|7272,7280|false|false|false|C1827465|Infusion route|infusion
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7272,7280|false|false|false|C0574032|Infusion procedures|infusion
Event|Event|SIMPLE_SEGMENT|7286,7297|false|false|false|||appropriate
Event|Event|SIMPLE_SEGMENT|7303,7312|false|false|false|||perfusion
Finding|Functional Concept|SIMPLE_SEGMENT|7303,7312|false|false|false|C4281794;C4723760|Perfusion (biological);Perfusion route|perfusion
Finding|Organism Function|SIMPLE_SEGMENT|7303,7312|false|false|false|C4281794;C4723760|Perfusion (biological);Perfusion route|perfusion
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7303,7312|false|false|false|C0031001;C4721534|Chemotherapeutic Perfusion;Perfusion (procedure)|perfusion
Event|Event|SIMPLE_SEGMENT|7313,7318|false|false|false|||study
Finding|Intellectual Product|SIMPLE_SEGMENT|7313,7318|false|false|false|C1705923|Study Object|study
Procedure|Research Activity|SIMPLE_SEGMENT|7313,7318|false|false|false|C0008972;C0947630;C2603343|Clinical Research;Scientific Study;Study|study
Event|Event|SIMPLE_SEGMENT|7323,7329|false|false|false|||normal
Event|Event|SIMPLE_SEGMENT|7335,7343|false|false|false|||interval
Finding|Intellectual Product|SIMPLE_SEGMENT|7335,7343|false|false|false|C1552654|Parameterized Data Type - Interval|interval
Event|Event|SIMPLE_SEGMENT|7345,7358|false|false|false|||normalization
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7368,7371|false|false|false|C2987138|Methylcytosine Dioxygenase TET1|LCx
Drug|Enzyme|SIMPLE_SEGMENT|7368,7371|false|false|false|C2987138|Methylcytosine Dioxygenase TET1|LCx
Finding|Gene or Genome|SIMPLE_SEGMENT|7368,7371|false|false|false|C1428863;C2987137|TET1 gene;TET1 wt Allele|LCx
Event|Event|SIMPLE_SEGMENT|7382,7391|false|false|false|||perfusion
Finding|Functional Concept|SIMPLE_SEGMENT|7382,7391|false|false|false|C4281794;C4723760|Perfusion (biological);Perfusion route|perfusion
Finding|Organism Function|SIMPLE_SEGMENT|7382,7391|false|false|false|C4281794;C4723760|Perfusion (biological);Perfusion route|perfusion
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7382,7391|false|false|false|C0031001;C4721534|Chemotherapeutic Perfusion;Perfusion (procedure)|perfusion
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7392,7398|false|false|false|C1861101|THYROID HORMONE PLASMA MEMBRANE TRANSPORT DEFECT|defect
Event|Event|SIMPLE_SEGMENT|7392,7398|false|false|false|||defect
Finding|Functional Concept|SIMPLE_SEGMENT|7392,7398|false|false|false|C1457869|Defect|defect
Event|Event|SIMPLE_SEGMENT|7400,7405|false|false|false|||Given
Event|Event|SIMPLE_SEGMENT|7420,7427|false|false|false|||quality
Event|Event|SIMPLE_SEGMENT|7432,7442|false|false|false|||tenderness
Finding|Mental Process|SIMPLE_SEGMENT|7432,7442|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|SIMPLE_SEGMENT|7432,7442|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Event|Event|SIMPLE_SEGMENT|7446,7455|false|false|false|||palpation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7446,7455|false|false|false|C0030247|Palpation|palpation
Event|Governmental or Regulatory Activity|SIMPLE_SEGMENT|7463,7467|false|false|false|C1510751|Academic Research Enhancement Awards|area
Event|Event|SIMPLE_SEGMENT|7472,7482|false|false|false|||discomfort
Finding|Sign or Symptom|SIMPLE_SEGMENT|7472,7482|false|false|false|C2364135|Discomfort|discomfort
Event|Event|SIMPLE_SEGMENT|7488,7496|false|false|false|||symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|7488,7496|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|7488,7496|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Idea or Concept|SIMPLE_SEGMENT|7502,7513|false|false|false|C0750501|most likely|most likely
Finding|Finding|SIMPLE_SEGMENT|7507,7513|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|7507,7513|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Drug|Organic Chemical|SIMPLE_SEGMENT|7514,7521|false|true|false|C0163712|Relate - vinyl resin|related
Event|Event|SIMPLE_SEGMENT|7514,7521|false|false|false|||related
Finding|Finding|SIMPLE_SEGMENT|7514,7521|false|true|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Finding|Functional Concept|SIMPLE_SEGMENT|7514,7521|false|true|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7526,7541|false|false|false|C0040213;C5779793|Costal chondritis;Tietze's Syndrome|costochondritis
Event|Event|SIMPLE_SEGMENT|7526,7541|false|false|false|||costochondritis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7551,7566|false|false|false|C2707260||musculoskeletal
Finding|Functional Concept|SIMPLE_SEGMENT|7551,7566|false|false|false|C0497254|Musculoskeletal|musculoskeletal
Event|Event|SIMPLE_SEGMENT|7567,7573|false|false|false|||causes
Finding|Functional Concept|SIMPLE_SEGMENT|7567,7573|false|false|false|C0015127;C1314792|Etiology;Etiology aspects|causes
Event|Event|SIMPLE_SEGMENT|7583,7590|false|false|false|||started
Drug|Organic Chemical|SIMPLE_SEGMENT|7595,7602|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7595,7602|false|false|false|C0004057|aspirin|aspirin
Event|Event|SIMPLE_SEGMENT|7595,7602|false|false|false|||aspirin
Event|Event|SIMPLE_SEGMENT|7628,7633|false|false|false|||trial
Procedure|Research Activity|SIMPLE_SEGMENT|7628,7633|false|false|false|C0008976|Clinical Trials|trial
Event|Event|SIMPLE_SEGMENT|7650,7658|false|false|false|||continue
Finding|Intellectual Product|SIMPLE_SEGMENT|7671,7675|false|false|false|C1561540|Transaction counts and value totals - week|week
Event|Event|SIMPLE_SEGMENT|7679,7687|false|false|false|||symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|7679,7687|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|7679,7687|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|SIMPLE_SEGMENT|7688,7695|false|false|false|||improve
Event|Event|SIMPLE_SEGMENT|7698,7705|false|false|false|||Chronic
Finding|Intellectual Product|SIMPLE_SEGMENT|7698,7705|false|false|false|C1547296|Chronic - Admission Level of Care Code|Chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|7698,7705|false|false|false|C1555457|Provision of recurring care for chronic illness|Chronic
Finding|Functional Concept|SIMPLE_SEGMENT|7706,7713|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Idea or Concept|SIMPLE_SEGMENT|7706,7713|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Intellectual Product|SIMPLE_SEGMENT|7706,7713|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|7706,7713|false|false|false|C0199168|Medical service|medical
Event|Event|SIMPLE_SEGMENT|7714,7722|false|false|false|||problems
Finding|Idea or Concept|SIMPLE_SEGMENT|7714,7722|false|false|false|C1546466|Problems - What subject filter|problems
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7726,7734|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|Diabetes
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7726,7743|false|false|false|C0011849|Diabetes Mellitus|Diabetes mellitus
Event|Event|SIMPLE_SEGMENT|7735,7743|false|false|false|||mellitus
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7755,7762|false|false|false|C1314782|Levemir|levemir
Drug|Hormone|SIMPLE_SEGMENT|7755,7762|false|false|false|C1314782|Levemir|levemir
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7755,7762|false|false|false|C1314782|Levemir|levemir
Event|Event|SIMPLE_SEGMENT|7755,7762|false|false|false|||levemir
Event|Event|SIMPLE_SEGMENT|7771,7779|false|false|false|||switched
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7794,7799|false|false|false|C0222045|Integumentary scale|scale
Event|Activity|SIMPLE_SEGMENT|7794,7799|false|false|false|C1947916|Scaling|scale
Event|Event|SIMPLE_SEGMENT|7794,7799|false|false|false|||scale
Finding|Conceptual Entity|SIMPLE_SEGMENT|7794,7799|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|scale
Finding|Intellectual Product|SIMPLE_SEGMENT|7794,7799|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|scale
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7803,7810|false|false|false|C0528249|Humalog|Humalog
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7803,7810|false|false|false|C0528249|Humalog|Humalog
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7814,7826|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|SIMPLE_SEGMENT|7814,7826|false|false|false|||Hypertension
Drug|Organic Chemical|SIMPLE_SEGMENT|7828,7836|false|false|false|C0126174|losartan|Losartan
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7828,7836|false|false|false|C0126174|losartan|Losartan
Event|Event|SIMPLE_SEGMENT|7828,7836|false|false|false|||Losartan
Event|Event|SIMPLE_SEGMENT|7841,7845|false|false|false|||held
Finding|Idea or Concept|SIMPLE_SEGMENT|7849,7854|false|false|false|C1552828|Table Frame - above|above
Event|Event|SIMPLE_SEGMENT|7862,7873|false|false|false|||hypotension
Finding|Finding|SIMPLE_SEGMENT|7862,7873|false|false|false|C0020649|Hypotension|hypotension
Finding|Intellectual Product|SIMPLE_SEGMENT|7879,7883|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Organic Chemical|SIMPLE_SEGMENT|7890,7900|false|false|false|C0022251|isosorbide|isosorbide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7890,7900|false|false|false|C0022251|isosorbide|isosorbide
Drug|Organic Chemical|SIMPLE_SEGMENT|7890,7912|false|false|false|C0064079|isosorbide mononitrate|isosorbide mononitrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7890,7912|false|false|false|C0064079|isosorbide mononitrate|isosorbide mononitrate
Event|Event|SIMPLE_SEGMENT|7901,7912|false|false|false|||mononitrate
Event|Event|SIMPLE_SEGMENT|7917,7925|false|false|false|||switched
Drug|Organic Chemical|SIMPLE_SEGMENT|7942,7952|false|false|false|C0022251|isosorbide|isosorbide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7942,7952|false|false|false|C0022251|isosorbide|isosorbide
Drug|Organic Chemical|SIMPLE_SEGMENT|7942,7962|false|false|false|C0022252|isosorbide dinitrate|isosorbide dinitrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7942,7962|false|false|false|C0022252|isosorbide dinitrate|isosorbide dinitrate
Event|Event|SIMPLE_SEGMENT|7963,7966|false|false|false|||TID
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7979,7993|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|hyperlipidemia
Event|Event|SIMPLE_SEGMENT|7979,7993|false|false|false|||hyperlipidemia
Finding|Finding|SIMPLE_SEGMENT|7979,7993|false|false|false|C0428465|Serum lipids high (finding)|hyperlipidemia
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7995,7999|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7995,7999|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|SIMPLE_SEGMENT|7995,7999|false|false|false|||COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|7995,7999|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8004,8008|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Event|Event|SIMPLE_SEGMENT|8004,8008|false|false|false|||GERD
Finding|Idea or Concept|SIMPLE_SEGMENT|8014,8018|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|8014,8018|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|8014,8018|false|false|false|C1553498|home health encounter|home
Event|Event|SIMPLE_SEGMENT|8019,8027|false|false|false|||regimens
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8019,8027|false|false|false|C0040808|Treatment Protocols|regimens
Event|Event|SIMPLE_SEGMENT|8034,8043|false|false|false|||continued
Finding|Idea or Concept|SIMPLE_SEGMENT|8048,8060|false|false|false|C1548597|Marketing basis - Transitional|TRANSITIONAL
Event|Event|SIMPLE_SEGMENT|8061,8067|false|false|false|||ISSUES
Finding|Body Substance|SIMPLE_SEGMENT|8071,8078|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|8071,8078|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|8071,8078|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Finding|SIMPLE_SEGMENT|8083,8086|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|SIMPLE_SEGMENT|8083,8086|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Finding|SIMPLE_SEGMENT|8083,8102|false|false|false|C0020649|Hypotension|low blood pressures
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8087,8092|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|8087,8092|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|8087,8092|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Finding|SIMPLE_SEGMENT|8087,8102|false|false|false|C1272641|Systemic arterial pressure|blood pressures
Event|Event|SIMPLE_SEGMENT|8093,8102|false|false|false|||pressures
Finding|Finding|SIMPLE_SEGMENT|8093,8102|false|false|false|C0460139|Pressure (finding)|pressures
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|8093,8102|false|false|false|C0033095||pressures
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|8120,8128|false|false|false|C0039155|Systole|systolic
Event|Event|SIMPLE_SEGMENT|8138,8145|false|false|false|||benefit
Finding|Finding|SIMPLE_SEGMENT|8151,8156|false|false|false|C0587267;C3810854|Close;Closed|close
Finding|Functional Concept|SIMPLE_SEGMENT|8151,8156|false|false|false|C0587267;C3810854|Close;Closed|close
Event|Activity|SIMPLE_SEGMENT|8157,8167|false|false|false|C1283169||monitoring
Event|Event|SIMPLE_SEGMENT|8157,8167|false|false|false|||monitoring
Procedure|Health Care Activity|SIMPLE_SEGMENT|8157,8167|false|false|false|C0150369|Preventive monitoring|monitoring
Event|Event|SIMPLE_SEGMENT|8172,8181|false|false|false|||titration
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8172,8181|false|false|true|C0162621|Titration Method|titration
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8185,8190|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|8185,8190|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|8185,8190|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Finding|SIMPLE_SEGMENT|8192,8200|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|SIMPLE_SEGMENT|8192,8200|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|8192,8200|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|8192,8200|false|false|false|C0033095||pressure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8201,8212|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8201,8212|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|8201,8212|false|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|8201,8212|false|false|false|C4284232|Medications|medications
Event|Event|SIMPLE_SEGMENT|8219,8229|false|false|false|||outpatient
Finding|Classification|SIMPLE_SEGMENT|8219,8229|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|8219,8229|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|SIMPLE_SEGMENT|8240,8251|false|false|false|||hypokalemic
Event|Event|SIMPLE_SEGMENT|8267,8276|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|8267,8276|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Drug|Organic Chemical|SIMPLE_SEGMENT|8292,8302|false|false|false|C0016860|furosemide|furosemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8292,8302|false|false|false|C0016860|furosemide|furosemide
Event|Event|SIMPLE_SEGMENT|8292,8302|false|false|false|||furosemide
Event|Event|SIMPLE_SEGMENT|8311,8315|false|false|false|||held
Event|Event|SIMPLE_SEGMENT|8325,8332|false|false|false|||recheck
Event|Event|SIMPLE_SEGMENT|8333,8337|false|false|false|||CHEM
Finding|Functional Concept|SIMPLE_SEGMENT|8333,8337|false|false|false|C0079107|chemical aspects|CHEM
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8333,8337|false|false|false|C0201682|Chemical procedure|CHEM
Event|Event|SIMPLE_SEGMENT|8353,8358|false|false|false|||visit
Finding|Social Behavior|SIMPLE_SEGMENT|8353,8358|false|false|false|C0545082|Visit|visit
Event|Event|SIMPLE_SEGMENT|8369,8378|false|false|false|||determine
Event|Event|SIMPLE_SEGMENT|8397,8404|false|false|false|||benefit
Event|Event|SIMPLE_SEGMENT|8413,8428|false|false|false|||supplementation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8413,8428|false|false|false|C0242297|Dietary Supplementation|supplementation
Event|Event|SIMPLE_SEGMENT|8434,8442|false|false|false|||elevated
Event|Event|SIMPLE_SEGMENT|8453,8462|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|8453,8462|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|8453,8462|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|8453,8462|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|8453,8462|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|SIMPLE_SEGMENT|8500,8507|false|false|false|||recheck
Finding|Idea or Concept|SIMPLE_SEGMENT|8515,8521|false|false|false|C1549636|Address type - Office|office
Event|Event|SIMPLE_SEGMENT|8536,8540|false|false|false|||code
Event|Occupational Activity|SIMPLE_SEGMENT|8536,8540|false|false|false|C0009219|Coding|code
Finding|Intellectual Product|SIMPLE_SEGMENT|8536,8540|false|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|code
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8543,8554|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8543,8554|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|8543,8554|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|8543,8554|false|false|false|C4284232|Medications|Medications
Finding|Finding|SIMPLE_SEGMENT|8543,8567|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|SIMPLE_SEGMENT|8558,8567|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|8558,8567|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8586,8596|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|8586,8596|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|8586,8601|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|SIMPLE_SEGMENT|8597,8601|false|false|false|||list
Finding|Intellectual Product|SIMPLE_SEGMENT|8597,8601|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|SIMPLE_SEGMENT|8605,8613|false|false|false|||accurate
Drug|Organic Chemical|SIMPLE_SEGMENT|8618,8626|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8618,8626|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|SIMPLE_SEGMENT|8618,8626|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|SIMPLE_SEGMENT|8618,8626|false|false|false|||complete
Finding|Functional Concept|SIMPLE_SEGMENT|8618,8626|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|SIMPLE_SEGMENT|8618,8626|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Organic Chemical|SIMPLE_SEGMENT|8631,8640|false|false|false|C0030049|oxycodone|Oxycodone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8631,8640|false|false|false|C0030049|oxycodone|Oxycodone
Event|Event|SIMPLE_SEGMENT|8631,8640|false|false|false|||Oxycodone
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8631,8640|false|false|false|C0524222|Oxycodone measurement|Oxycodone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8631,8654|false|false|false|C0717368|acetaminophen / oxycodone|Oxycodone-Acetaminophen
Drug|Organic Chemical|SIMPLE_SEGMENT|8641,8654|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8641,8654|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|SIMPLE_SEGMENT|8641,8654|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8641,8654|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8669,8672|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|SIMPLE_SEGMENT|8669,8672|false|false|false|||TAB
Event|Event|SIMPLE_SEGMENT|8676,8679|false|false|false|||Q8H
Finding|Gene or Genome|SIMPLE_SEGMENT|8680,8683|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8684,8688|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|8684,8688|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|8684,8688|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|8684,8688|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|SIMPLE_SEGMENT|8693,8706|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8693,8706|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Event|Event|SIMPLE_SEGMENT|8693,8706|false|false|false|||Nitroglycerin
Finding|Gene or Genome|SIMPLE_SEGMENT|8726,8729|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8730,8734|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|8730,8734|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|8730,8734|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|8730,8734|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|SIMPLE_SEGMENT|8739,8749|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8739,8749|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Organic Chemical|SIMPLE_SEGMENT|8739,8759|false|false|false|C0724633|metoprolol succinate|Metoprolol Succinate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8739,8759|false|false|false|C0724633|metoprolol succinate|Metoprolol Succinate
Drug|Organic Chemical|SIMPLE_SEGMENT|8750,8759|false|false|false|C0038617;C0220918|Succinates;succinate|Succinate
Event|Event|SIMPLE_SEGMENT|8750,8759|false|false|false|||Succinate
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8783,8790|false|false|false|C1314782|Levemir|Levemir
Drug|Hormone|SIMPLE_SEGMENT|8783,8790|false|false|false|C1314782|Levemir|Levemir
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8783,8790|false|false|false|C1314782|Levemir|Levemir
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8800,8807|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|SIMPLE_SEGMENT|8800,8807|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8800,8807|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|SIMPLE_SEGMENT|8800,8807|false|false|false|||insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|8800,8807|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8800,8807|false|false|false|C0202098|Insulin measurement|insulin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8800,8815|false|false|false|C0537270|insulin detemir|insulin detemir
Drug|Hormone|SIMPLE_SEGMENT|8800,8815|false|false|false|C0537270|insulin detemir|insulin detemir
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8800,8815|false|false|false|C0537270|insulin detemir|insulin detemir
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8808,8815|false|false|false|C0537270|insulin detemir|detemir
Drug|Hormone|SIMPLE_SEGMENT|8808,8815|false|false|false|C0537270|insulin detemir|detemir
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8808,8815|false|false|false|C0537270|insulin detemir|detemir
Event|Event|SIMPLE_SEGMENT|8808,8815|false|false|false|||detemir
Finding|Functional Concept|SIMPLE_SEGMENT|8826,8838|false|false|false|C1522438|Subcutaneous Route of Administration|subcutaneous
Drug|Organic Chemical|SIMPLE_SEGMENT|8859,8868|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8859,8868|false|false|false|C0001927|albuterol|albuterol
Event|Event|SIMPLE_SEGMENT|8859,8868|false|false|false|||albuterol
Drug|Organic Chemical|SIMPLE_SEGMENT|8859,8876|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8859,8876|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|8869,8876|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Inorganic Chemical|SIMPLE_SEGMENT|8869,8876|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8869,8876|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Event|Event|SIMPLE_SEGMENT|8869,8876|false|false|false|||sulfate
Finding|Functional Concept|SIMPLE_SEGMENT|8894,8904|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Finding|Organism Function|SIMPLE_SEGMENT|8894,8904|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Event|Event|SIMPLE_SEGMENT|8905,8910|false|false|false|||q4hrs
Event|Event|SIMPLE_SEGMENT|8911,8919|false|false|false|||wheezing
Finding|Sign or Symptom|SIMPLE_SEGMENT|8911,8919|false|false|false|C0043144|Wheezing|wheezing
Drug|Organic Chemical|SIMPLE_SEGMENT|8924,8931|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8924,8931|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|SIMPLE_SEGMENT|8924,8931|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|SIMPLE_SEGMENT|8924,8933|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|SIMPLE_SEGMENT|8924,8933|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8924,8933|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|SIMPLE_SEGMENT|8924,8933|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8924,8933|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Event|Event|SIMPLE_SEGMENT|8939,8943|false|false|false|||UNIT
Drug|Organic Chemical|SIMPLE_SEGMENT|8957,8966|false|false|false|C0040805|trazodone|TraZODone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8957,8966|false|false|false|C0040805|trazodone|TraZODone
Event|Event|SIMPLE_SEGMENT|8957,8966|false|false|false|||TraZODone
Drug|Organic Chemical|SIMPLE_SEGMENT|8984,8994|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8984,8994|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Organic Chemical|SIMPLE_SEGMENT|8984,9006|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8984,9006|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Event|Event|SIMPLE_SEGMENT|8995,9006|false|false|false|||Mononitrate
Finding|Finding|SIMPLE_SEGMENT|9008,9016|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|SIMPLE_SEGMENT|9008,9016|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|SIMPLE_SEGMENT|9017,9024|false|false|false|||Release
Finding|Functional Concept|SIMPLE_SEGMENT|9017,9024|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|9017,9024|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9017,9024|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|SIMPLE_SEGMENT|9046,9053|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9046,9053|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|SIMPLE_SEGMENT|9075,9087|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9075,9087|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|SIMPLE_SEGMENT|9105,9116|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9105,9116|false|false|false|C0082607|fluticasone|Fluticasone
Event|Event|SIMPLE_SEGMENT|9105,9116|false|false|false|||Fluticasone
Drug|Organic Chemical|SIMPLE_SEGMENT|9105,9127|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9105,9127|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Organic Chemical|SIMPLE_SEGMENT|9117,9127|false|false|false|C0033474;C0392214|Propionates;propionate|Propionate
Event|Event|SIMPLE_SEGMENT|9137,9141|false|false|false|||PUFF
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|9145,9148|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9145,9148|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9145,9148|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|9145,9148|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|9145,9148|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|9154,9166|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9154,9166|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Organic Chemical|SIMPLE_SEGMENT|9186,9196|false|false|false|C0244821|ropinirole|Ropinirole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9186,9196|false|false|false|C0244821|ropinirole|Ropinirole
Event|Event|SIMPLE_SEGMENT|9207,9210|false|false|false|||QPM
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9216,9223|false|false|false|C0528249|Humalog|HumaLOG
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9216,9223|false|false|false|C0528249|Humalog|HumaLOG
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9233,9240|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|SIMPLE_SEGMENT|9233,9240|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9233,9240|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|SIMPLE_SEGMENT|9233,9240|false|false|false|||insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|9233,9240|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9233,9240|false|false|false|C0202098|Insulin measurement|insulin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9233,9247|false|false|false|C0293359|insulin lispro|insulin lispro
Drug|Hormone|SIMPLE_SEGMENT|9233,9247|false|false|false|C0293359|insulin lispro|insulin lispro
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9233,9247|false|false|false|C0293359|insulin lispro|insulin lispro
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9241,9247|false|false|false|C0293359|insulin lispro|lispro
Drug|Hormone|SIMPLE_SEGMENT|9241,9247|false|false|false|C0293359|insulin lispro|lispro
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9241,9247|false|false|false|C0293359|insulin lispro|lispro
Event|Event|SIMPLE_SEGMENT|9241,9247|false|false|false|||lispro
Finding|Functional Concept|SIMPLE_SEGMENT|9253,9265|false|false|false|C1522438|Subcutaneous Route of Administration|SUBCUTANEOUS
Drug|Organic Chemical|SIMPLE_SEGMENT|9284,9293|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9284,9293|false|false|false|C0001927|albuterol|Albuterol
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9301,9304|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9301,9304|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9301,9304|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Finding|Cell Function|SIMPLE_SEGMENT|9301,9304|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Finding|Gene or Genome|SIMPLE_SEGMENT|9301,9304|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9312,9315|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9312,9315|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9312,9315|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Event|Event|SIMPLE_SEGMENT|9312,9315|false|false|false|||NEB
Finding|Cell Function|SIMPLE_SEGMENT|9312,9315|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|SIMPLE_SEGMENT|9312,9315|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|SIMPLE_SEGMENT|9323,9326|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|SIMPLE_SEGMENT|9327,9333|false|false|false|||wheeze
Finding|Sign or Symptom|SIMPLE_SEGMENT|9327,9333|false|false|false|C0043144|Wheezing|wheeze
Drug|Organic Chemical|SIMPLE_SEGMENT|9339,9352|false|false|false|C0025659|methocarbamol|Methocarbamol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9339,9352|false|false|false|C0025659|methocarbamol|Methocarbamol
Event|Event|SIMPLE_SEGMENT|9363,9366|false|false|false|||TID
Finding|Gene or Genome|SIMPLE_SEGMENT|9367,9370|false|false|false|C1422467|CIAO3 gene|PRN
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9371,9377|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Anatomy|Tissue|SIMPLE_SEGMENT|9371,9377|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Finding|Sign or Symptom|SIMPLE_SEGMENT|9371,9382|false|false|false|C0231528|Myalgia|muscle pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9378,9382|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|9378,9382|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|9378,9382|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|9378,9382|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|SIMPLE_SEGMENT|9388,9396|false|false|false|C0126174|losartan|Losartan
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9388,9396|false|false|false|C0126174|losartan|Losartan
Event|Event|SIMPLE_SEGMENT|9388,9396|false|false|false|||Losartan
Drug|Organic Chemical|SIMPLE_SEGMENT|9388,9406|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9388,9406|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9397,9406|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|9397,9406|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Food|SIMPLE_SEGMENT|9397,9406|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|9397,9406|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9397,9406|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Event|Event|SIMPLE_SEGMENT|9397,9406|false|false|false|||Potassium
Finding|Physiologic Function|SIMPLE_SEGMENT|9397,9406|false|false|false|C4553027|Potassium metabolic function|Potassium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9397,9406|false|false|false|C0202194|Potassium measurement|Potassium
Drug|Organic Chemical|SIMPLE_SEGMENT|9427,9437|false|false|false|C0016860|furosemide|Furosemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9427,9437|false|false|false|C0016860|furosemide|Furosemide
Drug|Organic Chemical|SIMPLE_SEGMENT|9458,9468|false|false|false|C0012091|diclofenac|diclofenac
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9458,9468|false|false|false|C0012091|diclofenac|diclofenac
Event|Event|SIMPLE_SEGMENT|9458,9468|false|false|false|||diclofenac
Drug|Organic Chemical|SIMPLE_SEGMENT|9458,9475|false|false|false|C0700583|diclofenac sodium|diclofenac sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9458,9475|false|false|false|C0700583|diclofenac sodium|diclofenac sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9469,9475|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|9469,9475|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9469,9475|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Event|Event|SIMPLE_SEGMENT|9469,9475|false|false|false|||sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|9469,9475|false|false|false|C4553025|Sodium metabolic function|sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9469,9475|false|false|false|C0337443|Sodium measurement|sodium
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9480,9487|false|false|false|C1710439|Topical Dosage Form|topical
Finding|Functional Concept|SIMPLE_SEGMENT|9480,9487|false|false|false|C1522168|Topical Route of Administration|topical
Event|Event|SIMPLE_SEGMENT|9488,9491|false|false|false|||TID
Finding|Gene or Genome|SIMPLE_SEGMENT|9492,9495|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9496,9500|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|9496,9500|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|9496,9500|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|9496,9500|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|9503,9512|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|9503,9512|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|9503,9512|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|9503,9512|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|9503,9512|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|9503,9524|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9513,9524|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9513,9524|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|9513,9524|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|9513,9524|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|SIMPLE_SEGMENT|9529,9538|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9529,9538|false|false|false|C0001927|albuterol|Albuterol
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9546,9549|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9546,9549|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9546,9549|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Finding|Cell Function|SIMPLE_SEGMENT|9546,9549|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Finding|Gene or Genome|SIMPLE_SEGMENT|9546,9549|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9557,9560|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9557,9560|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9557,9560|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Event|Event|SIMPLE_SEGMENT|9557,9560|false|false|false|||NEB
Finding|Cell Function|SIMPLE_SEGMENT|9557,9560|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|SIMPLE_SEGMENT|9557,9560|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|SIMPLE_SEGMENT|9568,9571|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|SIMPLE_SEGMENT|9572,9578|false|false|false|||wheeze
Finding|Sign or Symptom|SIMPLE_SEGMENT|9572,9578|false|false|false|C0043144|Wheezing|wheeze
Drug|Organic Chemical|SIMPLE_SEGMENT|9583,9595|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9583,9595|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|SIMPLE_SEGMENT|9612,9623|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9612,9623|false|false|false|C0082607|fluticasone|Fluticasone
Event|Event|SIMPLE_SEGMENT|9612,9623|false|false|false|||Fluticasone
Drug|Organic Chemical|SIMPLE_SEGMENT|9612,9634|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9612,9634|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Organic Chemical|SIMPLE_SEGMENT|9624,9634|false|false|false|C0033474;C0392214|Propionates;propionate|Propionate
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|9652,9655|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9652,9655|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9652,9655|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|9652,9655|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|9652,9655|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|9660,9673|false|false|false|C0025659|methocarbamol|Methocarbamol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9660,9673|false|false|false|C0025659|methocarbamol|Methocarbamol
Event|Event|SIMPLE_SEGMENT|9684,9687|false|false|false|||TID
Finding|Gene or Genome|SIMPLE_SEGMENT|9688,9691|false|false|false|C1422467|CIAO3 gene|PRN
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9692,9698|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Anatomy|Tissue|SIMPLE_SEGMENT|9692,9698|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Finding|Sign or Symptom|SIMPLE_SEGMENT|9692,9703|false|false|false|C0231528|Myalgia|muscle pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9699,9703|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|9699,9703|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|9699,9703|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|9699,9703|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|SIMPLE_SEGMENT|9708,9721|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9708,9721|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Event|Event|SIMPLE_SEGMENT|9708,9721|false|false|false|||Nitroglycerin
Finding|Gene or Genome|SIMPLE_SEGMENT|9741,9744|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9745,9749|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|9745,9749|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|9745,9749|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|9745,9749|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|SIMPLE_SEGMENT|9754,9766|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9754,9766|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Organic Chemical|SIMPLE_SEGMENT|9785,9795|false|false|false|C0244821|ropinirole|Ropinirole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9785,9795|false|false|false|C0244821|ropinirole|Ropinirole
Event|Event|SIMPLE_SEGMENT|9806,9809|false|false|false|||QPM
Drug|Organic Chemical|SIMPLE_SEGMENT|9814,9823|false|false|false|C0040805|trazodone|TraZODone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9814,9823|false|false|false|C0040805|trazodone|TraZODone
Drug|Organic Chemical|SIMPLE_SEGMENT|9841,9848|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9841,9848|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|SIMPLE_SEGMENT|9841,9848|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|SIMPLE_SEGMENT|9841,9850|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|SIMPLE_SEGMENT|9841,9850|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9841,9850|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|SIMPLE_SEGMENT|9841,9850|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9841,9850|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Event|Event|SIMPLE_SEGMENT|9849,9850|false|false|false|||D
Event|Event|SIMPLE_SEGMENT|9856,9860|false|false|false|||UNIT
Drug|Organic Chemical|SIMPLE_SEGMENT|9875,9884|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9875,9884|false|false|false|C0001927|albuterol|albuterol
Event|Event|SIMPLE_SEGMENT|9875,9884|false|false|false|||albuterol
Drug|Organic Chemical|SIMPLE_SEGMENT|9875,9892|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9875,9892|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|9885,9892|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Inorganic Chemical|SIMPLE_SEGMENT|9885,9892|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9885,9892|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Event|Event|SIMPLE_SEGMENT|9885,9892|false|false|false|||sulfate
Finding|Functional Concept|SIMPLE_SEGMENT|9910,9920|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|INHALATION
Finding|Organism Function|SIMPLE_SEGMENT|9910,9920|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|INHALATION
Event|Event|SIMPLE_SEGMENT|9927,9935|false|false|false|||wheezing
Finding|Sign or Symptom|SIMPLE_SEGMENT|9927,9935|false|false|false|C0043144|Wheezing|wheezing
Drug|Organic Chemical|SIMPLE_SEGMENT|9940,9950|false|false|false|C0012091|diclofenac|diclofenac
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9940,9950|false|false|false|C0012091|diclofenac|diclofenac
Event|Event|SIMPLE_SEGMENT|9940,9950|false|false|false|||diclofenac
Drug|Organic Chemical|SIMPLE_SEGMENT|9940,9957|false|false|false|C0700583|diclofenac sodium|diclofenac sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9940,9957|false|false|false|C0700583|diclofenac sodium|diclofenac sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9951,9957|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|9951,9957|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9951,9957|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Event|Event|SIMPLE_SEGMENT|9951,9957|false|false|false|||sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|9951,9957|false|false|false|C4553025|Sodium metabolic function|sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9951,9957|false|false|false|C0337443|Sodium measurement|sodium
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9962,9969|false|false|false|C1710439|Topical Dosage Form|topical
Finding|Functional Concept|SIMPLE_SEGMENT|9962,9969|false|false|false|C1522168|Topical Route of Administration|topical
Event|Event|SIMPLE_SEGMENT|9970,9973|false|false|false|||TID
Finding|Gene or Genome|SIMPLE_SEGMENT|9974,9977|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9978,9982|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|9978,9982|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|9978,9982|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|9978,9982|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|SIMPLE_SEGMENT|9988,9998|false|false|false|C0016860|furosemide|Furosemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9988,9998|false|false|false|C0016860|furosemide|Furosemide
Drug|Organic Chemical|SIMPLE_SEGMENT|10019,10029|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10019,10029|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Organic Chemical|SIMPLE_SEGMENT|10019,10041|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10019,10041|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Event|Event|SIMPLE_SEGMENT|10030,10041|false|false|false|||Mononitrate
Finding|Finding|SIMPLE_SEGMENT|10043,10051|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|SIMPLE_SEGMENT|10043,10051|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|SIMPLE_SEGMENT|10052,10059|false|false|false|||Release
Finding|Functional Concept|SIMPLE_SEGMENT|10052,10059|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|10052,10059|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10052,10059|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|SIMPLE_SEGMENT|10082,10092|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10082,10092|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Organic Chemical|SIMPLE_SEGMENT|10082,10102|false|false|false|C0724633|metoprolol succinate|Metoprolol Succinate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10082,10102|false|false|false|C0724633|metoprolol succinate|Metoprolol Succinate
Drug|Organic Chemical|SIMPLE_SEGMENT|10093,10102|false|false|false|C0038617;C0220918|Succinates;succinate|Succinate
Event|Event|SIMPLE_SEGMENT|10093,10102|false|false|false|||Succinate
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10127,10134|false|false|false|C0528249|Humalog|HumaLOG
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10127,10134|false|false|false|C0528249|Humalog|HumaLOG
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10144,10151|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|SIMPLE_SEGMENT|10144,10151|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10144,10151|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|SIMPLE_SEGMENT|10144,10151|false|false|false|||insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|10144,10151|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10144,10151|false|false|false|C0202098|Insulin measurement|insulin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10144,10158|false|false|false|C0293359|insulin lispro|insulin lispro
Drug|Hormone|SIMPLE_SEGMENT|10144,10158|false|false|false|C0293359|insulin lispro|insulin lispro
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10144,10158|false|false|false|C0293359|insulin lispro|insulin lispro
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10152,10158|false|false|false|C0293359|insulin lispro|lispro
Drug|Hormone|SIMPLE_SEGMENT|10152,10158|false|false|false|C0293359|insulin lispro|lispro
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10152,10158|false|false|false|C0293359|insulin lispro|lispro
Event|Event|SIMPLE_SEGMENT|10152,10158|false|false|false|||lispro
Finding|Functional Concept|SIMPLE_SEGMENT|10164,10176|false|false|false|C1522438|Subcutaneous Route of Administration|SUBCUTANEOUS
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10195,10202|false|false|false|C1314782|Levemir|Levemir
Drug|Hormone|SIMPLE_SEGMENT|10195,10202|false|false|false|C1314782|Levemir|Levemir
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10195,10202|false|false|false|C1314782|Levemir|Levemir
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10212,10219|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|SIMPLE_SEGMENT|10212,10219|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10212,10219|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|SIMPLE_SEGMENT|10212,10219|false|false|false|||insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|10212,10219|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10212,10219|false|false|false|C0202098|Insulin measurement|insulin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10212,10227|false|false|false|C0537270|insulin detemir|insulin detemir
Drug|Hormone|SIMPLE_SEGMENT|10212,10227|false|false|false|C0537270|insulin detemir|insulin detemir
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10212,10227|false|false|false|C0537270|insulin detemir|insulin detemir
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10220,10227|false|false|false|C0537270|insulin detemir|detemir
Drug|Hormone|SIMPLE_SEGMENT|10220,10227|false|false|false|C0537270|insulin detemir|detemir
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10220,10227|false|false|false|C0537270|insulin detemir|detemir
Event|Event|SIMPLE_SEGMENT|10220,10227|false|false|false|||detemir
Finding|Functional Concept|SIMPLE_SEGMENT|10238,10250|false|false|false|C1522438|Subcutaneous Route of Administration|subcutaneous
Drug|Organic Chemical|SIMPLE_SEGMENT|10272,10280|false|false|false|C0126174|losartan|Losartan
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10272,10280|false|false|false|C0126174|losartan|Losartan
Event|Event|SIMPLE_SEGMENT|10272,10280|false|false|false|||Losartan
Drug|Organic Chemical|SIMPLE_SEGMENT|10272,10290|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10272,10290|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|10281,10290|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|10281,10290|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Food|SIMPLE_SEGMENT|10281,10290|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|10281,10290|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10281,10290|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Event|Event|SIMPLE_SEGMENT|10281,10290|false|false|false|||Potassium
Finding|Physiologic Function|SIMPLE_SEGMENT|10281,10290|false|false|false|C4553027|Potassium metabolic function|Potassium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10281,10290|false|false|false|C0202194|Potassium measurement|Potassium
Drug|Organic Chemical|SIMPLE_SEGMENT|10311,10320|false|false|false|C0030049|oxycodone|Oxycodone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10311,10320|false|false|false|C0030049|oxycodone|Oxycodone
Event|Event|SIMPLE_SEGMENT|10311,10320|false|false|false|||Oxycodone
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10311,10320|false|false|false|C0524222|Oxycodone measurement|Oxycodone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10311,10334|false|false|false|C0717368|acetaminophen / oxycodone|Oxycodone-Acetaminophen
Drug|Organic Chemical|SIMPLE_SEGMENT|10321,10334|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10321,10334|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|SIMPLE_SEGMENT|10321,10334|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10321,10334|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10349,10352|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|SIMPLE_SEGMENT|10349,10352|false|false|false|||TAB
Event|Event|SIMPLE_SEGMENT|10356,10359|false|false|false|||Q8H
Finding|Gene or Genome|SIMPLE_SEGMENT|10360,10363|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10364,10368|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|10364,10368|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|10364,10368|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|10364,10368|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|SIMPLE_SEGMENT|10374,10381|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10374,10381|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|SIMPLE_SEGMENT|10401,10408|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10401,10408|false|false|false|C0004057|aspirin|aspirin
Event|Event|SIMPLE_SEGMENT|10401,10408|false|false|false|||aspirin
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10418,10424|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|SIMPLE_SEGMENT|10428,10436|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|10431,10436|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|10431,10436|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Event|Event|SIMPLE_SEGMENT|10457,10461|false|false|false|||Disp
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10468,10474|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|10475,10482|false|false|false|||Refills
Finding|Idea or Concept|SIMPLE_SEGMENT|10475,10482|false|false|false|C0807726|refill|Refills
Event|Event|SIMPLE_SEGMENT|10488,10497|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|10488,10497|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|10488,10497|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|10488,10497|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|10488,10497|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10488,10509|false|false|false|C4019243||Discharge Disposition
Finding|Finding|SIMPLE_SEGMENT|10488,10509|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10498,10509|false|false|false|C2926604||Disposition
Event|Event|SIMPLE_SEGMENT|10498,10509|false|false|false|||Disposition
Procedure|Health Care Activity|SIMPLE_SEGMENT|10498,10509|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|SIMPLE_SEGMENT|10511,10515|false|false|false|||Home
Finding|Idea or Concept|SIMPLE_SEGMENT|10511,10515|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|SIMPLE_SEGMENT|10511,10515|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|SIMPLE_SEGMENT|10511,10515|false|false|false|C1553498|home health encounter|Home
Event|Event|SIMPLE_SEGMENT|10518,10527|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|10518,10527|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|10518,10527|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|10518,10527|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|10518,10527|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|10518,10537|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10528,10537|false|false|false|C0945731||Diagnosis
Event|Event|SIMPLE_SEGMENT|10528,10537|false|false|false|||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|10528,10537|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|10528,10537|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10528,10537|false|false|false|C0011900|Diagnosis|Diagnosis
Anatomy|Body Location or Region|SIMPLE_SEGMENT|10541,10546|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|SIMPLE_SEGMENT|10541,10546|false|false|false|C0741025|Chest problem|Chest
Anatomy|Body Location or Region|SIMPLE_SEGMENT|10541,10551|false|false|false|C0205076;C4266615|Chest wall structure;Chest>Chest wall|Chest wall
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10541,10551|false|false|false|C0205076;C4266615|Chest wall structure;Chest>Chest wall|Chest wall
Finding|Sign or Symptom|SIMPLE_SEGMENT|10541,10556|false|false|false|C0008035;C0476280|Chest wall pain;Musculoskeletal chest pain|Chest wall pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10552,10556|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|10552,10556|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|10552,10556|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|10552,10556|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|10557,10565|false|false|false|||atypical
Finding|Finding|SIMPLE_SEGMENT|10557,10565|false|false|false|C0741302|atypia morphology|atypical
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10570,10576|false|false|false|C2926611||angina
Event|Event|SIMPLE_SEGMENT|10570,10576|false|false|false|||angina
Finding|Finding|SIMPLE_SEGMENT|10570,10576|false|false|false|C0002962;C2024883|Angina Pectoris|angina
Finding|Sign or Symptom|SIMPLE_SEGMENT|10570,10576|false|false|false|C0002962;C2024883|Angina Pectoris|angina
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10579,10594|false|false|false|C2707260||Musculoskeletal
Finding|Functional Concept|SIMPLE_SEGMENT|10579,10594|false|false|false|C0497254|Musculoskeletal|Musculoskeletal
Finding|Finding|SIMPLE_SEGMENT|10579,10599|false|false|false|C0026858|Musculoskeletal Pain|Musculoskeletal pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10595,10599|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|10595,10599|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|10595,10599|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|10595,10599|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Functional Concept|SIMPLE_SEGMENT|10608,10614|false|false|false|C0302891|Native (qualifier value)|native
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10615,10623|false|false|false|C0018787|Heart|coronary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10615,10630|false|false|false|C0205042|Coronary artery|coronary artery
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10624,10630|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|SIMPLE_SEGMENT|10624,10630|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10635,10641|false|false|false|C0813207|Creation of shunt|bypass
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10635,10647|false|false|false|C0185098|Bypass graft|bypass graft
Anatomy|Tissue|SIMPLE_SEGMENT|10642,10647|false|false|false|C0332835|Transplanted tissue|graft
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10642,10647|false|false|false|C0181074;C1705210|Graft Dosage Form;Graft material|graft
Finding|Intellectual Product|SIMPLE_SEGMENT|10642,10647|false|false|false|C1546653|Graft - Specimen Source Codes|graft
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10642,10647|false|false|false|C1961139;C3683798|Graft Procedures on the Head;Grafting procedure|graft
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10648,10655|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|10648,10655|false|false|false|||disease
Finding|Gene or Genome|SIMPLE_SEGMENT|10658,10662|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|Type
Finding|Intellectual Product|SIMPLE_SEGMENT|10658,10662|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|Type
Finding|Classification|SIMPLE_SEGMENT|10658,10664|false|false|false|C0441730|Type 2|Type 2
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10658,10673|false|false|false|C0011860|Diabetes Mellitus, Non-Insulin-Dependent|Type 2 Diabetes
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10658,10682|false|false|false|C0011860|Diabetes Mellitus, Non-Insulin-Dependent|Type 2 Diabetes mellitus
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10665,10673|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|Diabetes
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10665,10682|false|false|false|C0011849|Diabetes Mellitus|Diabetes mellitus
Event|Event|SIMPLE_SEGMENT|10674,10682|false|false|false|||mellitus
Event|Event|SIMPLE_SEGMENT|10691,10698|false|false|false|||Chronic
Finding|Intellectual Product|SIMPLE_SEGMENT|10691,10698|false|false|false|C1547296|Chronic - Admission Level of Care Code|Chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|10691,10698|false|false|false|C1555457|Provision of recurring care for chronic illness|Chronic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10691,10713|false|false|false|C1561643|Chronic Kidney Diseases|Chronic kidney disease
Finding|Classification|SIMPLE_SEGMENT|10691,10720|false|false|false|C2074731|chronic kidney disease stage|Chronic kidney disease, stage
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10691,10722|false|false|false|C2316787|Chronic kidney disease stage 3|Chronic kidney disease, stage 3
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10699,10705|false|false|false|C0022646;C0227665|Both kidneys;Kidney|kidney
Disorder|Neoplastic Process|SIMPLE_SEGMENT|10699,10705|false|false|false|C0496892;C0496927|Benign neoplasm of kidney;Neoplasm of uncertain or unknown behavior of kidney|kidney
Finding|Sign or Symptom|SIMPLE_SEGMENT|10699,10705|false|false|false|C0812426|Kidney problem|kidney
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10699,10705|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10699,10705|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10699,10713|false|true|false|C0022658|Kidney Diseases|kidney disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10706,10713|false|true|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|10706,10713|false|false|false|||disease
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10715,10720|false|false|false|C1300072|Tumor stage|stage
Finding|Intellectual Product|SIMPLE_SEGMENT|10715,10722|false|false|false|C0441771|Stage level 3|stage 3
Finding|Intellectual Product|SIMPLE_SEGMENT|10725,10730|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|Acute
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10725,10744|false|false|false|C0022660;C2609414|Acute kidney injury;Kidney Failure, Acute|Acute kidney injury
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|10725,10744|false|false|false|C0022660;C2609414|Acute kidney injury;Kidney Failure, Acute|Acute kidney injury
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10731,10737|false|false|false|C0022646;C0227665|Both kidneys;Kidney|kidney
Disorder|Neoplastic Process|SIMPLE_SEGMENT|10731,10737|false|false|false|C0496892;C0496927|Benign neoplasm of kidney;Neoplasm of uncertain or unknown behavior of kidney|kidney
Finding|Sign or Symptom|SIMPLE_SEGMENT|10731,10737|false|false|false|C0812426|Kidney problem|kidney
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10731,10737|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10731,10737|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|10731,10744|false|false|false|C0160420|Injury of kidney|kidney injury
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|10738,10744|false|false|false|C3263722;C3263723|Traumatic AND/OR non-traumatic injury;Traumatic injury|injury
Event|Event|SIMPLE_SEGMENT|10738,10744|false|false|false|||injury
Event|Event|SIMPLE_SEGMENT|10747,10754|false|false|false|||Chronic
Finding|Intellectual Product|SIMPLE_SEGMENT|10747,10754|false|false|false|C1547296|Chronic - Admission Level of Care Code|Chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|10747,10754|false|false|false|C1555457|Provision of recurring care for chronic illness|Chronic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10747,10784|false|false|false|C0024117|Chronic Obstructive Airway Disease|Chronic obstructive pulmonary disease
Finding|Functional Concept|SIMPLE_SEGMENT|10755,10766|false|false|false|C0549186|Obstructed|obstructive
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10755,10784|false|false|false|C0600260|Lung Diseases, Obstructive|obstructive pulmonary disease
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10767,10776|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10767,10776|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|10767,10776|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10767,10784|false|false|false|C0024115|Lung diseases|pulmonary disease
Finding|Finding|SIMPLE_SEGMENT|10767,10784|false|false|false|C0455540|History of - respiratory disease|pulmonary disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10777,10784|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|10777,10784|false|false|false|||disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10787,10799|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|SIMPLE_SEGMENT|10787,10799|false|false|false|||Hypertension
Event|Event|SIMPLE_SEGMENT|10802,10813|false|false|false|||Hypotension
Finding|Finding|SIMPLE_SEGMENT|10802,10813|false|false|false|C0020649|Hypotension|Hypotension
Event|Event|SIMPLE_SEGMENT|10816,10827|false|false|false|||Hypokalemia
Finding|Finding|SIMPLE_SEGMENT|10816,10827|false|false|false|C0020621|Hypokalemia|Hypokalemia
Finding|Intellectual Product|SIMPLE_SEGMENT|10830,10837|false|false|false|C1547296|Chronic - Admission Level of Care Code|Chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|10830,10837|false|false|false|C1555457|Provision of recurring care for chronic illness|Chronic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10830,10851|false|false|false|C0748678|shoulder pain chronic|Chronic shoulder pain
Anatomy|Body Location or Region|SIMPLE_SEGMENT|10838,10846|false|false|false|C0037004;C4299050|Shoulder;Upper extremity>Shoulder|shoulder
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10838,10846|false|false|false|C0221590;C0869975|Examination of shoulder(s);Procedures on Shoulder|shoulder
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10838,10846|false|false|false|C0221590;C0869975|Examination of shoulder(s);Procedures on Shoulder|shoulder
Finding|Sign or Symptom|SIMPLE_SEGMENT|10838,10851|false|false|false|C0037011|Shoulder Pain|shoulder pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10847,10851|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|10847,10851|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|10847,10851|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|10847,10851|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|10855,10864|false|false|false|C0027415|Narcotics|narcotics
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10855,10864|false|false|false|C0027415|Narcotics|narcotics
Event|Event|SIMPLE_SEGMENT|10855,10864|false|false|false|||narcotics
Finding|Functional Concept|SIMPLE_SEGMENT|10867,10878|false|false|false|C0549186|Obstructed|Obstructive
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10867,10890|false|false|false|C0520679|Sleep Apnea, Obstructive|Obstructive sleep apnea
Drug|Organic Chemical|SIMPLE_SEGMENT|10879,10884|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10879,10884|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Finding|Organism Function|SIMPLE_SEGMENT|10879,10884|false|false|false|C0037313|Sleep|sleep
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10879,10890|false|false|false|C0037315|Sleep Apnea Syndromes|sleep apnea
Event|Event|SIMPLE_SEGMENT|10885,10890|false|false|false|||apnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|10885,10890|false|false|false|C0003578|Apnea|apnea
Finding|Pathologic Function|SIMPLE_SEGMENT|10910,10916|false|false|false|C0232483|Reflux|reflux
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10917,10924|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|10917,10924|false|false|false|||disease
Event|Event|SIMPLE_SEGMENT|10927,10936|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|10927,10936|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|10927,10936|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|10927,10936|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|10927,10936|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10937,10946|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10937,10946|false|false|false|C0012634|Disease|Condition
Event|Event|SIMPLE_SEGMENT|10937,10946|false|false|false|||Condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|10937,10946|false|false|false|C1705253|Logical Condition|Condition
Finding|Mental Process|SIMPLE_SEGMENT|10948,10954|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10948,10961|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|SIMPLE_SEGMENT|10948,10961|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10955,10961|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|10955,10961|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|10963,10968|false|false|false|||Clear
Finding|Idea or Concept|SIMPLE_SEGMENT|10963,10968|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|SIMPLE_SEGMENT|10973,10981|false|false|false|||coherent
Finding|Finding|SIMPLE_SEGMENT|10973,10981|false|false|false|C4068804|Coherent|coherent
Event|Event|SIMPLE_SEGMENT|10983,10988|false|false|false|||Level
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10983,11005|false|false|false|C4050479||Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|10983,11005|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|SIMPLE_SEGMENT|10992,11005|false|false|false|||Consciousness
Finding|Finding|SIMPLE_SEGMENT|10992,11005|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|SIMPLE_SEGMENT|10992,11005|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11007,11012|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|11007,11012|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11007,11012|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|SIMPLE_SEGMENT|11007,11012|false|false|false|||Alert
Finding|Finding|SIMPLE_SEGMENT|11007,11012|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|11007,11012|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|11007,11012|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|SIMPLE_SEGMENT|11017,11028|false|false|false|||interactive
Finding|Functional Concept|SIMPLE_SEGMENT|11017,11028|false|false|false|C1704675|Interaction|interactive
Event|Activity|SIMPLE_SEGMENT|11030,11038|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|11030,11038|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|SIMPLE_SEGMENT|11030,11038|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11039,11045|false|false|false|C5889824||Status
Event|Event|SIMPLE_SEGMENT|11039,11045|false|false|false|||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|11039,11045|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|11047,11057|false|false|false|||Ambulatory
Finding|Functional Concept|SIMPLE_SEGMENT|11047,11057|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|SIMPLE_SEGMENT|11047,11057|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|SIMPLE_SEGMENT|11047,11057|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|SIMPLE_SEGMENT|11047,11057|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|SIMPLE_SEGMENT|11060,11071|false|false|false|||Independent
Finding|Finding|SIMPLE_SEGMENT|11060,11071|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|SIMPLE_SEGMENT|11060,11071|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Event|Event|SIMPLE_SEGMENT|11076,11085|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|11076,11085|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|11076,11085|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|11076,11085|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|11076,11085|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11076,11098|false|false|false|C3669312||Discharge Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|11076,11098|false|false|false|C4282220|Discharge instructions|Discharge Instructions
Procedure|Health Care Activity|SIMPLE_SEGMENT|11076,11098|false|false|false|C2266673|hospital discharge instructions (treatment)|Discharge Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11086,11098|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|11086,11098|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|11086,11098|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Finding|Gene or Genome|SIMPLE_SEGMENT|11100,11104|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Event|Event|SIMPLE_SEGMENT|11125,11133|false|false|false|||pleasure
Finding|Intellectual Product|SIMPLE_SEGMENT|11125,11133|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|SIMPLE_SEGMENT|11125,11133|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|SIMPLE_SEGMENT|11156,11160|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|11156,11160|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|11156,11160|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|11156,11160|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Event|Event|SIMPLE_SEGMENT|11184,11192|false|false|false|||admitted
Finding|Finding|SIMPLE_SEGMENT|11198,11204|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|SIMPLE_SEGMENT|11198,11204|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Anatomy|Body Location or Region|SIMPLE_SEGMENT|11205,11210|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|11205,11210|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11205,11215|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|11205,11215|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11211,11215|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|11211,11215|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|11211,11215|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|11211,11215|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11233,11239|false|false|false|C1718621|W stress|stress
Drug|Organic Chemical|SIMPLE_SEGMENT|11233,11239|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11233,11239|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Event|Event|SIMPLE_SEGMENT|11233,11239|false|false|false|||stress
Finding|Finding|SIMPLE_SEGMENT|11233,11239|false|false|false|C0038435|Stress|stress
Anatomy|Body Location or Region|SIMPLE_SEGMENT|11241,11245|false|false|false|C4318744|Test - temporal region|test
Event|Event|SIMPLE_SEGMENT|11241,11245|false|false|false|||test
Finding|Functional Concept|SIMPLE_SEGMENT|11241,11245|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Finding|Intellectual Product|SIMPLE_SEGMENT|11241,11245|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|11241,11245|false|false|false|C0456984|Test Result|test
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|11241,11245|false|false|false|C0022885|Laboratory Procedures|test
Event|Event|SIMPLE_SEGMENT|11251,11257|false|false|false|||showed
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11262,11266|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|11262,11266|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|11262,11266|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|11262,11266|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|11270,11278|false|false|false|||unlikely
Finding|Finding|SIMPLE_SEGMENT|11270,11278|false|false|false|C0750558|Unlikely|unlikely
Event|Event|SIMPLE_SEGMENT|11290,11298|false|false|false|||blockage
Finding|Finding|SIMPLE_SEGMENT|11290,11298|false|false|false|C1706968;C1879887;C2237319|Blockage (obstruction - finding);Partial Blockage within Medical Device|blockage
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11307,11315|false|false|false|C0003842;C0226004|Arterial system;Arteries|arteries
Anatomy|Body System|SIMPLE_SEGMENT|11307,11315|false|false|false|C0003842;C0226004|Arterial system;Arteries|arteries
Procedure|Health Care Activity|SIMPLE_SEGMENT|11307,11315|false|false|false|C0397581|Procedure on artery|arteries
Event|Event|SIMPLE_SEGMENT|11321,11325|false|false|false|||feed
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11331,11336|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|11331,11336|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Event|Event|SIMPLE_SEGMENT|11331,11336|false|false|false|||heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|11331,11336|false|false|false|C0795691|HEART PROBLEM|heart
Finding|Gene or Genome|SIMPLE_SEGMENT|11343,11346|true|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|lab
Finding|Intellectual Product|SIMPLE_SEGMENT|11343,11346|true|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|lab
Event|Event|SIMPLE_SEGMENT|11347,11351|true|false|false|||work
Event|Occupational Activity|SIMPLE_SEGMENT|11347,11351|true|false|false|C0043227|Work|work
Event|Event|SIMPLE_SEGMENT|11366,11373|true|false|false|||suggest
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|11374,11380|true|false|false|C3263722;C3263723|Traumatic AND/OR non-traumatic injury;Traumatic injury|injury
Event|Event|SIMPLE_SEGMENT|11374,11380|true|false|false|||injury
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11388,11393|true|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|11388,11393|true|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Event|Event|SIMPLE_SEGMENT|11388,11393|true|false|false|||heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|11388,11393|true|false|false|C0795691|HEART PROBLEM|heart
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11400,11404|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|11400,11404|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|11400,11404|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|11400,11404|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Idea or Concept|SIMPLE_SEGMENT|11429,11440|false|false|false|C0750501|most likely|most likely
Finding|Finding|SIMPLE_SEGMENT|11434,11440|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|11434,11440|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11441,11456|false|false|false|C2707260||musculoskeletal
Event|Event|SIMPLE_SEGMENT|11441,11456|false|false|false|||musculoskeletal
Finding|Functional Concept|SIMPLE_SEGMENT|11441,11456|false|false|false|C0497254|Musculoskeletal|musculoskeletal
Event|Event|SIMPLE_SEGMENT|11479,11486|false|false|false|||improve
Finding|Conceptual Entity|SIMPLE_SEGMENT|11492,11502|false|false|false|C1521721|Supportive assistance|supportive
Event|Event|SIMPLE_SEGMENT|11503,11511|false|false|false|||measures
Finding|Functional Concept|SIMPLE_SEGMENT|11503,11511|false|false|false|C1879489|Measures (attribute)|measures
Drug|Organic Chemical|SIMPLE_SEGMENT|11521,11528|false|false|false|C0699142|Tylenol|Tylenol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11521,11528|false|false|false|C0699142|Tylenol|Tylenol
Finding|Idea or Concept|SIMPLE_SEGMENT|11550,11553|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|11550,11553|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Finding|SIMPLE_SEGMENT|11559,11563|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|11559,11563|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|11559,11563|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|SIMPLE_SEGMENT|11583,11593|false|false|false|||prescribed
Finding|Finding|SIMPLE_SEGMENT|11594,11598|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|SIMPLE_SEGMENT|11594,11598|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|SIMPLE_SEGMENT|11594,11598|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Drug|Organic Chemical|SIMPLE_SEGMENT|11604,11611|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11604,11611|false|false|false|C0004057|aspirin|aspirin
Event|Event|SIMPLE_SEGMENT|11604,11611|false|false|false|||aspirin
Event|Event|SIMPLE_SEGMENT|11667,11678|false|false|false|||improvement
Finding|Conceptual Entity|SIMPLE_SEGMENT|11667,11678|false|false|false|C2986411|Improvement|improvement
Finding|Functional Concept|SIMPLE_SEGMENT|11687,11695|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|11687,11695|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|SIMPLE_SEGMENT|11696,11704|false|false|false|||continue
Finding|Intellectual Product|SIMPLE_SEGMENT|11717,11721|false|false|false|C1561540|Transaction counts and value totals - week|week
Event|Event|SIMPLE_SEGMENT|11733,11741|false|false|false|||symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|11733,11741|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|11733,11741|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|SIMPLE_SEGMENT|11742,11748|false|false|false|||worsen
Event|Event|SIMPLE_SEGMENT|11762,11771|true|false|false|||shortness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11762,11781|true|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|SIMPLE_SEGMENT|11762,11781|true|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|SIMPLE_SEGMENT|11775,11781|true|false|false|C0225386|Breath|breath
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11807,11814|true|false|false|C3854129||symptom
Event|Event|SIMPLE_SEGMENT|11807,11814|true|false|false|||symptom
Finding|Sign or Symptom|SIMPLE_SEGMENT|11807,11814|true|false|false|C1457887|Symptoms|symptom
Event|Event|SIMPLE_SEGMENT|11823,11826|true|false|false|||let
Finding|Intellectual Product|SIMPLE_SEGMENT|11832,11838|false|false|false|C2348314|Doctor - Title|doctor
Event|Event|SIMPLE_SEGMENT|11844,11849|false|false|false|||right
Finding|Functional Concept|SIMPLE_SEGMENT|11844,11849|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Event|Event|SIMPLE_SEGMENT|11876,11884|false|false|false|||pleasure
Finding|Intellectual Product|SIMPLE_SEGMENT|11876,11884|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|SIMPLE_SEGMENT|11876,11884|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|SIMPLE_SEGMENT|11907,11911|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|11907,11911|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|11907,11911|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|11907,11911|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Anatomy|Body System|SIMPLE_SEGMENT|11949,11959|false|false|false|C0007226|Cardiovascular system|Cardiology
Procedure|Health Care Activity|SIMPLE_SEGMENT|11967,11975|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11976,11988|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|11976,11988|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|11976,11988|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

