 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Procedure|Health Care Activity|SIMPLE_SEGMENT|42,51|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|42,56|false|false|false|C2598112||Admission Date
Finding|Body Substance|SIMPLE_SEGMENT|76,85|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|76,85|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|76,85|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|76,85|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|76,90|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|108,113|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|108,113|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|108,113|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|132,135|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|143,150|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|143,150|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|152,160|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Drug|Indicator, Reagent, or Diagnostic Aid|Allergies|178,181|false|false|false|C0013343|Dyes|Dye
Drug|Biologically Active Substance|Allergies|183,189|false|false|false|C0021968;C0885449|Iodine, Homeopathic preparation;iodine|Iodine
Drug|Element, Ion, or Isotope|Allergies|183,189|false|false|false|C0021968;C0885449|Iodine, Homeopathic preparation;iodine|Iodine
Drug|Pharmacologic Substance|Allergies|183,189|false|false|false|C0021968;C0885449|Iodine, Homeopathic preparation;iodine|Iodine
Event|Activity|Allergies|190,200|false|false|false|C2700400|Contain (action)|Containing
Finding|Functional Concept|Allergies|190,200|false|false|false|C0332256|Containing (qualifier value)|Containing
Drug|Indicator, Reagent, or Diagnostic Aid|Allergies|201,209|false|false|false|C0009924|Contrast Media|Contrast
Drug|Indicator, Reagent, or Diagnostic Aid|Allergies|201,215|false|false|false|C0009924|Contrast Media|Contrast Media
Anatomy|Tissue|Allergies|210,215|false|false|false|C0162867;C1254021|Media layer;Tunica Media|Media
Finding|Intellectual Product|Allergies|210,215|false|false|false|C0009458;C0677540|Communications Media;PAMS Media|Media
Drug|Organic Chemical|Allergies|218,227|false|false|false|C0030049|oxycodone|Oxycodone
Drug|Pharmacologic Substance|Allergies|218,227|false|false|false|C0030049|oxycodone|Oxycodone
Procedure|Laboratory Procedure|Allergies|218,227|false|false|false|C0524222|Oxycodone measurement|Oxycodone
Drug|Organic Chemical|Allergies|231,241|false|false|false|C0055729|cilostazol|cilostazol
Drug|Pharmacologic Substance|Allergies|231,241|false|false|false|C0055729|cilostazol|cilostazol
Drug|Organic Chemical|Allergies|244,255|false|false|false|C1569608|varenicline|Varenicline
Drug|Pharmacologic Substance|Allergies|244,255|false|false|false|C1569608|varenicline|Varenicline
Finding|Functional Concept|Allergies|258,267|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|Chief Complaint|292,299|false|false|false|C0013404;C2024878|Dyspnea|Dyspnea
Finding|Sign or Symptom|Chief Complaint|292,299|false|false|false|C0013404;C2024878|Dyspnea|Dyspnea
Anatomy|Body Part, Organ, or Organ Component|Chief Complaint|301,307|false|false|false|C0018792|Heart Atrium|Atrial
Attribute|Clinical Attribute|Chief Complaint|301,320|false|false|false|C2926591||Atrial Fibrillation
Disorder|Disease or Syndrome|Chief Complaint|301,320|false|false|false|C0004238|Atrial Fibrillation|Atrial Fibrillation
Lab|Laboratory or Test Result|Chief Complaint|301,320|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Atrial Fibrillation
Disorder|Disease or Syndrome|Chief Complaint|308,320|false|false|false|C0232197|Fibrillation|Fibrillation
Finding|Classification|Chief Complaint|323,328|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|329,337|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|329,337|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|341,359|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|350,359|false|false|false|C0945766||Procedure
Event|Occupational Activity|Chief Complaint|350,359|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|350,359|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|350,359|false|false|false|C0184661|Interventional procedure|Procedure
Disorder|Disease or Syndrome|History of Present Illness|416,420|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|History of Present Illness|416,420|false|false|false|C1647218|COPD pharmacologic substance|COPD
Finding|Gene or Genome|History of Present Illness|416,420|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|History of Present Illness|437,440|false|false|false|C0020538|Hypertensive disease|htn
Disorder|Disease or Syndrome|History of Present Illness|442,446|false|false|false|C0004238|Atrial Fibrillation|afib
Lab|Laboratory or Test Result|History of Present Illness|442,446|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|afib
Finding|Finding|History of Present Illness|466,473|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|History of Present Illness|466,473|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Disorder|Disease or Syndrome|History of Present Illness|503,507|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|History of Present Illness|503,507|false|false|false|C1647218|COPD pharmacologic substance|COPD
Finding|Gene or Genome|History of Present Illness|503,507|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|History of Present Illness|526,530|false|false|false|C0004238|Atrial Fibrillation|Afib
Lab|Laboratory or Test Result|History of Present Illness|526,530|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Afib
Finding|Finding|History of Present Illness|536,539|false|false|false|C1417822;C3540498;C4050414|NR1D2 gene;NR1D2 wt Allele;Rapid Virologic Response|RVR
Finding|Gene or Genome|History of Present Illness|536,539|false|false|false|C1417822;C3540498;C4050414|NR1D2 gene;NR1D2 wt Allele;Rapid Virologic Response|RVR
Finding|Body Substance|History of Present Illness|548,555|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|548,555|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|548,555|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Disorder|Disease or Syndrome|History of Present Illness|604,608|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|History of Present Illness|604,608|false|false|false|C1647218|COPD pharmacologic substance|COPD
Finding|Gene or Genome|History of Present Illness|604,608|false|false|false|C1412502|ARCN1 gene|COPD
Finding|Finding|History of Present Illness|609,614|false|false|false|C1517205;C3540542|Exacerbation of cGVHD;Flare|flare
Finding|Sign or Symptom|History of Present Illness|609,614|false|false|false|C1517205;C3540542|Exacerbation of cGVHD;Flare|flare
Drug|Hormone|History of Present Illness|642,652|false|false|false|C0032952|prednisone|prednisone
Drug|Organic Chemical|History of Present Illness|642,652|false|false|false|C0032952|prednisone|prednisone
Drug|Pharmacologic Substance|History of Present Illness|642,652|false|false|false|C0032952|prednisone|prednisone
Procedure|Health Care Activity|History of Present Illness|653,658|false|false|false|C0441640||taper
Drug|Antibiotic|History of Present Illness|684,696|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Clinical Drug|History of Present Illness|684,696|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Organic Chemical|History of Present Illness|684,696|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Finding|Finding|History of Present Illness|726,730|false|false|false|C5575035|Well (answer to question)|well
Finding|Intellectual Product|History of Present Illness|732,736|false|false|false|C1720594|Then - dosing instruction fragment|then
Finding|Finding|History of Present Illness|747,754|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|History of Present Illness|747,754|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Finding|History of Present Illness|747,762|false|false|false|C0743330|Rest Dyspnea|dyspnea at rest
Finding|Functional Concept|History of Present Illness|755,762|false|false|false|C0443144|At rest (qualifier value)|at rest
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|758,762|false|false|false|C1742913|REST protein, human|rest
Drug|Biologically Active Substance|History of Present Illness|758,762|false|false|false|C1742913|REST protein, human|rest
Finding|Daily or Recreational Activity|History of Present Illness|758,762|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Gene or Genome|History of Present Illness|758,762|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Molecular Function|History of Present Illness|758,762|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Organism Function|History of Present Illness|779,787|false|false|false|C0015264|Exertion|exertion
Finding|Sign or Symptom|History of Present Illness|816,819|false|false|false|C0013404|Dyspnea|SOB
Finding|Functional Concept|History of Present Illness|841,849|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|History of Present Illness|841,849|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Idea or Concept|History of Present Illness|856,866|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|History of Present Illness|856,871|false|false|false|C0332290|Consistent with|consistent with
Disorder|Disease or Syndrome|History of Present Illness|876,880|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|History of Present Illness|876,880|false|false|false|C1647218|COPD pharmacologic substance|COPD
Finding|Gene or Genome|History of Present Illness|876,880|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|History of Present Illness|894,897|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|894,897|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|History of Present Illness|894,897|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|894,897|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|History of Present Illness|894,897|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|History of Present Illness|894,897|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|History of Present Illness|894,897|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|History of Present Illness|894,897|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Finding|Gene or Genome|History of Present Illness|894,897|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|History of Present Illness|894,897|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Disorder|Disease or Syndrome|History of Present Illness|948,952|false|false|false|C0004238|Atrial Fibrillation|Afib
Lab|Laboratory or Test Result|History of Present Illness|948,952|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Afib
Finding|Finding|History of Present Illness|956,959|false|false|false|C1417822;C3540498;C4050414|NR1D2 gene;NR1D2 wt Allele;Rapid Virologic Response|RVR
Finding|Gene or Genome|History of Present Illness|956,959|false|false|false|C1417822;C3540498;C4050414|NR1D2 gene;NR1D2 wt Allele;Rapid Virologic Response|RVR
Event|Activity|History of Present Illness|961,965|false|false|false|C0871208|Rating (action)|rate
Finding|Idea or Concept|History of Present Illness|961,965|false|false|false|C1549480|Amount type - Rate|rate
Finding|Conceptual Entity|History of Present Illness|993,1000|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|993,1000|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|History of Present Illness|993,1000|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|993,1003|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|History of Present Illness|1004,1008|false|false|false|C0004238|Atrial Fibrillation|afib
Lab|Laboratory or Test Result|History of Present Illness|1004,1008|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|afib
Finding|Sign or Symptom|History of Present Illness|1052,1055|false|false|false|C0013404|Dyspnea|SOB
Disorder|Disease or Syndrome|History of Present Illness|1060,1064|false|false|false|C0004238|Atrial Fibrillation|afib
Lab|Laboratory or Test Result|History of Present Illness|1060,1064|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|afib
Finding|Finding|History of Present Illness|1070,1073|false|false|false|C1417822;C3540498;C4050414|NR1D2 gene;NR1D2 wt Allele;Rapid Virologic Response|RVR
Finding|Gene or Genome|History of Present Illness|1070,1073|false|false|false|C1417822;C3540498;C4050414|NR1D2 gene;NR1D2 wt Allele;Rapid Virologic Response|RVR
Finding|Individual Behavior|History of Present Illness|1096,1105|false|false|false|C1321605|Compliance behavior|compliant
Drug|Biomedical or Dental Material|History of Present Illness|1111,1115|false|false|false|C1300458|Nebulizer solution|nebs
Drug|Organic Chemical|History of Present Illness|1120,1127|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Drug|Pharmacologic Substance|History of Present Illness|1120,1127|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Finding|Intellectual Product|History of Present Illness|1136,1143|false|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1136,1143|false|false|false|C0040808|Treatment Protocols|regimen
Attribute|Clinical Attribute|History of Present Illness|1165,1170|false|false|false|C1717255||edema
Finding|Pathologic Function|History of Present Illness|1165,1170|false|false|false|C0013604|Edema|edema
Finding|Finding|History of Present Illness|1172,1181|false|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Finding|Sign or Symptom|History of Present Illness|1172,1181|false|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Finding|Daily or Recreational Activity|History of Present Illness|1201,1207|true|false|false|C0040802|travel|travel
Procedure|Health Care Activity|History of Present Illness|1201,1207|true|false|false|C1555670|travel charge|travel
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1209,1218|false|false|false|C0543467|Operative Surgical Procedures|surgeries
Anatomy|Body Location or Region|History of Present Illness|1243,1248|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|1243,1248|false|false|false|C0741025|Chest problem|chest
Finding|Sign or Symptom|History of Present Illness|1243,1258|false|false|false|C0232292|Chest tightness|chest tightness
Disorder|Disease or Syndrome|History of Present Illness|1287,1291|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|History of Present Illness|1287,1291|false|false|false|C1647218|COPD pharmacologic substance|COPD
Finding|Gene or Genome|History of Present Illness|1287,1291|false|false|false|C1412502|ARCN1 gene|COPD
Finding|Sign or Symptom|History of Present Illness|1307,1313|true|false|false|C0015967|Fever|fevers
Finding|Sign or Symptom|History of Present Illness|1317,1325|true|false|false|C0010200|Coughing|coughing
Event|Occupational Activity|History of Present Illness|1329,1339|false|false|false|C0033268|production|production
Finding|Intellectual Product|History of Present Illness|1329,1339|false|false|false|C1548180|Production Processing ID|production
Finding|Body Substance|History of Present Illness|1343,1349|false|false|false|C0038056;C1546789;C1576419|Specimen Type - Sputum;Sputum|sputum
Finding|Intellectual Product|History of Present Illness|1343,1349|false|false|false|C0038056;C1546789;C1576419|Specimen Type - Sputum;Sputum|sputum
Disorder|Disease or Syndrome|Past Medical History|1391,1397|false|false|false|C0004096|Asthma|ASTHMA
Disorder|Disease or Syndrome|Past Medical History|1398,1402|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Past Medical History|1398,1402|false|false|false|C1647218|COPD pharmacologic substance|COPD
Finding|Gene or Genome|Past Medical History|1398,1402|false|false|false|C1412502|ARCN1 gene|COPD
Finding|Finding|Past Medical History|1406,1414|false|false|false|C0741302|atypia morphology|ATYPICAL
Finding|Sign or Symptom|Past Medical History|1406,1425|false|false|false|C0262384|Atypical chest pain|ATYPICAL CHEST PAIN
Anatomy|Body Location or Region|Past Medical History|1415,1420|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|CHEST
Finding|Finding|Past Medical History|1415,1420|false|false|false|C0741025|Chest problem|CHEST
Attribute|Clinical Attribute|Past Medical History|1415,1425|false|false|false|C2926613||CHEST PAIN
Finding|Sign or Symptom|Past Medical History|1415,1425|false|false|false|C0008031|Chest Pain|CHEST PAIN
Attribute|Clinical Attribute|Past Medical History|1421,1425|false|true|false|C2598155||PAIN
Finding|Functional Concept|Past Medical History|1421,1425|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|PAIN
Finding|Sign or Symptom|Past Medical History|1421,1425|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|PAIN
Anatomy|Body Location or Region|Past Medical History|1429,1437|false|false|false|C0027530|Neck|CERVICAL
Disorder|Disease or Syndrome|Past Medical History|1429,1449|false|false|false|C0263884|Cervical radiculitis|CERVICAL RADICULITIS
Disorder|Disease or Syndrome|Past Medical History|1438,1449|false|false|false|C0034544|Radiculitis|RADICULITIS
Anatomy|Body Location or Region|Past Medical History|1453,1461|false|false|false|C0027530|Neck|CERVICAL
Disorder|Disease or Syndrome|Past Medical History|1453,1473|false|false|false|C0158241;C1384641|Cervical spondylosis;Cervical spondylosis without myelopathy|CERVICAL SPONDYLOSIS
Disorder|Disease or Syndrome|Past Medical History|1462,1473|false|false|false|C0038019|Spondylosis|SPONDYLOSIS
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1477,1485|false|false|false|C0018787|Heart|CORONARY
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1477,1492|false|false|false|C0205042|Coronary artery|CORONARY ARTERY
Disorder|Disease or Syndrome|Past Medical History|1477,1500|false|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|CORONARY ARTERY DISEASE
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1486,1492|false|false|false|C0003842;C0226004|Arterial system;Arteries|ARTERY
Anatomy|Body System|Past Medical History|1486,1492|false|false|false|C0003842;C0226004|Arterial system;Arteries|ARTERY
Disorder|Disease or Syndrome|Past Medical History|1486,1500|false|false|false|C0852949|Arteriopathic disease|ARTERY DISEASE
Disorder|Disease or Syndrome|Past Medical History|1493,1500|false|false|false|C0012634|Disease|DISEASE
Finding|Sign or Symptom|Past Medical History|1504,1512|false|false|false|C0018681|Headache|HEADACHE
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1516,1519|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|HIP
Drug|Amino Acid, Peptide, or Protein|Past Medical History|1516,1519|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|HIP
Drug|Biologically Active Substance|Past Medical History|1516,1519|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|HIP
Drug|Pharmacologic Substance|Past Medical History|1516,1519|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|HIP
Finding|Gene or Genome|Past Medical History|1516,1519|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|HIP
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1516,1519|false|false|false|C1292890|Procedure on hip|HIP
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1516,1531|false|false|false|C0392806|Prosthetic arthroplasty of hip (procedure)|HIP REPLACEMENT
Finding|Functional Concept|Past Medical History|1520,1531|false|false|false|C0559956|Replacement|REPLACEMENT
Procedure|Health Care Activity|Past Medical History|1520,1531|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|REPLACEMENT
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1520,1531|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|REPLACEMENT
Disorder|Disease or Syndrome|Past Medical History|1535,1549|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|HYPERLIPIDEMIA
Finding|Finding|Past Medical History|1535,1549|false|false|false|C0428465|Serum lipids high (finding)|HYPERLIPIDEMIA
Disorder|Disease or Syndrome|Past Medical History|1553,1565|false|false|false|C0020538|Hypertensive disease|HYPERTENSION
Disorder|Disease or Syndrome|Past Medical History|1569,1583|false|false|false|C0029408|Degenerative polyarthritis|OSTEOARTHRITIS
Disorder|Disease or Syndrome|Past Medical History|1587,1593|false|false|false|C0019340;C0854331|Herpes simplex dermatitis|HERPES
Disorder|Disease or Syndrome|Past Medical History|1587,1600|false|false|false|C0019360;C0042338|Herpes zoster (disorder);herpesvirus 3, human|HERPES ZOSTER
Disorder|Virus|Past Medical History|1587,1600|false|false|false|C0019360;C0042338|Herpes zoster (disorder);herpesvirus 3, human|HERPES ZOSTER
Disorder|Disease or Syndrome|Past Medical History|1594,1600|false|false|false|C0019360|Herpes zoster (disorder)|ZOSTER
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1604,1610|false|false|false|C0018792|Heart Atrium|ATRIAL
Attribute|Clinical Attribute|Past Medical History|1604,1623|false|false|false|C2926591||ATRIAL FIBRILLATION
Disorder|Disease or Syndrome|Past Medical History|1604,1623|false|false|false|C0004238|Atrial Fibrillation|ATRIAL FIBRILLATION
Lab|Laboratory or Test Result|Past Medical History|1604,1623|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|ATRIAL FIBRILLATION
Disorder|Disease or Syndrome|Past Medical History|1611,1623|false|false|false|C0232197|Fibrillation|FIBRILLATION
Disorder|Mental or Behavioral Dysfunction|Past Medical History|1627,1634|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|ANXIETY
Finding|Sign or Symptom|Past Medical History|1627,1634|false|false|false|C0860603|Anxiety symptoms|ANXIETY
Finding|Intellectual Product|Past Medical History|1638,1654|false|false|false|C1314977|Gastrointestinal attachment|GASTROINTESTINAL
Finding|Pathologic Function|Past Medical History|1638,1663|false|false|false|C0017181|Gastrointestinal Hemorrhage|GASTROINTESTINAL BLEEDING
Finding|Pathologic Function|Past Medical History|1655,1663|false|false|false|C0019080|Hemorrhage|BLEEDING
Disorder|Disease or Syndrome|Past Medical History|1667,1681|false|false|false|C0029408|Degenerative polyarthritis|OSTEOARTHRITIS
Finding|Functional Concept|Past Medical History|1685,1700|false|false|false|C0333482|atherosclerotic|ATHEROSCLEROTIC
Disorder|Disease or Syndrome|Past Medical History|1685,1723|false|false|false|C0004153|Atherosclerosis|ATHEROSCLEROTIC CARDIOVASCULAR DISEASE
Anatomy|Body System|Past Medical History|1701,1715|false|false|false|C0007226;C3887460|Cardiovascular;Cardiovascular system|CARDIOVASCULAR
Disorder|Disease or Syndrome|Past Medical History|1701,1723|false|false|false|C0007222|Cardiovascular Diseases|CARDIOVASCULAR DISEASE
Disorder|Disease or Syndrome|Past Medical History|1716,1723|false|false|false|C0012634|Disease|DISEASE
Disorder|Disease or Syndrome|Past Medical History|1727,1754|false|false|false|C0085096|Peripheral Vascular Diseases|PERIPHERAL VASCULAR DISEASE
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1738,1746|false|false|false|C0005847|Blood Vessel|VASCULAR
Disorder|Disease or Syndrome|Past Medical History|1738,1754|false|false|false|C0042373|Vascular Diseases|VASCULAR DISEASE
Disorder|Disease or Syndrome|Past Medical History|1747,1754|false|false|false|C0012634|Disease|DISEASE
Finding|Idea or Concept|Family Medical History|1793,1799|false|false|false|C1546508|Relationship - Mother|Mother
Disorder|Disease or Syndrome|Family Medical History|1806,1809|false|false|false|C0020538|Hypertensive disease|HTN
Finding|Conceptual Entity|Family Medical History|1812,1818|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Idea or Concept|Family Medical History|1812,1818|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Conceptual Entity|Family Medical History|1829,1836|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Finding|Idea or Concept|Family Medical History|1829,1836|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Finding|Conceptual Entity|Family Medical History|1844,1851|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Finding|Idea or Concept|Family Medical History|1844,1851|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Finding|Finding|Family Medical History|1860,1868|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|Family Medical History|1860,1868|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|Family Medical History|1860,1868|false|false|false|C0031809|Physical Examination|Physical
Procedure|Health Care Activity|Family Medical History|1874,1883|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Finding|Finding|Family Medical History|1884,1892|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|Family Medical History|1884,1892|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|Family Medical History|1884,1892|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|Family Medical History|1884,1897|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAM
Procedure|Health Care Activity|Family Medical History|1884,1897|false|false|false|C0031809|Physical Examination|PHYSICAL EXAM
Finding|Functional Concept|Family Medical History|1893,1897|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|Family Medical History|1893,1897|false|false|false|C0582103|Medical Examination|EXAM
Finding|Classification|Family Medical History|1932,1939|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|Family Medical History|1932,1939|false|false|false|C3812897|General medical service|GENERAL
Finding|Finding|Family Medical History|1941,1945|false|false|false|C5575035|Well (answer to question)|Well
Disorder|Disease or Syndrome|Family Medical History|1957,1960|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|Family Medical History|1957,1960|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|Family Medical History|1957,1960|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Family Medical History|1957,1960|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|Family Medical History|1957,1960|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Finding|Finding|Family Medical History|1957,1960|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Disorder|Congenital Abnormality|Family Medical History|1965,1981|true|false|false|C0158784|Accessory skeletal muscle|accessory muscle
Finding|Finding|Family Medical History|1965,1985|true|false|false|C1821466|Use of accessory muscles|accessory muscle use
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1975,1981|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Anatomy|Tissue|Family Medical History|1975,1981|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Finding|Functional Concept|Family Medical History|1982,1985|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|Family Medical History|1982,1985|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Anatomy|Body Location or Region|Family Medical History|1990,1995|false|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2003,2009|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|Family Medical History|2003,2009|false|false|false|C0036412|Scleral Diseases|Sclera
Procedure|Health Care Activity|Family Medical History|2003,2009|false|false|false|C2228481|examination of sclera|Sclera
Finding|Finding|Family Medical History|2010,2019|false|false|false|C0205180|Anicteric|anicteric
Finding|Finding|Family Medical History|2021,2026|false|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Anatomy|Body Location or Region|Family Medical History|2037,2041|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|Family Medical History|2037,2041|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|Family Medical History|2037,2041|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Finding|Finding|Family Medical History|2046,2049|true|false|false|C0425687|Jugular venous engorgement|JVD
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2053,2060|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|Family Medical History|2053,2060|false|false|false|C1314974|Cardiac attachment|CARDIAC
Finding|Finding|Family Medical History|2072,2078|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|Family Medical History|2072,2078|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Event|Activity|Family Medical History|2087,2091|false|false|false|C0871208|Rating (action)|rate
Finding|Idea or Concept|Family Medical History|2087,2091|false|false|false|C1549480|Amount type - Rate|rate
Finding|Finding|Family Medical History|2112,2119|false|false|false|C0018808|Heart murmur|murmurs
Finding|Finding|Family Medical History|2120,2124|false|false|false|C0232267|Pericardial friction rub|rubs
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2137,2142|false|false|false|C0024109|Lung|LUNGS
Drug|Inorganic Chemical|Family Medical History|2151,2154|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|Family Medical History|2151,2154|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|Family Medical History|2151,2154|false|false|false|C0001861;C3536832|Air (substance);air|air
Finding|Finding|Family Medical History|2151,2154|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|Family Medical History|2151,2154|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|Family Medical History|2151,2154|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Finding|Family Medical History|2155,2159|false|false|false|C5575035|Well (answer to question)|well
Finding|Functional Concept|Family Medical History|2173,2178|false|false|false|C1883002|Sequence Chromatogram|Trace
Finding|Organism Function|Family Medical History|2179,2190|false|false|false|C0004048|Inspiration (function)|inspiratory
Finding|Sign or Symptom|Family Medical History|2179,2199|false|false|false|C0231874|Inspiratory wheezing|inspiratory wheezing
Finding|Sign or Symptom|Family Medical History|2191,2199|false|false|false|C0043144|Wheezing|wheezing
Finding|Organism Function|Family Medical History|2212,2222|false|false|false|C0231800|Expiration, Respiratory|expiratory
Finding|Sign or Symptom|Family Medical History|2212,2231|false|false|false|C0231875|Expiratory wheezing|expiratory wheezing
Finding|Sign or Symptom|Family Medical History|2223,2231|false|false|false|C0043144|Wheezing|wheezing
Anatomy|Body Location or Region|Family Medical History|2239,2243|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2239,2243|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Family Medical History|2239,2243|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Family Medical History|2239,2243|false|false|false|C0740941|Lung Problem|lung
Finding|Finding|Family Medical History|2256,2264|false|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Finding|Finding|Family Medical History|2265,2272|false|false|false|C0035508|Rhonchi|rhonchi
Anatomy|Body Location or Region|Family Medical History|2277,2284|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|Family Medical History|2277,2284|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Finding|Finding|Family Medical History|2277,2284|false|false|false|C0941288|Abdomen problem|ABDOMEN
Disorder|Disease or Syndrome|Family Medical History|2286,2290|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Finding|Gene or Genome|Family Medical History|2301,2304|true|false|false|C1537594|LRRC4B gene|HSM
Finding|Mental Process|Family Medical History|2308,2318|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|Family Medical History|2308,2318|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2323,2334|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2349,2356|false|false|false|C0015811|Femur|femoral
Finding|Finding|Family Medical History|2357,2363|true|false|false|C0006318|Bruit|bruits
Finding|Body Substance|Family Medical History|2368,2377|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|Family Medical History|2368,2377|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|Family Medical History|2368,2377|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|Family Medical History|2368,2377|false|false|false|C0030685|Patient Discharge|DISCHARGE
Finding|Finding|Family Medical History|2378,2386|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|Family Medical History|2378,2386|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|Family Medical History|2378,2386|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|Family Medical History|2378,2391|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAM
Procedure|Health Care Activity|Family Medical History|2378,2391|false|false|false|C0031809|Physical Examination|PHYSICAL EXAM
Finding|Functional Concept|Family Medical History|2387,2391|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|Family Medical History|2387,2391|false|false|false|C0582103|Medical Examination|EXAM
Finding|Classification|Family Medical History|2420,2427|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|Family Medical History|2420,2427|false|false|false|C3812897|General medical service|GENERAL
Disorder|Disease or Syndrome|Family Medical History|2429,2432|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|Family Medical History|2429,2432|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|Family Medical History|2429,2432|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Family Medical History|2429,2432|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|Family Medical History|2429,2432|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Finding|Finding|Family Medical History|2429,2432|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Location or Region|Family Medical History|2433,2438|false|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2446,2452|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|Family Medical History|2446,2452|false|false|false|C0036412|Scleral Diseases|Sclera
Procedure|Health Care Activity|Family Medical History|2446,2452|false|false|false|C2228481|examination of sclera|Sclera
Finding|Finding|Family Medical History|2453,2462|false|false|false|C0205180|Anicteric|anicteric
Finding|Idea or Concept|Family Medical History|2494,2499|false|false|false|C1550016|Remote control command - Clear|clear
Anatomy|Body Location or Region|Family Medical History|2501,2505|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|Family Medical History|2501,2505|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|Family Medical History|2501,2505|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Finding|Finding|Family Medical History|2510,2513|true|false|false|C0425687|Jugular venous engorgement|JVD
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2516,2523|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|Family Medical History|2516,2523|false|false|false|C1314974|Cardiac attachment|CARDIAC
Finding|Finding|Family Medical History|2548,2555|true|false|false|C0018808|Heart murmur|murmurs
Finding|Finding|Family Medical History|2556,2560|true|false|false|C0232267|Pericardial friction rub|rubs
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2572,2577|false|false|false|C0024109|Lung|LUNGS
Drug|Inorganic Chemical|Family Medical History|2594,2597|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|Family Medical History|2594,2597|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|Family Medical History|2594,2597|false|false|false|C0001861;C3536832|Air (substance);air|air
Finding|Finding|Family Medical History|2594,2597|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|Family Medical History|2594,2597|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|Family Medical History|2594,2597|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Phenomenon|Natural Phenomenon or Process|Family Medical History|2594,2606|false|false|false|C0001868|Air Movements|air movement
Finding|Organism Function|Family Medical History|2598,2606|false|false|false|C0026649|Movement|movement
Finding|Idea or Concept|Family Medical History|2608,2619|false|false|false|C0750502|Significant|significant
Finding|Sign or Symptom|Family Medical History|2620,2628|false|false|false|C0043144|Wheezing|wheezing
Finding|Finding|Family Medical History|2644,2651|false|false|false|C0035508|Rhonchi|rhonchi
Finding|Finding|Family Medical History|2656,2664|true|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Anatomy|Body Location or Region|Family Medical History|2667,2674|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|Family Medical History|2667,2674|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Finding|Finding|Family Medical History|2667,2674|false|false|false|C0941288|Abdomen problem|ABDOMEN
Disorder|Disease or Syndrome|Family Medical History|2676,2680|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Finding|Gene or Genome|Family Medical History|2691,2694|true|false|false|C1537594|LRRC4B gene|HSM
Finding|Mental Process|Family Medical History|2698,2708|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|Family Medical History|2698,2708|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2712,2723|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Procedure|Health Care Activity|Family Medical History|2757,2766|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Lab|Laboratory or Test Result|Family Medical History|2767,2771|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|Family Medical History|2785,2790|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|Family Medical History|2785,2790|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|Family Medical History|2791,2794|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|Family Medical History|2799,2802|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|Family Medical History|2799,2802|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|Family Medical History|2799,2802|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|Family Medical History|2808,2811|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|Family Medical History|2808,2811|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|Family Medical History|2808,2811|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|Family Medical History|2808,2811|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|Family Medical History|2817,2820|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|Family Medical History|2817,2820|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|Family Medical History|2828,2831|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|Family Medical History|2828,2831|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|Family Medical History|2828,2831|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|Family Medical History|2828,2831|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|Family Medical History|2836,2839|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|Family Medical History|2836,2839|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|Family Medical History|2836,2839|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|Family Medical History|2836,2839|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|Family Medical History|2836,2839|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|Family Medical History|2846,2850|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|Family Medical History|2879,2882|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|Family Medical History|2899,2904|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|Family Medical History|2899,2904|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Finding|Body Substance|Family Medical History|2917,2923|false|false|false|C0024202|Lymph|Lymphs
Drug|Antibiotic|Family Medical History|2929,2934|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|Family Medical History|2929,2934|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|Family Medical History|2929,2934|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|Family Medical History|2941,2944|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|Eos
Finding|Gene or Genome|Family Medical History|2941,2944|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|Eos
Disorder|Disease or Syndrome|Family Medical History|3049,3054|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|Family Medical History|3049,3054|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|Family Medical History|3059,3062|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Procedure|Laboratory Procedure|Family Medical History|3059,3062|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|Family Medical History|3084,3089|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|Family Medical History|3084,3089|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|Family Medical History|3084,3097|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|Family Medical History|3084,3097|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|Family Medical History|3084,3097|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|Family Medical History|3090,3097|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|Family Medical History|3090,3097|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|Family Medical History|3090,3097|false|false|false|C0017725|glucose|Glucose
Lab|Laboratory or Test Result|Family Medical History|3090,3097|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|Family Medical History|3090,3097|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|Family Medical History|3143,3147|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|Family Medical History|3143,3147|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|Family Medical History|3143,3147|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|Family Medical History|3172,3177|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|Family Medical History|3172,3177|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|Family Medical History|3172,3185|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|Family Medical History|3178,3185|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|Family Medical History|3178,3185|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|Family Medical History|3178,3185|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|Family Medical History|3178,3185|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|Family Medical History|3178,3185|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Finding|Physiologic Function|Family Medical History|3178,3185|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|Family Medical History|3178,3185|false|false|false|C0201925|Calcium measurement|Calcium
Lab|Laboratory or Test Result|Family Medical History|3217,3221|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|Family Medical History|3235,3240|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|Family Medical History|3235,3240|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|Family Medical History|3267,3272|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|Family Medical History|3267,3272|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|Family Medical History|3273,3278|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|Family Medical History|3273,3278|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|Family Medical History|3273,3278|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|Family Medical History|3273,3278|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Disorder|Disease or Syndrome|Family Medical History|3307,3312|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|Family Medical History|3307,3312|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|Family Medical History|3336,3339|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Drug|Biologically Active Substance|Family Medical History|3336,3339|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Drug|Hormone|Family Medical History|3336,3339|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Drug|Pharmacologic Substance|Family Medical History|3336,3339|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Finding|Gene or Genome|Family Medical History|3336,3339|false|false|false|C1334121;C1336604;C1705002|IL5 gene;TERF1 gene;TERF1 wt Allele|TRF
Disorder|Disease or Syndrome|Family Medical History|3356,3361|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|Family Medical History|3356,3361|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Attribute|Clinical Attribute|Family Medical History|3362,3365|false|false|false|C2708739||TSH
Drug|Amino Acid, Peptide, or Protein|Family Medical History|3362,3365|false|false|false|C0040160|thyrotropin|TSH
Drug|Hormone|Family Medical History|3362,3365|false|false|false|C0040160|thyrotropin|TSH
Drug|Pharmacologic Substance|Family Medical History|3362,3365|false|false|false|C0040160|thyrotropin|TSH
Procedure|Laboratory Procedure|Family Medical History|3362,3365|false|false|false|C0202230|Thyroid stimulating hormone measurement|TSH
Disorder|Disease or Syndrome|Family Medical History|3383,3388|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|Family Medical History|3383,3388|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Finding|Classification|Family Medical History|3393,3396|false|false|false|C0391840;C4521535|Partial pressure of Oxygen;US Military enlisted E5|pO2
Finding|Molecular Function|Family Medical History|3393,3396|false|false|false|C0391840;C4521535|Partial pressure of Oxygen;US Military enlisted E5|pO2
Procedure|Laboratory Procedure|Family Medical History|3393,3396|false|false|false|C1283004|PO2 measurement|pO2
Lab|Laboratory or Test Result|Family Medical History|3401,3405|false|false|false|C0391839|Carbon dioxide, partial pressure|pCO2
Procedure|Laboratory Procedure|Family Medical History|3401,3405|false|false|false|C0201931|Carbon dioxide measurement, partial pressure|pCO2
Anatomy|Body Location or Region|Family Medical History|3431,3435|false|false|false|C2987514|Anatomical base|Base
Drug|Biomedical or Dental Material|Family Medical History|3431,3435|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|Base
Drug|Chemical Viewed Functionally|Family Medical History|3431,3435|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|Base
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Family Medical History|3431,3435|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|Base
Finding|Gene or Genome|Family Medical History|3431,3435|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|Base
Finding|Idea or Concept|Family Medical History|3431,3435|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|Base
Disorder|Disease or Syndrome|Family Medical History|3458,3463|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|Family Medical History|3458,3463|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Finding|Functional Concept|Family Medical History|3468,3472|false|false|false|C0332296|Free of (attribute)|FREE
Finding|Intellectual Product|Family Medical History|3474,3480|false|false|false|C1552596;C3244286|Direct - PostalAddressUse;direct address|DIRECT
Finding|Functional Concept|Family Medical History|3481,3489|false|false|false|C4723631|Dialysis Method of Administration|DIALYSIS
Phenomenon|Natural Phenomenon or Process|Family Medical History|3481,3489|false|false|false|C0011945|Physical Dialysis|DIALYSIS
Procedure|Therapeutic or Preventive Procedure|Family Medical History|3481,3489|false|false|false|C0011946;C4551529|Dialysis procedure;Renal Dialysis|DIALYSIS
Anatomy|Body Location or Region|Family Medical History|3490,3494|false|false|false|C4318744|Test - temporal region|Test
Finding|Functional Concept|Family Medical History|3490,3494|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|Test
Finding|Intellectual Product|Family Medical History|3490,3494|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|Test
Lab|Laboratory or Test Result|Family Medical History|3490,3494|false|false|false|C0456984|Test Result|Test
Procedure|Laboratory Procedure|Family Medical History|3490,3494|false|false|false|C0022885|Laboratory Procedures|Test
Finding|Body Substance|Family Medical History|3498,3507|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|Family Medical History|3498,3507|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|Family Medical History|3498,3507|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|Family Medical History|3498,3507|false|false|false|C0030685|Patient Discharge|DISCHARGE
Lab|Laboratory or Test Result|Family Medical History|3508,3512|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|Family Medical History|3530,3535|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|Family Medical History|3530,3535|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|Family Medical History|3536,3539|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|Family Medical History|3546,3549|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|Family Medical History|3546,3549|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|Family Medical History|3546,3549|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|Family Medical History|3555,3558|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|Family Medical History|3555,3558|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|Family Medical History|3555,3558|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|Family Medical History|3555,3558|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|Family Medical History|3564,3567|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|Family Medical History|3564,3567|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|Family Medical History|3575,3578|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|Family Medical History|3575,3578|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|Family Medical History|3575,3578|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|Family Medical History|3575,3578|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|Family Medical History|3583,3586|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|Family Medical History|3583,3586|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|Family Medical History|3583,3586|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|Family Medical History|3583,3586|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|Family Medical History|3583,3586|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|Family Medical History|3593,3597|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|Family Medical History|3626,3629|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|Family Medical History|3646,3651|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|Family Medical History|3646,3651|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|Family Medical History|3646,3659|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|Family Medical History|3646,3659|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|Family Medical History|3646,3659|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|Family Medical History|3652,3659|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|Family Medical History|3652,3659|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|Family Medical History|3652,3659|false|false|false|C0017725|glucose|Glucose
Lab|Laboratory or Test Result|Family Medical History|3652,3659|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|Family Medical History|3652,3659|false|false|false|C0337438|Glucose measurement|Glucose
Disorder|Disease or Syndrome|Family Medical History|3733,3738|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|Family Medical History|3733,3738|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|Family Medical History|3733,3746|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|Family Medical History|3739,3746|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|Family Medical History|3739,3746|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|Family Medical History|3739,3746|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|Family Medical History|3739,3746|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|Family Medical History|3739,3746|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Finding|Physiologic Function|Family Medical History|3739,3746|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|Family Medical History|3739,3746|false|false|false|C0201925|Calcium measurement|Calcium
Finding|Finding|Family Medical History|3768,3775|false|false|false|C0740845|Imaging problem|IMAGING
Procedure|Diagnostic Procedure|Family Medical History|3768,3775|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|IMAGING
Anatomy|Body Location or Region|Family Medical History|3781,3786|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|Family Medical History|3781,3786|false|false|false|C0741025|Chest problem|Chest
Procedure|Diagnostic Procedure|Family Medical History|3781,3792|false|false|false|C0039985|Plain chest X-ray|Chest X ray
Phenomenon|Natural Phenomenon or Process|Family Medical History|3787,3792|false|false|false|C0043309|Roentgen Rays|X ray
Procedure|Diagnostic Procedure|Family Medical History|3787,3792|false|false|false|C1306645;C1962945|Plain x-ray;Radiographic imaging procedure|X ray
Finding|Gene or Genome|Family Medical History|3789,3792|false|false|false|C1428870;C5444437|RAB35 wt Allele;SH3YL1 gene|ray
Phenomenon|Natural Phenomenon or Process|Family Medical History|3789,3792|false|false|false|C0851346|Radiation|ray
Attribute|Clinical Attribute|Family Medical History|3794,3802|false|false|false|C3172260||Relative
Finding|Idea or Concept|Family Medical History|3794,3802|false|false|false|C1546849|Living Arrangement - Relative|Relative
Finding|Functional Concept|Family Medical History|3803,3811|false|false|false|C0442805|Increase|increase
Finding|Finding|Family Medical History|3815,3822|false|false|false|C0029053;C1265876|Abnormally opaque structure (morphologic abnormality);Decreased translucency|opacity
Finding|Pathologic Function|Family Medical History|3815,3822|false|false|false|C0029053;C1265876|Abnormally opaque structure (morphologic abnormality);Decreased translucency|opacity
Anatomy|Body Location or Region|Family Medical History|3832,3836|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|3832,3836|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Family Medical History|3832,3836|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Family Medical History|3832,3836|false|false|false|C0740941|Lung Problem|lung
Drug|Chemical Viewed Functionally|Family Medical History|3838,3843|false|false|false|C0178499|Base|bases
Disorder|Disease or Syndrome|Family Medical History|3878,3882|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Anatomy|Body Location or Region|Family Medical History|3878,3889|false|false|false|C0225317;C4532079|Neck+Chest>Soft tissue;soft tissue|soft tissue
Anatomy|Tissue|Family Medical History|3878,3889|false|false|false|C0225317;C4532079|Neck+Chest>Soft tissue;soft tissue|soft tissue
Anatomy|Tissue|Family Medical History|3883,3889|false|false|false|C0040300|Body tissue|tissue
Finding|Intellectual Product|Family Medical History|3883,3889|false|true|false|C1547928|Tissue Specimen Code|tissue
Disorder|Disease or Syndrome|Family Medical History|3903,3916|false|false|false|C0521530|Lung consolidation|consolidation
Finding|Finding|Family Medical History|3951,3963|false|false|false|C0750484;C1611825|Confirmation;confirmation - ResponseLevel|confirmation
Finding|Intellectual Product|Family Medical History|3951,3963|false|false|false|C0750484;C1611825|Confirmation;confirmation - ResponseLevel|confirmation
Anatomy|Body Location or Region|Family Medical History|3970,3975|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|Family Medical History|3970,3975|false|false|false|C0741025|Chest problem|Chest
Procedure|Diagnostic Procedure|Family Medical History|3970,3981|false|false|false|C0039985|Plain chest X-ray|Chest X ray
Phenomenon|Natural Phenomenon or Process|Family Medical History|3976,3981|false|false|false|C0043309|Roentgen Rays|X ray
Procedure|Diagnostic Procedure|Family Medical History|3976,3981|false|false|false|C1306645;C1962945|Plain x-ray;Radiographic imaging procedure|X ray
Finding|Gene or Genome|Family Medical History|3978,3981|false|false|false|C1428870;C5444437|RAB35 wt Allele;SH3YL1 gene|ray
Phenomenon|Natural Phenomenon or Process|Family Medical History|3978,3981|false|false|false|C0851346|Radiation|ray
Disorder|Anatomical Abnormality|Family Medical History|3992,4006|false|false|false|C0020449|Hyperdistention|hyperinflation
Disorder|Disease or Syndrome|Family Medical History|4022,4034|false|false|false|C0032326|Pneumothorax|pneumothorax
Finding|Body Substance|Family Medical History|4036,4044|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|Family Medical History|4036,4044|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|Family Medical History|4036,4044|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Disorder|Disease or Syndrome|Family Medical History|4046,4059|false|false|false|C0521530|Lung consolidation|consolidation
Anatomy|Body Space or Junction|Family Medical History|4063,4066|false|false|false|C0262212|Choroidal fissure|CHF
Disorder|Disease or Syndrome|Family Medical History|4063,4066|false|false|false|C0018802|Congestive heart failure|CHF
Finding|Finding|Family Medical History|4078,4086|false|false|false|C0332148|Probable diagnosis|probable
Disorder|Disease or Syndrome|Family Medical History|4088,4098|false|false|false|C0029453|Osteopenia|osteopenia
Finding|Conceptual Entity|Hospital Course|4145,4152|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|4145,4152|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Hospital Course|4145,4152|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|4145,4155|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|Hospital Course|4156,4159|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Hospital Course|4156,4159|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Hospital Course|4156,4159|false|false|false|C1504769|DFFB protein, human|CAD
Finding|Gene or Genome|Hospital Course|4156,4159|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Hospital Course|4156,4159|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Hospital Course|4156,4159|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4156,4159|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Disorder|Disease or Syndrome|Hospital Course|4161,4164|false|false|false|C0085096|Peripheral Vascular Diseases|PVD
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4161,4164|false|false|false|C4521226|Pomalidomide/Bortezomib/Dexamethasone Regimen|PVD
Disorder|Disease or Syndrome|Hospital Course|4171,4175|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Hospital Course|4171,4175|false|false|false|C1647218|COPD pharmacologic substance|COPD
Finding|Gene or Genome|Hospital Course|4171,4175|false|false|false|C1412502|ARCN1 gene|COPD
Finding|Conceptual Entity|Hospital Course|4180,4187|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|4180,4187|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Hospital Course|4180,4187|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|4180,4190|false|false|false|C0262926|Medical History|history of
Anatomy|Body Location or Region|Hospital Course|4201,4206|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Hospital Course|4201,4206|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Hospital Course|4201,4211|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|Hospital Course|4201,4211|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Hospital Course|4207,4211|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|4207,4211|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|4207,4211|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Disorder|Disease or Syndrome|Hospital Course|4231,4235|false|false|false|C0004238|Atrial Fibrillation|afib
Lab|Laboratory or Test Result|Hospital Course|4231,4235|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|afib
Finding|Finding|Hospital Course|4242,4245|false|false|false|C1417822;C3540498;C4050414|NR1D2 gene;NR1D2 wt Allele;Rapid Virologic Response|RVR
Finding|Gene or Genome|Hospital Course|4242,4245|false|false|false|C1417822;C3540498;C4050414|NR1D2 gene;NR1D2 wt Allele;Rapid Virologic Response|RVR
Disorder|Disease or Syndrome|Hospital Course|4250,4254|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Hospital Course|4250,4254|false|false|false|C1647218|COPD pharmacologic substance|COPD
Finding|Gene or Genome|Hospital Course|4250,4254|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|Hospital Course|4250,4267|false|false|false|C0740304|COPD exacerbation|COPD exacerbation
Finding|Finding|Hospital Course|4255,4267|false|false|false|C4086268|Exacerbation|exacerbation
Finding|Intellectual Product|Hospital Course|4273,4278|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|ACUTE
Finding|Idea or Concept|Hospital Course|4279,4287|false|false|false|C1546466|Problems - What subject filter|PROBLEMS
Disorder|Disease or Syndrome|Hospital Course|4291,4295|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Hospital Course|4291,4295|false|false|false|C1647218|COPD pharmacologic substance|COPD
Finding|Gene or Genome|Hospital Course|4291,4295|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|Hospital Course|4291,4308|false|false|false|C0740304|COPD exacerbation|COPD exacerbation
Finding|Finding|Hospital Course|4296,4308|false|false|false|C4086268|Exacerbation|exacerbation
Finding|Social Behavior|Hospital Course|4340,4346|false|false|false|C0545082|Visit|visits
Procedure|Health Care Activity|Hospital Course|4340,4346|false|false|false|C1512346|Patient Visit|visits
Disorder|Disease or Syndrome|Hospital Course|4352,4356|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Hospital Course|4352,4356|false|false|false|C1647218|COPD pharmacologic substance|COPD
Finding|Gene or Genome|Hospital Course|4352,4356|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|Hospital Course|4352,4369|false|false|false|C0740304|COPD exacerbation|COPD exacerbation
Finding|Finding|Hospital Course|4357,4369|false|false|false|C4086268|Exacerbation|exacerbation
Drug|Hormone|Hospital Course|4414,4424|false|false|false|C0032952|prednisone|prednisone
Drug|Organic Chemical|Hospital Course|4414,4424|false|false|false|C0032952|prednisone|prednisone
Drug|Pharmacologic Substance|Hospital Course|4414,4424|false|false|false|C0032952|prednisone|prednisone
Disorder|Disease or Syndrome|Hospital Course|4453,4456|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|Hospital Course|4453,4456|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|Hospital Course|4453,4456|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|Hospital Course|4453,4456|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|Hospital Course|4453,4456|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|Hospital Course|4453,4456|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|Hospital Course|4453,4456|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|Hospital Course|4453,4456|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Finding|Gene or Genome|Hospital Course|4453,4456|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|Hospital Course|4453,4456|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Idea or Concept|Hospital Course|4459,4465|false|false|false|C1549636|Address type - Office|office
Finding|Finding|Hospital Course|4482,4489|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|Hospital Course|4482,4489|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Finding|Hospital Course|4503,4510|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|Hospital Course|4503,4510|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4503,4510|false|false|false|C0087111|Therapeutic procedure|therapy
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4540,4545|false|false|false|C0028429||nasal
Drug|Biomedical or Dental Material|Hospital Course|4540,4545|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Organic Chemical|Hospital Course|4540,4545|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Pharmacologic Substance|Hospital Course|4540,4545|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Finding|Finding|Hospital Course|4540,4545|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Functional Concept|Hospital Course|4540,4545|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Sign or Symptom|Hospital Course|4540,4556|false|false|false|C0027424|Nasal congestion (finding)|nasal congestion
Finding|Pathologic Function|Hospital Course|4546,4556|false|false|false|C0700148|Congestion|congestion
Finding|Functional Concept|Hospital Course|4571,4576|false|false|false|C0521026|Viral|viral
Disorder|Disease or Syndrome|Hospital Course|4577,4580|false|false|false|C0041912|Upper Respiratory Infections|URI
Finding|Gene or Genome|Hospital Course|4577,4580|false|false|false|C1421895;C1548524;C3272713|URI1 gene;URI1 wt Allele;Uniform Resource Identifier|URI
Finding|Intellectual Product|Hospital Course|4577,4580|false|false|false|C1421895;C1548524;C3272713|URI1 gene;URI1 wt Allele;Uniform Resource Identifier|URI
Attribute|Clinical Attribute|Hospital Course|4581,4588|false|false|false|C0032930|Precipitating Factors|trigger
Disorder|Disease or Syndrome|Hospital Course|4629,4633|false|false|false|C0004238|Atrial Fibrillation|afib
Lab|Laboratory or Test Result|Hospital Course|4629,4633|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|afib
Finding|Finding|Hospital Course|4639,4642|false|false|false|C1417822;C3540498;C4050414|NR1D2 gene;NR1D2 wt Allele;Rapid Virologic Response|RVR
Finding|Gene or Genome|Hospital Course|4639,4642|false|false|false|C1417822;C3540498;C4050414|NR1D2 gene;NR1D2 wt Allele;Rapid Virologic Response|RVR
Drug|Organic Chemical|Hospital Course|4699,4706|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Pharmacologic Substance|Hospital Course|4699,4706|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Substance|Hospital Course|4699,4706|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Finding|Conceptual Entity|Hospital Course|4699,4706|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Functional Concept|Hospital Course|4699,4706|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Idea or Concept|Hospital Course|4699,4706|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4714,4719|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Hospital Course|4714,4719|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Hospital Course|4714,4719|false|false|false|C0795691|HEART PROBLEM|heart
Attribute|Clinical Attribute|Hospital Course|4714,4724|false|false|false|C0018810;C0488794|heart rate|heart rate
Finding|Finding|Hospital Course|4714,4724|false|false|false|C2041121||heart rate
Procedure|Health Care Activity|Hospital Course|4714,4724|false|false|false|C2197023|examination of heart rate|heart rate
Event|Activity|Hospital Course|4720,4724|false|false|false|C0871208|Rating (action)|rate
Finding|Idea or Concept|Hospital Course|4720,4724|false|false|false|C1549480|Amount type - Rate|rate
Procedure|Health Care Activity|Hospital Course|4742,4751|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Anatomy|Anatomical Structure|Hospital Course|4759,4764|false|false|false|C3714591|Floor (anatomic)|floor
Finding|Sign or Symptom|Hospital Course|4789,4797|false|false|false|C0043144|Wheezing|wheezing
Finding|Finding|Hospital Course|4799,4808|false|false|false|C0442805;C5236002|Increase;Increased (finding)|increased
Finding|Functional Concept|Hospital Course|4799,4808|false|false|false|C0442805;C5236002|Increase;Increased (finding)|increased
Finding|Sign or Symptom|Hospital Course|4799,4826|false|false|false|C0859927|Increased work of breathing|increased work of breathing
Event|Occupational Activity|Hospital Course|4809,4813|false|false|false|C0043227|Work|work
Finding|Organ or Tissue Function|Hospital Course|4809,4826|false|false|false|C0043229|Work of Breathing|work of breathing
Attribute|Clinical Attribute|Hospital Course|4817,4826|false|false|false|C5885990||breathing
Finding|Finding|Hospital Course|4817,4826|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|Hospital Course|4817,4826|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|Hospital Course|4817,4826|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|Hospital Course|4817,4826|false|false|false|C1160636|respiratory system process|breathing
Finding|Intellectual Product|Hospital Course|4832,4836|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|poor
Drug|Inorganic Chemical|Hospital Course|4837,4840|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|Hospital Course|4837,4840|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|Hospital Course|4837,4840|false|false|false|C0001861;C3536832|Air (substance);air|air
Finding|Finding|Hospital Course|4837,4840|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|Hospital Course|4837,4840|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|Hospital Course|4837,4840|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Phenomenon|Natural Phenomenon or Process|Hospital Course|4837,4849|false|false|false|C0001868|Air Movements|air movement
Finding|Organism Function|Hospital Course|4841,4849|false|false|false|C0026649|Movement|movement
Drug|Organic Chemical|Hospital Course|4880,4890|false|false|false|C0701466|Solu-Medrol|solumedrol
Drug|Pharmacologic Substance|Hospital Course|4880,4890|false|false|false|C0701466|Solu-Medrol|solumedrol
Drug|Hormone|Hospital Course|4919,4929|false|false|false|C0032952|prednisone|prednisone
Drug|Organic Chemical|Hospital Course|4919,4929|false|false|false|C0032952|prednisone|prednisone
Drug|Pharmacologic Substance|Hospital Course|4919,4929|false|false|false|C0032952|prednisone|prednisone
Finding|Idea or Concept|Hospital Course|4941,4945|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|4941,4945|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|4941,4945|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Hospital Course|4946,4958|false|false|false|C0039771|theophylline|theophylline
Drug|Pharmacologic Substance|Hospital Course|4946,4958|false|false|false|C0039771|theophylline|theophylline
Procedure|Laboratory Procedure|Hospital Course|4946,4958|false|false|false|C0039773|Assay of theophylline|theophylline
Disorder|Mental or Behavioral Dysfunction|Hospital Course|4986,4989|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|4986,4989|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|4986,4989|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|4986,4989|false|false|false|C1332410|BID gene|BID
Disorder|Mental or Behavioral Dysfunction|Hospital Course|5000,5003|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5000,5003|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|5000,5003|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|5000,5003|false|false|false|C1332410|BID gene|BID
Finding|Finding|Hospital Course|5048,5063|false|false|false|C0080203|Tachyarrhythmia|tachyarrhythmia
Drug|Organic Chemical|Hospital Course|5083,5094|false|false|false|C0027235|ipratropium|ipratropium
Drug|Pharmacologic Substance|Hospital Course|5083,5094|false|false|false|C0027235|ipratropium|ipratropium
Drug|Biomedical or Dental Material|Hospital Course|5095,5099|false|false|false|C1300458|Nebulizer solution|nebs
Drug|Organic Chemical|Hospital Course|5106,5115|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|Hospital Course|5106,5115|false|false|false|C0001927|albuterol|albuterol
Drug|Biomedical or Dental Material|Hospital Course|5116,5120|false|false|false|C1300458|Nebulizer solution|nebs
Drug|Organic Chemical|Hospital Course|5130,5141|false|false|false|C0082607|fluticasone|fluticasone
Drug|Pharmacologic Substance|Hospital Course|5130,5141|false|false|false|C0082607|fluticasone|fluticasone
Drug|Pharmacologic Substance|Hospital Course|5130,5152|false|false|false|C0939232|fluticasone / salmeterol|fluticasone-salmeterol
Drug|Organic Chemical|Hospital Course|5142,5152|false|false|false|C0073992|salmeterol|salmeterol
Drug|Pharmacologic Substance|Hospital Course|5142,5152|false|false|false|C0073992|salmeterol|salmeterol
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5154,5163|false|false|false|C0024109|Lung|Pulmonary
Attribute|Clinical Attribute|Hospital Course|5154,5163|false|false|false|C2707265||Pulmonary
Finding|Finding|Hospital Course|5154,5163|false|false|false|C4522268|Pulmonary (intended site)|Pulmonary
Procedure|Research Activity|Hospital Course|5197,5202|false|false|false|C0008976|Clinical Trials|trial
Finding|Organ or Tissue Function|Hospital Course|5206,5214|false|false|false|C0012797|Diuresis|diuresis
Drug|Organic Chemical|Hospital Course|5241,5246|false|false|false|C0699992|Lasix|Lasix
Drug|Pharmacologic Substance|Hospital Course|5241,5246|false|false|false|C0699992|Lasix|Lasix
Finding|Finding|Hospital Course|5250,5254|false|false|false|C5575035|Well (answer to question)|well
Drug|Antibiotic|Hospital Course|5256,5268|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|Azithromycin
Drug|Clinical Drug|Hospital Course|5256,5268|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|Azithromycin
Drug|Organic Chemical|Hospital Course|5256,5268|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|Azithromycin
Drug|Organic Chemical|Hospital Course|5325,5337|false|false|false|C0039771|theophylline|theophylline
Drug|Pharmacologic Substance|Hospital Course|5325,5337|false|false|false|C0039771|theophylline|theophylline
Procedure|Laboratory Procedure|Hospital Course|5325,5337|false|false|false|C0039773|Assay of theophylline|theophylline
Drug|Organic Chemical|Hospital Course|5342,5352|false|false|false|C0002598|amiodarone|amiodarone
Drug|Pharmacologic Substance|Hospital Course|5342,5352|false|false|false|C0002598|amiodarone|amiodarone
Procedure|Laboratory Procedure|Hospital Course|5342,5352|false|false|false|C5399868|Drug assay amiodarone|amiodarone
Finding|Idea or Concept|Hospital Course|5392,5395|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|5392,5395|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Antibiotic|Hospital Course|5406,5417|false|false|false|C0007561|ceftriaxone|ceftriaxone
Drug|Organic Chemical|Hospital Course|5406,5417|false|false|false|C0007561|ceftriaxone|ceftriaxone
Drug|Antibiotic|Hospital Course|5469,5480|false|false|false|C0055011|cefpodoxime|cefpodoxime
Drug|Organic Chemical|Hospital Course|5469,5480|false|false|false|C0055011|cefpodoxime|cefpodoxime
Drug|Hormone|Hospital Course|5509,5519|false|false|false|C0032952|prednisone|prednisone
Drug|Organic Chemical|Hospital Course|5509,5519|false|false|false|C0032952|prednisone|prednisone
Drug|Pharmacologic Substance|Hospital Course|5509,5519|false|false|false|C0032952|prednisone|prednisone
Procedure|Health Care Activity|Hospital Course|5520,5525|false|false|false|C0441640||taper
Finding|Intellectual Product|Hospital Course|5563,5567|false|false|false|C1720594|Then - dosing instruction fragment|then
Procedure|Health Care Activity|Hospital Course|5588,5592|false|false|false|C1315068|Pulmonary ventilator management|pulm
Finding|Functional Concept|Hospital Course|5593,5599|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|Hospital Course|5593,5599|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|Hospital Course|5593,5602|false|false|false|C0589120|Follow-up status|follow up
Procedure|Health Care Activity|Hospital Course|5593,5602|false|false|false|C1522577|follow-up|follow up
Finding|Finding|Hospital Course|5607,5611|false|false|false|C5575035|Well (answer to question)|well
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5631,5640|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Hospital Course|5631,5640|false|false|false|C2707265||pulmonary
Finding|Finding|Hospital Course|5631,5640|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5641,5646|false|false|false|C0034991|Rehabilitation therapy|rehab
Finding|Functional Concept|Hospital Course|5738,5750|false|false|false|C2348609|Supplement|supplemental
Disorder|Disease or Syndrome|Hospital Course|5772,5777|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5782,5788|false|false|false|C0018792|Heart Atrium|Atrial
Attribute|Clinical Attribute|Hospital Course|5782,5801|false|false|false|C2926591||Atrial fibrillation
Disorder|Disease or Syndrome|Hospital Course|5782,5801|false|false|false|C0004238|Atrial Fibrillation|Atrial fibrillation
Lab|Laboratory or Test Result|Hospital Course|5782,5801|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Atrial fibrillation
Disorder|Disease or Syndrome|Hospital Course|5789,5801|false|false|false|C0232197|Fibrillation|fibrillation
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5821,5827|false|false|false|C0018792|Heart Atrium|atrial
Disorder|Disease or Syndrome|Hospital Course|5829,5841|false|false|false|C0232197|Fibrillation|fibrillation
Drug|Organic Chemical|Hospital Course|5863,5873|false|false|false|C0002598|amiodarone|amiodarone
Drug|Pharmacologic Substance|Hospital Course|5863,5873|false|false|false|C0002598|amiodarone|amiodarone
Procedure|Laboratory Procedure|Hospital Course|5863,5873|false|false|false|C5399868|Drug assay amiodarone|amiodarone
Drug|Organic Chemical|Hospital Course|5878,5886|false|false|false|C1831808|apixaban|apixaban
Drug|Pharmacologic Substance|Hospital Course|5878,5886|false|false|false|C1831808|apixaban|apixaban
Disorder|Disease or Syndrome|Hospital Course|5932,5935|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|Hospital Course|5932,5935|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|Hospital Course|5932,5935|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5932,5935|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|Hospital Course|5932,5935|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|Hospital Course|5932,5935|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|Hospital Course|5932,5935|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|Hospital Course|5932,5935|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Finding|Gene or Genome|Hospital Course|5932,5935|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|Hospital Course|5932,5935|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Idea or Concept|Hospital Course|5938,5944|false|false|false|C1549636|Address type - Office|office
Finding|Functional Concept|Hospital Course|5946,5955|false|false|false|C0871157|Prompting|prompting
Procedure|Health Care Activity|Hospital Course|5961,5969|false|false|false|C0034927|Patient referral|referral
Procedure|Health Care Activity|Hospital Course|5961,5972|false|false|false|C2585021|Referral to|referral to
Disorder|Disease or Syndrome|Hospital Course|5985,5989|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Hospital Course|5985,5989|false|false|false|C1647218|COPD pharmacologic substance|COPD
Finding|Gene or Genome|Hospital Course|5985,5989|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|Hospital Course|5985,6002|false|false|false|C0740304|COPD exacerbation|COPD exacerbation
Finding|Finding|Hospital Course|5990,6002|false|false|false|C4086268|Exacerbation|exacerbation
Finding|Finding|Hospital Course|6011,6017|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Hospital Course|6011,6017|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Attribute|Clinical Attribute|Hospital Course|6037,6048|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Hospital Course|6037,6048|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|Hospital Course|6037,6048|false|false|false|C4284232|Medications|medications
Finding|Finding|Hospital Course|6054,6062|false|false|false|C0332149|Possible|possibly
Drug|Organic Chemical|Hospital Course|6091,6103|false|false|false|C0039771|theophylline|theophylline
Drug|Pharmacologic Substance|Hospital Course|6091,6103|false|false|false|C0039771|theophylline|theophylline
Procedure|Laboratory Procedure|Hospital Course|6091,6103|false|false|false|C0039773|Assay of theophylline|theophylline
Drug|Organic Chemical|Hospital Course|6126,6135|false|false|false|C0012373|diltiazem|diltiazem
Drug|Pharmacologic Substance|Hospital Course|6126,6135|false|false|false|C0012373|diltiazem|diltiazem
Disorder|Neoplastic Process|Hospital Course|6136,6139|false|false|false|C1135868|Gestational Trophoblastic Neoplasms|gtt
Drug|Biomedical or Dental Material|Hospital Course|6136,6139|false|false|false|C0991568|Drops - Drug Form|gtt
Procedure|Laboratory Procedure|Hospital Course|6136,6139|false|false|false|C0017741|Glucose tolerance test|gtt
Drug|Organic Chemical|Hospital Course|6193,6202|false|false|false|C0012373|diltiazem|diltiazem
Drug|Pharmacologic Substance|Hospital Course|6193,6202|false|false|false|C0012373|diltiazem|diltiazem
Event|Activity|Hospital Course|6221,6228|false|false|false|C1706079||arrival
Finding|Functional Concept|Hospital Course|6221,6228|false|false|false|C1555577|arrival - ActRelationshipType|arrival
Anatomy|Anatomical Structure|Hospital Course|6236,6241|false|false|false|C3714591|Floor (anatomic)|floor
Drug|Organic Chemical|Hospital Course|6279,6289|false|false|false|C0002598|amiodarone|amiodarone
Drug|Pharmacologic Substance|Hospital Course|6279,6289|false|false|false|C0002598|amiodarone|amiodarone
Procedure|Laboratory Procedure|Hospital Course|6279,6289|false|false|false|C5399868|Drug assay amiodarone|amiodarone
Drug|Organic Chemical|Hospital Course|6294,6302|false|false|false|C1831808|apixaban|apixaban
Drug|Pharmacologic Substance|Hospital Course|6294,6302|false|false|false|C1831808|apixaban|apixaban
Drug|Organic Chemical|Hospital Course|6323,6335|false|false|false|C0039771|theophylline|theophylline
Drug|Pharmacologic Substance|Hospital Course|6323,6335|false|false|false|C0039771|theophylline|theophylline
Procedure|Laboratory Procedure|Hospital Course|6323,6335|false|false|false|C0039773|Assay of theophylline|theophylline
Disorder|Mental or Behavioral Dysfunction|Hospital Course|6361,6364|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6361,6364|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|6361,6364|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|6361,6364|false|false|false|C1332410|BID gene|BID
Disorder|Mental or Behavioral Dysfunction|Hospital Course|6377,6380|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6377,6380|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|6377,6380|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|6377,6380|false|false|false|C1332410|BID gene|BID
Drug|Biologically Active Substance|Hospital Course|6384,6388|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Drug|Element, Ion, or Isotope|Hospital Course|6384,6388|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Drug|Pharmacologic Substance|Hospital Course|6384,6388|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Procedure|Laboratory Procedure|Hospital Course|6384,6388|false|false|false|C0337439|Iron measurement|Iron
Disorder|Disease or Syndrome|Hospital Course|6384,6399|false|false|false|C0162316;C0240066|Iron deficiency;Iron deficiency anemia|Iron deficiency
Disorder|Disease or Syndrome|Hospital Course|6384,6406|false|false|false|C0162316|Iron deficiency anemia|Iron deficiency anemia
Disorder|Disease or Syndrome|Hospital Course|6389,6399|false|false|false|C0162429|Malnutrition|deficiency
Finding|Functional Concept|Hospital Course|6389,6399|false|false|false|C0011155|Deficiency|deficiency
Disorder|Disease or Syndrome|Hospital Course|6389,6406|false|false|false|C0041782|Deficiency anemias|deficiency anemia
Disorder|Disease or Syndrome|Hospital Course|6400,6406|false|false|false|C0002871|Anemia|anemia
Finding|Body Substance|Hospital Course|6408,6415|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|6408,6415|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|6408,6415|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Finding|Hospital Course|6434,6444|false|false|false|C0302870|microcytic|microcytic
Disorder|Disease or Syndrome|Hospital Course|6446,6452|false|false|false|C0002871|Anemia|anemia
Finding|Finding|Hospital Course|6458,6461|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|Hospital Course|6458,6461|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Finding|Hospital Course|6458,6466|false|false|false|C0860975|Iron low|low iron
Drug|Biologically Active Substance|Hospital Course|6462,6466|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Element, Ion, or Isotope|Hospital Course|6462,6466|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Pharmacologic Substance|Hospital Course|6462,6466|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Procedure|Laboratory Procedure|Hospital Course|6462,6466|false|false|false|C0337439|Iron measurement|iron
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6471,6479|false|false|false|C0015879|Ferritin|ferritin
Drug|Biologically Active Substance|Hospital Course|6471,6479|false|false|false|C0015879|Ferritin|ferritin
Drug|Pharmacologic Substance|Hospital Course|6471,6479|false|false|false|C0015879|Ferritin|ferritin
Procedure|Laboratory Procedure|Hospital Course|6471,6479|false|false|false|C0373607|Ferritin measurement|ferritin
Finding|Finding|Hospital Course|6497,6502|false|false|false|C3714655|On IV|on IV
Drug|Element, Ion, or Isotope|Hospital Course|6500,6507|false|false|false|C0082568|ferryl iron|IV iron
Drug|Biologically Active Substance|Hospital Course|6503,6507|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Element, Ion, or Isotope|Hospital Course|6503,6507|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Pharmacologic Substance|Hospital Course|6503,6507|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Procedure|Laboratory Procedure|Hospital Course|6503,6507|false|false|false|C0337439|Iron measurement|iron
Drug|Inorganic Chemical|Hospital Course|6516,6522|false|false|false|C3848561|ferric cation|ferric
Drug|Pharmacologic Substance|Hospital Course|6516,6522|false|false|false|C3848561|ferric cation|ferric
Drug|Organic Chemical|Hospital Course|6516,6532|false|false|false|C0060235|ferric gluconate|ferric gluconate
Drug|Pharmacologic Substance|Hospital Course|6516,6532|false|false|false|C0060235|ferric gluconate|ferric gluconate
Drug|Biologically Active Substance|Hospital Course|6523,6532|false|false|false|C0017714;C0220836|Gluconates;gluconate|gluconate
Drug|Organic Chemical|Hospital Course|6523,6532|false|false|false|C0017714;C0220836|Gluconates;gluconate|gluconate
Drug|Pharmacologic Substance|Hospital Course|6523,6532|false|false|false|C0017714;C0220836|Gluconates;gluconate|gluconate
Drug|Biologically Active Substance|Hospital Course|6566,6570|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Element, Ion, or Isotope|Hospital Course|6566,6570|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Pharmacologic Substance|Hospital Course|6566,6570|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Procedure|Laboratory Procedure|Hospital Course|6566,6570|false|false|false|C0337439|Iron measurement|iron
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6579,6584|false|false|false|C0021853|Intestines|bowel
Procedure|Health Care Activity|Hospital Course|6579,6592|false|false|false|C5979615|Bowel Regimen|bowel regimen
Finding|Intellectual Product|Hospital Course|6585,6592|false|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6585,6592|false|false|false|C0040808|Treatment Protocols|regimen
Finding|Intellectual Product|Hospital Course|6606,6612|false|false|false|C1547311|Patient Condition Code - Stable|stable
Finding|Idea or Concept|Hospital Course|6656,6664|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Hospital Course|6656,6667|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Finding|Pathologic Function|Hospital Course|6668,6676|true|false|false|C0019080|Hemorrhage|bleeding
Finding|Idea or Concept|Hospital Course|6679,6691|false|false|false|C1548597|Marketing basis - Transitional|Transitional
Finding|Body Substance|Hospital Course|6702,6709|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|6702,6709|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|6702,6709|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Hormone|Hospital Course|6724,6734|false|false|false|C0032952|prednisone|prednisone
Drug|Organic Chemical|Hospital Course|6724,6734|false|false|false|C0032952|prednisone|prednisone
Drug|Pharmacologic Substance|Hospital Course|6724,6734|false|false|false|C0032952|prednisone|prednisone
Procedure|Health Care Activity|Hospital Course|6735,6740|false|false|false|C0441640||taper
Finding|Finding|Hospital Course|6742,6750|false|false|false|C0392756|Reduced|decrease
Finding|Intellectual Product|Hospital Course|6790,6794|false|false|false|C1720594|Then - dosing instruction fragment|then
Finding|Body Substance|Hospital Course|6838,6845|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|6838,6845|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|6838,6845|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Disorder|Disease or Syndrome|Hospital Course|6862,6866|false|false|false|C0270724|Infantile Neuroaxonal Dystrophy|plan
Finding|Functional Concept|Hospital Course|6862,6866|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Intellectual Product|Hospital Course|6862,6866|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Mental Process|Hospital Course|6862,6866|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6902,6911|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Hospital Course|6902,6911|false|false|false|C2707265||pulmonary
Finding|Finding|Hospital Course|6902,6911|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6912,6917|false|false|false|C0034991|Rehabilitation therapy|rehab
Event|Activity|Hospital Course|6944,6955|false|false|false|C0003629|Appointments|appointment
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6962,6971|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Hospital Course|6962,6971|false|false|false|C2707265||pulmonary
Finding|Finding|Hospital Course|6962,6971|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6972,6977|false|false|false|C0034991|Rehabilitation therapy|rehab
Finding|Body Substance|Hospital Course|6981,6988|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|6981,6988|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|6981,6988|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Antibiotic|Hospital Course|7018,7029|false|false|false|C0055011|cefpodoxime|cefpodoxime
Drug|Organic Chemical|Hospital Course|7018,7029|false|false|false|C0055011|cefpodoxime|cefpodoxime
Drug|Organic Chemical|Hospital Course|7033,7041|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|Hospital Course|7033,7041|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|Hospital Course|7033,7041|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Finding|Functional Concept|Hospital Course|7033,7041|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|Hospital Course|7033,7041|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|Hospital Course|7045,7048|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|7045,7048|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Antibiotic|Hospital Course|7059,7070|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Finding|Finding|Hospital Course|7075,7081|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|Hospital Course|7075,7081|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Disorder|Disease or Syndrome|Hospital Course|7082,7086|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Hospital Course|7082,7086|false|false|false|C1647218|COPD pharmacologic substance|COPD
Finding|Gene or Genome|Hospital Course|7082,7086|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|Hospital Course|7082,7099|false|false|false|C0740304|COPD exacerbation|COPD exacerbation
Finding|Finding|Hospital Course|7087,7099|false|false|false|C4086268|Exacerbation|exacerbation
Finding|Body Substance|Hospital Course|7102,7109|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|7102,7109|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|7102,7109|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|7146,7156|false|false|false|C0549178|Continuous|continuous
Finding|Idea or Concept|Hospital Course|7157,7161|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|7157,7161|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|7157,7161|false|false|false|C1553498|home health encounter|home
Finding|Body Substance|Hospital Course|7167,7174|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|7167,7174|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|7167,7174|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Organic Chemical|Hospital Course|7177,7189|false|false|false|C0039771|theophylline|theophylline
Drug|Pharmacologic Substance|Hospital Course|7177,7189|false|false|false|C0039771|theophylline|theophylline
Procedure|Laboratory Procedure|Hospital Course|7177,7189|false|false|false|C0039773|Assay of theophylline|theophylline
Disorder|Mental or Behavioral Dysfunction|Hospital Course|7212,7215|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7212,7215|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|7212,7215|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|7212,7215|false|false|false|C1332410|BID gene|BID
Disorder|Mental or Behavioral Dysfunction|Hospital Course|7226,7229|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7226,7229|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|7226,7229|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|7226,7229|false|false|false|C1332410|BID gene|BID
Disorder|Disease or Syndrome|Hospital Course|7242,7246|false|false|false|C0004238|Atrial Fibrillation|afib
Lab|Laboratory or Test Result|Hospital Course|7242,7246|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|afib
Finding|Finding|Hospital Course|7252,7255|false|false|false|C1417822;C3540498;C4050414|NR1D2 gene;NR1D2 wt Allele;Rapid Virologic Response|RVR
Finding|Gene or Genome|Hospital Course|7252,7255|false|false|false|C1417822;C3540498;C4050414|NR1D2 gene;NR1D2 wt Allele;Rapid Virologic Response|RVR
Drug|Organic Chemical|Hospital Course|7287,7299|false|false|false|C0039771|theophylline|theophylline
Drug|Pharmacologic Substance|Hospital Course|7287,7299|false|false|false|C0039771|theophylline|theophylline
Procedure|Laboratory Procedure|Hospital Course|7287,7299|false|false|false|C0039773|Assay of theophylline|theophylline
Finding|Finding|Hospital Course|7300,7304|false|false|false|C0043084|Weaning|wean
Finding|Functional Concept|Hospital Course|7310,7318|false|false|false|C0332287;C1883712|Add - instruction imperative;In addition to|addition
Drug|Antibiotic|Hospital Course|7322,7334|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Clinical Drug|Hospital Course|7322,7334|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Organic Chemical|Hospital Course|7322,7334|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Finding|Body Substance|Hospital Course|7360,7367|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|7360,7367|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|7360,7367|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Organic Chemical|Hospital Course|7376,7386|false|false|false|C0002598|amiodarone|amiodarone
Drug|Pharmacologic Substance|Hospital Course|7376,7386|false|false|false|C0002598|amiodarone|amiodarone
Procedure|Laboratory Procedure|Hospital Course|7376,7386|false|false|false|C5399868|Drug assay amiodarone|amiodarone
Drug|Organic Chemical|Hospital Course|7396,7407|false|false|false|C0965618|roflumilast|roflumilast
Drug|Pharmacologic Substance|Hospital Course|7396,7407|false|false|false|C0965618|roflumilast|roflumilast
Finding|Finding|Hospital Course|7409,7416|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|Hospital Course|7409,7416|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7409,7416|false|false|false|C0087111|Therapeutic procedure|therapy
Finding|Body Substance|Hospital Course|7419,7426|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|7419,7426|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|7419,7426|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Biologically Active Substance|Hospital Course|7439,7443|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Element, Ion, or Isotope|Hospital Course|7439,7443|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Pharmacologic Substance|Hospital Course|7439,7443|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Procedure|Laboratory Procedure|Hospital Course|7439,7443|false|false|false|C0337439|Iron measurement|iron
Finding|Functional Concept|Hospital Course|7444,7453|false|false|false|C0011155|Deficiency|deficient
Finding|Finding|Hospital Course|7463,7468|false|false|false|C3714655|On IV|on IV
Drug|Element, Ion, or Isotope|Hospital Course|7466,7473|false|false|false|C0082568|ferryl iron|IV iron
Drug|Biologically Active Substance|Hospital Course|7469,7473|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Element, Ion, or Isotope|Hospital Course|7469,7473|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Pharmacologic Substance|Hospital Course|7469,7473|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Procedure|Laboratory Procedure|Hospital Course|7469,7473|false|false|false|C0337439|Iron measurement|iron
Drug|Biologically Active Substance|Hospital Course|7503,7507|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Element, Ion, or Isotope|Hospital Course|7503,7507|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Pharmacologic Substance|Hospital Course|7503,7507|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Procedure|Laboratory Procedure|Hospital Course|7503,7507|false|false|false|C0337439|Iron measurement|iron
Finding|Body Substance|Hospital Course|7510,7517|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|7510,7517|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|7510,7517|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Finding|Hospital Course|7532,7544|false|false|false|C0586553|Raised TSH level|elevated TSH
Attribute|Clinical Attribute|Hospital Course|7541,7544|false|false|false|C2708739||TSH
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7541,7544|false|false|false|C0040160|thyrotropin|TSH
Drug|Hormone|Hospital Course|7541,7544|false|false|false|C0040160|thyrotropin|TSH
Drug|Pharmacologic Substance|Hospital Course|7541,7544|false|false|false|C0040160|thyrotropin|TSH
Procedure|Laboratory Procedure|Hospital Course|7541,7544|false|false|false|C0202230|Thyroid stimulating hormone measurement|TSH
Finding|Functional Concept|Hospital Course|7563,7567|false|false|false|C0332296|Free of (attribute)|free
Procedure|Laboratory Procedure|Hospital Course|7563,7570|false|false|false|C0202225|T4 free measurement|free T4
Finding|Idea or Concept|Hospital Course|7582,7589|false|false|false|C1691786;C1704475|Pending - Allergy Clinical Status;Pending - referral status|pending
Finding|Body Substance|Hospital Course|7593,7602|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|7593,7602|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|7593,7602|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|7593,7602|false|false|false|C0030685|Patient Discharge|discharge
Event|Occupational Activity|Hospital Course|7605,7609|false|false|false|C0009219|Coding|Code
Finding|Intellectual Product|Hospital Course|7605,7609|false|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|Code
Finding|Finding|Hospital Course|7618,7627|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Finding|Idea or Concept|Hospital Course|7618,7627|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Finding|Intellectual Product|Hospital Course|7618,7627|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Finding|Pathologic Function|Hospital Course|7618,7627|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Phenomenon|Phenomenon or Process|Hospital Course|7618,7627|false|false|false|C0013956|Emergency Situation|Emergency
Procedure|Health Care Activity|Hospital Course|7618,7627|false|false|false|C1553500|emergency encounter|Emergency
Finding|Functional Concept|Hospital Course|7618,7635|false|false|false|C1552023|emergency contact|Emergency Contact
Event|Activity|Hospital Course|7628,7635|false|false|false|C3812666|Personal Contact|Contact
Finding|Functional Concept|Hospital Course|7628,7635|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|Contact
Finding|Idea or Concept|Hospital Course|7628,7635|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|Contact
Finding|Intellectual Product|Hospital Course|7628,7635|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|Contact
Phenomenon|Phenomenon or Process|Hospital Course|7628,7635|false|false|false|C0392367|Physical contact|Contact
Procedure|Health Care Activity|Hospital Course|7683,7692|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|Hospital Course|7711,7721|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|Hospital Course|7711,7721|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|Hospital Course|7711,7726|false|false|false|C0746470|MEDICATION LIST|Medication list
Finding|Intellectual Product|Hospital Course|7722,7726|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Drug|Organic Chemical|Hospital Course|7743,7751|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|Hospital Course|7743,7751|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|Hospital Course|7743,7751|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Finding|Functional Concept|Hospital Course|7743,7751|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|Hospital Course|7743,7751|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Organic Chemical|Hospital Course|7756,7769|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Hospital Course|7756,7769|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Procedure|Laboratory Procedure|Hospital Course|7756,7769|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|Hospital Course|7784,7787|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|7788,7792|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|7788,7792|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|7788,7792|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|Hospital Course|7797,7805|false|false|false|C1831808|apixaban|Apixaban
Drug|Pharmacologic Substance|Hospital Course|7797,7805|false|false|false|C1831808|apixaban|Apixaban
Disorder|Mental or Behavioral Dysfunction|Hospital Course|7814,7817|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7814,7817|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|7814,7817|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|7814,7817|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|7822,7831|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|Hospital Course|7822,7831|false|false|false|C0001927|albuterol|Albuterol
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7839,7842|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biologically Active Substance|Hospital Course|7839,7842|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biomedical or Dental Material|Hospital Course|7839,7842|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Finding|Cell Function|Hospital Course|7839,7842|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Finding|Gene or Genome|Hospital Course|7839,7842|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7850,7853|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biologically Active Substance|Hospital Course|7850,7853|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biomedical or Dental Material|Hospital Course|7850,7853|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Finding|Cell Function|Hospital Course|7850,7853|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|Hospital Course|7850,7853|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|Hospital Course|7861,7864|false|false|false|C1422467|CIAO3 gene|PRN
Finding|Body Substance|Hospital Course|7879,7885|false|false|false|C0225386|Breath|breath
Drug|Organic Chemical|Hospital Course|7890,7900|false|false|false|C0002598|amiodarone|Amiodarone
Drug|Pharmacologic Substance|Hospital Course|7890,7900|false|false|false|C0002598|amiodarone|Amiodarone
Procedure|Laboratory Procedure|Hospital Course|7890,7900|false|false|false|C5399868|Drug assay amiodarone|Amiodarone
Drug|Organic Chemical|Hospital Course|7921,7933|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|Hospital Course|7921,7933|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|Hospital Course|7951,7967|false|false|false|C0003921;C2608262;C3853661|Artificial Tears;Lubricant Eye Drops;artificial tears (medication)|Artificial Tears
Finding|Body Substance|Hospital Course|7962,7967|false|false|false|C0039409;C1547924;C1611838|Tears (substance);Tears specimen|Tears
Finding|Intellectual Product|Hospital Course|7962,7967|false|false|false|C0039409;C1547924;C1611838|Tears (substance);Tears specimen|Tears
Drug|Biomedical or Dental Material|Hospital Course|7972,7976|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|Hospital Course|7972,7976|false|false|false|C1705648|Dropping|DROP
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7977,7986|false|false|false|C0229118|Structure of both eyes|BOTH EYES
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7982,7986|false|false|false|C0015392|Eye|EYES
Attribute|Clinical Attribute|Hospital Course|7982,7986|false|false|false|C5848506||EYES
Finding|Gene or Genome|Hospital Course|7987,7990|false|false|false|C1422467|CIAO3 gene|PRN
Finding|Intellectual Product|Hospital Course|7991,8001|false|false|false|C1706307;C2700617;C5575347|Have Vulvar Irritation question;Irritability - emotion;Irritation (finding)|irritation
Finding|Mental Process|Hospital Course|7991,8001|false|false|false|C1706307;C2700617;C5575347|Have Vulvar Irritation question;Irritability - emotion;Irritation (finding)|irritation
Finding|Pathologic Function|Hospital Course|7991,8001|false|false|false|C1706307;C2700617;C5575347|Have Vulvar Irritation question;Irritability - emotion;Irritation (finding)|irritation
Phenomenon|Phenomenon or Process|Hospital Course|7991,8001|false|false|false|C0441723|Irritation|irritation
Drug|Organic Chemical|Hospital Course|8006,8017|false|false|false|C0090306|latanoprost|Latanoprost
Drug|Pharmacologic Substance|Hospital Course|8006,8017|false|false|false|C0090306|latanoprost|Latanoprost
Finding|Functional Concept|Hospital Course|8025,8030|false|false|false|C1522230|Ophthalmic Route of Administration|Ophth
Drug|Biomedical or Dental Material|Hospital Course|8040,8044|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|Hospital Course|8040,8044|false|false|false|C1705648|Dropping|DROP
Finding|Functional Concept|Hospital Course|8045,8049|false|false|false|C1552822|Table Cell Horizontal Align - left|LEFT
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8045,8053|false|false|false|C0229090|Left eye structure|LEFT EYE
Procedure|Diagnostic Procedure|Hospital Course|8045,8053|false|false|false|C2141124|examination of left eye|LEFT EYE
Anatomy|Body Location or Region|Hospital Course|8050,8053|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|EYE
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8050,8053|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|EYE
Disorder|Disease or Syndrome|Hospital Course|8050,8053|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|EYE
Disorder|Neoplastic Process|Hospital Course|8050,8053|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|EYE
Finding|Body Substance|Hospital Course|8050,8053|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|EYE
Finding|Finding|Hospital Course|8050,8053|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|EYE
Finding|Intellectual Product|Hospital Course|8050,8053|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|EYE
Drug|Organic Chemical|Hospital Course|8062,8071|false|false|false|C0012373|diltiazem|Diltiazem
Drug|Pharmacologic Substance|Hospital Course|8062,8071|false|false|false|C0012373|diltiazem|Diltiazem
Finding|Finding|Hospital Course|8072,8080|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|8072,8080|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|8081,8088|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|8081,8088|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8081,8088|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8099,8102|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8099,8102|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|8099,8102|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|8099,8102|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|8107,8118|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Hospital Course|8107,8118|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Organic Chemical|Hospital Course|8107,8129|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Pharmacologic Substance|Hospital Course|8107,8129|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Organic Chemical|Hospital Course|8119,8129|false|false|false|C0033474;C0392214|Propionates;propionate|Propionate
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8130,8135|false|false|false|C0028429||NASAL
Drug|Biomedical or Dental Material|Hospital Course|8130,8135|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Drug|Organic Chemical|Hospital Course|8130,8135|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Drug|Pharmacologic Substance|Hospital Course|8130,8135|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Finding|Finding|Hospital Course|8130,8135|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|NASAL
Finding|Functional Concept|Hospital Course|8130,8135|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|NASAL
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8146,8149|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8146,8149|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|8146,8149|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|8146,8149|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|8155,8166|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Hospital Course|8155,8166|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Hospital Course|8155,8177|false|false|false|C0939232|fluticasone / salmeterol|Fluticasone-Salmeterol
Drug|Organic Chemical|Hospital Course|8155,8184|false|false|false|C4762496|Fluticasone-Salmeterol Diskus|Fluticasone-Salmeterol Diskus
Drug|Pharmacologic Substance|Hospital Course|8155,8184|false|false|false|C4762496|Fluticasone-Salmeterol Diskus|Fluticasone-Salmeterol Diskus
Drug|Organic Chemical|Hospital Course|8167,8177|false|false|false|C0073992|salmeterol|Salmeterol
Drug|Pharmacologic Substance|Hospital Course|8167,8177|false|false|false|C0073992|salmeterol|Salmeterol
Drug|Biomedical or Dental Material|Hospital Course|8197,8200|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Organic Chemical|Hospital Course|8197,8200|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Pharmacologic Substance|Hospital Course|8197,8200|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Finding|Functional Concept|Hospital Course|8197,8200|false|false|false|C0205535|Inhalation Route of Administration|INH
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8204,8207|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8204,8207|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|8204,8207|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|8204,8207|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|8213,8232|false|false|false|C0020261|hydrochlorothiazide|Hydrochlorothiazide
Drug|Pharmacologic Substance|Hospital Course|8213,8232|false|false|false|C0020261|hydrochlorothiazide|Hydrochlorothiazide
Drug|Organic Chemical|Hospital Course|8253,8263|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Pharmacologic Substance|Hospital Course|8253,8263|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Organic Chemical|Hospital Course|8253,8275|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Drug|Pharmacologic Substance|Hospital Course|8253,8275|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Finding|Finding|Hospital Course|8277,8285|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|8277,8285|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|8286,8293|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|8286,8293|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8286,8293|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|Hospital Course|8316,8325|false|false|false|C0024002|lorazepam|Lorazepam
Drug|Pharmacologic Substance|Hospital Course|8316,8325|false|false|false|C0024002|lorazepam|Lorazepam
Finding|Gene or Genome|Hospital Course|8340,8343|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Pharmacologic Substance|Hospital Course|8344,8352|false|false|false|C1950154|Insomnia homeopathic medication|insomnia
Finding|Sign or Symptom|Hospital Course|8344,8352|false|false|false|C0917801|Sleeplessness|insomnia
Drug|Organic Chemical|Hospital Course|8358,8370|false|false|false|C0039771|theophylline|Theophylline
Drug|Pharmacologic Substance|Hospital Course|8358,8370|false|false|false|C0039771|theophylline|Theophylline
Procedure|Laboratory Procedure|Hospital Course|8358,8370|false|false|false|C0039773|Assay of theophylline|Theophylline
Drug|Organic Chemical|Hospital Course|8358,8373|false|false|false|C2241157|Theophylline ER|Theophylline ER
Drug|Pharmacologic Substance|Hospital Course|8358,8373|false|false|false|C2241157|Theophylline ER|Theophylline ER
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8384,8387|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8384,8387|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|8384,8387|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|8384,8387|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|8393,8403|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Pharmacologic Substance|Hospital Course|8393,8403|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Organic Chemical|Hospital Course|8425,8435|false|false|false|C0213771|tiotropium|Tiotropium
Drug|Pharmacologic Substance|Hospital Course|8425,8435|false|false|false|C0213771|tiotropium|Tiotropium
Drug|Organic Chemical|Hospital Course|8425,8443|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Pharmacologic Substance|Hospital Course|8425,8443|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Inorganic Chemical|Hospital Course|8436,8443|false|false|false|C0006222|Bromides|Bromide
Procedure|Laboratory Procedure|Hospital Course|8436,8443|false|false|false|C0202341|Bromides measurement|Bromide
Disorder|Congenital Abnormality|Hospital Course|8446,8449|false|false|false|C1855179|CATARACT, ANTERIOR POLAR|CAP
Drug|Biomedical or Dental Material|Hospital Course|8446,8449|false|false|false|C0006935|capsule (pharmacologic)|CAP
Finding|Gene or Genome|Hospital Course|8446,8449|false|false|false|C1416891;C1418551;C1419093;C1422073;C1422760;C2985259;C4522312|BRD4 gene;BRD4 wt Allele;CAP1 gene;HACD1 gene;LNPEP gene;SERPINB6 gene;SORBS1 gene|CAP
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8446,8449|false|false|false|C0278651;C0280547;C1879916|CAP Regimen;cisplatin/cyclophosphamide/doxorubicin protocol;cyclophosphamide/doxorubicin/prednisone protocol|CAP
Drug|Organic Chemical|Hospital Course|8464,8477|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|Hospital Course|8464,8477|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|Hospital Course|8464,8477|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Inorganic Chemical|Hospital Course|8480,8488|false|false|false|C0026162|Minerals|minerals
Drug|Biomedical or Dental Material|Hospital Course|8491,8494|false|false|false|C0039225|Tablet Dosage Form|TAB
Drug|Organic Chemical|Hospital Course|8509,8516|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|Hospital Course|8509,8516|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|Hospital Course|8537,8548|false|false|false|C0165590|dorzolamide|Dorzolamide
Drug|Pharmacologic Substance|Hospital Course|8537,8548|false|false|false|C0165590|dorzolamide|Dorzolamide
Finding|Functional Concept|Hospital Course|8552,8557|false|false|false|C1522230|Ophthalmic Route of Administration|Ophth
Drug|Biomedical or Dental Material|Hospital Course|8567,8571|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|Hospital Course|8567,8571|false|false|false|C1705648|Dropping|DROP
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8572,8581|false|false|false|C0229118|Structure of both eyes|BOTH EYES
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8577,8581|false|false|false|C0015392|Eye|EYES
Attribute|Clinical Attribute|Hospital Course|8577,8581|false|false|false|C5848506||EYES
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8582,8585|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8582,8585|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|8582,8585|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|8582,8585|false|false|false|C1332410|BID gene|BID
Finding|Body Substance|Hospital Course|8590,8599|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|8590,8599|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|8590,8599|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|8590,8599|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|8590,8611|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|8600,8611|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|8600,8611|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|Hospital Course|8600,8611|false|false|false|C4284232|Medications|Medications
Finding|Idea or Concept|Hospital Course|8616,8620|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|8616,8620|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|8616,8620|false|false|false|C1553498|home health encounter|Home
Finding|Idea or Concept|Hospital Course|8633,8643|false|false|false|C0549178|Continuous|continuous
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8644,8649|false|false|false|C0028429||nasal
Drug|Biomedical or Dental Material|Hospital Course|8644,8649|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Organic Chemical|Hospital Course|8644,8649|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Pharmacologic Substance|Hospital Course|8644,8649|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Finding|Finding|Hospital Course|8644,8649|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Functional Concept|Hospital Course|8644,8649|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8650,8657|false|false|false|C1550232|Body Parts - Cannula|cannula
Finding|Body Substance|Hospital Course|8650,8657|false|false|false|C1546577;C1550622|Specimen Type - Cannula|cannula
Finding|Intellectual Product|Hospital Course|8650,8657|false|false|false|C1546577;C1550622|Specimen Type - Cannula|cannula
Finding|Organism Function|Hospital Course|8663,8671|false|false|false|C0015264|Exertion|exertion
Attribute|Clinical Attribute|Hospital Course|8672,8681|false|false|false|C0945731||Diagnosis
Finding|Classification|Hospital Course|8672,8681|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|8672,8681|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|8672,8681|false|false|false|C0011900|Diagnosis|Diagnosis
Finding|Intellectual Product|Hospital Course|8683,8690|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|Hospital Course|8683,8690|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Disorder|Disease or Syndrome|Hospital Course|8683,8720|false|false|false|C0024117|Chronic Obstructive Airway Disease|chronic obstructive pulmonary disease
Finding|Functional Concept|Hospital Course|8691,8702|false|false|false|C0549186|Obstructed|obstructive
Disorder|Disease or Syndrome|Hospital Course|8691,8720|false|false|false|C0600260|Lung Diseases, Obstructive|obstructive pulmonary disease
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8703,8712|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Hospital Course|8703,8712|false|false|false|C2707265||pulmonary
Finding|Finding|Hospital Course|8703,8712|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Disorder|Disease or Syndrome|Hospital Course|8703,8720|false|false|false|C0024115|Lung diseases|pulmonary disease
Finding|Finding|Hospital Course|8703,8720|false|false|false|C0455540|History of - respiratory disease|pulmonary disease
Disorder|Disease or Syndrome|Hospital Course|8713,8720|false|false|false|C0012634|Disease|disease
Finding|Functional Concept|Hospital Course|8739,8744|false|false|false|C0686904|Patient need for (contextual qualifier)|Needs
Finding|Idea or Concept|Hospital Course|8746,8753|false|false|false|C0549178|Continuous|ongoing
Drug|Organic Chemical|Hospital Course|8765,8778|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Hospital Course|8765,8778|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Procedure|Laboratory Procedure|Hospital Course|8765,8778|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|Hospital Course|8793,8796|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|8797,8801|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|8797,8801|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|8797,8801|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|Hospital Course|8806,8816|false|false|false|C0002598|amiodarone|Amiodarone
Drug|Pharmacologic Substance|Hospital Course|8806,8816|false|false|false|C0002598|amiodarone|Amiodarone
Procedure|Laboratory Procedure|Hospital Course|8806,8816|false|false|false|C5399868|Drug assay amiodarone|Amiodarone
Drug|Organic Chemical|Hospital Course|8837,8845|false|false|false|C1831808|apixaban|Apixaban
Drug|Pharmacologic Substance|Hospital Course|8837,8845|false|false|false|C1831808|apixaban|Apixaban
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8854,8857|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8854,8857|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|8854,8857|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|8854,8857|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|8862,8871|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|Hospital Course|8862,8871|false|false|false|C0001927|albuterol|Albuterol
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8879,8882|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biologically Active Substance|Hospital Course|8879,8882|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biomedical or Dental Material|Hospital Course|8879,8882|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Finding|Cell Function|Hospital Course|8879,8882|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Finding|Gene or Genome|Hospital Course|8879,8882|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8890,8893|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biologically Active Substance|Hospital Course|8890,8893|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biomedical or Dental Material|Hospital Course|8890,8893|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Finding|Cell Function|Hospital Course|8890,8893|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|Hospital Course|8890,8893|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|Hospital Course|8901,8904|false|false|false|C1422467|CIAO3 gene|PRN
Finding|Body Substance|Hospital Course|8919,8925|false|false|false|C0225386|Breath|breath
Drug|Pharmacologic Substance|Hospital Course|8930,8946|false|false|false|C0003921;C2608262;C3853661|Artificial Tears;Lubricant Eye Drops;artificial tears (medication)|Artificial Tears
Finding|Body Substance|Hospital Course|8941,8946|false|false|false|C0039409;C1547924;C1611838|Tears (substance);Tears specimen|Tears
Finding|Intellectual Product|Hospital Course|8941,8946|false|false|false|C0039409;C1547924;C1611838|Tears (substance);Tears specimen|Tears
Drug|Biomedical or Dental Material|Hospital Course|8951,8955|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|Hospital Course|8951,8955|false|false|false|C1705648|Dropping|DROP
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8956,8965|false|false|false|C0229118|Structure of both eyes|BOTH EYES
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8961,8965|false|false|false|C0015392|Eye|EYES
Attribute|Clinical Attribute|Hospital Course|8961,8965|false|false|false|C5848506||EYES
Finding|Gene or Genome|Hospital Course|8966,8969|false|false|false|C1422467|CIAO3 gene|PRN
Finding|Intellectual Product|Hospital Course|8970,8980|false|false|false|C1706307;C2700617;C5575347|Have Vulvar Irritation question;Irritability - emotion;Irritation (finding)|irritation
Finding|Mental Process|Hospital Course|8970,8980|false|false|false|C1706307;C2700617;C5575347|Have Vulvar Irritation question;Irritability - emotion;Irritation (finding)|irritation
Finding|Pathologic Function|Hospital Course|8970,8980|false|false|false|C1706307;C2700617;C5575347|Have Vulvar Irritation question;Irritability - emotion;Irritation (finding)|irritation
Phenomenon|Phenomenon or Process|Hospital Course|8970,8980|false|false|false|C0441723|Irritation|irritation
Drug|Organic Chemical|Hospital Course|8985,8992|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|Hospital Course|8985,8992|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|Hospital Course|9012,9024|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|Hospital Course|9012,9024|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|Hospital Course|9042,9051|false|false|false|C0012373|diltiazem|Diltiazem
Drug|Pharmacologic Substance|Hospital Course|9042,9051|false|false|false|C0012373|diltiazem|Diltiazem
Finding|Finding|Hospital Course|9052,9060|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|9052,9060|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|9061,9068|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|9061,9068|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9061,9068|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9079,9082|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9079,9082|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|9079,9082|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|9079,9082|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|9088,9099|false|false|false|C0165590|dorzolamide|Dorzolamide
Drug|Pharmacologic Substance|Hospital Course|9088,9099|false|false|false|C0165590|dorzolamide|Dorzolamide
Finding|Functional Concept|Hospital Course|9103,9108|false|false|false|C1522230|Ophthalmic Route of Administration|Ophth
Drug|Biomedical or Dental Material|Hospital Course|9118,9122|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|Hospital Course|9118,9122|false|false|false|C1705648|Dropping|DROP
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9123,9132|false|false|false|C0229118|Structure of both eyes|BOTH EYES
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9128,9132|false|false|false|C0015392|Eye|EYES
Attribute|Clinical Attribute|Hospital Course|9128,9132|false|false|false|C5848506||EYES
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9133,9136|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9133,9136|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|9133,9136|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|9133,9136|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|9142,9153|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Hospital Course|9142,9153|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Organic Chemical|Hospital Course|9142,9164|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Pharmacologic Substance|Hospital Course|9142,9164|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Organic Chemical|Hospital Course|9154,9164|false|false|false|C0033474;C0392214|Propionates;propionate|Propionate
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9165,9170|false|false|false|C0028429||NASAL
Drug|Biomedical or Dental Material|Hospital Course|9165,9170|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Drug|Organic Chemical|Hospital Course|9165,9170|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Drug|Pharmacologic Substance|Hospital Course|9165,9170|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Finding|Finding|Hospital Course|9165,9170|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|NASAL
Finding|Functional Concept|Hospital Course|9165,9170|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|NASAL
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9181,9184|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9181,9184|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|9181,9184|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|9181,9184|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|9190,9201|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Hospital Course|9190,9201|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Hospital Course|9190,9212|false|false|false|C0939232|fluticasone / salmeterol|Fluticasone-Salmeterol
Drug|Organic Chemical|Hospital Course|9190,9219|false|false|false|C4762496|Fluticasone-Salmeterol Diskus|Fluticasone-Salmeterol Diskus
Drug|Pharmacologic Substance|Hospital Course|9190,9219|false|false|false|C4762496|Fluticasone-Salmeterol Diskus|Fluticasone-Salmeterol Diskus
Drug|Organic Chemical|Hospital Course|9202,9212|false|false|false|C0073992|salmeterol|Salmeterol
Drug|Pharmacologic Substance|Hospital Course|9202,9212|false|false|false|C0073992|salmeterol|Salmeterol
Drug|Biomedical or Dental Material|Hospital Course|9232,9235|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Organic Chemical|Hospital Course|9232,9235|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Pharmacologic Substance|Hospital Course|9232,9235|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Finding|Functional Concept|Hospital Course|9232,9235|false|false|false|C0205535|Inhalation Route of Administration|INH
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9239,9242|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9239,9242|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|9239,9242|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|9239,9242|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|9248,9267|false|false|false|C0020261|hydrochlorothiazide|Hydrochlorothiazide
Drug|Pharmacologic Substance|Hospital Course|9248,9267|false|false|false|C0020261|hydrochlorothiazide|Hydrochlorothiazide
Drug|Organic Chemical|Hospital Course|9288,9298|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Pharmacologic Substance|Hospital Course|9288,9298|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Organic Chemical|Hospital Course|9288,9310|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Drug|Pharmacologic Substance|Hospital Course|9288,9310|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Finding|Finding|Hospital Course|9312,9320|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|9312,9320|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|9321,9328|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|9321,9328|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9321,9328|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|Hospital Course|9351,9362|false|false|false|C0090306|latanoprost|Latanoprost
Drug|Pharmacologic Substance|Hospital Course|9351,9362|false|false|false|C0090306|latanoprost|Latanoprost
Finding|Functional Concept|Hospital Course|9370,9375|false|false|false|C1522230|Ophthalmic Route of Administration|Ophth
Drug|Biomedical or Dental Material|Hospital Course|9385,9389|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|Hospital Course|9385,9389|false|false|false|C1705648|Dropping|DROP
Finding|Functional Concept|Hospital Course|9390,9394|false|false|false|C1552822|Table Cell Horizontal Align - left|LEFT
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9390,9398|false|false|false|C0229090|Left eye structure|LEFT EYE
Procedure|Diagnostic Procedure|Hospital Course|9390,9398|false|false|false|C2141124|examination of left eye|LEFT EYE
Anatomy|Body Location or Region|Hospital Course|9395,9398|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|EYE
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9395,9398|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|EYE
Disorder|Disease or Syndrome|Hospital Course|9395,9398|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|EYE
Disorder|Neoplastic Process|Hospital Course|9395,9398|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|EYE
Finding|Body Substance|Hospital Course|9395,9398|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|EYE
Finding|Finding|Hospital Course|9395,9398|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|EYE
Finding|Intellectual Product|Hospital Course|9395,9398|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|EYE
Drug|Organic Chemical|Hospital Course|9408,9417|false|false|false|C0024002|lorazepam|Lorazepam
Drug|Pharmacologic Substance|Hospital Course|9408,9417|false|false|false|C0024002|lorazepam|Lorazepam
Finding|Gene or Genome|Hospital Course|9432,9435|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Pharmacologic Substance|Hospital Course|9436,9444|false|false|false|C1950154|Insomnia homeopathic medication|insomnia
Finding|Sign or Symptom|Hospital Course|9436,9444|false|false|false|C0917801|Sleeplessness|insomnia
Drug|Organic Chemical|Hospital Course|9450,9463|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|Hospital Course|9450,9463|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|Hospital Course|9450,9463|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Inorganic Chemical|Hospital Course|9466,9474|false|false|false|C0026162|Minerals|minerals
Drug|Biomedical or Dental Material|Hospital Course|9477,9480|false|false|false|C0039225|Tablet Dosage Form|TAB
Drug|Organic Chemical|Hospital Course|9495,9505|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Pharmacologic Substance|Hospital Course|9495,9505|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Organic Chemical|Hospital Course|9527,9537|false|false|false|C0213771|tiotropium|Tiotropium
Drug|Pharmacologic Substance|Hospital Course|9527,9537|false|false|false|C0213771|tiotropium|Tiotropium
Drug|Organic Chemical|Hospital Course|9527,9545|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Pharmacologic Substance|Hospital Course|9527,9545|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Inorganic Chemical|Hospital Course|9538,9545|false|false|false|C0006222|Bromides|Bromide
Procedure|Laboratory Procedure|Hospital Course|9538,9545|false|false|false|C0202341|Bromides measurement|Bromide
Disorder|Congenital Abnormality|Hospital Course|9548,9551|false|false|false|C1855179|CATARACT, ANTERIOR POLAR|CAP
Drug|Biomedical or Dental Material|Hospital Course|9548,9551|false|false|false|C0006935|capsule (pharmacologic)|CAP
Finding|Gene or Genome|Hospital Course|9548,9551|false|false|false|C1416891;C1418551;C1419093;C1422073;C1422760;C2985259;C4522312|BRD4 gene;BRD4 wt Allele;CAP1 gene;HACD1 gene;LNPEP gene;SERPINB6 gene;SORBS1 gene|CAP
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9548,9551|false|false|false|C0278651;C0280547;C1879916|CAP Regimen;cisplatin/cyclophosphamide/doxorubicin protocol;cyclophosphamide/doxorubicin/prednisone protocol|CAP
Drug|Organic Chemical|Hospital Course|9566,9578|false|false|false|C0039771|theophylline|Theophylline
Drug|Pharmacologic Substance|Hospital Course|9566,9578|false|false|false|C0039771|theophylline|Theophylline
Procedure|Laboratory Procedure|Hospital Course|9566,9578|false|false|false|C0039773|Assay of theophylline|Theophylline
Drug|Organic Chemical|Hospital Course|9566,9581|false|false|false|C0939729|Theophylline SR|Theophylline SR
Drug|Pharmacologic Substance|Hospital Course|9566,9581|false|false|false|C0939729|Theophylline SR|Theophylline SR
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9592,9595|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9592,9595|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|9592,9595|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|9592,9595|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|9601,9613|false|false|false|C0039771|theophylline|theophylline
Drug|Pharmacologic Substance|Hospital Course|9601,9613|false|false|false|C0039771|theophylline|theophylline
Procedure|Laboratory Procedure|Hospital Course|9601,9613|false|false|false|C0039773|Assay of theophylline|theophylline
Drug|Biomedical or Dental Material|Hospital Course|9623,9629|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|Hospital Course|9633,9641|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|9636,9641|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|9636,9641|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Idea or Concept|Hospital Course|9650,9653|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|9650,9653|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Activity|Hospital Course|9654,9658|false|false|false|C1880359|Dispense (activity)|Disp
Finding|Gene or Genome|Hospital Course|9654,9658|false|false|false|C2828567|PRSS30P gene|Disp
Drug|Biomedical or Dental Material|Hospital Course|9665,9671|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|Hospital Course|9672,9679|false|false|false|C0807726|refill|Refills
Drug|Antibiotic|Hospital Course|9687,9698|false|false|false|C0055011|cefpodoxime|Cefpodoxime
Drug|Organic Chemical|Hospital Course|9687,9698|false|false|false|C0055011|cefpodoxime|Cefpodoxime
Drug|Antibiotic|Hospital Course|9687,9707|false|false|false|C0108938|cefpodoxime proxetil|Cefpodoxime Proxetil
Drug|Organic Chemical|Hospital Course|9687,9707|false|false|false|C0108938|cefpodoxime proxetil|Cefpodoxime Proxetil
Drug|Pharmacologic Substance|Hospital Course|9723,9731|false|false|false|C0720099|Duration brand of oxymetazoline|Duration
Drug|Antibiotic|Hospital Course|9745,9756|false|false|false|C0055011|cefpodoxime|cefpodoxime
Drug|Organic Chemical|Hospital Course|9745,9756|false|false|false|C0055011|cefpodoxime|cefpodoxime
Drug|Biomedical or Dental Material|Hospital Course|9766,9772|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|Hospital Course|9776,9784|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|9779,9784|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|9779,9784|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Idea or Concept|Hospital Course|9793,9796|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|9793,9796|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Biomedical or Dental Material|Hospital Course|9807,9813|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|Hospital Course|9814,9821|false|false|false|C0807726|refill|Refills
Drug|Element, Ion, or Isotope|Hospital Course|9829,9836|false|false|false|C2346592|Ferrous|Ferrous
Drug|Inorganic Chemical|Hospital Course|9829,9844|false|false|false|C0060282|ferrous sulfate|Ferrous Sulfate
Drug|Pharmacologic Substance|Hospital Course|9829,9844|false|false|false|C0060282|ferrous sulfate|Ferrous Sulfate
Drug|Element, Ion, or Isotope|Hospital Course|9837,9844|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Inorganic Chemical|Hospital Course|9837,9844|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Pharmacologic Substance|Hospital Course|9837,9844|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Element, Ion, or Isotope|Hospital Course|9866,9873|false|false|false|C2346592|Ferrous|ferrous
Drug|Inorganic Chemical|Hospital Course|9866,9881|false|false|false|C0060282|ferrous sulfate|ferrous sulfate
Drug|Pharmacologic Substance|Hospital Course|9866,9881|false|false|false|C0060282|ferrous sulfate|ferrous sulfate
Drug|Element, Ion, or Isotope|Hospital Course|9874,9881|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Inorganic Chemical|Hospital Course|9874,9881|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Pharmacologic Substance|Hospital Course|9874,9881|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Biologically Active Substance|Hospital Course|9896,9900|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Element, Ion, or Isotope|Hospital Course|9896,9900|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Pharmacologic Substance|Hospital Course|9896,9900|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Procedure|Laboratory Procedure|Hospital Course|9896,9900|false|false|false|C0337439|Iron measurement|iron
Drug|Biomedical or Dental Material|Hospital Course|9904,9910|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|Hospital Course|9914,9922|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|9917,9922|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|9917,9922|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Biomedical or Dental Material|Hospital Course|9940,9946|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|Hospital Course|9947,9954|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|9962,9970|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|Hospital Course|9962,9970|false|false|false|C1692318|docusate|Docusate
Drug|Organic Chemical|Hospital Course|9962,9977|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|Hospital Course|9962,9977|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|Hospital Course|9971,9977|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|9971,9977|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|9971,9977|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Finding|Physiologic Function|Hospital Course|9971,9977|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|9971,9977|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9988,9991|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9988,9991|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|9988,9991|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|9988,9991|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|9997,10005|false|false|false|C1692318|docusate|docusate
Drug|Pharmacologic Substance|Hospital Course|9997,10005|false|false|false|C1692318|docusate|docusate
Drug|Organic Chemical|Hospital Course|9997,10012|false|false|false|C0243237|docusate sodium|docusate sodium
Drug|Pharmacologic Substance|Hospital Course|9997,10012|false|false|false|C0243237|docusate sodium|docusate sodium
Drug|Biologically Active Substance|Hospital Course|10006,10012|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Element, Ion, or Isotope|Hospital Course|10006,10012|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Pharmacologic Substance|Hospital Course|10006,10012|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Finding|Physiologic Function|Hospital Course|10006,10012|false|false|false|C4553025|Sodium metabolic function|sodium
Procedure|Laboratory Procedure|Hospital Course|10006,10012|false|false|false|C0337443|Sodium measurement|sodium
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10022,10029|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Anatomy|Cell Component|Hospital Course|10022,10029|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Drug|Biomedical or Dental Material|Hospital Course|10022,10029|false|false|false|C0006935|capsule (pharmacologic)|capsule
Finding|Functional Concept|Hospital Course|10033,10041|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|10036,10041|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|10036,10041|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Idea or Concept|Hospital Course|10050,10053|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|10050,10053|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10065,10072|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|10065,10072|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|10065,10072|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Finding|Idea or Concept|Hospital Course|10073,10080|false|false|false|C0807726|refill|Refills
Drug|Biomedical or Dental Material|Hospital Course|10088,10100|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|Polyethylene
Drug|Organic Chemical|Hospital Course|10088,10100|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|Polyethylene
Drug|Organic Chemical|Hospital Course|10088,10107|false|false|false|C0032483|polyethylene glycols|Polyethylene Glycol
Drug|Pharmacologic Substance|Hospital Course|10088,10107|false|false|false|C0032483|polyethylene glycols|Polyethylene Glycol
Drug|Hazardous or Poisonous Substance|Hospital Course|10101,10107|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|Glycol
Drug|Organic Chemical|Hospital Course|10101,10107|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|Glycol
Drug|Biomedical or Dental Material|Hospital Course|10127,10139|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|polyethylene
Drug|Organic Chemical|Hospital Course|10127,10139|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|polyethylene
Drug|Organic Chemical|Hospital Course|10127,10146|false|false|false|C0032483|polyethylene glycols|polyethylene glycol
Drug|Pharmacologic Substance|Hospital Course|10127,10146|false|false|false|C0032483|polyethylene glycols|polyethylene glycol
Drug|Organic Chemical|Hospital Course|10127,10151|false|false|false|C0724672|polyethylene glycol 3350|polyethylene glycol 3350
Drug|Pharmacologic Substance|Hospital Course|10127,10151|false|false|false|C0724672|polyethylene glycol 3350|polyethylene glycol 3350
Drug|Hazardous or Poisonous Substance|Hospital Course|10140,10146|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|glycol
Drug|Organic Chemical|Hospital Course|10140,10146|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|glycol
Drug|Biomedical or Dental Material|Hospital Course|10167,10173|false|false|false|C0032861;C1382110|Powder dose form;powder physical state|powder
Drug|Substance|Hospital Course|10167,10173|false|false|false|C0032861;C1382110|Powder dose form;powder physical state|powder
Finding|Functional Concept|Hospital Course|10177,10185|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|10180,10185|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|10180,10185|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Idea or Concept|Hospital Course|10193,10200|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|10208,10219|false|false|false|C0027235|ipratropium|Ipratropium
Drug|Pharmacologic Substance|Hospital Course|10208,10219|false|false|false|C0027235|ipratropium|Ipratropium
Drug|Organic Chemical|Hospital Course|10208,10227|false|false|false|C0700580|ipratropium bromide|Ipratropium Bromide
Drug|Pharmacologic Substance|Hospital Course|10208,10227|false|false|false|C0700580|ipratropium bromide|Ipratropium Bromide
Drug|Inorganic Chemical|Hospital Course|10220,10227|false|false|false|C0006222|Bromides|Bromide
Procedure|Laboratory Procedure|Hospital Course|10220,10227|false|false|false|C0202341|Bromides measurement|Bromide
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10228,10231|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biologically Active Substance|Hospital Course|10228,10231|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biomedical or Dental Material|Hospital Course|10228,10231|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Finding|Cell Function|Hospital Course|10228,10231|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Finding|Gene or Genome|Hospital Course|10228,10231|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10234,10237|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biologically Active Substance|Hospital Course|10234,10237|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biomedical or Dental Material|Hospital Course|10234,10237|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Finding|Cell Function|Hospital Course|10234,10237|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|Hospital Course|10234,10237|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|Hospital Course|10245,10248|false|false|false|C1422467|CIAO3 gene|PRN
Finding|Finding|Hospital Course|10249,10256|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|Hospital Course|10249,10256|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|Hospital Course|10258,10266|false|false|false|C0043144|Wheezing|wheezing
Drug|Organic Chemical|Hospital Course|10272,10283|false|false|false|C0027235|ipratropium|ipratropium
Drug|Pharmacologic Substance|Hospital Course|10272,10283|false|false|false|C0027235|ipratropium|ipratropium
Drug|Organic Chemical|Hospital Course|10272,10291|false|false|false|C0700580|ipratropium bromide|ipratropium bromide
Drug|Pharmacologic Substance|Hospital Course|10272,10291|false|false|false|C0700580|ipratropium bromide|ipratropium bromide
Drug|Inorganic Chemical|Hospital Course|10284,10291|false|false|false|C0006222|Bromides|bromide
Procedure|Laboratory Procedure|Hospital Course|10284,10291|false|false|false|C0202341|Bromides measurement|bromide
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10314,10317|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|neb
Drug|Biologically Active Substance|Hospital Course|10314,10317|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|neb
Drug|Biomedical or Dental Material|Hospital Course|10314,10317|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|neb
Finding|Cell Function|Hospital Course|10314,10317|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|neb
Finding|Gene or Genome|Hospital Course|10314,10317|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|neb
Drug|Biomedical or Dental Material|Hospital Course|10318,10321|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Organic Chemical|Hospital Course|10318,10321|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Pharmacologic Substance|Hospital Course|10318,10321|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Finding|Functional Concept|Hospital Course|10318,10321|false|false|false|C0205535|Inhalation Route of Administration|INH
Finding|Intellectual Product|Hospital Course|10322,10327|false|false|false|C1720374|Every - dosing instruction fragment|Every
Finding|Idea or Concept|Hospital Course|10356,10363|false|false|false|C0807726|refill|Refills
Drug|Hormone|Hospital Course|10371,10381|false|false|false|C0032952|prednisone|PredniSONE
Drug|Organic Chemical|Hospital Course|10371,10381|false|false|false|C0032952|prednisone|PredniSONE
Drug|Pharmacologic Substance|Hospital Course|10371,10381|false|false|false|C0032952|prednisone|PredniSONE
Finding|Intellectual Product|Hospital Course|10409,10413|false|false|false|C1720594|Then - dosing instruction fragment|then
Finding|Intellectual Product|Hospital Course|10426,10430|false|false|false|C1720594|Then - dosing instruction fragment|then
Finding|Intellectual Product|Hospital Course|10442,10446|false|false|false|C1720594|Then - dosing instruction fragment|then
Finding|Intellectual Product|Hospital Course|10458,10462|false|false|false|C1720594|Then - dosing instruction fragment|then
Finding|Idea or Concept|Hospital Course|10469,10476|false|false|false|C0549178|Continuous|ongoing
Procedure|Health Care Activity|Hospital Course|10478,10485|false|false|false|C0441640||Tapered
Drug|Hormone|Hospital Course|10503,10513|false|false|false|C0032952|prednisone|prednisone
Drug|Organic Chemical|Hospital Course|10503,10513|false|false|false|C0032952|prednisone|prednisone
Drug|Pharmacologic Substance|Hospital Course|10503,10513|false|false|false|C0032952|prednisone|prednisone
Drug|Biomedical or Dental Material|Hospital Course|10527,10533|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|Hospital Course|10537,10545|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|10540,10545|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|10540,10545|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Biomedical or Dental Material|Hospital Course|10569,10575|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|Hospital Course|10576,10583|false|false|false|C0807726|refill|Refills
Finding|Body Substance|Hospital Course|10590,10599|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|10590,10599|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|10590,10599|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|10590,10599|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|10590,10611|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|10590,10611|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|10600,10611|false|false|false|C2926604||Disposition
Procedure|Health Care Activity|Hospital Course|10600,10611|false|false|false|C0184758|Patient disposition|Disposition
Finding|Idea or Concept|Hospital Course|10613,10617|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|10613,10617|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|10613,10617|false|false|false|C1553498|home health encounter|Home
Event|Occupational Activity|Hospital Course|10623,10630|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|Hospital Course|10623,10630|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Finding|Intellectual Product|Hospital Course|10633,10641|false|false|false|C4695111|ADMIN.FACILITY|Facility
Finding|Body Substance|Hospital Course|10649,10658|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|10649,10658|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|10649,10658|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|10649,10658|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|10649,10668|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|10659,10668|false|false|false|C0945731||Diagnosis
Finding|Classification|Hospital Course|10659,10668|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|10659,10668|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|10659,10668|false|false|false|C0011900|Diagnosis|Diagnosis
Finding|Intellectual Product|Principle Diagnosis|10689,10696|false|false|false|C1547296|Chronic - Admission Level of Care Code|Chronic
Procedure|Health Care Activity|Principle Diagnosis|10689,10696|false|false|false|C1555457|Provision of recurring care for chronic illness|Chronic
Disorder|Disease or Syndrome|Principle Diagnosis|10689,10726|false|false|false|C0024117|Chronic Obstructive Airway Disease|Chronic obstructive pulmonary disease
Finding|Functional Concept|Principle Diagnosis|10697,10708|false|false|false|C0549186|Obstructed|obstructive
Disorder|Disease or Syndrome|Principle Diagnosis|10697,10726|false|false|false|C0600260|Lung Diseases, Obstructive|obstructive pulmonary disease
Anatomy|Body Part, Organ, or Organ Component|Principle Diagnosis|10709,10718|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Principle Diagnosis|10709,10718|false|false|false|C2707265||pulmonary
Finding|Finding|Principle Diagnosis|10709,10718|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Disorder|Disease or Syndrome|Principle Diagnosis|10709,10726|false|false|false|C0024115|Lung diseases|pulmonary disease
Finding|Finding|Principle Diagnosis|10709,10726|false|false|false|C0455540|History of - respiratory disease|pulmonary disease
Disorder|Disease or Syndrome|Principle Diagnosis|10719,10726|false|true|false|C0012634|Disease|disease
Anatomy|Body Part, Organ, or Organ Component|Principle Diagnosis|10727,10733|false|false|false|C0018792|Heart Atrium|Atrial
Attribute|Clinical Attribute|Principle Diagnosis|10727,10746|false|false|false|C2926591||Atrial fibrillation
Disorder|Disease or Syndrome|Principle Diagnosis|10727,10746|false|false|false|C0004238|Atrial Fibrillation|Atrial fibrillation
Lab|Laboratory or Test Result|Principle Diagnosis|10727,10746|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Atrial fibrillation
Disorder|Disease or Syndrome|Principle Diagnosis|10727,10778|false|false|false|C1142306|Atrial fibrillation with rapid ventricular response|Atrial fibrillation with rapid ventricular response
Procedure|Diagnostic Procedure|Principle Diagnosis|10727,10778|false|false|false|C3853730|continuous electrocardiogram monitoring atrial fibrillation with rapid ventricular response|Atrial fibrillation with rapid ventricular response
Disorder|Disease or Syndrome|Principle Diagnosis|10734,10746|false|false|false|C0232197|Fibrillation|fibrillation
Disorder|Disease or Syndrome|Principle Diagnosis|10752,10778|false|false|false|C0748243|rapid ventricular response|rapid ventricular response
Anatomy|Body Part, Organ, or Organ Component|Principle Diagnosis|10758,10769|false|false|false|C0018827|Heart Ventricle|ventricular
Finding|Finding|Principle Diagnosis|10770,10778|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Intellectual Product|Principle Diagnosis|10770,10778|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Mental Process|Principle Diagnosis|10770,10778|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Disorder|Neoplastic Process|Principle Diagnosis|10780,10789|false|false|false|C0027627|Neoplasm Metastasis|Secondary
Finding|Functional Concept|Principle Diagnosis|10780,10789|false|false|false|C1522484|metastatic qualifier|Secondary
Procedure|Diagnostic Procedure|Principle Diagnosis|10790,10799|false|false|false|C0011900|Diagnosis|diagnoses
Disorder|Disease or Syndrome|Principle Diagnosis|10801,10813|false|false|false|C0020538|Hypertensive disease|Hypertension
Anatomy|Body Part, Organ, or Organ Component|Principle Diagnosis|10814,10822|false|false|false|C0018787|Heart|Coronary
Anatomy|Body Part, Organ, or Organ Component|Principle Diagnosis|10814,10829|false|false|false|C0205042|Coronary artery|Coronary artery
Disorder|Disease or Syndrome|Principle Diagnosis|10814,10837|false|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|Coronary artery disease
Anatomy|Body Part, Organ, or Organ Component|Principle Diagnosis|10823,10829|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|Principle Diagnosis|10823,10829|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Disorder|Disease or Syndrome|Principle Diagnosis|10823,10837|false|false|false|C0852949|Arteriopathic disease|artery disease
Disorder|Disease or Syndrome|Principle Diagnosis|10830,10837|false|false|false|C0012634|Disease|disease
Disorder|Disease or Syndrome|Principle Diagnosis|10838,10865|false|false|false|C0085096|Peripheral Vascular Diseases|Peripheral vascular disease
Anatomy|Body Part, Organ, or Organ Component|Principle Diagnosis|10849,10857|false|false|false|C0005847|Blood Vessel|vascular
Disorder|Disease or Syndrome|Principle Diagnosis|10849,10865|false|false|false|C0042373|Vascular Diseases|vascular disease
Disorder|Disease or Syndrome|Principle Diagnosis|10858,10865|false|false|false|C0012634|Disease|disease
Finding|Mental Process|Discharge Condition|10890,10896|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|10890,10903|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|10890,10903|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|10897,10903|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|10897,10903|false|false|false|C1546481|What subject filter - Status|Status
Finding|Idea or Concept|Discharge Condition|10905,10910|false|false|false|C1550016|Remote control command - Clear|Clear
Finding|Finding|Discharge Condition|10915,10923|false|false|false|C4068804|Coherent|coherent
Attribute|Clinical Attribute|Discharge Condition|10925,10947|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|10925,10947|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Finding|Finding|Discharge Condition|10934,10947|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|10934,10947|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|10949,10954|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|10949,10954|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|10949,10954|false|false|false|C0718338|Alert brand of caffeine|Alert
Finding|Finding|Discharge Condition|10949,10954|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|10949,10954|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|10949,10954|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|10959,10970|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|10972,10980|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|10972,10980|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|10972,10980|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|10981,10987|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|10981,10987|false|false|false|C1546481|What subject filter - Status|Status
Finding|Functional Concept|Discharge Condition|10989,10999|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|Discharge Condition|10989,10999|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|Discharge Condition|10989,10999|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|Discharge Condition|10989,10999|false|false|false|C1561560|ambulatory encounter|Ambulatory
Finding|Finding|Discharge Condition|11002,11013|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|Discharge Condition|11002,11013|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Gene or Genome|Discharge Instructions|11042,11046|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Finding|Finding|Discharge Instructions|11111,11121|false|false|false|C1299586|Has difficulty doing (qualifier value)|difficulty
Finding|Sign or Symptom|Discharge Instructions|11111,11131|false|false|false|C0013404;C0476273|Dyspnea;Respiratory distress|difficulty breathing
Attribute|Clinical Attribute|Discharge Instructions|11122,11131|false|false|false|C5885990||breathing
Finding|Finding|Discharge Instructions|11122,11131|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|Discharge Instructions|11122,11131|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|Discharge Instructions|11122,11131|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|Discharge Instructions|11122,11131|false|false|false|C1160636|respiratory system process|breathing
Finding|Finding|Discharge Instructions|11168,11172|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|fast
Finding|Gene or Genome|Discharge Instructions|11168,11172|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|fast
Finding|Molecular Function|Discharge Instructions|11168,11172|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|fast
Finding|Finding|Discharge Instructions|11168,11183|false|false|false|C0039231|Tachycardia|fast heart rate
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|11173,11178|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Discharge Instructions|11173,11178|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Discharge Instructions|11173,11178|false|false|false|C0795691|HEART PROBLEM|heart
Attribute|Clinical Attribute|Discharge Instructions|11173,11183|false|false|false|C0018810;C0488794|heart rate|heart rate
Finding|Finding|Discharge Instructions|11173,11183|false|false|false|C2041121||heart rate
Procedure|Health Care Activity|Discharge Instructions|11173,11183|false|false|false|C2197023|examination of heart rate|heart rate
Event|Activity|Discharge Instructions|11179,11183|false|false|false|C0871208|Rating (action)|rate
Finding|Idea or Concept|Discharge Instructions|11179,11183|false|false|false|C1549480|Amount type - Rate|rate
Finding|Finding|Discharge Instructions|11190,11200|false|false|false|C1299586|Has difficulty doing (qualifier value)|difficulty
Finding|Sign or Symptom|Discharge Instructions|11190,11210|false|false|false|C0013404;C0476273|Dyspnea;Respiratory distress|difficulty breathing
Attribute|Clinical Attribute|Discharge Instructions|11201,11210|false|false|false|C5885990||breathing
Finding|Finding|Discharge Instructions|11201,11210|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|Discharge Instructions|11201,11210|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|Discharge Instructions|11201,11210|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|Discharge Instructions|11201,11210|false|false|false|C1160636|respiratory system process|breathing
Disorder|Disease or Syndrome|Discharge Instructions|11228,11232|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Discharge Instructions|11228,11232|false|false|false|C1647218|COPD pharmacologic substance|COPD
Finding|Gene or Genome|Discharge Instructions|11228,11232|false|false|false|C1412502|ARCN1 gene|COPD
Finding|Finding|Discharge Instructions|11247,11251|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|fast
Finding|Gene or Genome|Discharge Instructions|11247,11251|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|fast
Finding|Molecular Function|Discharge Instructions|11247,11251|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|fast
Finding|Finding|Discharge Instructions|11247,11262|false|false|false|C0039231|Tachycardia|fast heart rate
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|11252,11257|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Discharge Instructions|11252,11257|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Discharge Instructions|11252,11257|false|false|false|C0795691|HEART PROBLEM|heart
Attribute|Clinical Attribute|Discharge Instructions|11252,11262|false|false|false|C0018810;C0488794|heart rate|heart rate
Finding|Finding|Discharge Instructions|11252,11262|false|false|false|C2041121||heart rate
Procedure|Health Care Activity|Discharge Instructions|11252,11262|false|false|false|C2197023|examination of heart rate|heart rate
Event|Activity|Discharge Instructions|11258,11262|false|false|false|C0871208|Rating (action)|rate
Finding|Idea or Concept|Discharge Instructions|11258,11262|false|false|false|C1549480|Amount type - Rate|rate
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|11280,11286|false|false|false|C0018792|Heart Atrium|atrial
Attribute|Clinical Attribute|Discharge Instructions|11280,11299|false|false|false|C2926591||atrial fibrillation
Disorder|Disease or Syndrome|Discharge Instructions|11280,11299|false|false|false|C0004238|Atrial Fibrillation|atrial fibrillation
Lab|Laboratory or Test Result|Discharge Instructions|11280,11299|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|atrial fibrillation
Disorder|Disease or Syndrome|Discharge Instructions|11287,11299|false|false|false|C0232197|Fibrillation|fibrillation
Finding|Finding|Discharge Instructions|11313,11333|false|false|false|C0237314|Irregular heart beat|irregular heart rate
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|11323,11328|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Discharge Instructions|11323,11328|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Discharge Instructions|11323,11328|false|false|false|C0795691|HEART PROBLEM|heart
Attribute|Clinical Attribute|Discharge Instructions|11323,11333|false|false|false|C0018810;C0488794|heart rate|heart rate
Finding|Finding|Discharge Instructions|11323,11333|false|false|false|C2041121||heart rate
Procedure|Health Care Activity|Discharge Instructions|11323,11333|false|false|false|C2197023|examination of heart rate|heart rate
Event|Activity|Discharge Instructions|11329,11333|false|false|false|C0871208|Rating (action)|rate
Finding|Idea or Concept|Discharge Instructions|11329,11333|false|false|false|C1549480|Amount type - Rate|rate
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|11364,11369|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Discharge Instructions|11364,11369|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Discharge Instructions|11364,11369|false|false|false|C0795691|HEART PROBLEM|heart
Attribute|Clinical Attribute|Discharge Instructions|11392,11403|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Discharge Instructions|11392,11403|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|Discharge Instructions|11392,11403|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Discharge Instructions|11435,11447|false|false|false|C0039771|theophylline|theophylline
Drug|Pharmacologic Substance|Discharge Instructions|11435,11447|false|false|false|C0039771|theophylline|theophylline
Procedure|Laboratory Procedure|Discharge Instructions|11435,11447|false|false|false|C0039773|Assay of theophylline|theophylline
Finding|Finding|Discharge Instructions|11454,11460|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Discharge Instructions|11454,11460|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|11481,11486|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Discharge Instructions|11481,11486|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Discharge Instructions|11481,11486|false|false|false|C0795691|HEART PROBLEM|heart
Attribute|Clinical Attribute|Discharge Instructions|11481,11491|false|false|false|C0018810;C0488794|heart rate|heart rate
Finding|Finding|Discharge Instructions|11481,11491|false|false|false|C2041121||heart rate
Procedure|Health Care Activity|Discharge Instructions|11481,11491|false|false|false|C2197023|examination of heart rate|heart rate
Event|Activity|Discharge Instructions|11487,11491|false|false|false|C0871208|Rating (action)|rate
Finding|Idea or Concept|Discharge Instructions|11487,11491|false|false|false|C1549480|Amount type - Rate|rate
Drug|Pharmacologic Substance|Discharge Instructions|11519,11529|false|false|false|C0013227|Pharmaceutical Preparations|medication
Finding|Intellectual Product|Discharge Instructions|11519,11529|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Finding|Finding|Discharge Instructions|11545,11552|false|false|false|C4534363|At home|at home
Finding|Idea or Concept|Discharge Instructions|11548,11552|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Discharge Instructions|11548,11552|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Discharge Instructions|11548,11552|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Discharge Instructions|11554,11563|false|false|false|C0012373|diltiazem|diltiazem
Drug|Pharmacologic Substance|Discharge Instructions|11554,11563|false|false|false|C0012373|diltiazem|diltiazem
Disorder|Disease or Syndrome|Discharge Instructions|11595,11599|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Discharge Instructions|11595,11599|false|false|false|C1647218|COPD pharmacologic substance|COPD
Finding|Gene or Genome|Discharge Instructions|11595,11599|false|false|false|C1412502|ARCN1 gene|COPD
Finding|Finding|Discharge Instructions|11604,11610|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Discharge Instructions|11604,11610|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Disorder|Disease or Syndrome|Discharge Instructions|11633,11637|false|false|false|C0009443;C0024117|Chronic Obstructive Airway Disease;Common Cold|cold
Drug|Organic Chemical|Discharge Instructions|11633,11637|false|false|false|C0719425|Cold brand of chlorpheniramine-phenylpropanolamine|cold
Drug|Pharmacologic Substance|Discharge Instructions|11633,11637|false|false|false|C0719425|Cold brand of chlorpheniramine-phenylpropanolamine|cold
Finding|Organism Function|Discharge Instructions|11633,11637|false|false|false|C0234192|Cold Sensation|cold
Phenomenon|Natural Phenomenon or Process|Discharge Instructions|11633,11637|false|false|false|C0009264|Cold Temperature|cold
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|11633,11637|false|false|false|C0010412|Cold Therapy|cold
Finding|Finding|Discharge Instructions|11654,11659|false|false|false|C1517205;C3540542|Exacerbation of cGVHD;Flare|flare
Finding|Sign or Symptom|Discharge Instructions|11654,11659|false|false|false|C1517205;C3540542|Exacerbation of cGVHD;Flare|flare
Finding|Finding|Discharge Instructions|11669,11676|false|false|false|C1551395;C1552745;C1561576|Alert level - Serious;Device Alert Level - Serious;Equipment Alert Level - Serious|serious
Finding|Idea or Concept|Discharge Instructions|11669,11676|false|false|false|C1551395;C1552745;C1561576|Alert level - Serious;Device Alert Level - Serious;Equipment Alert Level - Serious|serious
Drug|Organic Chemical|Discharge Instructions|11690,11698|false|false|false|C0038317|Steroids|steroids
Drug|Pharmacologic Substance|Discharge Instructions|11690,11698|false|false|false|C0038317|Steroids|steroids
Finding|Organism Function|Discharge Instructions|11708,11715|false|false|false|C0004048|Inspiration (function)|inhaled
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|11717,11727|false|false|false|C0087111|Therapeutic procedure|treatments
Anatomy|Body Location or Region|Discharge Instructions|11759,11763|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|11759,11763|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Discharge Instructions|11759,11763|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Discharge Instructions|11759,11763|false|false|false|C0740941|Lung Problem|lung
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|11788,11797|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Discharge Instructions|11788,11797|false|false|false|C2707265||pulmonary
Finding|Finding|Discharge Instructions|11788,11797|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|11798,11803|false|false|false|C0034991|Rehabilitation therapy|rehab
Finding|Intellectual Product|Discharge Instructions|11812,11816|false|false|false|C4724437|SURE Test|sure
Anatomy|Body Location or Region|Discharge Instructions|11822,11826|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|11822,11826|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Discharge Instructions|11822,11826|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Discharge Instructions|11822,11826|false|false|false|C0740941|Lung Problem|lung
Disorder|Disease or Syndrome|Discharge Instructions|11822,11834|false|false|false|C0024115|Lung diseases|lung disease
Disorder|Disease or Syndrome|Discharge Instructions|11827,11834|false|false|false|C0012634|Disease|disease
Finding|Finding|Discharge Instructions|11856,11860|false|false|false|C5575035|Well (answer to question)|well
Finding|Finding|Discharge Instructions|11864,11872|false|false|false|C0332149|Possible|possible
Finding|Idea or Concept|Discharge Instructions|11910,11918|false|false|false|C1547192|Organization unit type - Hospital|hospital
Finding|Intellectual Product|Discharge Instructions|11922,11927|false|false|false|C4050225|Often - answer to question|often
Event|Activity|Discharge Instructions|11961,11972|false|false|false|C0003629|Appointments|appointment
Finding|Intellectual Product|Discharge Instructions|11994,12002|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|Discharge Instructions|11994,12002|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|Discharge Instructions|12025,12029|false|false|false|C1947933|care activity|care
Finding|Finding|Discharge Instructions|12025,12029|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|12025,12029|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Disorder|Disease or Syndrome|Discharge Instructions|12052,12056|false|false|false|C0339510|Vitelliform Macular Dystrophy|best
Finding|Gene or Genome|Discharge Instructions|12052,12056|false|false|false|C1826421;C5781213|BEST1 gene;BEST1 wt Allele|best
Procedure|Health Care Activity|Discharge Instructions|12101,12109|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|12110,12122|false|false|false|C3263700||Instructions
Finding|Intellectual Product|Discharge Instructions|12110,12122|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

