CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Pharmaceutical Preparations|Drug|false|false||MEDICINEnull|Medicine|Title|false|false||MEDICINEnull|INJECTION, MEROPENEM, 100 MG ADMINISTERED|Drug|false|false||meropenem
null|meropenem|Drug|false|false||meropenem
null|meropenem|Drug|false|false||meropenemnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Complaint (finding)|Finding|false|false||Complaintnull|null|Attribute|false|false||Complaintnull|Respiratory Failure|Disorder|false|false||Respiratory Failurenull|Respiratory attachment|Finding|false|false||Respiratory
null|respiratory|Finding|false|false||Respiratory
null|null|Finding|false|false||Respiratory
null|Respiratory specimen|Finding|false|false||Respiratorynull|Respiratory rate|Attribute|false|false||Respiratorynull|Failure (biologic function)|Finding|false|false||Failure
null|Failure|Finding|false|false||Failure
null|Personal failure|Finding|false|false||Failurenull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|mechanical method|Finding|false|false||Mechanicalnull|Mechanical Treatments|Procedure|false|false||Mechanicalnull|Intubation (procedure)|Procedure|false|false||Intubationnull|Arteries|Anatomy|false|false||Arterialnull|Arterial|Modifier|false|false||Arterialnull|Line Specimen|Drug|false|false||Line
null|Long Interspersed Elements|Drug|false|false||Line
null|Long Interspersed Elements|Drug|false|false||Linenull|line source specimen code|Finding|false|false||Linenull|Intravascular line|Device|false|false||Linenull|Linear|Modifier|false|false||Linenull|Line Unit of Length|LabModifier|false|false||Linenull|central venous|Modifier|false|false||Central Venousnull|Central brand of multivitamin with minerals|Drug|false|false||Central
null|Central brand of multivitamin with minerals|Drug|false|false||Centralnull|Central Minus|Procedure|false|false||Centralnull|Central|Modifier|false|false||Centralnull|venous access|Device|false|false||Venous Accessnull|Veins|Anatomy|false|false||Venousnull|Venous|Modifier|false|false||Venousnull|Role Class - access|Finding|false|false||Accessnull|Access|Modifier|false|false||Accessnull|Line Specimen|Drug|false|false||Line
null|Long Interspersed Elements|Drug|false|false||Line
null|Long Interspersed Elements|Drug|false|false||Linenull|line source specimen code|Finding|false|false||Linenull|Intravascular line|Device|false|false||Linenull|Linear|Modifier|false|false||Linenull|Line Unit of Length|LabModifier|false|false||Linenull|Transaction counts and value totals - year|Finding|false|false||year
null|Precision - year|Finding|false|false||yearnull|year|Time|false|false||yearnull|Old|Time|false|false||oldnull|Woman|Subject|false|false||woman
null|Human, Female adult|Subject|false|false||womannull|Recent|Time|false|false||recentlynull|Sepsis|Disorder|false|false||sepsis
null|Septicemia|Disorder|false|false||sepsisnull|Sepsis <Sepsidae>|Entity|false|false||sepsisnull|Shock|Finding|false|false||shocknull|Readmission|Procedure|false|false||readmissionnull|Hypoxia, CTCAE|Finding|false|false||hypoxia
null|Hypoxia|Finding|false|false||hypoxianull|Hypercapnia|Finding|false|false||hypercarbianull|Respiratory attachment|Finding|false|false||respiratory
null|respiratory|Finding|false|false||respiratory
null|null|Finding|false|false||respiratory
null|Respiratory specimen|Finding|false|false||respiratorynull|Respiratory rate|Attribute|false|false||respiratorynull|Emotional distress|Finding|false|false||distress
null|Distress|Finding|false|false||distressnull|Respiratory Failure|Disorder|false|false||respiratory failurenull|Respiratory attachment|Finding|false|false||respiratory
null|respiratory|Finding|false|false||respiratory
null|null|Finding|false|false||respiratory
null|Respiratory specimen|Finding|false|false||respiratorynull|Respiratory rate|Attribute|false|false||respiratorynull|Failure (biologic function)|Finding|false|false||failure
null|Failure|Finding|false|false||failure
null|Personal failure|Finding|false|false||failurenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Rehabilitation therapy|Procedure|false|false||rehabnull|Depressed mood|Disorder|false|false||depressednull|Mental state|Finding|false|false||mental statusnull|null|Attribute|false|false||mental status
null|null|Attribute|false|false||mental statusnull|Psyche structure|Finding|false|false||mentalnull|What subject filter - Status|Finding|false|false||statusnull|null|Attribute|false|false||statusnull|Social status|Modifier|false|false||status
null|Status|Modifier|false|false||statusnull|Tachypnea|Finding|false|false||tachypneanull|null|Finding|false|false||dyspnea
null|Dyspnea|Finding|false|false||dyspneanull|Ethyl Methanesulfonate|Drug|false|false||EMS
null|Ethyl Methanesulfonate|Drug|false|false||EMS
null|Ethyl Methanesulfonate|Drug|false|false||EMSnull|EMSLR gene|Finding|false|false||EMSnull|Emergency Medical Services|Procedure|false|false||EMSnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Intubation (procedure)|Procedure|false|false||intubationnull|Airway structure|Anatomy|false|false||airway
null|Chest>Airway|Anatomy|false|false||airwaynull|Artificial Airways|Device|false|false||airwaynull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Certification patient type - Emergency|Finding|false|false||emergency
null|Consent Non-Disclosure Reason - Emergency|Finding|false|false||emergency
null|Admission Type - Emergency|Finding|false|false||emergency
null|Referral category - Emergency|Finding|false|false||emergency
null|Emergencies [Disease/Finding]|Finding|false|false||emergency
null|Consent Bypass Reason - Emergency|Finding|false|false||emergency
null|Level of Care - Emergency|Finding|false|false||emergency
null|Encounter Admission Source - emergency|Finding|false|false||emergency
null|Patient Class - Emergency|Finding|false|false||emergency
null|Visit Priority Code - Emergency|Finding|false|false||emergencynull|emergency encounter|Procedure|false|false||emergencynull|Emergency Situation|Phenomenon|false|false||emergencynull|Specialty Type - Emergency|Title|false|false||emergencynull|Bale out|Time|false|false||emergencynull|Department - No suggested values defined|Finding|false|false||department
null|Organization Unit Type - Department|Finding|false|false||department
null|Department - Charge type|Finding|false|false||departmentnull|Department|Entity|false|false||departmentnull|Patient location type - Department|Modifier|false|false||department
null|Department - Person location type|Modifier|false|false||departmentnull|Report (document)|Finding|true|false||reportsnull|Reporting|Procedure|true|false||reportsnull|Increasing frequency of cough|Finding|true|false||increased coughingnull|Increased (finding)|Finding|true|false||increased
null|Increase|Finding|true|false||increasednull|Increased|LabModifier|false|false||increasednull|Coughing|Finding|true|false||coughingnull|Has patient|Finding|false|false||patient hasnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Complicated|Finding|false|false||complicatednull|Medical referral type|Finding|false|false||medical
null|Medical|Finding|false|false||medical
null|Medical school type|Finding|false|false||medicalnull|Medical service|Procedure|false|false||medicalnull|Course|Time|false|false||coursenull|Transaction counts and value totals - month|Finding|false|false||month
null|Precision - month|Finding|false|false||monthnull|month|Time|false|false||month
null|Monthly (qualifier value)|Time|false|false||monthnull|BRIEF Health Literacy Screening Tool|Finding|false|false||brief
null|Behavior Rating Inventory of Executive Function|Finding|false|false||briefnull|Brief|Time|false|false||briefnull|Shortened|Modifier|false|false||briefnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Initially|Time|false|false||initiallynull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Clostridium difficile colitis|Disorder|false|false||c.diff colitisnull|Colitis|Disorder|false|false||colitisnull|Sepsis|Disorder|false|false||sepsis
null|Septicemia|Disorder|false|false||sepsisnull|Sepsis <Sepsidae>|Entity|false|false||sepsisnull|Respiratory Failure|Disorder|false|false||respiratory failurenull|Respiratory attachment|Finding|false|false||respiratory
null|respiratory|Finding|false|false||respiratory
null|null|Finding|false|false||respiratory
null|Respiratory specimen|Finding|false|false||respiratorynull|Respiratory rate|Attribute|false|false||respiratorynull|Failure (biologic function)|Finding|false|false||failure
null|Failure|Finding|false|false||failure
null|Personal failure|Finding|false|false||failurenull|Intubation (procedure)|Procedure|false|false||intubationnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Dyspnea|Finding|false|false||SOBnull|A1BG gene|Finding|false|false||ABGnull|Analysis of arterial blood gases and pH|Procedure|false|false||ABGnull|Biphasic Continuous Positive Airway Pressure|Procedure|false|false||biPAPnull|HDAC1 protein, human|Drug|false|false||HD1
null|HDAC1 protein, human|Drug|false|false||HD1null|HDAC1 wt Allele|Finding|false|false||HD1
null|HDAC1 gene|Finding|false|false||HD1
null|PLEC wt Allele|Finding|false|false||HD1null|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygennull|Oxygen Therapy Care|Procedure|false|false||oxygennull|Oxygen Equipment Location|Modifier|false|false||oxygennull|Requirement|Finding|false|false||requirementnull|Science of Etiology|Finding|false|false||etiology
null|Etiology aspects|Finding|false|false||etiology
null|Etiology|Finding|false|false||etiologynull|Respiratory attachment|Finding|false|false||respiratory
null|respiratory|Finding|false|false||respiratory
null|null|Finding|false|false||respiratory
null|Respiratory specimen|Finding|false|false||respiratorynull|Respiratory rate|Attribute|false|false||respiratorynull|Failure (biologic function)|Finding|false|false||failure
null|Failure|Finding|false|false||failure
null|Personal failure|Finding|false|false||failurenull|Hypoventilation|Finding|false|false||hypoventilationnull|Somnolence|Disorder|false|false||somnolencenull|Drowsiness|Finding|false|false||somnolencenull|Relate - vinyl resin|Drug|false|false||relatednull|Role Link Type - related|Finding|false|false||related
null|Related (finding)|Finding|false|false||relatednull|Definitely Related to Intervention|Modifier|false|false||related
null|Relationships|Modifier|false|false||relatednull|Oversedation|Finding|false|false||oversedationnull|Zyprexa|Drug|false|false||zyprexa
null|Zyprexa|Drug|false|false||zyprexanull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Cancer/Testis Antigen|Drug|false|false||CTAnull|PCYT1A wt Allele|Finding|false|false||CTA
null|CERNA3 gene|Finding|false|false||CTAnull|Cardiac Computerized Tomographic Angiography|Procedure|false|false||CTAnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Negative|Finding|false|false||negative fornull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Remote control command - Clear|Finding|false|false||clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|Evidence of (contextual qualifier)|Finding|false|false||evidence ofnull|Evidence|Finding|false|false||evidencenull|Pneumonia|Disorder|false|false||pneumonianull|Initially|Time|false|false||initiallynull|SMC3 protein, human|Drug|false|false||HCAP
null|SMC3 protein, human|Drug|false|false||HCAPnull|SMC3 wt Allele|Finding|false|false||HCAP
null|RNGTT gene|Finding|false|false||HCAP
null|SMC3 gene|Finding|false|false||HCAP
null|DCD gene|Finding|false|false||HCAPnull|Cyclophosphamide/Altretamine/Doxorubicin/Cisplatin Regimen|Procedure|false|false||HCAPnull|Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE|Drug|false|false||antibiotics
null|Antibiotics|Drug|false|false||antibiotics
null|Antibiotics, ophthalmologic|Drug|false|false||antibiotics
null|Antibiotics, Gynecological|Drug|false|false||antibiotics
null|antibiotics, intestinal|Drug|false|false||antibiotics
null|Antibiotic throat preparations|Drug|false|false||antibiotics
null|Antibiotics, Antitubercular|Drug|false|false||antibiotics
null|Antibiotics for systemic use|Drug|false|false||antibiotics
null|Antifungal Antibiotics, Topical|Drug|false|false||antibioticsnull|cefepime|Drug|false|false||cefepime
null|cefepime|Drug|false|false||cefepimenull|null|Time|false|false||priornull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Culture (Anthropological)|Finding|false|false||culturesnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Lung consolidation|Disorder|true|false||consolidationnull|Consolidation|Modifier|false|false||consolidationnull|Imaging problem|Finding|false|false||imagingnull|Diagnostic Imaging|Procedure|false|false||imaging
null|Imaging Techniques|Procedure|false|false||imagingnull|Imaging Technology|Title|false|false||imagingnull|Initial (abbreviation)|Finding|false|false||initialnull|Initially|Time|false|false||initialnull|Firstly|Modifier|false|false||initialnull|Systole|Finding|false|false||systolicnull|Respiratory, thoracic and mediastinal disorders|Disorder|false|false||Respnull|Respiratory rate|Attribute|false|false||Respnull|Spontaneous respiration|Finding|false|false||spontaneous respirationsnull|Respiration|Finding|false|false||respirationsnull|SAT1 protein, human|Drug|false|false||Sat
null|SAT1 protein, human|Drug|false|false||Satnull|College Entrance Examination Board Scholastic Aptitude Test|Finding|false|false||Sat
null|SAT1 wt Allele|Finding|false|false||Sat
null|SAT1 gene|Finding|false|false||Satnull|Santali language|Entity|false|false||Satnull|Initial (abbreviation)|Finding|false|false||Initialnull|Initially|Time|false|false||Initialnull|Firstly|Modifier|false|false||Initialnull|Laboratory test finding|Lab|false|false||labsnull|Hemopoietic stem cell transplant|Procedure|false|false||hct
null|Hematocrit Measurement|Procedure|false|false||hctnull|Leukocytes|Anatomy|false|false||wbcnull|creatinine|Drug|false|false||creatinine
null|creatinine|Drug|false|false||creatininenull|Creatinine metabolic function|Finding|false|false||creatininenull|Creatinine measurement|Procedure|false|false||creatininenull|Edo Language|Entity|false|false||BINnull|Bin|LabModifier|false|false||BINnull|lipase|Drug|false|false||lipase
null|lipase|Drug|false|false||lipase
null|lipase|Drug|false|false||lipasenull|Lipase measurement|Procedure|false|false||lipasenull|lactate|Drug|false|false||lactate
null|lactate|Drug|false|false||lactate
null|Lactates|Drug|false|false||lactatenull|Lactic acid measurement|Procedure|false|false||lactatenull|Plain chest X-ray|Procedure|false|false||cxrnull|Bilateral|Modifier|false|false||bilateralnull|Pleural Diseases|Disorder|false|false||pleuralnull|Pleura|Anatomy|false|false||pleuralnull|Pleural|Modifier|false|false||pleuralnull|effusion|Finding|false|false||effusionsnull|LARGE1 wt Allele|Finding|false|false||large
null|LARGE1 gene|Finding|false|false||largenull|Large|LabModifier|false|false||largenull|BRAF Gene Rearrangement|Disorder|false|false||positivenull|Rh Positive Blood Group|Finding|false|false||positive
null|Positive Finding|Finding|false|false||positive
null|Positive|Finding|false|false||positivenull|Positive Charge|Modifier|false|false||positivenull|Positive Number|LabModifier|false|false||positivenull|Nitrites|Drug|false|false||nitrites
null|Nitrites|Drug|false|false||nitrites
null|Nitrites|Drug|false|false||nitritesnull|Leukocytes|Anatomy|false|false||wbcnull|Respiratory Failure|Disorder|false|false||respiratory failurenull|Respiratory attachment|Finding|false|false||respiratory
null|respiratory|Finding|false|false||respiratory
null|null|Finding|false|false||respiratory
null|Respiratory specimen|Finding|false|false||respiratorynull|Respiratory rate|Attribute|false|false||respiratorynull|Failure (biologic function)|Finding|false|false||failure
null|Failure|Finding|false|false||failure
null|Personal failure|Finding|false|false||failurenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Intubated|Finding|false|false||intubatednull|Initial (abbreviation)|Finding|false|false||initialnull|Initially|Time|false|false||initialnull|Firstly|Modifier|false|false||initialnull|A1BG gene|Finding|false|false||ABGnull|Analysis of arterial blood gases and pH|Procedure|false|false||ABGnull|SLC35G1 gene|Finding|false|false||post
null|DESI1 gene|Finding|false|false||postnull|Post Device|Device|false|false||postnull|Post|Time|false|false||postnull|Intubation (procedure)|Procedure|false|false||intubationnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|vancomycin|Drug|false|false||vancomycin
null|vancomycin|Drug|false|false||vancomycinnull|Vancomycin measurement|Procedure|false|false||vancomycinnull|cefepime|Drug|false|false||cefepime
null|cefepime|Drug|false|false||cefepimenull|coverage - HL7PublishingDomain|Finding|false|false||coverage
null|null|Finding|false|false||coverage
null|coverage - financial contract|Finding|false|false||coveragenull|Urinary tract|Anatomy|false|false||urinarynull|urinary|Modifier|false|false||urinarynull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Source (property) (qualifier value)|Finding|false|false||source
null|Term Source|Finding|false|false||source
null|Source|Finding|false|false||sourcenull|Intubation (procedure)|Procedure|false|false||intubationnull|Levophed|Drug|false|false||levophed
null|Levophed|Drug|false|false||levophednull|phenylephrine|Drug|false|false||phenylephrine
null|phenylephrine|Drug|false|false||phenylephrinenull|Peripherally inserted central catheter (physical object)|Device|false|false||PICC linenull|Peripherally Inserted Central Catheter Line Insertion|Procedure|false|false||PICCnull|Peripherally inserted central catheter (physical object)|Device|false|false||PICCnull|Line Specimen|Drug|false|false||line
null|Long Interspersed Elements|Drug|false|false||line
null|Long Interspersed Elements|Drug|false|false||linenull|line source specimen code|Finding|false|false||linenull|Intravascular line|Device|false|false||linenull|Linear|Modifier|false|false||linenull|Line Unit of Length|LabModifier|false|false||linenull|Changing|Finding|false|false||alterednull|Mental state|Finding|false|false||mental statusnull|null|Attribute|false|false||mental status
null|null|Attribute|false|false||mental statusnull|Psyche structure|Finding|false|false||mentalnull|What subject filter - Status|Finding|false|false||statusnull|null|Attribute|false|false||statusnull|Social status|Modifier|false|false||status
null|Status|Modifier|false|false||statusnull|arrival - ActRelationshipType|Finding|false|false||arrivalnull|null|Event|false|false||arrivalnull|CAT scan of head|Procedure|false|false||head CTnull|Problems with head|Disorder|false|false||headnull|Procedure on head|Procedure|false|false||headnull|Structure of head of caudate nucleus|Anatomy|false|false||head
null|Head|Anatomy|false|false||headnull|Head Device|Device|false|false||headnull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|findings aspects|Finding|false|false||findingsnull|null|Attribute|false|false||findingsnull|Transfer - product ownership|Finding|false|false||transfer
null|Transfer Technique|Finding|false|false||transfer
null|ActClass - transfer|Finding|false|false||transfer
null|null|Finding|false|false||transfernull|Transfer (immobility management)|Procedure|false|false||transfernull|Settings (qualitative concept)|Modifier|false|false||settingsnull|Fraction of inspired oxygen|Finding|false|false||fio2null|fraction of inspired oxygen (FiO2) (treatment)|Procedure|false|false||fio2
null|Inspired Oxygen Fraction Test|Procedure|false|false||fio2null|null|Attribute|false|false||fio2null|Positive end expiratory pressure (finding)|Finding|false|false||peepnull|Positive End-Expiratory Pressure|Procedure|false|false||peepnull|Sedation|Finding|false|false||Sedation
null|Sedated state|Finding|false|false||Sedationnull|Sedation procedure|Procedure|false|false||Sedationnull|midazolam|Drug|false|false||midazolam
null|midazolam|Drug|false|false||midazolamnull|fentanyl|Drug|false|false||fentanyl
null|fentanyl|Drug|false|false||fentanylnull|Fentanyl measurement|Procedure|false|false||fentanylnull|Levophed|Drug|false|false||levophed
null|Levophed|Drug|false|false||levophednull|Living Alone|Finding|false|false||alonenull|alone - group size|Subject|false|false||alonenull|Singular|LabModifier|false|false||alonenull|Microtubule-Associated Proteins|Drug|false|false||MAPs
null|Microtubule-Associated Proteins|Drug|false|false||MAPsnull|C3orf62 gene|Finding|false|false||MAPs
null|Map|Finding|false|false||MAPsnull|arrival - ActRelationshipType|Finding|false|false||arrivalnull|null|Event|false|false||arrivalnull|Fraction of inspired oxygen|Finding|false|false||FiO2null|fraction of inspired oxygen (FiO2) (treatment)|Procedure|false|false||FiO2
null|Inspired Oxygen Fraction Test|Procedure|false|false||FiO2null|null|Attribute|false|false||FiO2null|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Levophed|Drug|false|false||levophed
null|Levophed|Drug|false|false||levophednull|Sedated state|Finding|false|false||sedatednull|Confusional Arousals|Disorder|false|false||unresponsivenull|Unresponsive to Treatment|Finding|false|false||unresponsive
null|unresponsive behavior|Finding|false|false||unresponsivenull|Participation Mode - verbal|Finding|false|false||verbalnull|Consent Mode - Verbal|Procedure|false|false||verbalnull|Verbal|Modifier|false|false||verbalnull|Pain|Finding|false|false||painfulnull|Stimulus|Phenomenon|false|false||stimulinull|Thought|Finding|false|false||thought
null|null|Finding|false|false||thoughtnull|Behavior Rating Inventory of Executive Function|Finding|false|false||brief
null|BRIEF Health Literacy Screening Tool|Finding|false|false||briefnull|Brief|Time|false|false||briefnull|Shortened|Modifier|false|false||briefnull|Episode of|Time|false|false||episode ofnull|Episode of|Time|false|false||episodenull|Decerebrate Posturing|Finding|false|false||decerebrate posturing
null|Decerebrate State|Finding|false|false||decerebrate posturingnull|Posturing|Disorder|false|false||posturingnull|Upper Extremity|Anatomy|false|false||upper extremitiesnull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|All extremities|Anatomy|false|false||extremities
null|Limb structure|Anatomy|false|false||extremitiesnull|Review of systems (procedure)|Procedure|false|false||Review of systemsnull|null|Attribute|false|false||Review of systems
null|null|Attribute|false|false||Review of systemsnull|Review of|Finding|false|false||Review ofnull|Review (Publication Type)|Finding|false|false||Review
null|Act Class - review|Finding|false|false||Reviewnull|System|Finding|false|false||systemsnull|Unable|Finding|false|false||Unablenull|Obtain|Finding|false|false||Obtainnull|Acquisition (action)|Event|false|false||Obtainnull|Anemia|Disorder|false|false||Anemianull|Anemia <Anemiaceae>|Entity|false|false||Anemianull|borderline cholesterol|Lab|false|false||Borderline cholesterolnull|Borderline|Modifier|false|false||Borderlinenull|cholesterol|Drug|false|false||cholesterol
null|cholesterol|Drug|false|false||cholesterolnull|Cholesterol measurement|Procedure|false|false||cholesterolnull|Recurrent|Time|false|false||Recurrent
null|Episodic|Time|false|false||Recurrentnull|Flatulence|Finding|false|false||Flatulencenull|Heart murmur|Finding|false|false||Heart Murmurnull|Malignant neoplasm of heart|Disorder|false|false||Heart
null|benign neoplasm of heart|Disorder|false|false||Heartnull|HEART PROBLEM|Finding|false|false||Heartnull|Chest>Heart|Anatomy|false|false||Heart
null|Heart|Anatomy|false|false||Heartnull|Heart murmur|Finding|false|false||Murmurnull|Hypertensive disease|Disorder|false|false||Hypertensionnull|Hypothyroidism|Disorder|false|false||Hypothyroidismnull|Mitral Valve Insufficiency|Disorder|false|false||Mitral Regurgitationnull|mitral|Modifier|false|false||Mitralnull|Regurgitation|Finding|false|false||Regurgitation
null|Regurgitates after swallowing|Finding|false|false||Regurgitationnull|Regurgitation - mechanism|Phenomenon|false|false||Regurgitationnull|Osteoporosis|Disorder|false|false||Osteoporosisnull|Encounter due to family history of osteoporosis|Finding|false|false||Osteoporosisnull|Pneumonia|Disorder|false|false||Pneumonianull|Sinusitis|Disorder|false|false||Sinusitisnull|Long Variable|Modifier|false|false||Long
null|Long|Modifier|false|false||Longnull|null|Finding|false|false||history of hypertensionnull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Hypertensive disease|Disorder|false|false||hypertensionnull|ErbB Receptors|Drug|false|false||her family
null|ErbB Receptors|Drug|false|false||her familynull|ErbB Receptors|Finding|false|false||her familynull|Entity Name Part Type - family|Finding|false|false||family
null|Last Name|Finding|false|false||family
null|Living Arrangement - Family|Finding|false|false||family
null|Family (taxonomic)|Finding|false|false||family
null|Family Collection|Finding|false|false||familynull|Family|Subject|false|false||familynull|Indirect exposure mechanism - Father|Finding|false|false||Father
null|Relationship - Father|Finding|false|false||Father
null|Father - courtesy title|Finding|false|false||Fathernull|Father (person)|Subject|false|false||Fathernull|Entity Name Part Type - family|Finding|false|false||family
null|Last Name|Finding|false|false||family
null|Living Arrangement - Family|Finding|false|false||family
null|Family (taxonomic)|Finding|false|false||family
null|Family Collection|Finding|false|false||familynull|Family|Subject|false|false||familynull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Numerous|LabModifier|false|false||multiplenull|Malignant Neoplasms|Disorder|false|false||cancersnull|Grandfather|Subject|false|false||grandfathernull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Malignant neoplasm of stomach|Disorder|false|false||stomach cancer
null|Stomach Carcinoma|Disorder|false|false||stomach cancernull|Neoplasm of uncertain or unknown behavior of stomach|Disorder|false|false||stomach
null|Stomach Diseases|Disorder|false|false||stomach
null|Benign neoplasm of stomach|Disorder|false|false||stomach
null|Carcinoma in situ of stomach|Disorder|false|false||stomachnull|Stomach problem|Finding|false|false||stomachnull|Procedure on stomach|Procedure|false|false||stomachnull|Stomach structure|Anatomy|false|false||stomach
null|Abdomen>Stomach|Anatomy|false|false||stomach
null|Stomach|Anatomy|false|false||stomachnull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Uncle|Subject|false|false||unclenull|Medical History|Finding|false|true||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Throat Homeopathic Medication|Drug|false|true||throatnull|Specimen Type - Throat|Finding|false|true||throat
null|null|Finding|false|true||throatnull|Anterior portion of neck|Anatomy|false|false||throat
null|Throat|Anatomy|false|false||throat
null|Pharyngeal structure|Anatomy|false|false||throatnull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Medical History|Finding|true|false||history ofnull|History of present illness (finding)|Finding|true|false||history
null|History of previous events|Finding|true|false||history
null|Historical aspects qualifier|Finding|true|false||history
null|Medical History|Finding|true|false||history
null|Concept History|Finding|true|false||historynull|History|Subject|false|false||historynull|Malignant tumor of colon|Disorder|true|false||colon cancersnull|Neoplasm of uncertain or unknown behavior of colon|Disorder|true|false||colon
null|Colonic Diseases|Disorder|true|false||colon
null|Carcinoma in situ of colon|Disorder|true|false||colonnull|COLON PROBLEM|Finding|true|false||colonnull|Colon structure (body structure)|Anatomy|false|false||colon
null|Abdomen+Pelvis>Colon|Anatomy|false|false||colonnull|TUBE,COLON,22FR,RADIOPAQUE RUBBER B#7370|Device|true|false||colonnull|Colon <Coloninae>|Entity|true|false||colonnull|Malignant Neoplasms|Disorder|true|false||cancersnull|Indirect exposure mechanism - Father|Finding|false|false||Father
null|Relationship - Father|Finding|false|false||Father
null|Father - courtesy title|Finding|false|false||Fathernull|Father (person)|Subject|false|false||Fathernull|Cerebrovascular accident|Disorder|false|false||strokenull|Stroke (heart beat)|Finding|false|false||strokenull|Entity Name Part Type - family|Finding|false|false||family
null|Last Name|Finding|false|false||family
null|Living Arrangement - Family|Finding|false|false||family
null|Family (taxonomic)|Finding|false|false||family
null|Family Collection|Finding|false|false||familynull|Family|Subject|false|false||familynull|Relationship - Mother|Finding|false|false||Mothernull|Mother (person)|Subject|false|false||Mothernull|null|Anatomy|false|false||heart valve
null|Heart Valves|Anatomy|false|false||heart valvenull|Malignant neoplasm of heart|Disorder|false|false||heart
null|benign neoplasm of heart|Disorder|false|false||heartnull|HEART PROBLEM|Finding|false|false||heartnull|Chest>Heart|Anatomy|false|false||heart
null|Heart|Anatomy|false|false||heartnull|Anatomical valve|Anatomy|false|false||valvenull|Valve (physical object)|Device|false|false||valve
null|Valve Device|Device|false|false||valve
null|medical valve|Device|false|false||valvenull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|physical examination (physical finding)|Finding|false|false||PHYSICAL EXAMnull|Physical Examination|Procedure|false|false||PHYSICAL EXAMnull|physical examination (physical finding)|Finding|false|false||PHYSICAL
null|Physical|Finding|false|false||PHYSICALnull|Physical Examination|Procedure|false|false||PHYSICALnull|Exam|Finding|false|false||EXAMnull|Medical Examination|Procedure|false|false||EXAMnull|Fraction of inspired oxygen|Finding|false|false||FiO2null|fraction of inspired oxygen (FiO2) (treatment)|Procedure|false|false||FiO2
null|Inspired Oxygen Fraction Test|Procedure|false|false||FiO2null|null|Attribute|false|false||FiO2null|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||Generalnull|General medical service|Procedure|false|false||Generalnull|Generalized|Modifier|false|false||Generalnull|Intubated|Finding|false|false||Intubatednull|Confusional Arousals|Disorder|false|false||unresponsivenull|Unresponsive to Treatment|Finding|false|false||unresponsive
null|unresponsive behavior|Finding|false|false||unresponsivenull|Acute limbic encephalitis following transplant|Disorder|false|false||palenull|Body pale (finding)|Finding|false|false||pale
null|Pallor of skin|Finding|false|false||palenull|Pale color saturation|Modifier|false|false||pale
null|Pale color|Modifier|false|false||palenull|Very|Modifier|false|false||verynull|Thin (qualifier value)|Modifier|false|false||thinnull|HEENT|Anatomy|false|false||HEENTnull|Scleral Diseases|Disorder|false|false||Scleranull|examination of sclera|Procedure|false|false||Scleranull|Sclera|Anatomy|false|false||Scleranull|Anicteric|Finding|false|false||anictericnull|Myelofibrosis|Disorder|false|false||MMMnull|Medial part of medial mammillary nucleus|Anatomy|false|false||MMMnull|Oropharyngeal|Anatomy|false|false||oropharynxnull|Remote control command - Clear|Finding|false|false||clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|Pupil|Anatomy|false|false||pupilsnull|Constricting sensation quality|Finding|false|false||constrictednull|Sluggish|Finding|false|false||sluggishnull|Present|Finding|false|false||present
null|Presentation|Finding|false|false||presentnull|Passive joint movement of neck (finding)|Finding|false|false||Neck
null|Neck problem|Finding|false|false||Necknull|dendritic spine neck|Anatomy|false|false||Neck
null|Neck|Anatomy|false|false||Necknull|Supple|Finding|false|false||supplenull|Jugular venous pressure|Finding|false|false||JVPnull|Elevated|Modifier|false|false||elevated
null|High|Modifier|false|false||elevatednull|Leukocyte adhesion deficiency type 1|Disorder|true|false||LAD
null|Leukocyte adhesion deficiency|Disorder|true|false||LADnull|ITGB2 wt Allele|Finding|true|false||LAD
null|DLD gene|Finding|true|false||LADnull|Anterior descending branch of left coronary artery|Anatomy|true|false||LADnull|Ladino Language|Entity|true|false||LADnull|Regular|Modifier|false|false||Regularnull|Amount type - Rate|Finding|false|false||ratenull|Rating (action)|Event|false|false||ratenull|Rate|LabModifier|false|false||ratenull|Rhythm|Finding|false|false||rhythm
null|rhythmic process (biological)|Finding|false|false||rhythmnull|SYSTOLIC EJECTION MURMUR|Finding|false|false||SEMnull|Microscopes, Electron, Scanning|Device|false|false||SEMnull|Standard Error|LabModifier|false|false||SEMnull|Vitelliform Macular Dystrophy|Disorder|false|false||bestnull|BEST1 wt Allele|Finding|false|false||best
null|BEST1 gene|Finding|false|false||bestnull|best (quality)|Modifier|false|false||bestnull|midline catheter (treatment)|Procedure|false|false||midline catheternull|Midline catheter (device)|Device|false|false||midline catheternull|midline cell component|Anatomy|false|false||midlinenull|Midline (qualifier value)|Modifier|false|false||midlinenull|null|Finding|false|false||catheternull|catheter device|Device|false|false||catheter
null|XXX>Catheter|Device|false|false||catheternull|Present|Finding|false|false||present
null|Presentation|Finding|false|false||presentnull|Right arm|Anatomy|false|false||R armnull|Anorectal Malformations|Disorder|false|false||armnull|AKR1A1 wt Allele|Finding|false|false||arm
null|ARMC9 gene|Finding|false|false||armnull|Protocol Treatment Arm|Procedure|false|false||arm
null|Axillary Reverse Mapping|Procedure|false|false||arm
null|Study Arm|Procedure|false|false||armnull|Upper arm|Anatomy|false|false||arm
null|null|Anatomy|false|false||arm
null|Upper Extremity|Anatomy|false|false||armnull|Lung|Anatomy|false|false||Lungsnull|Bilateral|Modifier|false|false||Bilateralnull|Basilar Rales|Finding|false|false||crackles
null|Rales|Finding|false|false||cracklesnull|Spontaneous respiration|Finding|true|false||spontaneous respirationsnull|Spontaneous|Finding|true|false||spontaneousnull|Respiration|Finding|true|false||respirationsnull|Trophoblastic tumor, epithelioid|Disorder|false|false||ETTnull|Place - dosing instruction imperative|Finding|false|false||placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|Malignant neoplasm of abdomen|Disorder|false|false||Abdomennull|Abdomen problem|Finding|false|false||Abdomennull|Abdomen|Anatomy|false|false||Abdomen
null|Abdominal Cavity|Anatomy|false|false||Abdomennull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||softnull|Soft|Modifier|false|false||softnull|Bowel sounds|Finding|false|false||bowel soundsnull|Intestines|Anatomy|false|false||bowelnull|null|Device|false|false||soundsnull|null|Phenomenon|false|false||soundsnull|Present|Finding|false|false||present
null|Presentation|Finding|false|false||presentnull|Organomegaly|Finding|false|false||organomegalynull|Present|Finding|false|false||present
null|Presentation|Finding|false|false||presentnull|Candida|Entity|false|false||candidalnull|Eruption of skin (disorder)|Disorder|false|false||rashnull|Skin rash|Finding|false|false||rash
null|Eruptions|Finding|false|false||rash
null|Exanthema|Finding|false|false||rashnull|Pelvis>Groin|Anatomy|false|false||groin
null|Inguinal region|Anatomy|false|false||groin
null|Inguinal part of abdomen|Anatomy|false|false||groinnull|Academic Research Enhancement Awards|Event|false|false||areanull|Geographic Locations|Entity|false|false||areanull|Area|Modifier|false|false||areanull|powder physical state|Drug|false|false||powder
null|Powder dose form|Drug|false|false||powdernull|miconazole|Drug|false|false||miconazole
null|miconazole|Drug|false|false||miconazolenull|powder physical state|Drug|false|false||powder
null|Powder dose form|Drug|false|false||powdernull|Present|Finding|false|false||present
null|Presentation|Finding|false|false||presentnull|Distribution [PK]|Finding|false|false||distribution
null|Distribution|Finding|false|false||distributionnull|Spatial Distribution|Modifier|false|false||distributionnull|Hereditary Multiple Exostoses|Disorder|false|false||Extnull|EXT1 wt Allele|Finding|false|false||Ext
null|EXT1 gene|Finding|false|false||Extnull|Feels warm|Finding|false|false||warmnull|warming process|Phenomenon|false|false||warmnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false||pulsesnull|Clubbing|Disorder|true|false||clubbingnull|Cyanosis|Finding|true|false||cyanosisnull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Neurology speciality|Title|false|false||Neuronull|Neurologic (qualifier value)|Modifier|false|false||Neuronull|Unable|Finding|false|false||Unablenull|Unresponsiveness|Finding|false|false||unresponsivenessnull|Has patient|Finding|false|false||patient hasnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|All extremities|Anatomy|false|false||all extremitiesnull|All extremities|Anatomy|false|false||extremities
null|Limb structure|Anatomy|false|false||extremitiesnull|Decerebration procedure|Procedure|false|false||decerebrationnull|Upper Extremity|Anatomy|false|false||upper extremitiesnull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|All extremities|Anatomy|false|false||extremities
null|Limb structure|Anatomy|false|false||extremitiesnull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|physical examination (physical finding)|Finding|false|false||PHYSICAL EXAMnull|Physical Examination|Procedure|false|false||PHYSICAL EXAMnull|physical examination (physical finding)|Finding|false|false||PHYSICAL
null|Physical|Finding|false|false||PHYSICALnull|Physical Examination|Procedure|false|false||PHYSICALnull|Exam|Finding|false|false||EXAMnull|Medical Examination|Procedure|false|false||EXAMnull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|Laboratory test finding|Lab|false|false||LABSnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Creatine Kinase|Drug|false|false||CPK
null|Creatine Kinase|Drug|false|false||CPKnull|PIK3C2A gene|Finding|false|false||CPKnull|Creatine kinase measurement|Procedure|false|false||CPKnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|lipase|Drug|false|false||Lipase
null|lipase|Drug|false|false||Lipase
null|lipase|Drug|false|false||Lipasenull|Lipase measurement|Procedure|false|false||Lipasenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MB
null|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MBnull|creatine kinase activity|Finding|false|false||CK-MBnull|Serum creatine phosphokinase MB isoenzyme measurement|Procedure|false|false||CK-MB
null|Creatine kinase MB measurement|Procedure|false|false||CK-MBnull|MB-6|Drug|false|false||MB-6null|Blood calcium measurement|Procedure|false|false||BLOOD Calciumnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Iron Drug Class|Drug|false|false||Iron
null|iron|Drug|false|false||Iron
null|iron|Drug|false|false||Iron
null|iron|Drug|false|false||Iron
null|Ferrum metallicum, Homeopathic preparation|Drug|false|false||Ironnull|Iron measurement|Procedure|false|false||Ironnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|folate|Drug|false|false||Folate
null|folate|Drug|false|false||Folate
null|folate|Drug|false|false||Folatenull|Folic acid measurement|Procedure|false|false||Folatenull|Thyrotropin-Releasing Hormone, human|Drug|false|false||TRF
null|IL5 protein, human|Drug|false|false||TRF
null|IL5 protein, human|Drug|false|false||TRF
null|thyrotropin-releasing hormone|Drug|false|false||TRF
null|thyrotropin-releasing hormone|Drug|false|false||TRF
null|thyrotropin-releasing hormone|Drug|false|false||TRF
null|Tocotrienol-rich Fraction|Drug|false|false||TRF
null|Thyrotropin-Releasing Hormone, human|Drug|false|false||TRFnull|TERF1 wt Allele|Finding|false|false||TRF
null|TERF1 gene|Finding|false|false||TRF
null|IL5 gene|Finding|false|false||TRFnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Arylsulfatase A, human|Drug|false|false||ASA
null|Arylsulfatase A, human|Drug|false|false||ASA
null|aspirin|Drug|false|false||ASA
null|aspirin|Drug|false|false||ASAnull|ARSA gene|Finding|false|false||ASAnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|CNS depressants ethanol|Drug|false|false||Ethanol
null|CNS depressants ethanol|Drug|false|false||Ethanol
null|antiseptics ethanol|Drug|false|false||Ethanol
null|antiseptics ethanol|Drug|false|false||Ethanol
null|ethanol|Drug|false|false||Ethanol
null|ethanol|Drug|false|false||Ethanolnull|Toxic effect of ethyl alcohol|Disorder|false|false||Ethanolnull|Ethanol measurement|Procedure|false|false||Ethanolnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Partial pressure of Oxygen|Finding|false|false||pO2
null|US Military enlisted E5|Finding|false|false||pO2null|PO2 measurement|Procedure|false|false||pO2null|Carbon dioxide measurement, partial pressure|Procedure|false|false||pCO2null|Carbon dioxide, partial pressure|Lab|false|false||pCO2null|nitrogenous base|Drug|false|false||Base
null|Base|Drug|false|false||Base
null|Dental Base|Drug|false|false||Base
null|base - RoleClass|Drug|false|false||Basenull|Base - General Qualifier|Finding|false|false||Base
null|BPIFA4P gene|Finding|false|false||Base
null|Base - RX Component Type|Finding|false|false||Basenull|Anatomical base|Anatomy|false|false||Basenull|Base - unit of product usage|LabModifier|false|false||Basenull|Published Comment|Finding|false|false||Comment
null|Comment|Finding|false|false||Commentnull|Green color|Modifier|false|false||GREENnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|lactate|Drug|false|false||Lactate
null|lactate|Drug|false|false||Lactate
null|Lactates|Drug|false|false||Lactatenull|Lactic acid measurement|Procedure|false|false||Lactatenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|SAT1 protein, human|Drug|false|false||Sat
null|SAT1 protein, human|Drug|false|false||Satnull|College Entrance Examination Board Scholastic Aptitude Test|Finding|false|false||Sat
null|SAT1 wt Allele|Finding|false|false||Sat
null|SAT1 gene|Finding|false|false||Satnull|Santali language|Entity|false|false||Satnull|Color of urine|Finding|false|false||URINE Colornull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|color additive|Drug|false|false||Color
null|Coloring Excipient|Drug|false|false||Colornull|color - solid dosage form|Modifier|false|false||Color
null|Color|Modifier|false|false||Colornull|Color quantity|LabModifier|false|false||Colornull|Yellow color|Modifier|false|false||Yellownull|Cloudy|Modifier|false|false||Hazynull|Mandibular right first molar mesial prosthesis|Device|false|false||30PMnull|Hematuria|Disorder|false|false||URINE Bloodnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Blood and lymphatic system disorders|Disorder|false|false||Bloodnull|peripheral blood|Finding|false|false||Blood
null|Blood|Finding|false|false||Blood
null|In Blood|Finding|false|false||Bloodnull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||MODnull|nitrite ion|Drug|false|false||Nitrite
null|Nitrites|Drug|false|false||Nitrite
null|Nitrites|Drug|false|false||Nitrite
null|Nitrites|Drug|false|false||Nitrite
null|nitrite ion|Drug|false|false||Nitrite
null|nitrite ion|Drug|false|false||Nitritenull|Health Maintenance Organization Point of Service Plan|Finding|false|false||POSnull|Structure of parieto-occipital fissure|Anatomy|false|false||POSnull|Point-of-service (POS) plan|Entity|false|false||POS
null|Local - Managed care POS|Entity|false|false||POSnull|Proteins|Drug|false|false||Protein
null|Proteins|Drug|false|false||Proteinnull|Protein Info|Finding|false|false||Proteinnull|Protein measurement|Procedure|false|false||Proteinnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Ketones|Drug|false|false||Ketonenull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Mandibular right first molar mesial prosthesis|Device|false|false||30PMnull|null|Lab|false|false||URINE RBC
null|Red blood cells urine positive|Lab|false|false||URINE RBCnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Leukocytes|Anatomy|false|false||WBCnull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||MODnull|Yeast, Dried|Drug|false|false||Yeast
null|Candida albicans allergenic extract|Drug|false|false||Yeast
null|Candida albicans allergenic extract|Drug|false|false||Yeast
null|Candida albicans allergenic extract|Drug|false|false||Yeastnull|Saccharomyces cerevisiae|Entity|false|false||Yeast
null|Yeasts|Entity|false|false||Yeastnull|Tissue Factor Pathway Inhibitor, human|Drug|false|false||Epi
null|epinephrine|Drug|false|false||Epi
null|epinephrine|Drug|false|false||Epi
null|epinephrine|Drug|false|false||Epi
null|Tissue Factor Pathway Inhibitor, human|Drug|false|false||Epinull|Exocrine pancreatic insufficiency|Disorder|false|false||Epinull|Eysenck personality inventory|Finding|false|false||Epi
null|TFPI wt Allele|Finding|false|false||Epi
null|TFPI gene|Finding|false|false||Epinull|Electronic Portal Imaging|Procedure|false|false||Epi
null|Echo-Planar Imaging|Procedure|false|false||Epinull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Mandibular right first molar mesial prosthesis|Device|false|false||30PMnull|Mucus in urine (finding)|Finding|false|false||URINE Mucousnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Mucus (substance)|Finding|false|false||Mucous
null|mucus layer|Finding|false|false||Mucousnull|Mucous appearance|Modifier|false|false||Mucousnull|Retinoic Acid Response Element|Finding|false|false||RAREnull|Infrequent|Time|false|false||RAREnull|Rare|Modifier|false|false||RAREnull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|Laboratory test finding|Lab|false|false||LABSnull|Microbiology Diagnostic Service Section ID|Finding|false|false||MICROBIOLOGY
null|Microbiological|Finding|false|false||MICROBIOLOGY
null|Microbiology - Laboratory Class|Finding|false|false||MICROBIOLOGYnull|Microbiology procedure|Procedure|false|false||MICROBIOLOGYnull|Science of Microbiology|Title|false|false||MICROBIOLOGYnull|Urine culture|Procedure|false|false||Urine culturenull|Portion of urine|Finding|false|false||Urine
null|null|Finding|false|false||Urine
null|Urine|Finding|false|false||Urine
null|In Urine|Finding|false|false||Urine
null|Urine specimen|Finding|false|false||Urinenull|Culture Dose Form|Drug|false|false||culturenull|Culture (Anthropological)|Finding|false|false||culture
null|Cultural aspects|Finding|false|false||culturenull|Microbial culture (procedure)|Procedure|false|false||culture
null|Laboratory culture|Procedure|false|false||culturenull|Pseudomonas aeruginosa infection|Disorder|false|false||PSEUDOMONAS AERUGINOSAnull|Pseudomonas aeruginosa|Entity|false|false||PSEUDOMONAS AERUGINOSAnull|Pseudomonas Infections|Disorder|false|false||PSEUDOMONASnull|Pseudomonas|Entity|false|false||PSEUDOMONASnull|organisms/mL|LabModifier|false|false||ORGANISMS/MLnull|Organism|Entity|false|false||ORGANISMSnull|per milliliter|LabModifier|false|false||/MLnull|Antimicrobial susceptibility|Finding|false|false||SENSITIVITIESnull|methyl isocyanate|Drug|false|false||MIC
null|methyl isocyanate|Drug|false|false||MICnull|Ductal Carcinoma In Situ with Microinvasion|Disorder|false|false||MICnull|cisplatin/ifosfamide/mitomycin protocol|Procedure|false|false||MIC
null|Minimum Inhibitory Concentration Test|Procedure|false|false||MICnull|Micmac language|Entity|false|false||MICnull|Microgram per Milliliter|LabModifier|false|false||MCG/MLnull|microgram|LabModifier|false|false||MCGnull|per milliliter|LabModifier|false|false||/MLnull|amikacin|Drug|false|false||AMIKACIN
null|amikacin|Drug|false|false||AMIKACINnull|Amikacin measurement|Procedure|false|false||AMIKACINnull|cefepime|Drug|false|false||CEFEPIME
null|cefepime|Drug|false|false||CEFEPIMEnull|ceftazidime|Drug|false|false||CEFTAZIDIME
null|ceftazidime|Drug|false|false||CEFTAZIDIMEnull|ciprofloxacin|Drug|false|false||CIPROFLOXACIN
null|ciprofloxacin|Drug|false|false||CIPROFLOXACINnull|gentamicin|Drug|false|false||GENTAMICIN
null|gentamicin|Drug|false|false||GENTAMICINnull|Gentamicin measurement|Procedure|false|false||GENTAMICINnull|INJECTION, MEROPENEM, 100 MG ADMINISTERED|Drug|false|false||MEROPENEM
null|meropenem|Drug|false|false||MEROPENEM
null|meropenem|Drug|false|false||MEROPENEMnull|piperacillin|Drug|false|false||PIPERACILLIN
null|piperacillin|Drug|false|false||PIPERACILLINnull|tazobactam|Drug|false|false||TAZO
null|tazobactam|Drug|false|false||TAZOnull|tobramycin|Drug|false|false||TOBRAMYCIN
null|tobramycin|Drug|false|false||TOBRAMYCINnull|Tobramycin measurement|Procedure|false|false||TOBRAMYCINnull|Blood culture|Procedure|false|false||Blood culturenull|Blood and lymphatic system disorders|Disorder|false|false||Bloodnull|peripheral blood|Finding|false|false||Blood
null|Blood|Finding|false|false||Blood
null|In Blood|Finding|false|false||Bloodnull|Culture Dose Form|Drug|false|false||culturenull|Culture (Anthropological)|Finding|false|false||culture
null|Cultural aspects|Finding|false|false||culturenull|Microbial culture (procedure)|Procedure|false|false||culture
null|Laboratory culture|Procedure|false|false||culturenull|Lactobacillus species|Entity|false|false||LACTOBACILLUS SPECIES
null|Lactobacillus|Entity|false|false||LACTOBACILLUS SPECIESnull|Lactobacillus|Entity|false|false||LACTOBACILLUSnull|Species - Nature of Abnormal Testing|Finding|false|false||SPECIES
null|Species|Finding|false|false||SPECIESnull|SET protein, human|Drug|false|false||set
null|SET protein, human|Drug|false|false||setnull|Parameterized Data Type - Set|Finding|false|false||set
null|Set scale|Finding|false|false||set
null|Set (Psychology)|Finding|false|false||set
null|SET gene|Finding|false|false||set
null|set (group)|Finding|false|false||setnull|Act Relationship Subset - previous|Time|false|false||previous
null|Previous|Time|false|false||previousnull|day|Time|false|false||daysnull|Antimicrobial susceptibility|Finding|false|false||SENSITIVITIESnull|methyl isocyanate|Drug|false|false||MIC
null|methyl isocyanate|Drug|false|false||MICnull|Ductal Carcinoma In Situ with Microinvasion|Disorder|false|false||MICnull|cisplatin/ifosfamide/mitomycin protocol|Procedure|false|false||MIC
null|Minimum Inhibitory Concentration Test|Procedure|false|false||MICnull|Micmac language|Entity|false|false||MICnull|Microgram per Milliliter|LabModifier|false|false||MCG/MLnull|microgram|LabModifier|false|false||MCGnull|per milliliter|LabModifier|false|false||/MLnull|ampicillin|Drug|false|false||AMPICILLIN
null|ampicillins|Drug|false|false||AMPICILLIN
null|ampicillins|Drug|false|false||AMPICILLIN
null|ampicillin|Drug|false|false||AMPICILLINnull|gentamicin|Drug|false|false||GENTAMICIN
null|gentamicin|Drug|false|false||GENTAMICINnull|Gentamicin measurement|Procedure|false|false||GENTAMICINnull|penicillin G|Drug|false|false||PENICILLIN G
null|penicillin G|Drug|false|false||PENICILLIN Gnull|penicillins|Drug|false|false||PENICILLIN
null|penicillins|Drug|false|false||PENICILLINnull|Microbial culture of sputum|Procedure|false|false||Sputum culturenull|Specimen Type - Sputum|Finding|false|false||Sputum
null|null|Finding|false|false||Sputum
null|Sputum|Finding|false|false||Sputumnull|Culture Dose Form|Drug|false|false||culturenull|Culture (Anthropological)|Finding|false|false||culture
null|Cultural aspects|Finding|false|false||culturenull|Microbial culture (procedure)|Procedure|false|false||culture
null|Laboratory culture|Procedure|false|false||culturenull|endotracheal|Modifier|false|false||endotrachealnull|Source (property) (qualifier value)|Finding|false|false||source
null|Term Source|Finding|false|false||source
null|Source|Finding|false|false||sourcenull|Gram's stain|Drug|false|false||GRAM STAIN
null|Gram's stain|Drug|false|false||GRAM STAINnull|Bacterial stain, routine|Procedure|false|false||GRAM STAINnull|gram|LabModifier|false|false||GRAMnull|Stains|Drug|false|false||STAINnull|Staining method|Procedure|false|false||STAINnull|Epithelial Cells|Anatomy|false|false||epithelial cellsnull|Epithelial|Modifier|false|false||epithelialnull|Cells|Anatomy|false|false||cellsnull|Per 100x Field|LabModifier|false|false||/100X fieldnull|Knowledge Field|Finding|false|false||field
null|Force Field|Finding|false|false||field
null|Field|Finding|false|false||fieldnull|field - patient encounter|Procedure|false|false||fieldnull|Knowledge Field|Finding|false|false||FIELD
null|Force Field|Finding|false|false||FIELD
null|Field|Finding|false|false||FIELDnull|field - patient encounter|Procedure|false|false||FIELDnull|Saccharomycetales|Entity|false|false||BUDDING YEASTnull|Cell budding|Finding|false|false||BUDDINGnull|Yeast, Dried|Drug|false|false||YEAST
null|Candida albicans allergenic extract|Drug|false|false||YEAST
null|Candida albicans allergenic extract|Drug|false|false||YEAST
null|Candida albicans allergenic extract|Drug|false|false||YEASTnull|Saccharomyces cerevisiae|Entity|false|false||YEAST
null|Yeasts|Entity|false|false||YEASTnull|pseudohyphae|Entity|false|false||PSEUDOHYPHAEnull|Knowledge Field|Finding|false|false||FIELD
null|Force Field|Finding|false|false||FIELD
null|Field|Finding|false|false||FIELDnull|field - patient encounter|Procedure|false|false||FIELDnull|Gram-Positive Cocci|Entity|false|false||GRAM POSITIVE COCCInull|gram|LabModifier|false|false||GRAMnull|BRAF Gene Rearrangement|Disorder|false|false||POSITIVEnull|Rh Positive Blood Group|Finding|false|false||POSITIVE
null|Positive Finding|Finding|false|false||POSITIVE
null|Positive|Finding|false|false||POSITIVEnull|Positive Charge|Modifier|false|false||POSITIVEnull|Positive Number|LabModifier|false|false||POSITIVEnull|Cocci bacteria|Entity|false|false||COCCInull|Respiratory culture|Procedure|false|false||RESPIRATORY CULTUREnull|Respiratory attachment|Finding|false|false||RESPIRATORY
null|respiratory|Finding|false|false||RESPIRATORY
null|null|Finding|false|false||RESPIRATORY
null|Respiratory specimen|Finding|false|false||RESPIRATORYnull|Respiratory rate|Attribute|false|false||RESPIRATORYnull|Culture Dose Form|Drug|false|false||CULTUREnull|Culture (Anthropological)|Finding|false|false||CULTURE
null|Cultural aspects|Finding|false|false||CULTUREnull|Microbial culture (procedure)|Procedure|false|false||CULTURE
null|Laboratory culture|Procedure|false|false||CULTUREnull|Diagnosis Type - Final|Finding|false|false||Finalnull|Final|Time|false|false||Finalnull|End-stage|Modifier|false|false||Finalnull|Moderate growth|Modifier|false|false||MODERATE GROWTHnull|Moderate - Severity of Illness Code|Finding|false|false||MODERATE
null|Moderate|Finding|false|false||MODERATEnull|Moderate (severity modifier)|Modifier|false|false||MODERATE
null|Moderate - Allergy Severity|Modifier|false|false||MODERATE
null|Moderation|Modifier|false|false||MODERATEnull|Growth & development aspects|Finding|false|false||GROWTH
null|Tissue Growth|Finding|false|false||GROWTH
null|Growth|Finding|false|false||GROWTH
null|growth aspects|Finding|false|false||GROWTHnull|Growth action|Phenomenon|false|false||GROWTHnull|Symbiotic|Finding|false|false||Commensalnull|Commensal parasite|Entity|false|false||Commensalnull|Pharyngeal/Respiratory Flora|Entity|false|false||Respiratory Floranull|Respiratory attachment|Finding|false|false||Respiratory
null|respiratory|Finding|false|false||Respiratory
null|null|Finding|false|false||Respiratory
null|Respiratory specimen|Finding|false|false||Respiratorynull|Respiratory rate|Attribute|false|false||Respiratorynull|Yeast, Dried|Drug|false|false||YEAST
null|Candida albicans allergenic extract|Drug|false|false||YEAST
null|Candida albicans allergenic extract|Drug|false|false||YEAST
null|Candida albicans allergenic extract|Drug|false|false||YEASTnull|Saccharomyces cerevisiae|Entity|false|false||YEAST
null|Yeasts|Entity|false|false||YEASTnull|Growth & development aspects|Finding|false|false||GROWTH
null|Tissue Growth|Finding|false|false||GROWTH
null|Growth|Finding|false|false||GROWTH
null|growth aspects|Finding|false|false||GROWTHnull|Growth action|Phenomenon|false|false||GROWTHnull|Legionella culture|Procedure|false|false||LEGIONELLA CULTUREnull|Legionella|Entity|false|false||LEGIONELLAnull|Culture Dose Form|Drug|false|false||CULTUREnull|Culture (Anthropological)|Finding|false|false||CULTURE
null|Cultural aspects|Finding|false|false||CULTUREnull|Microbial culture (procedure)|Procedure|false|false||CULTURE
null|Laboratory culture|Procedure|false|false||CULTUREnull|Preliminary|Time|false|false||Preliminarynull|Legionella|Entity|true|false||LEGIONELLAnull|Urine culture|Procedure|false|false||Urine culturenull|Portion of urine|Finding|false|false||Urine
null|null|Finding|false|false||Urine
null|Urine|Finding|false|false||Urine
null|In Urine|Finding|false|false||Urine
null|Urine specimen|Finding|false|false||Urinenull|Culture Dose Form|Drug|false|false||culturenull|Culture (Anthropological)|Finding|false|false||culture
null|Cultural aspects|Finding|false|false||culturenull|Microbial culture (procedure)|Procedure|false|false||culture
null|Laboratory culture|Procedure|false|false||culturenull|Yeast, Dried|Drug|false|false||YEAST
null|Candida albicans allergenic extract|Drug|false|false||YEAST
null|Candida albicans allergenic extract|Drug|false|false||YEAST
null|Candida albicans allergenic extract|Drug|false|false||YEASTnull|Saccharomyces cerevisiae|Entity|false|false||YEAST
null|Yeasts|Entity|false|false||YEASTnull|organisms/mL|LabModifier|false|false||ORGANISMS/MLnull|Organism|Entity|false|false||ORGANISMSnull|per milliliter|LabModifier|false|false||/MLnull|Blood culture|Procedure|false|false||Blood culturenull|Blood and lymphatic system disorders|Disorder|false|false||Bloodnull|peripheral blood|Finding|false|false||Blood
null|Blood|Finding|false|false||Blood
null|In Blood|Finding|false|false||Bloodnull|Culture Dose Form|Drug|false|false||culturenull|Culture (Anthropological)|Finding|false|false||culture
null|Cultural aspects|Finding|false|false||culturenull|Microbial culture (procedure)|Procedure|false|false||culture
null|Laboratory culture|Procedure|false|false||culturenull|Diagnosis Type - Final|Finding|false|false||finalnull|Final|Time|false|false||finalnull|End-stage|Modifier|false|false||finalnull|Rh Negative Blood Group|Finding|false|false||NEGATIVE
null|Negative|Finding|false|false||NEGATIVE
null|Negative Finding|Finding|false|false||NEGATIVEnull|Expression Negative|Lab|false|false||NEGATIVEnull|Negative - qualifier|Modifier|false|false||NEGATIVE
null|Negative Charge|Modifier|false|false||NEGATIVEnull|Negative Number|LabModifier|false|false||NEGATIVEnull|Blood culture|Procedure|false|false||Blood culturenull|Blood and lymphatic system disorders|Disorder|false|false||Bloodnull|peripheral blood|Finding|false|false||Blood
null|Blood|Finding|false|false||Blood
null|In Blood|Finding|false|false||Bloodnull|Culture Dose Form|Drug|false|false||culturenull|Culture (Anthropological)|Finding|false|false||culture
null|Cultural aspects|Finding|false|false||culturenull|Microbial culture (procedure)|Procedure|false|false||culture
null|Laboratory culture|Procedure|false|false||culturenull|Diagnosis Type - Final|Finding|false|false||finalnull|Final|Time|false|false||finalnull|End-stage|Modifier|false|false||finalnull|Rh Negative Blood Group|Finding|false|false||NEGATIVE
null|Negative|Finding|false|false||NEGATIVE
null|Negative Finding|Finding|false|false||NEGATIVEnull|Expression Negative|Lab|false|false||NEGATIVEnull|Negative - qualifier|Modifier|false|false||NEGATIVE
null|Negative Charge|Modifier|false|false||NEGATIVEnull|Negative Number|LabModifier|false|false||NEGATIVEnull|Blood culture|Procedure|false|false||Blood culturenull|Blood and lymphatic system disorders|Disorder|false|false||Bloodnull|peripheral blood|Finding|false|false||Blood
null|Blood|Finding|false|false||Blood
null|In Blood|Finding|false|false||Bloodnull|Culture Dose Form|Drug|false|false||culturenull|Culture (Anthropological)|Finding|false|false||culture
null|Cultural aspects|Finding|false|false||culturenull|Microbial culture (procedure)|Procedure|false|false||culture
null|Laboratory culture|Procedure|false|false||culturenull|Pending - Allergy Clinical Status|Finding|false|false||pending
null|Pending - referral status|Finding|false|false||pendingnull|Pending - status|Time|false|false||pendingnull|pending - ManagedParticipationStatus|Modifier|false|false||pending
null|pending - RoleStatus|Modifier|false|false||pending
null|Pending - Day type|Modifier|false|false||pendingnull|Growth & development aspects|Finding|true|false||GROWTH
null|Tissue Growth|Finding|true|false||GROWTH
null|Growth|Finding|true|false||GROWTH
null|growth aspects|Finding|true|false||GROWTHnull|Growth action|Phenomenon|true|false||GROWTHnull|Plain chest X-ray|Procedure|false|false||CHEST X-RAYnull|Chest problem|Finding|false|false||CHESTnull|Chest|Anatomy|false|false||CHEST
null|Anterior thoracic region|Anatomy|false|false||CHESTnull|ActClaimAttachmentCategoryCode - x-ray|Finding|false|false||X-RAY
null|roentgenographic|Finding|false|false||X-RAYnull|Plain x-ray|Procedure|false|false||X-RAY
null|Diagnostic radiologic examination|Procedure|false|false||X-RAY
null|Radiographic imaging procedure|Procedure|false|false||X-RAYnull|Roentgen Rays|Phenomenon|false|false||X-RAYnull|Bilateral pleural effusion|Disorder|false|false||Bilateral pleural effusionnull|Bilateral|Modifier|false|false||Bilateralnull|Pleural effusion (disorder)|Finding|false|false||pleural effusion
null|Pleural effusion fluid|Finding|false|false||pleural effusion
null|null|Finding|false|false||pleural effusionnull|Pleural Diseases|Disorder|false|false||pleuralnull|Pleura|Anatomy|false|false||pleuralnull|Pleural|Modifier|false|false||pleuralnull|Effusion (substance)|Finding|false|false||effusion
null|null|Finding|false|false||effusion
null|effusion|Finding|false|false||effusionnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Greater Than|LabModifier|false|false||greater thannull|Greater|LabModifier|false|false||greaternull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Underlying|Finding|false|false||Underlyingnull|Lung consolidation|Disorder|false|false||consolidationnull|Consolidation|Modifier|false|false||consolidationnull|Completely - dosing instruction fragment|Finding|false|false||completelynull|Complete|Modifier|false|false||completelynull|Endotracheal tube|Device|false|false||Endotracheal tubenull|endotracheal|Modifier|false|false||Endotrachealnull|Unspecified tube|Finding|false|false||tube
null|TUBE1 gene|Finding|false|false||tubenull|biomedical tube device|Device|false|false||tube
null|Packaging Tube|Device|false|false||tubenull|tube|Modifier|false|false||tubenull|Tube (unit of presentation)|LabModifier|false|false||tube
null|Tube Dosing Unit|LabModifier|false|false||tubenull|Structure of carina|Anatomy|false|false||carina
null|Keel structure|Anatomy|false|false||carinanull|Recommendation|Finding|false|false||Recommendnull|Repositioning (procedure)|Procedure|false|false||repositioningnull|Unspecified tube|Finding|false|false||tube
null|TUBE1 gene|Finding|false|false||tubenull|biomedical tube device|Device|false|false||tube
null|Packaging Tube|Device|false|false||tubenull|tube|Modifier|false|false||tubenull|Tube (unit of presentation)|LabModifier|false|false||tube
null|Tube Dosing Unit|LabModifier|false|false||tubenull|Neoplasm of uncertain or unknown behavior of stomach|Disorder|false|false||stomach
null|Stomach Diseases|Disorder|false|false||stomach
null|Benign neoplasm of stomach|Disorder|false|false||stomach
null|Carcinoma in situ of stomach|Disorder|false|false||stomachnull|Stomach problem|Finding|false|false||stomachnull|Procedure on stomach|Procedure|false|false||stomachnull|Stomach structure|Anatomy|false|false||stomach
null|Abdomen>Stomach|Anatomy|false|false||stomach
null|Stomach|Anatomy|false|false||stomachnull|Distal Resection Margin|Attribute|false|false||distalnull|Distal (qualifier value)|Modifier|false|false||distalnull|Carcinoma in situ of esophagus|Disorder|false|false||esophagus
null|Esophageal Diseases|Disorder|false|false||esophagus
null|Benign neoplasm of esophagus|Disorder|false|false||esophagusnull|Esophagus problem|Finding|false|false||esophagusnull|Procedures on the esophagus|Procedure|false|false||esophagusnull|Chest>Esophagus|Anatomy|false|false||esophagus
null|Esophagus|Anatomy|false|false||esophagusnull|Table Cell Horizontal Align - right|Finding|false|false||Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|Peripherally Inserted Central Catheter Line Insertion|Procedure|false|false||PICCnull|Peripherally inserted central catheter (physical object)|Device|false|false||PICCnull|Axilla|Anatomy|false|false||axillanull|CAT scan of head|Procedure|false|false||CT HEADnull|null|Attribute|false|false||CT HEADnull|Problems with head|Disorder|false|false||HEADnull|Procedure on head|Procedure|false|false||HEADnull|Structure of head of caudate nucleus|Anatomy|false|false||HEAD
null|Head|Anatomy|false|false||HEADnull|Head Device|Device|false|false||HEADnull|Contrast Media|Drug|true|false||CONTRASTnull|Contrast|Modifier|false|false||CONTRASTnull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Hemorrhage|Finding|false|false||hemorrhagenull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Infarction|Finding|false|false||infarctionnull|Mass Effect|Finding|false|false||mass effectnull|Mass of body structure|Finding|false|false||mass
null|Morphology, Attenuation, Size, and Structure Criteria|Finding|false|false||mass
null|null|Finding|false|false||mass
null|FBN1 wt Allele|Finding|false|false||mass
null|FBN1 gene|Finding|false|false||mass
null|Mass of body region|Finding|false|false||massnull|Mass, a measure of quantity of matter|LabModifier|false|false||mass
null|Molecular Mass|LabModifier|false|false||massnull|Effect, Appearance|Modifier|false|false||effect
null|Effect|Modifier|false|false||effectnull|Heart Ventricle|Anatomy|false|false||ventriclesnull|Prominent|Modifier|false|false||prominentnull|Glycation End Products, Advanced|Drug|false|false||age
null|Glycation End Products, Advanced|Drug|false|false||agenull|null|Attribute|false|false||agenull|Age|Subject|false|false||agenull|Relate - vinyl resin|Drug|false|false||relatednull|Role Link Type - related|Finding|false|false||related
null|Related (finding)|Finding|false|false||relatednull|Definitely Related to Intervention|Modifier|false|false||related
null|Relationships|Modifier|false|false||relatednull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|Atrophic|Finding|false|false||atrophynull|Periventricular white matter hypodensities|Finding|false|false||Periventricular white matter hypodensitiesnull|Periventricular white matter|Anatomy|false|false||Periventricular white matternull|Periventricular|Modifier|false|false||Periventricularnull|White matter|Anatomy|false|false||white matternull|White (population group)|Subject|false|false||white
null|Caucasian|Subject|false|false||white
null|Caucasians|Subject|false|false||whitenull|White color|Modifier|false|false||whitenull|Consistent with|Finding|false|false||compatible withnull|Compatible|Modifier|false|false||compatible withnull|Consistent with|Finding|false|false||compatiblenull|Compatible|Modifier|false|false||compatiblenull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Structure of small blood vessel (organ)|Anatomy|false|false||small vesselnull|Small|LabModifier|false|false||smallnull|Vessel Positions|Anatomy|false|false||vessel
null|Blood Vessel|Anatomy|false|false||vesselnull|Vessel (unit of presentation)|LabModifier|false|false||vesselnull|Ischemic|Finding|false|false||ischemicnull|Disease|Disorder|false|false||diseasenull|Basal|Modifier|false|false||Basalnull|Cistern|Anatomy|false|false||cisternsnull|Legal patent|Finding|false|false||patentnull|Open|Modifier|false|false||patentnull|Preservation Technique|Procedure|false|false||preservation
null|Biologic Preservation|Procedure|false|false||preservationnull|Gray color|Modifier|false|false||graynull|Gray unit of radiation dose|LabModifier|false|false||graynull|White (population group)|Subject|false|false||white
null|Caucasian|Subject|false|false||white
null|Caucasians|Subject|false|false||whitenull|White color|Modifier|false|false||whitenull|Cell Differentiation process|Finding|false|false||differentiation
null|Differentiation|Finding|false|false||differentiationnull|Cellular Differentiation Qualifier|Attribute|false|false||differentiationnull|Fracture|Disorder|true|false||fracturenull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Malignant neoplasm of nasal cavity|Disorder|false|false||nasal cavitynull|examination of nasal cavity|Procedure|false|false||nasal cavitynull|Nasal cavity|Anatomy|false|false||nasal cavitynull|Nasal brand of oxymetazoline|Drug|false|false||nasal
null|Nasal brand of oxymetazoline|Drug|false|false||nasal
null|Nasal dosage form|Drug|false|false||nasalnull|Nasal Route of Administration|Finding|false|false||nasal
null|Nasal (intended site)|Finding|false|false||nasalnull|null|Anatomy|false|false||nasalnull|Dental caries|Disorder|false|false||cavity
null|Cavitation|Disorder|false|false||cavitynull|Body cavities|Anatomy|false|false||cavitynull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Secondary to|Modifier|false|false||secondary tonull|Neoplasm Metastasis|Disorder|false|false||secondarynull|metastatic qualifier|Finding|false|false||secondarynull|Secondary to|Modifier|false|false||secondarynull|second (number)|LabModifier|false|false||secondarynull|Intubated|Finding|false|false||intubatednull|State|Finding|false|false||statenull|Geographic state|Entity|false|false||state
null|US State|Entity|false|false||statenull|atherosclerotic|Finding|false|false||Atheroscleroticnull|Mural|Modifier|false|false||muralnull|Pathologic calcification, calcified structure|Finding|false|false||calcifications
null|Physiologic calcification|Finding|false|false||calcificationsnull|Calcified (qualifier value)|Modifier|false|false||calcificationsnull|Code System Type - Internal|Modifier|false|false||internal
null|Internal Surface|Modifier|false|false||internal
null|Internal|Modifier|false|false||internalnull|Carotid Arteries|Anatomy|false|false||carotid arteries
null|Head+Neck>Carotid artery|Anatomy|false|false||carotid arteriesnull|Carotid Arteries|Anatomy|false|false||carotidnull|Procedure on artery|Procedure|false|false||arteriesnull|Arteries|Anatomy|false|false||arteries
null|Arterial system|Anatomy|false|false||arteriesnull|Present|Finding|false|false||present
null|Presentation|Finding|false|false||presentnull|Nasal sinus|Anatomy|false|false||paranasal sinusesnull|pathologic fistula|Disorder|false|false||sinusesnull|Head>Sinuses|Anatomy|false|false||sinuses
null|Nasal sinus|Anatomy|false|false||sinusesnull|Pneumatic mastoid cell|Anatomy|false|false||mastoid air cellsnull|examination of mastoid region|Procedure|false|false||mastoidnull|Mastoid process|Anatomy|false|false||mastoid
null|null|Anatomy|false|false||mastoid
null|Head>Mastoid|Anatomy|false|false||mastoidnull|Air (substance)|Drug|false|false||air
null|air|Drug|false|false||air
null|air|Drug|false|false||airnull|ACUTE INSULIN RESPONSE|Finding|false|false||air
null|AIRN gene|Finding|false|false||air
null|AI/RHEUM|Finding|false|false||airnull|Cells|Anatomy|false|false||cellsnull|Malignant neoplasm of middle ear|Disorder|false|false||middle ear
null|Disorder of middle ear|Disorder|false|false||middle earnull|examination of middle ear|Procedure|false|false||middle earnull|middle ear|Anatomy|false|false||middle earnull|Table Cell Vertical Align - middle|Finding|false|false||middlenull|Middle|Modifier|false|false||middle
null|Midline (qualifier value)|Modifier|false|false||middlenull|Ear and labyrinth disorders|Disorder|false|false||earnull|SpecimenType - Ear|Finding|false|false||ear
null|null|Finding|false|false||earnull|Ear structure|Anatomy|false|false||ear
null|null|Anatomy|false|false||earnull|Dental caries|Disorder|false|false||cavities
null|Cavitation|Disorder|false|false||cavitiesnull|Body cavities|Anatomy|false|false||cavitiesnull|Remote control command - Clear|Finding|false|false||clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|Bilateral|Modifier|false|false||Bilateralnull|Ocular (intended site)|Finding|false|false||ocular
null|Vision|Finding|false|false||ocular
null|Ocular (qualifier)|Finding|false|false||ocularnull|Orbital region|Anatomy|false|false||ocular
null|Eye|Anatomy|false|false||ocularnull|Lens Device|Device|false|false||lensesnull|impression (attitude)|Finding|false|false||IMPRESSION
null|EKG impression|Finding|false|false||IMPRESSIONnull|Intracranial Hemorrhage|Finding|false|false||intracranial hemorrhagenull|Intracranial Route of Administration|Finding|false|false||intracranialnull|Intracranial|Anatomy|false|false||intracranialnull|Hemorrhage|Finding|false|false||hemorrhagenull|Mass Effect|Finding|false|false||mass effectnull|Mass of body structure|Finding|false|false||mass
null|Morphology, Attenuation, Size, and Structure Criteria|Finding|false|false||mass
null|null|Finding|false|false||mass
null|FBN1 wt Allele|Finding|false|false||mass
null|FBN1 gene|Finding|false|false||mass
null|Mass of body region|Finding|false|false||massnull|Mass, a measure of quantity of matter|LabModifier|false|false||mass
null|Molecular Mass|LabModifier|false|false||massnull|Effect, Appearance|Modifier|false|false||effect
null|Effect|Modifier|false|false||effectnull|Transthoracic echocardiography|Procedure|false|false||TTEnull|Left atrial structure|Anatomy|false|false||left atriumnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Heart Atrium|Anatomy|false|false||atriumnull|size|Modifier|false|false||sizenull|size - solid dosage form|LabModifier|false|false||sizenull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Focal hypertrophy|Finding|false|false||focal hypertrophynull|Focal|Modifier|false|false||focalnull|Hypertrophy|Finding|false|false||hypertrophynull|Basal|Modifier|false|false||basalnull|Septum of telencephalon|Anatomy|false|false||septum
null|Cell septum|Anatomy|false|false||septum
null|Septum - general anatomical term|Anatomy|false|false||septumnull|Left ventricular cavity size|Attribute|false|false||left ventricular cavity sizenull|Cavity of left ventricle|Anatomy|false|false||left ventricular cavitynull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Cavity of ventricle|Anatomy|false|false||ventricular cavitynull|Heart Ventricle|Anatomy|false|false||ventricularnull|Ventricular|Modifier|false|false||ventricularnull|Dental caries|Disorder|false|false||cavity
null|Cavitation|Disorder|false|false||cavitynull|Body cavities|Anatomy|false|false||cavitynull|size|Modifier|false|false||sizenull|size - solid dosage form|LabModifier|false|false||sizenull|Table Cell Horizontal Align - left|Finding|false|false||Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|Heart Ventricle|Anatomy|false|false||ventricularnull|Ventricular|Modifier|false|false||ventricularnull|Systole|Finding|false|false||systolicnull|Function (attribute)|Finding|false|false||function
null|physiological aspects|Finding|false|false||function
null|Mathematical Operator|Finding|false|false||function
null|Functional Status|Finding|false|false||functionnull|Function Axis|Subject|false|false||functionnull|Table Cell Horizontal Align - right|Finding|false|false||Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|Heart Ventricle|Anatomy|false|false||ventricularnull|Ventricular|Modifier|false|false||ventricularnull|chamber [body part]|Anatomy|false|false||chambernull|Chamber (physical object)|Device|false|false||chambernull|size|Modifier|false|false||sizenull|size - solid dosage form|LabModifier|false|false||sizenull|Free of (attribute)|Finding|false|false||freenull|Empty (qualifier)|Modifier|false|false||freenull|Wall motion|Attribute|false|false||wall motionnull|Walls of a building|Device|false|false||wallnull|Motion|Phenomenon|false|false||motionnull|Aortic valve structure|Anatomy|false|false||aortic valve
null|Chest>Aortic valve|Anatomy|false|false||aortic valvenull|Aorta|Anatomy|false|false||aorticnull|Anatomical valve|Anatomy|false|false||valvenull|Valve (physical object)|Device|false|false||valve
null|Valve Device|Device|false|false||valve
null|medical valve|Device|false|false||valvenull|MILDLY|Modifier|false|false||mildly
null|Mild (qualifier value)|Modifier|false|false||mildlynull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Aortic valve structure|Anatomy|false|false||aortic valve
null|Chest>Aortic valve|Anatomy|false|false||aortic valvenull|Aorta|Anatomy|false|false||aorticnull|Anatomical valve|Anatomy|false|false||valvenull|Valve (physical object)|Device|false|false||valve
null|Valve Device|Device|false|false||valve
null|medical valve|Device|false|false||valvenull|Stenosis|Finding|false|false||stenosisnull|Stenosis <Pimeliinae>|Entity|false|false||stenosisnull|Stenosis Morphology|Modifier|false|false||stenosisnull|Valve Area|Finding|false|false||valve areanull|Anatomical valve|Anatomy|false|false||valvenull|Valve (physical object)|Device|false|false||valve
null|Valve Device|Device|false|false||valve
null|medical valve|Device|false|false||valvenull|Academic Research Enhancement Awards|Event|false|false||areanull|Geographic Locations|Entity|false|false||areanull|Area|Modifier|false|false||areanull|Chiari malformation type II|Disorder|false|false||cm2null|sq. cm|LabModifier|false|false||cm2null|Sequence Chromatogram|Finding|false|false||Tracenull|Trace Dosing Unit|LabModifier|false|false||Trace
null|trace amount|LabModifier|false|false||Trace
null|unknown - trace|LabModifier|false|false||Tracenull|Aortic Valve Insufficiency|Disorder|false|false||aortic regurgitationnull|Aorta|Anatomy|false|false||aorticnull|Regurgitation|Finding|false|false||regurgitation
null|Regurgitates after swallowing|Finding|false|false||regurgitationnull|Regurgitation - mechanism|Phenomenon|false|false||regurgitationnull|Mitral Valve|Anatomy|false|false||mitral valvenull|mitral|Modifier|false|false||mitralnull|Anatomical valve|Anatomy|false|false||valvenull|Valve (physical object)|Device|false|false||valve
null|Valve Device|Device|false|false||valve
null|medical valve|Device|false|false||valvenull|MILDLY|Modifier|false|false||mildly
null|Mild (qualifier value)|Modifier|false|false||mildlynull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Mitral valve annular calcification|Disorder|false|false||mitral annular calcificationnull|Premature calcification of mitral annulus|Finding|false|false||mitral annular calcificationnull|mitral|Modifier|false|false||mitralnull|Annular shape|Modifier|false|false||annularnull|Physiologic calcification|Finding|false|false||calcification
null|Calcification|Finding|false|false||calcification
null|Calcinosis|Finding|false|false||calcificationnull|Calcified (qualifier value)|Modifier|false|false||calcificationnull|Moderate - Severity of Illness Code|Finding|false|false||Moderate
null|Moderate|Finding|false|false||Moderatenull|Moderate (severity modifier)|Modifier|false|false||Moderate
null|Moderate - Allergy Severity|Modifier|false|false||Moderate
null|Moderation|Modifier|false|false||Moderatenull|mitral|Modifier|false|false||mitralnull|Regurgitation|Finding|false|false||regurgitation
null|Regurgitates after swallowing|Finding|false|false||regurgitationnull|Regurgitation - mechanism|Phenomenon|false|false||regurgitationnull|Acoustic shadowing|Finding|false|false||acoustic shadowingnull|Acoustics|Phenomenon|false|false||acousticnull|Shadowing (regime/therapy)|Procedure|false|false||shadowing
null|Shadowing (Histology)|Procedure|false|false||shadowingnull|With intensity|Modifier|false|false||severity
null|Severities|Modifier|false|false||severitynull|Mitral Valve Insufficiency|Disorder|false|false||mitral regurgitationnull|mitral|Modifier|false|false||mitralnull|Regurgitation|Finding|false|false||regurgitation
null|Regurgitates after swallowing|Finding|false|false||regurgitationnull|Regurgitation - mechanism|Phenomenon|false|false||regurgitationnull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Pulmonary artery structure|Anatomy|false|false||pulmonary arterynull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Arterial system|Anatomy|false|false||artery
null|Arteries|Anatomy|false|false||arterynull|Systolic Hypertension|Disorder|false|false||systolic hypertensionnull|Systole|Finding|false|false||systolicnull|Hypertensive disease|Disorder|false|false||hypertensionnull|Pericardial effusion|Disorder|true|false||pericardial effusionnull|Pericardial effusion body substance|Finding|true|false||pericardial effusionnull|Pericardial (qualifier value)|Anatomy|false|false||pericardial
null|Pericardial sac structure|Anatomy|false|false||pericardialnull|Effusion (substance)|Finding|true|false||effusion
null|null|Finding|true|false||effusion
null|effusion|Finding|true|false||effusionnull|null|Time|false|false||priornull|Study Object|Finding|false|false||studynull|Scientific Study|Procedure|false|false||study
null|Study|Procedure|false|false||study
null|Clinical Research|Procedure|false|false||studynull|Room of building - Study|Device|false|false||studynull|Similarity|Modifier|false|false||similarnull|Special Handling Code - Upright|Finding|false|false||UPRIGHTnull|Entity Handling - upright|Phenomenon|false|false||UPRIGHTnull|Upright|Modifier|false|false||UPRIGHTnull|Plain chest X-ray|Procedure|false|false||CHEST X-RAYnull|Chest problem|Finding|false|false||CHESTnull|Chest|Anatomy|false|false||CHEST
null|Anterior thoracic region|Anatomy|false|false||CHESTnull|ActClaimAttachmentCategoryCode - x-ray|Finding|false|false||X-RAY
null|roentgenographic|Finding|false|false||X-RAYnull|Plain x-ray|Procedure|false|false||X-RAY
null|Diagnostic radiologic examination|Procedure|false|false||X-RAY
null|Radiographic imaging procedure|Procedure|false|false||X-RAYnull|Roentgen Rays|Phenomenon|false|false||X-RAYnull|Most Recent|Time|false|false||most recentnull|Recent|Time|false|false||recentnull|Study Object|Finding|false|false||studynull|Scientific Study|Procedure|false|false||study
null|Study|Procedure|false|false||study
null|Clinical Research|Procedure|false|false||studynull|Room of building - Study|Device|false|false||studynull|Improvement|Finding|false|false||improvementnull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Pulmonary Edema|Finding|false|false||pulmonary edemanull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Reduced|Finding|false|false||decreasenull|Decrease|LabModifier|false|false||decreasenull|Small|LabModifier|false|false||smallnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Pleural effusion (disorder)|Finding|false|false||pleural effusion
null|Pleural effusion fluid|Finding|false|false||pleural effusion
null|null|Finding|false|false||pleural effusionnull|Pleural Diseases|Disorder|false|false||pleuralnull|Pleura|Anatomy|false|false||pleuralnull|Pleural|Modifier|false|false||pleuralnull|Effusion (substance)|Finding|false|false||effusion
null|null|Finding|false|false||effusion
null|effusion|Finding|false|false||effusionnull|Moderate - Severity of Illness Code|Finding|false|false||Moderate
null|Moderate|Finding|false|false||Moderatenull|Moderate (severity modifier)|Modifier|false|false||Moderate
null|Moderate - Allergy Severity|Modifier|false|false||Moderate
null|Moderation|Modifier|false|false||Moderatenull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Pleural effusion (disorder)|Finding|false|false||pleural effusion
null|Pleural effusion fluid|Finding|false|false||pleural effusion
null|null|Finding|false|false||pleural effusionnull|Pleural Diseases|Disorder|false|false||pleuralnull|Pleura|Anatomy|false|false||pleuralnull|Pleural|Modifier|false|false||pleuralnull|Effusion (substance)|Finding|false|false||effusion
null|null|Finding|false|false||effusion
null|effusion|Finding|false|false||effusionnull|Atelectasis|Finding|false|false||atelectasisnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Special Handling Code - Upright|Finding|false|false||UPRIGHTnull|Entity Handling - upright|Phenomenon|false|false||UPRIGHTnull|Upright|Modifier|false|false||UPRIGHTnull|Plain chest X-ray|Procedure|false|false||CHEST X-RAYnull|Chest problem|Finding|false|false||CHESTnull|Chest|Anatomy|false|false||CHEST
null|Anterior thoracic region|Anatomy|false|false||CHESTnull|ActClaimAttachmentCategoryCode - x-ray|Finding|false|false||X-RAY
null|roentgenographic|Finding|false|false||X-RAYnull|Plain x-ray|Procedure|false|false||X-RAY
null|Diagnostic radiologic examination|Procedure|false|false||X-RAY
null|Radiographic imaging procedure|Procedure|false|false||X-RAYnull|Roentgen Rays|Phenomenon|false|false||X-RAYnull|Cardiac attachment|Finding|false|false||Cardiacnull|Heart|Anatomy|false|false||Cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||Cardiacnull|size|Modifier|false|false||sizenull|size - solid dosage form|LabModifier|false|false||sizenull|Long Interspersed Elements|Drug|false|false||Lines
null|Long Interspersed Elements|Drug|false|false||Linesnull|Lines Quantity Limit Request|Finding|false|false||Linesnull|Lines - QueryQuantityUnit|Modifier|false|false||Lines
null|Linear|Modifier|false|false||Linesnull|null|Finding|false|false||tubesnull|biomedical tube device|Device|false|false||tubesnull|Tube Dosing Unit|LabModifier|false|false||tubesnull|Type of Agreement - Standard|Finding|false|false||standard
null|Standard (document)|Finding|false|false||standardnull|Standard base excess calculation technique|Procedure|false|false||standardnull|Standard (qualifier)|Modifier|false|false||standardnull|Position of phenotypic abnormality|Modifier|false|false||position
null|Positioning (attribute)|Modifier|false|false||positionnull|LARGE1 wt Allele|Finding|false|false||Large
null|LARGE1 gene|Finding|false|false||Largenull|Large|LabModifier|false|false||Largenull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Moderate - Severity of Illness Code|Finding|false|false||moderate
null|Moderate|Finding|false|false||moderatenull|Moderate (severity modifier)|Modifier|false|false||moderate
null|Moderate - Allergy Severity|Modifier|false|false||moderate
null|Moderation|Modifier|false|false||moderatenull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Pleural effusion (disorder)|Finding|false|false||pleural effusionsnull|Pleural Diseases|Disorder|false|false||pleuralnull|Pleura|Anatomy|false|false||pleuralnull|Pleural|Modifier|false|false||pleuralnull|effusion|Finding|false|false||effusionsnull|null|Finding|false|false||unchangednull|About The Same|Modifier|false|false||unchangednull|Positioning patient (procedure)|Procedure|false|false||positioning
null|Positioning - therapy|Procedure|false|false||positioningnull|Positioning (attribute)|Modifier|false|false||positioningnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Structure of right upper lobe of lung|Anatomy|false|false||Right upper lobenull|Table Cell Horizontal Align - right|Finding|false|false||Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|Structure of upper lobe of lung|Anatomy|false|false||upper lobenull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|AKT1S1 wt Allele|Finding|false|false||lobe
null|AKT1S1 gene|Finding|false|false||lobenull|lobe|Anatomy|false|false||lobenull|Abnormally opaque structure (morphologic abnormality)|Finding|false|false||opacity
null|Decreased translucency|Finding|false|false||opacitynull|Consistent with|Finding|false|false||consistent withnull|Compatible|Modifier|false|false||consistent withnull|Consistent with|Finding|false|false||consistentnull|Atelectasis|Finding|false|false||atelectasisnull|Pleural effusion (disorder)|Finding|false|false||Pleural effusionsnull|Pleural Diseases|Disorder|false|false||Pleuralnull|Pleura|Anatomy|false|false||Pleuralnull|Pleural|Modifier|false|false||Pleuralnull|effusion|Finding|false|false||effusionsnull|Atelectasis|Finding|false|false||atelectasisnull|Greater|LabModifier|false|false||larger
null|Large|LabModifier|false|false||largernull|RIGHT SIDE (USED TO IDENTIFY PROCEDURES PERFORMED ON THE RIGHT SIDE OF THE BODY)|Modifier|false|false||right side
null|Right|Modifier|false|false||right sidenull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Side|Modifier|false|false||sidenull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Blood Vessel|Anatomy|false|false||vascularnull|Vascular|Modifier|false|false||vascularnull|Congestion|Finding|false|false||congestionnull|Transaction counts and value totals - year|Finding|false|false||year
null|Precision - year|Finding|false|false||yearnull|year|Time|false|false||yearnull|Old|Time|false|false||oldnull|Woman|Subject|false|false||woman
null|Human, Female adult|Subject|false|false||womannull|Recent|Time|false|false||recentlynull|Sepsis|Disorder|false|false||sepsis
null|Septicemia|Disorder|false|false||sepsisnull|Sepsis <Sepsidae>|Entity|false|false||sepsisnull|Shock|Finding|false|false||shocknull|Readmission|Procedure|false|false||readmissionnull|Hypoxia, CTCAE|Finding|false|false||hypoxia
null|Hypoxia|Finding|false|false||hypoxianull|Hypercapnia|Finding|false|false||hypercarbianull|Respiratory attachment|Finding|false|false||respiratory
null|respiratory|Finding|false|false||respiratory
null|null|Finding|false|false||respiratory
null|Respiratory specimen|Finding|false|false||respiratorynull|Respiratory rate|Attribute|false|false||respiratorynull|Failure (biologic function)|Finding|false|false||failure
null|Failure|Finding|false|false||failure
null|Personal failure|Finding|false|false||failurenull|Urinary tract infection|Disorder|false|false||urinary tract infectionnull|Urinary tract|Anatomy|false|false||urinary tract
null|Urinary system|Anatomy|false|false||urinary tractnull|Urinary tract|Anatomy|false|false||urinarynull|urinary|Modifier|false|false||urinarynull|Tract|Anatomy|false|false||tractnull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|Respiratory Failure|Disorder|false|false||Respiratory Failurenull|Respiratory attachment|Finding|false|false||Respiratory
null|respiratory|Finding|false|false||Respiratory
null|null|Finding|false|false||Respiratory
null|Respiratory specimen|Finding|false|false||Respiratorynull|Respiratory rate|Attribute|false|false||Respiratorynull|Failure (biologic function)|Finding|false|false||Failure
null|Failure|Finding|false|false||Failure
null|Personal failure|Finding|false|false||Failurenull|Science of Etiology|Finding|false|false||Etiology
null|Etiology aspects|Finding|false|false||Etiology
null|Etiology|Finding|false|false||Etiologynull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Multifactorial|Finding|false|false||multifactorialnull|Respiratory insufficiency due to muscle weakness|Finding|false|false||respiratory muscle weakness
null|Respiratory muscle weakness|Finding|false|false||respiratory muscle weaknessnull|Respiratory Muscles|Anatomy|false|false||respiratory musclenull|Respiratory attachment|Finding|false|false||respiratory
null|respiratory|Finding|false|false||respiratory
null|null|Finding|false|false||respiratory
null|Respiratory specimen|Finding|false|false||respiratorynull|Respiratory rate|Attribute|false|false||respiratorynull|Paresis|Disorder|false|false||muscle weaknessnull|Muscle Weakness|Finding|false|false||muscle weaknessnull|Muscle (organ)|Anatomy|false|false||muscle
null|Muscle Tissue|Anatomy|false|false||musclenull|Weakness|Finding|false|false||weakness
null|Asthenia|Finding|false|false||weaknessnull|Pulmonary ventilator management|Procedure|false|false||pulmnull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Pleural effusion (disorder)|Finding|false|false||pleural effusionsnull|Pleural Diseases|Disorder|false|false||pleuralnull|Pleura|Anatomy|false|false||pleuralnull|Pleural|Modifier|false|false||pleuralnull|effusion|Finding|false|false||effusionsnull|On admission|Time|false|false||on admissionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|ActClaimAttachmentCategoryCode - x-ray|Finding|false|false||x-ray
null|roentgenographic|Finding|false|false||x-raynull|Plain x-ray|Procedure|false|false||x-ray
null|Diagnostic radiologic examination|Procedure|false|false||x-ray
null|Radiographic imaging procedure|Procedure|false|false||x-raynull|Roentgen Rays|Phenomenon|false|false||x-raynull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|mitral|Modifier|false|false||mitralnull|Intubated|Finding|false|false||intubatednull|Pulmonary Edema|Finding|false|false||pulmonary edemanull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Respiratory Muscles|Anatomy|false|false||respiratory musclenull|Respiratory attachment|Finding|false|false||respiratory
null|respiratory|Finding|false|false||respiratory
null|null|Finding|false|false||respiratory
null|Respiratory specimen|Finding|false|false||respiratorynull|Respiratory rate|Attribute|false|false||respiratorynull|Muscle (organ)|Anatomy|false|false||muscle
null|Muscle Tissue|Anatomy|false|false||musclenull|Weakness|Finding|false|false||weakness
null|Asthenia|Finding|false|false||weaknessnull|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group|Finding|false|false||poor
null|Patient Condition Code - Poor|Finding|false|false||poornull|Poverty|Subject|false|false||poornull|Language Proficiency - Poor|Modifier|false|false||poor
null|Specimen Quality - Poor|Modifier|false|false||poor
null|Poor - grade|Modifier|false|false||poor
null|Poor - qualifier|Modifier|false|false||poornull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Inspiratory force|Finding|false|false||inspiratory forcenull|Inspiration (function)|Finding|false|false||inspiratorynull|Mechanical force|Phenomenon|false|false||force
null|Force|Phenomenon|false|false||forcenull|Protein S100-A8|Drug|false|false||NIF
null|Protein S100-A8|Drug|false|false||NIF
null|Protein S100-A9|Drug|false|false||NIF
null|Protein S100-A9|Drug|false|false||NIFnull|S100A9 wt Allele|Finding|false|false||NIF
null|S100A8 wt Allele|Finding|false|false||NIF
null|S100A9 gene|Finding|false|false||NIFnull|Protein S100-A8|Drug|false|false||NIF
null|Protein S100-A8|Drug|false|false||NIF
null|Protein S100-A9|Drug|false|false||NIF
null|Protein S100-A9|Drug|false|false||NIFnull|S100A9 wt Allele|Finding|false|false||NIF
null|S100A8 wt Allele|Finding|false|false||NIF
null|S100A9 gene|Finding|false|false||NIFnull|Optimization|Event|false|false||optimizationnull|Nutrition (function)|Finding|false|false||nutrition
null|Nutritional status|Finding|false|false||nutrition
null|Nutrition outcomes|Finding|false|false||nutritionnull|Feeding and dietary regimes|Procedure|false|false||nutrition
null|Nutritional Study|Procedure|false|false||nutritionnull|Science of nutrition|Title|false|false||nutritionnull|Supportive care|Procedure|false|false||supportive care
null|Palliative Care|Procedure|false|false||supportive carenull|Supportive assistance|Finding|false|false||supportivenull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Pulmonary Edema|Finding|false|false||pulmonary edemanull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Precaution Code - Aggressive|Finding|false|false||aggressive
null|Aggressive behavior|Finding|false|false||aggressive
null|Risk Codes - Aggressive|Finding|false|false||aggressivenull|Aggressive course|Time|false|false||aggressivenull|Entity Risk - aggressive|Modifier|false|false||aggressivenull|Diuresis|Finding|false|false||diuresisnull|Lasix|Drug|false|false||Lasix
null|Lasix|Drug|false|false||Lasixnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Lasix|Drug|false|false||Lasix
null|Lasix|Drug|false|false||Lasixnull|Biomaterial Treatment|Finding|false|false||treatment
null|Treating|Finding|false|false||treatment
null|therapeutic aspects|Finding|false|false||treatmentnull|treatment - ActInformationManagementReason|Procedure|false|false||treatment
null|Administration (procedure)|Procedure|false|false||treatment
null|Therapeutic procedure|Procedure|false|false||treatmentnull|Able (qualifier value)|Finding|false|false||ablenull|Ability|Subject|false|false||ablenull|Oxygen nasal cannula|Device|false|false||nasal cannula
null|Nasal Cannula|Device|false|false||nasal cannulanull|Nasal brand of oxymetazoline|Drug|false|false||nasal
null|Nasal brand of oxymetazoline|Drug|false|false||nasal
null|Nasal dosage form|Drug|false|false||nasalnull|Nasal Route of Administration|Finding|false|false||nasal
null|Nasal (intended site)|Finding|false|false||nasalnull|null|Anatomy|false|false||nasalnull|Specimen Type - Cannula|Finding|false|false||cannula
null|null|Finding|false|false||cannulanull|Body Parts - Cannula|Anatomy|false|false||cannulanull|Cannula device|Device|false|false||cannulanull|Calamus <grasshoppers>|Entity|false|false||cannulanull|lisinopril|Drug|false|false||Lisinopril
null|lisinopril|Drug|false|false||Lisinoprilnull|Daily|Time|false|false||dailynull|Reduced|Finding|false|false||reductionnull|Reduction procedure|Procedure|false|false||reduction
null|Surgical reduction|Procedure|false|false||reductionnull|Reduction (chemical)|Phenomenon|false|false||reductionnull|contextual factors|Finding|false|false||settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Further|Modifier|false|false||furthernull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Dosage|LabModifier|false|false||dosesnull|Lasix|Drug|false|false||Lasix
null|Lasix|Drug|false|false||Lasixnull|Rehabilitation therapy|Procedure|false|false||rehabnull|Lasix|Drug|false|false||Lasix
null|Lasix|Drug|false|false||Lasixnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|lisinopril|Drug|false|false||lisinopril
null|lisinopril|Drug|false|false||lisinoprilnull|Observation Interpretation - better|Finding|false|false||betternull|Better|Modifier|false|false||betternull|Reduced|Finding|false|false||reductionnull|Reduction procedure|Procedure|false|false||reduction
null|Surgical reduction|Procedure|false|false||reductionnull|Reduction (chemical)|Phenomenon|false|false||reductionnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|Pseudomonas Infections|Disorder|false|false||Pseudomonasnull|Pseudomonas|Entity|false|false||Pseudomonasnull|urinastatin|Drug|false|false||UTI
null|urinastatin|Drug|false|false||UTInull|Urinary tract infection|Disorder|false|false||UTInull|AMBP wt Allele|Finding|false|false||UTI
null|AMBP gene|Finding|false|false||UTInull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Pseudomonas Infections|Disorder|false|false||Pseudomonasnull|Pseudomonas|Entity|false|false||Pseudomonasnull|Sensitive|Finding|false|false||sensitive tonull|Sensitive|Finding|false|false||sensitivenull|stimulus sensitivity|Modifier|false|false||sensitivenull|gentamicin|Drug|false|false||Gentamicin
null|gentamicin|Drug|false|false||Gentamicinnull|Gentamicin measurement|Procedure|false|false||Gentamicinnull|Urine culture|Procedure|false|false||urine culturenull|Portion of urine|Finding|false|false||urine
null|null|Finding|false|false||urine
null|Urine|Finding|false|false||urine
null|In Urine|Finding|false|false||urine
null|Urine specimen|Finding|false|false||urinenull|Culture Dose Form|Drug|false|false||culturenull|Culture (Anthropological)|Finding|false|false||culture
null|Cultural aspects|Finding|false|false||culturenull|Microbial culture (procedure)|Procedure|false|false||culture
null|Laboratory culture|Procedure|false|false||culturenull|Initially|Time|false|false||initiallynull|Double (qualifier value)|Finding|false|false||doublenull|Doubling|Event|false|false||doublenull|Double Value Type|Modifier|false|false||doublenull|coverage - HL7PublishingDomain|Finding|false|false||coverage
null|null|Finding|false|false||coverage
null|coverage - financial contract|Finding|false|false||coveragenull|Cipro|Drug|false|false||Cipro
null|Cipro|Drug|false|false||Cipronull|cefepime|Drug|false|false||Cefepime
null|cefepime|Drug|false|false||Cefepimenull|Culture (Anthropological)|Finding|false|false||culturesnull|Pending - Allergy Clinical Status|Finding|false|false||pending
null|Pending - referral status|Finding|false|false||pendingnull|Pending - status|Time|false|false||pendingnull|pending - ManagedParticipationStatus|Modifier|false|false||pending
null|pending - RoleStatus|Modifier|false|false||pending
null|Pending - Day type|Modifier|false|false||pendingnull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|cefepime|Drug|false|false||Cefepime
null|cefepime|Drug|false|false||Cefepimenull|Living Alone|Finding|false|false||alonenull|alone - group size|Subject|false|false||alonenull|Singular|LabModifier|false|false||alonenull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|Concern|Finding|false|false||concernnull|Drug Eruptions|Finding|false|false||drug rashnull|Pharmaceutical Preparations|Drug|false|false||drug
null|Pharmacologic Substance|Drug|false|false||drugnull|Drug problem|Finding|false|false||drugnull|Eruption of skin (disorder)|Disorder|false|false||rashnull|Skin rash|Finding|false|false||rash
null|Eruptions|Finding|false|false||rash
null|Exanthema|Finding|false|false||rashnull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|Zosyn|Drug|false|false||Zosyn
null|Zosyn|Drug|false|false||Zosynnull|Zosyn|Drug|false|false||Zosyn
null|Zosyn|Drug|false|false||Zosynnull|Course|Time|false|false||coursenull|Total|Modifier|false|false||totalnull|day|Time|false|false||daysnull|Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE|Drug|false|false||antibiotics
null|Antibiotics|Drug|false|false||antibiotics
null|Antibiotics, ophthalmologic|Drug|false|false||antibiotics
null|Antibiotics, Gynecological|Drug|false|false||antibiotics
null|antibiotics, intestinal|Drug|false|false||antibiotics
null|Antibiotic throat preparations|Drug|false|false||antibiotics
null|Antibiotics, Antitubercular|Drug|false|false||antibiotics
null|Antibiotics for systemic use|Drug|false|false||antibiotics
null|Antifungal Antibiotics, Topical|Drug|false|false||antibioticsnull|Complicated|Finding|false|false||complicatednull|urinastatin|Drug|false|false||UTI
null|urinastatin|Drug|false|false||UTInull|Urinary tract infection|Disorder|false|false||UTInull|AMBP wt Allele|Finding|false|false||UTI
null|AMBP gene|Finding|false|false||UTInull|Eruption of skin (disorder)|Disorder|false|false||RASHnull|Skin rash|Finding|false|false||RASH
null|Eruptions|Finding|false|false||RASH
null|Exanthema|Finding|false|false||RASHnull|DYRK3 gene|Finding|false|false||red
null|Redness|Finding|false|false||red
null|IK gene|Finding|false|false||rednull|Radiological Exposure Device|Device|false|false||rednull|Red color|Modifier|false|false||rednull|Macular rash|Finding|false|false||macular rashnull|macular|Modifier|false|false||macularnull|Eruption of skin (disorder)|Disorder|false|false||rashnull|Skin rash|Finding|false|false||rash
null|Eruptions|Finding|false|false||rash
null|Exanthema|Finding|false|false||rashnull|All extremities|Anatomy|false|false||extremities
null|Limb structure|Anatomy|false|false||extremitiesnull|Initially|Time|false|false||initiallynull|Drug Eruptions|Finding|false|false||drug rashnull|Pharmaceutical Preparations|Drug|false|false||drug
null|Pharmacologic Substance|Drug|false|false||drugnull|Drug problem|Finding|false|false||drugnull|Eruption of skin (disorder)|Disorder|false|false||rashnull|Skin rash|Finding|false|false||rash
null|Eruptions|Finding|false|false||rash
null|Exanthema|Finding|false|false||rashnull|Late|Time|false|false||laternull|More|LabModifier|false|false||morenull|Consistent with|Finding|false|false||consistent withnull|Compatible|Modifier|false|false||consistent withnull|Consistent with|Finding|false|false||consistentnull|Contact Dermatitis|Disorder|false|false||contact dermatitisnull|Contact with|Finding|false|false||contact
null|Contact - HL7 Attribution|Finding|false|false||contact
null|Communication Contact|Finding|false|false||contactnull|contact person|Subject|false|false||contactnull|Physical contact|Phenomenon|false|false||contactnull|Personal Contact|Event|false|false||contactnull|Dermatitis|Disorder|false|false||dermatitisnull|Eczema|Disorder|false|false||eczemanull|triamcinolone|Drug|false|false||Triamcinolone
null|triamcinolone|Drug|false|false||Triamcinolonenull|Emollient Cream|Drug|false|false||cream
null|Cream|Drug|false|false||cream
null|Dairy Cream|Drug|false|false||creamnull|Eruption of skin (disorder)|Disorder|false|false||rashnull|Skin rash|Finding|false|false||rash
null|Eruptions|Finding|false|false||rash
null|Exanthema|Finding|false|false||rashnull|Colitis|Disorder|false|false||Colitisnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Recent|Time|false|false||recentlynull|Colitis|Disorder|false|false||colitisnull|Sepsis|Disorder|false|false||sepsis
null|Septicemia|Disorder|false|false||sepsisnull|Sepsis <Sepsidae>|Entity|false|false||sepsisnull|Repeat Object|Finding|false|false||Repeat
null|Repeat|Finding|false|false||Repeatnull|Repeat Pattern|Time|false|false||Repeatnull|Residual Cancer Burden Class 0|Finding|false|false||PCR
null|Pathologic Complete Response|Finding|false|false||PCRnull|Probe with target amplification technique|Procedure|false|false||PCR
null|Polymerase Chain Reaction|Procedure|false|false||PCRnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Last|Modifier|false|false||lastnull|Hospitalization|Procedure|false|false||hospitalizationnull|vancomycin|Drug|false|false||vancomycin
null|vancomycin|Drug|false|false||vancomycinnull|Vancomycin measurement|Procedure|false|false||vancomycinnull|Course|Time|false|false||coursenull|vancomycin|Drug|false|false||vancomycin
null|vancomycin|Drug|false|false||vancomycinnull|Vancomycin measurement|Procedure|false|false||vancomycinnull|during hospitalization|Time|false|false||during hospitalizationnull|Hospitalization|Procedure|false|false||hospitalizationnull|Concurrent|Time|false|false||concurrentnull|Biomaterial Treatment|Finding|false|false||treatment
null|Treating|Finding|false|false||treatment
null|therapeutic aspects|Finding|false|false||treatmentnull|treatment - ActInformationManagementReason|Procedure|false|false||treatment
null|Administration (procedure)|Procedure|false|false||treatment
null|Therapeutic procedure|Procedure|false|false||treatmentnull|Widening|Modifier|false|false||broadnull|Spectrum|Finding|false|false||spectrumnull|Electromagnetic Spectrum|LabModifier|false|false||spectrumnull|Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE|Drug|false|false||antibiotics
null|Antibiotics|Drug|false|false||antibiotics
null|Antibiotics, ophthalmologic|Drug|false|false||antibiotics
null|Antibiotics, Gynecological|Drug|false|false||antibiotics
null|antibiotics, intestinal|Drug|false|false||antibiotics
null|Antibiotic throat preparations|Drug|false|false||antibiotics
null|Antibiotics, Antitubercular|Drug|false|false||antibiotics
null|Antibiotics for systemic use|Drug|false|false||antibiotics
null|Antifungal Antibiotics, Topical|Drug|false|false||antibioticsnull|Zosyn|Drug|false|false||zosyn
null|Zosyn|Drug|false|false||zosynnull|Pseudomonas Infections|Disorder|false|false||pseudomonasnull|Pseudomonas|Entity|false|false||pseudomonasnull|urinastatin|Drug|false|false||UTI
null|urinastatin|Drug|false|false||UTInull|Urinary tract infection|Disorder|false|false||UTInull|AMBP wt Allele|Finding|false|false||UTI
null|AMBP gene|Finding|false|false||UTInull|Zosyn|Drug|false|false||zosyn
null|Zosyn|Drug|false|false||zosynnull|vancomycin|Drug|false|false||vanco
null|vancomycin|Drug|false|false||vanconull|Anemia|Disorder|false|false||Anemianull|Anemia <Anemiaceae>|Entity|false|false||Anemianull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|null|Finding|false|false||guaiac positive stoolsnull|guaiac positive|Lab|false|false||guaiac positivenull|guaiac|Drug|false|false||guaiac
null|guaiac|Drug|false|false||guaiacnull|BRAF Gene Rearrangement|Disorder|false|false||positivenull|Rh Positive Blood Group|Finding|false|false||positive
null|Positive Finding|Finding|false|false||positive
null|Positive|Finding|false|false||positivenull|Positive Charge|Modifier|false|false||positivenull|Positive Number|LabModifier|false|false||positivenull|Feces|Finding|false|false||stoolsnull|null|Attribute|false|false||stoolsnull|Stool seat|Device|false|false||stoolsnull|Last|Modifier|false|false||lastnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Message Waiting Priority - High|Finding|false|false||high
null|high - ActExposureLevelCode|Finding|false|false||high
null|IPSS Risk Category High|Finding|false|false||high
null|IPSS-R Risk Category High|Finding|false|false||high
null|High (finding)|Finding|false|false||highnull|Observation Value - High|Modifier|false|false||high
null|High|Modifier|false|false||high
null|Abnormally high|Modifier|false|false||highnull|Hospitalization|Procedure|false|false||hospitalizationnull|Storage Unit|Device|false|false||unit
null|Unit device|Device|false|false||unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||unit
null|Unit of Measure|LabModifier|false|false||unit
null|Unit|LabModifier|false|false||unit
null|Enzyme Unit|LabModifier|false|false||unitnull|Colloids|Drug|false|false||colloidnull|Colloid, body substance|Finding|false|false||colloidnull|pressure support|Procedure|false|false||pressure supportnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|Support brand of multivitamin|Drug|false|false||support
null|Support brand of multivitamin|Drug|false|false||support
null|Support brand of multivitamin|Drug|false|false||supportnull|Supportive assistance|Finding|false|false||supportnull|Supportive care|Procedure|false|false||supportnull|Support - dental|Attribute|false|false||supportnull|null|Device|false|false||supportnull|Hypothyroidism|Disorder|false|false||Hypothyroidismnull|Synthetic Levothyroxine|Drug|false|false||levothyroxine
null|Synthetic Levothyroxine|Drug|false|false||levothyroxine
null|levothyroxine|Drug|false|false||levothyroxine
null|levothyroxine|Drug|false|false||levothyroxine
null|levothyroxine|Drug|false|false||levothyroxinenull|microgram|LabModifier|false|false||mcgnull|Daily|Time|false|false||dailynull|Gastroesophageal reflux disease|Disorder|false|false||GERDnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|omeprazole|Drug|false|false||omeprazole
null|omeprazole|Drug|false|false||omeprazolenull|Last|Modifier|false|false||lastnull|Hospitalization|Procedure|false|false||hospitalizationnull|BRAF Gene Rearrangement|Disorder|false|false||positivenull|Rh Positive Blood Group|Finding|false|false||positive
null|Positive Finding|Finding|false|false||positive
null|Positive|Finding|false|false||positivenull|Positive Charge|Modifier|false|false||positivenull|Positive Number|LabModifier|false|false||positivenull|Histamine H2 Antagonists|Drug|false|false||H2 blockernull|Prophylactic treatment|Procedure|false|false||prophylaxisnull|prevention & control|Modifier|false|false||prophylaxisnull|contextual factors|Finding|false|false||settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|Delirium|Disorder|false|false||deliriumnull|famotidine|Drug|false|false||Famotidine
null|famotidine|Drug|false|false||Famotidinenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Delirium|Disorder|false|false||deliriousnull|Electrocardiogram image|Finding|false|false||EKG
null|Electrocardiogram|Finding|false|false||EKGnull|Electrocardiography|Procedure|false|false||EKGnull|Changing|Finding|false|false||Changesnull|Changed status|LabModifier|false|false||Changesnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Lateral|Modifier|false|false||lateralnull|SULT1E1 wt Allele|Finding|false|false||STE
null|SULT1E1 gene|Finding|false|false||STEnull|MILDLY|Modifier|false|false||mildly
null|Mild (qualifier value)|Modifier|false|false||mildlynull|Elevated|Modifier|false|false||elevated
null|High|Modifier|false|false||elevatednull|Troponin|Drug|false|false||troponin
null|Troponin|Drug|false|false||troponinnull|Troponin measurement|Procedure|false|false||troponinnull|Per Megabase Pair|LabModifier|false|false||/MBnull|Residential flat|Device|false|false||flatnull|Flat shape|Modifier|false|false||flatnull|On admission|Time|false|false||on admissionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Blunt (object)|Device|false|false||bluntnull|Blunted|Modifier|false|false||bluntnull|Traumatic AND/OR non-traumatic injury|Disorder|false|false||injury
null|Traumatic injury|Disorder|false|false||injurynull|Compressed structure|Finding|false|false||compressionsnull|Compression|Phenomenon|false|false||compressionsnull|Ischemia co-occurrent and due to increased oxygen demand|Disorder|false|false||demand ischemianull|Economic demand|Finding|false|false||demandnull|Demand (clinical)|Procedure|false|false||demandnull|Ischemia|Finding|false|false||ischemianull|Ischemia Procedure|Procedure|false|false||ischemianull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Femur|Anatomy|false|false||femoralnull|contextual factors|Finding|false|false||settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|Hypotension|Finding|false|false||hypotensionnull|Inventory of Callous-Unemotional Traits|Finding|false|false||ICUnull|Structure of intraculminate fissure|Anatomy|false|false||ICUnull|intensive care unit|Device|false|false||ICUnull|intensive care unit|Entity|false|false||ICUnull|Peripherally Inserted Central Catheter Line Insertion|Procedure|false|false||PICCnull|Peripherally inserted central catheter (physical object)|Device|false|false||PICCnull|SET protein, human|Drug|false|false||set
null|SET protein, human|Drug|false|false||setnull|Parameterized Data Type - Set|Finding|false|false||set
null|Set scale|Finding|false|false||set
null|Set (Psychology)|Finding|false|false||set
null|SET gene|Finding|false|false||set
null|set (group)|Finding|false|false||setnull|Lactobacillus|Entity|false|false||Lactobacillusnull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false||skin
null|Skin and subcutaneous tissue disorders|Disorder|false|false||skinnull|Skin Specimen Source Code|Finding|false|false||skin
null|Skin Specimen|Finding|false|false||skinnull|Skin, Human|Anatomy|false|false||skin
null|Skin|Anatomy|false|false||skinnull|Contaminant|Drug|false|false||contaminantnull|surveillance aspects|Finding|false|false||surveillancenull|Medical Surveillance|Procedure|false|false||surveillancenull|legal surveillance|Event|false|false||surveillancenull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Marketing basis - Transitional|Finding|false|false||TRANSITIONALnull|Transitional cell morphology|Modifier|false|false||TRANSITIONALnull|MDF Attribute Type - Code|Finding|false|false||Code
null|A Codes|Finding|false|false||Code
null|Code|Finding|false|false||Codenull|Coding|Event|false|false||Codenull|Full|Modifier|false|false||Fullnull|Laboratory test finding|Lab|false|false||Labsnull|Daily|Time|false|false||dailynull|Basic metabolic panel|Procedure|false|false||chem 7null|chemical aspects|Finding|false|false||chemnull|Chemical procedure|Procedure|false|false||chemnull|Science of Chemistry|Subject|false|false||chemnull|Phos <Photinae>|Entity|false|false||phosnull|Nutrition (function)|Finding|false|false||Nutrition
null|Nutritional status|Finding|false|false||Nutrition
null|Nutrition outcomes|Finding|false|false||Nutritionnull|Feeding and dietary regimes|Procedure|false|false||Nutrition
null|Nutritional Study|Procedure|false|false||Nutritionnull|Science of nutrition|Title|false|false||Nutritionnull|Unspecified tube|Finding|false|false||Tube
null|TUBE1 gene|Finding|false|false||Tubenull|biomedical tube device|Device|false|false||Tube
null|Packaging Tube|Device|false|false||Tubenull|tube|Modifier|false|false||Tubenull|Tube (unit of presentation)|LabModifier|false|false||Tube
null|Tube Dosing Unit|LabModifier|false|false||Tubenull|Soft diet|Procedure|false|false||soft dietnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||softnull|Soft|Modifier|false|false||softnull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Thin (qualifier value)|Modifier|false|false||thinnull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|fluticasone|Drug|false|false||fluticasone
null|fluticasone|Drug|false|false||fluticasonenull|mcg/actuation|LabModifier|false|false||mcg/actuationnull|microgram|LabModifier|false|false||mcgnull|Actuation (unit of presentation)|LabModifier|false|false||actuationnull|SPRAY, SUSPENSION|Drug|false|false||Spray, Suspensionnull|Spray Dosage Form|Drug|false|false||Spraynull|Spray (administration method)|Finding|false|false||Spraynull|Spray (action)|Event|false|false||Spraynull|Spray Dosing Unit|LabModifier|false|false||Spraynull|Suspension substance|Drug|false|false||Suspension
null|Suspensions|Drug|false|false||Suspensionnull|Suspension (action)|Finding|false|false||Suspensionnull|Puff Dosing Unit|LabModifier|false|false||puffsnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Synthetic Levothyroxine|Drug|false|false||levothyroxine
null|Synthetic Levothyroxine|Drug|false|false||levothyroxine
null|levothyroxine|Drug|false|false||levothyroxine
null|levothyroxine|Drug|false|false||levothyroxine
null|levothyroxine|Drug|false|false||levothyroxinenull|microgram|LabModifier|false|false||mcgnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Daily|Time|false|false||DAILYnull|Acetaminophen [EPC]|Drug|false|false||acetaminophen
null|acetaminophen|Drug|false|false||acetaminophen
null|acetaminophen|Drug|false|false||acetaminophennull|Acetaminophen measurement|Procedure|false|false||acetaminophennull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletsnull|CIAO3 gene|Finding|false|false||prnnull|As required|Time|false|false||prn
null|Pro Re Nata|Time|false|false||prnnull|polyvinyl alcohol|Drug|false|false||polyvinyl alcoholnull|Polyvinyls|Drug|false|false||polyvinyl
null|Polyvinyls|Drug|false|false||polyvinylnull|Alcohols|Drug|false|false||alcohol
null|Alcohols|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcoholnull|Alcohol - Recreational Drug Use Code|Finding|false|false||alcoholnull|Drops - Drug Form|Drug|false|false||Dropsnull|Drop Dosing Unit|LabModifier|false|false||Dropsnull|Hour|Time|false|false||hoursnull|CIAO3 gene|Finding|false|false||prnnull|As required|Time|false|false||prn
null|Pro Re Nata|Time|false|false||prnnull|insulin lispro|Drug|true|false||insulin lispro
null|insulin lispro|Drug|true|false||insulin lispro
null|insulin lispro|Drug|true|false||insulin lispronull|insulin, regular, human|Drug|false|false||insulin
null|Insulin [EPC]|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulinnull|INS gene|Finding|false|false||insulinnull|Insulin measurement|Procedure|false|false||insulinnull|insulin lispro|Drug|false|false||lispro
null|insulin lispro|Drug|false|false||lispro
null|insulin lispro|Drug|false|false||lispronull|Unit per Milliliter|LabModifier|false|false||unit/mLnull|Storage Unit|Device|false|false||unit
null|Unit device|Device|false|false||unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||unit
null|Unit of Measure|LabModifier|false|false||unit
null|Unit|LabModifier|false|false||unit
null|Enzyme Unit|LabModifier|false|false||unitnull|per milliliter|LabModifier|false|false||/mLnull|Solution Dosage Form|Drug|false|false||Solution
null|Solutions|Drug|false|false||Solution
null|Pharmaceutical Solutions|Drug|false|false||Solutionnull|Resolution|Finding|false|false||Solutionnull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|sliding scale|Procedure|false|false||Sliding scalenull|Sliding|Finding|false|false||Slidingnull|Scale, LOINC Axis 5|Finding|false|false||scale
null|Base Number|Finding|false|false||scale
null|Scale - rank|Finding|false|false||scalenull|Integumentary scale|Anatomy|false|false||scalenull|Weight measurement scales|Device|false|false||scalenull|Scaling|Event|false|false||scalenull|Unit - NCI Thesaurus Property|LabModifier|false|false||units
null|Unit of Measure|LabModifier|false|false||units
null|Unit|LabModifier|false|false||unitsnull|Subcutaneous Route of Administration|Finding|false|false||Subcutaneousnull|subcutaneous|Modifier|false|false||Subcutaneousnull|Three times daily|Time|false|false||three times a daynull|Thrice|LabModifier|false|false||three timesnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Unit - NCI Thesaurus Property|LabModifier|false|false||units
null|Unit of Measure|LabModifier|false|false||units
null|Unit|LabModifier|false|false||unitsnull|Unit - NCI Thesaurus Property|LabModifier|false|false||units
null|Unit of Measure|LabModifier|false|false||units
null|Unit|LabModifier|false|false||unitsnull|Unit - NCI Thesaurus Property|LabModifier|false|false||units
null|Unit of Measure|LabModifier|false|false||units
null|Unit|LabModifier|false|false||unitsnull|Unit - NCI Thesaurus Property|LabModifier|false|false||units
null|Unit of Measure|LabModifier|false|false||units
null|Unit|LabModifier|false|false||unitsnull|Unit - NCI Thesaurus Property|LabModifier|false|false||units
null|Unit of Measure|LabModifier|false|false||units
null|Unit|LabModifier|false|false||unitsnull|Unit - NCI Thesaurus Property|LabModifier|false|false||units
null|Unit of Measure|LabModifier|false|false||units
null|Unit|LabModifier|false|false||unitsnull|Call - dosing instruction fragment|Finding|false|false||call
null|Call (Instruction)|Finding|false|false||call
null|Decision|Finding|false|false||call
null|CHL1 gene|Finding|false|false||callnull|miconazole nitrate|Drug|false|false||miconazole nitrate
null|miconazole nitrate|Drug|false|false||miconazole nitratenull|miconazole|Drug|false|false||miconazole
null|miconazole|Drug|false|false||miconazolenull|nitrate ion|Drug|false|false||nitrate
null|nitrate ion|Drug|false|false||nitrate
null|Nitrate|Drug|false|false||nitrate
null|Nitrates|Drug|false|false||nitratenull|powder physical state|Drug|false|false||Powder
null|Powder dose form|Drug|false|false||Powdernull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|CIAO3 gene|Finding|false|false||prnnull|As required|Time|false|false||prn
null|Pro Re Nata|Time|false|false||prnnull|Eruption of skin (disorder)|Disorder|false|false||rashnull|Skin rash|Finding|false|false||rash
null|Eruptions|Finding|false|false||rash
null|Exanthema|Finding|false|false||rashnull|vancomycin|Drug|false|false||vancomycin
null|vancomycin|Drug|false|false||vancomycinnull|Vancomycin measurement|Procedure|false|false||vancomycinnull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Every six hours|Time|false|false||Q6Hnull|7 days|Time|false|false||7 daysnull|day|Time|false|false||daysnull|heparin, porcine|Drug|false|false||heparin (porcine)
null|heparin, porcine|Drug|false|false||heparin (porcine)
null|heparin, porcine|Drug|false|false||heparin (porcine)null|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparinnull|Porcine prosthetic valve|Finding|false|false||porcinenull|Porcine species|Entity|false|false||porcine
null|Family suidae|Entity|false|false||porcinenull|Unit per Milliliter|LabModifier|false|false||unit/mLnull|Storage Unit|Device|false|false||unit
null|Unit device|Device|false|false||unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||unit
null|Unit of Measure|LabModifier|false|false||unit
null|Unit|LabModifier|false|false||unit
null|Enzyme Unit|LabModifier|false|false||unitnull|per milliliter|LabModifier|false|false||/mLnull|Solution Dosage Form|Drug|false|false||Solution
null|Solutions|Drug|false|false||Solution
null|Pharmaceutical Solutions|Drug|false|false||Solutionnull|Resolution|Finding|false|false||Solutionnull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|albuterol sulfate|Drug|false|false||albuterol sulfate
null|albuterol sulfate|Drug|false|false||albuterol sulfatenull|albuterol|Drug|false|false||albuterol
null|albuterol|Drug|false|false||albuterolnull|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||sulfate
null|Sulfates, Inorganic|Drug|false|false||sulfate
null|sulfate ion|Drug|false|false||sulfate
null|sulfate ion|Drug|false|false||sulfate
null|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||sulfatenull|Solution Dosage Form|Drug|false|false||Solution
null|Solutions|Drug|false|false||Solution
null|Pharmaceutical Solutions|Drug|false|false||Solutionnull|Resolution|Finding|false|false||Solutionnull|CIAO3 gene|Finding|false|false||prnnull|As required|Time|false|false||prn
null|Pro Re Nata|Time|false|false||prnnull|Dyspnea|Finding|false|false||SOBnull|ipratropium bromide|Drug|false|false||ipratropium bromide
null|ipratropium bromide|Drug|false|false||ipratropium bromidenull|ipratropium|Drug|false|false||ipratropium
null|ipratropium|Drug|false|false||ipratropiumnull|Bromides|Drug|false|false||bromidenull|Bromides measurement|Procedure|false|false||bromidenull|Solution Dosage Form|Drug|false|false||Solution
null|Solutions|Drug|false|false||Solution
null|Pharmaceutical Solutions|Drug|false|false||Solutionnull|Resolution|Finding|false|false||Solutionnull|CIAO3 gene|Finding|false|false||prnnull|As required|Time|false|false||prn
null|Pro Re Nata|Time|false|false||prnnull|Dyspnea|Finding|false|false||SOBnull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|null|Drug|false|false||Vancomycin Oralnull|vancomycin|Drug|false|false||Vancomycin
null|vancomycin|Drug|false|false||Vancomycinnull|Vancomycin measurement|Procedure|false|false||Vancomycinnull|Oral Liquid Product|Drug|false|false||Oral Liquidnull|Oral Dosage Form|Drug|false|false||Oralnull|Oral Route of Administration|Finding|false|false||Oral
null|Oral (intended site)|Finding|false|false||Oralnull|Oral cavity|Anatomy|false|false||Oralnull|Oral|Modifier|false|false||Oralnull|Liquid Dosage Form|Drug|false|false||Liquid
null|Liquid substance|Drug|false|false||Liquidnull|Liquid (finding)|Finding|false|false||Liquidnull|Liquid diet|Procedure|false|false||Liquidnull|Liquid (state of matter)|Modifier|false|false||Liquidnull|Every six hours|Time|false|false||Q6Hnull|Duration brand of oxymetazoline|Drug|false|false||Durationnull|Duration (temporal concept)|Time|false|false||Durationnull|day|Time|false|false||Daysnull|Last|Modifier|false|false||Lastnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|fluticasone propionate|Drug|false|false||Fluticasone Propionate
null|fluticasone propionate|Drug|false|false||Fluticasone Propionatenull|fluticasone|Drug|false|false||Fluticasone
null|fluticasone|Drug|false|false||Fluticasonenull|propionate|Drug|false|false||Propionate
null|Propionates|Drug|false|false||Propionatenull|Puff Dosing Unit|LabModifier|false|false||PUFF
null|Picofarad|LabModifier|false|false||PUFFnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|levothyroxine sodium|Drug|false|false||Levothyroxine Sodium
null|levothyroxine sodium|Drug|false|false||Levothyroxine Sodium
null|levothyroxine sodium|Drug|false|false||Levothyroxine Sodiumnull|Synthetic Levothyroxine|Drug|false|false||Levothyroxine
null|Synthetic Levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxinenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|microgram|LabModifier|false|false||mcgnull|Daily|Time|false|false||DAILYnull|triamcinolone acetonide|Drug|false|false||Triamcinolone Acetonide
null|triamcinolone acetonide|Drug|false|false||Triamcinolone Acetonidenull|triamcinolone|Drug|false|false||Triamcinolone
null|triamcinolone|Drug|false|false||Triamcinolonenull|Emollient Cream|Drug|false|false||Cream
null|Cream|Drug|false|false||Cream
null|Dairy Cream|Drug|false|false||Creamnull|APPL1 gene|Finding|false|false||Applnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Liposarcoma, Pleomorphic|Disorder|false|false||pls
null|Papillon-Lefevre Disease|Disorder|false|false||pls
null|Lateral Sclerosis|Disorder|false|false||plsnull|CTSC wt Allele|Finding|false|false||pls
null|CTSC gene|Finding|false|false||plsnull|Thin (qualifier value)|Modifier|false|false||thinnull|anatomical layer|Anatomy|false|false||layernull|Chicken laying egg for human food|Entity|false|false||layernull|Coating (film)|Modifier|false|false||layernull|Eruption of skin (disorder)|Disorder|false|false||rashnull|Skin rash|Finding|false|false||rash
null|Eruptions|Finding|false|false||rash
null|Exanthema|Finding|false|false||rashnull|miconazole|Drug|false|false||Miconazole
null|miconazole|Drug|false|false||Miconazolenull|powder physical state|Drug|false|false||Powder
null|Powder dose form|Drug|false|false||Powdernull|APPL1 gene|Finding|false|false||Applnull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|Rash of groin|Finding|false|false||groin rashnull|Pelvis>Groin|Anatomy|false|false||groin
null|Inguinal region|Anatomy|false|false||groin
null|Inguinal part of abdomen|Anatomy|false|false||groinnull|Eruption of skin (disorder)|Disorder|false|false||rashnull|Skin rash|Finding|false|false||rash
null|Eruptions|Finding|false|false||rash
null|Exanthema|Finding|false|false||rashnull|insulin, regular, human|Drug|false|false||Insulin
null|Insulin [EPC]|Drug|false|false||Insulin
null|INS protein, human|Drug|false|false||Insulin
null|INS protein, human|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Insulin Drug Class|Drug|false|false||Insulin
null|Insulin Drug Class|Drug|false|false||Insulin
null|insulin, regular, human|Drug|false|false||Insulin
null|insulin, regular, human|Drug|false|false||Insulinnull|INS gene|Finding|false|false||Insulinnull|Insulin measurement|Procedure|false|false||Insulinnull|sliding scale|Procedure|false|false||Sliding Scalenull|Sliding|Finding|false|false||Slidingnull|Scale, LOINC Axis 5|Finding|false|false||Scale
null|Base Number|Finding|false|false||Scale
null|Scale - rank|Finding|false|false||Scalenull|Integumentary scale|Anatomy|false|false||Scalenull|Weight measurement scales|Device|false|false||Scalenull|Scaling|Event|false|false||Scalenull|insulin, regular, human|Drug|false|false||Insulin
null|Insulin [EPC]|Drug|false|false||Insulin
null|INS protein, human|Drug|false|false||Insulin
null|INS protein, human|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Insulin Drug Class|Drug|false|false||Insulin
null|Insulin Drug Class|Drug|false|false||Insulin
null|insulin, regular, human|Drug|false|false||Insulin
null|insulin, regular, human|Drug|false|false||Insulinnull|INS gene|Finding|false|false||Insulinnull|Insulin measurement|Procedure|false|false||Insulinnull|sliding scale|Procedure|false|false||Sliding Scalenull|Sliding|Finding|false|false||Slidingnull|Scale, LOINC Axis 5|Finding|false|false||Scale
null|Base Number|Finding|false|false||Scale
null|Scale - rank|Finding|false|false||Scalenull|Integumentary scale|Anatomy|false|false||Scalenull|Weight measurement scales|Device|false|false||Scalenull|Scaling|Event|false|false||Scalenull|insulin lispro|Drug|false|false||lispro Insulin
null|insulin lispro|Drug|false|false||lispro Insulin
null|insulin lispro|Drug|false|false||lispro Insulinnull|insulin lispro|Drug|false|false||lispro
null|insulin lispro|Drug|false|false||lispro
null|insulin lispro|Drug|false|false||lispronull|insulin, regular, human|Drug|false|false||Insulin
null|Insulin [EPC]|Drug|false|false||Insulin
null|INS protein, human|Drug|false|false||Insulin
null|INS protein, human|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Insulin Drug Class|Drug|false|false||Insulin
null|Insulin Drug Class|Drug|false|false||Insulin
null|insulin, regular, human|Drug|false|false||Insulin
null|insulin, regular, human|Drug|false|false||Insulinnull|INS gene|Finding|false|false||Insulinnull|Insulin measurement|Procedure|false|false||Insulinnull|lisinopril|Drug|false|false||Lisinopril
null|lisinopril|Drug|false|false||Lisinoprilnull|Daily|Time|false|false||DAILYnull|Hold - dosing instruction fragment|Finding|false|false||HOLD
null|hold - Data Operation|Finding|false|false||HOLDnull|Hold (action)|Event|false|false||HOLDnull|Androgen Binding Protein|Drug|false|false||SBP
null|Androgen Binding Protein|Drug|false|false||SBPnull|CCHCR1 wt Allele|Finding|false|false||SBP
null|SHBG wt Allele|Finding|false|false||SBPnull|Systolic blood pressure measurement|Procedure|false|false||SBPnull|Systolic Pressure|Attribute|false|false||SBPnull|famotidine|Drug|false|false||Famotidine
null|famotidine|Drug|false|false||Famotidinenull|Every twelve hours|Time|false|false||Q12Hnull|heparin, porcine|Drug|false|false||Heparin
null|heparin, porcine|Drug|false|false||Heparin
null|heparin, porcine|Drug|false|false||Heparin
null|heparin|Drug|false|false||Heparin
null|heparin|Drug|false|false||Heparin
null|heparin|Drug|false|false||Heparinnull|Storage Unit|Device|false|false||UNIT
null|Unit device|Device|false|false||UNITnull|Unit - NCI Thesaurus Property|LabModifier|false|false||UNIT
null|Unit of Measure|LabModifier|false|false||UNIT
null|Unit|LabModifier|false|false||UNIT
null|Enzyme Unit|LabModifier|false|false||UNITnull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|polyvinyl alcohol|Drug|false|false||polyvinyl alcoholnull|Polyvinyls|Drug|false|false||polyvinyl
null|Polyvinyls|Drug|false|false||polyvinylnull|Alcohols|Drug|false|false||alcohol
null|Alcohols|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcoholnull|Alcohol - Recreational Drug Use Code|Finding|false|false||alcoholnull|Hour|Time|false|false||hoursnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Dry Eyes brand of ocular lubricant|Drug|false|false||dry eyesnull|Dry Eye Syndromes|Disorder|false|false||dry eyes
null|Keratoconjunctivitis Sicca|Disorder|false|false||dry eyesnull|Dryness of eye|Finding|false|false||dry eyesnull|Eye|Anatomy|false|false||eyesnull|null|Attribute|false|false||eyesnull|docusate sodium|Drug|false|false||Docusate Sodium
null|docusate sodium|Drug|false|false||Docusate Sodiumnull|docusate|Drug|false|false||Docusate
null|docusate|Drug|false|false||Docusatenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|Liquid Dosage Form|Drug|false|false||Liquid
null|Liquid substance|Drug|false|false||Liquidnull|Liquid (finding)|Finding|false|false||Liquidnull|Liquid diet|Procedure|false|false||Liquidnull|Liquid (state of matter)|Modifier|false|false||Liquidnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|furosemide|Drug|false|false||Furosemide
null|furosemide|Drug|false|false||Furosemidenull|Daily|Time|false|false||DAILYnull|Hypervolemia (finding)|Finding|false|false||volume overloadnull|Volume (publication)|Finding|false|false||volumenull|Volume|LabModifier|false|false||volumenull|Check|Finding|false|false||checknull|null|Event|false|false||checknull|Electrolytes|Drug|false|false||electrolytes
null|Electrolytes|Drug|false|false||electrolytes
null|Electrolyte [EPC]|Drug|false|false||electrolytesnull|albuterol|Drug|false|false||Albuterol
null|albuterol|Drug|false|false||Albuterolnull|NEB protein, human|Drug|false|false||Neb
null|NEB protein, human|Drug|false|false||Neb
null|Nebulizer solution|Drug|false|false||Nebnull|NEB gene|Finding|false|false||Neb
null|mitotic nuclear membrane disassembly|Finding|false|false||Nebnull|NEB protein, human|Drug|false|false||NEB
null|NEB protein, human|Drug|false|false||NEB
null|Nebulizer solution|Drug|false|false||NEBnull|NEB gene|Finding|false|false||NEB
null|mitotic nuclear membrane disassembly|Finding|false|false||NEBnull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Wheezing|Finding|false|false||wheezenull|ipratropium bromide|Drug|false|false||Ipratropium Bromide
null|ipratropium bromide|Drug|false|false||Ipratropium Bromidenull|ipratropium|Drug|false|false||Ipratropium
null|ipratropium|Drug|false|false||Ipratropiumnull|Bromides|Drug|false|false||Bromidenull|Bromides measurement|Procedure|false|false||Bromidenull|NEB protein, human|Drug|false|false||Neb
null|NEB protein, human|Drug|false|false||Neb
null|Nebulizer solution|Drug|false|false||Nebnull|NEB gene|Finding|false|false||Neb
null|mitotic nuclear membrane disassembly|Finding|false|false||Nebnull|NEB protein, human|Drug|false|false||NEB
null|NEB protein, human|Drug|false|false||NEB
null|Nebulizer solution|Drug|false|false||NEBnull|NEB gene|Finding|false|false||NEB
null|mitotic nuclear membrane disassembly|Finding|false|false||NEBnull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Wheezing|Finding|false|false||wheezenull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|long-term care|Procedure|false|false||Extended Carenull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|In care (finding)|Finding|false|false||Care
null|Continuity Assessment Record and Evaluation|Finding|false|false||Carenull|care activity|Event|false|false||Carenull|ADMIN.FACILITY|Finding|false|false||Facilitynull|Facility (object)|Device|false|false||Facilitynull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Admission Level of Care Code - Acute|Finding|false|false||ACUTE
null|Acute - Triage Code|Finding|false|false||ACUTEnull|acute|Time|false|false||ACUTEnull|Respiratory Failure|Disorder|false|false||respiratory failurenull|Respiratory attachment|Finding|false|false||respiratory
null|respiratory|Finding|false|false||respiratory
null|null|Finding|false|false||respiratory
null|Respiratory specimen|Finding|false|false||respiratorynull|Respiratory rate|Attribute|false|false||respiratorynull|Failure (biologic function)|Finding|false|false||failure
null|Failure|Finding|false|false||failure
null|Personal failure|Finding|false|false||failurenull|Sepsis|Disorder|false|false||Sepsis
null|Septicemia|Disorder|false|false||Sepsisnull|Sepsis <Sepsidae>|Entity|false|false||Sepsisnull|Urinary tract|Anatomy|false|false||urinarynull|urinary|Modifier|false|false||urinarynull|Source (property) (qualifier value)|Finding|false|false||source
null|Term Source|Finding|false|false||source
null|Source|Finding|false|false||sourcenull|Recurrent|Time|false|false||Recurrent
null|Episodic|Time|false|false||Recurrentnull|Colitis|Disorder|false|false||colitisnull|Chronic - Admission Level of Care Code|Finding|false|false||CHRONICnull|Provision of recurring care for chronic illness|Procedure|false|false||CHRONICnull|chronic|Time|false|false||CHRONICnull|Hypothyroidism|Disorder|false|false||Hypothyroidismnull|Chronic anemia|Disorder|false|false||Chronic anemianull|Chronic - Admission Level of Care Code|Finding|false|false||Chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||Chronicnull|chronic|Time|false|false||Chronicnull|Anemia|Disorder|false|false||anemianull|Anemia <Anemiaceae>|Entity|false|false||anemianull|Mitral Valve Insufficiency|Disorder|false|false||Mitral regurgitationnull|mitral|Modifier|false|false||Mitralnull|Regurgitation|Finding|false|false||regurgitation
null|Regurgitates after swallowing|Finding|false|false||regurgitationnull|Regurgitation - mechanism|Phenomenon|false|false||regurgitationnull|Osteoporosis|Disorder|false|false||Osteoporosisnull|Encounter due to family history of osteoporosis|Finding|false|false||Osteoporosisnull|Sjogren's Syndrome|Disorder|false|false||Sjogren syndromenull|Syndrome|Disorder|false|false||syndromenull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|BORNHOLM EYE DISEASE|Disorder|false|false||Bednull|Bachelor of Education|Finding|false|false||Bednull|Beds|Device|false|false||Bednull|Patient Location - Bed|Modifier|false|false||Bednull|Helping Behavior|Finding|false|false||assistancenull|Assisted (qualifier value)|Modifier|false|false||assistancenull|Chairs|Device|false|false||chairnull|Chairperson|Subject|false|false||chairnull|has wheelchair at home (history)|Finding|false|false||wheelchair
null|Wheelchair Usually Used|Finding|false|false||wheelchairnull|wheelchair|Device|false|false||wheelchairnull|FBXW7-AS1 gene|Finding|false|false||Dearnull|Production Class Code - Pleasure|Finding|false|false||pleasure
null|pleasurable emotion|Finding|false|false||pleasurenull|Pleasure - Animals raised for recreation|Entity|false|false||pleasurenull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Respiratory Failure|Disorder|false|false||respiratory failurenull|Respiratory attachment|Finding|false|false||respiratory
null|respiratory|Finding|false|false||respiratory
null|null|Finding|false|false||respiratory
null|Respiratory specimen|Finding|false|false||respiratorynull|Respiratory rate|Attribute|false|false||respiratorynull|Failure (biologic function)|Finding|false|false||failure
null|Failure|Finding|false|false||failure
null|Personal failure|Finding|false|false||failurenull|Intubation (procedure)|Procedure|false|false||intubationnull|mechanical method|Finding|false|false||mechanicalnull|Mechanical Treatments|Procedure|false|false||mechanicalnull|Ventilation, function (observable entity)|Finding|false|false||ventilation
null|Respiration|Finding|false|false||ventilationnull|Assisted breathing|Procedure|false|false||ventilationnull|Environmental air flow|Phenomenon|false|false||ventilationnull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|combination - answer to question|Finding|false|false||combinationnull|combination of objects|Entity|false|false||combinationnull|Combined|Modifier|false|false||combinationnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Weakness|Finding|false|false||weakness
null|Asthenia|Finding|false|false||weaknessnull|Chronic disease|Disorder|false|false||chronic illnessnull|Reported history of chronic illness|Finding|false|false||chronic illnessnull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Illness (finding)|Finding|false|false||illnessnull|Pleural effusion (disorder)|Finding|false|false||pleural effusionsnull|Pleural Diseases|Disorder|false|false||pleuralnull|Pleura|Anatomy|false|false||pleuralnull|Pleural|Modifier|false|false||pleuralnull|effusion|Finding|false|false||effusionsnull|Pulmonary Edema|Finding|false|false||pulmonary edemanull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Lung|Anatomy|false|false||lungsnull|Urinary tract infection|Disorder|false|false||urinary tract infectionnull|Urinary tract|Anatomy|false|false||urinary tract
null|Urinary system|Anatomy|false|false||urinary tractnull|Urinary tract|Anatomy|false|false||urinarynull|urinary|Modifier|false|false||urinarynull|Tract|Anatomy|false|false||tractnull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|Sepsis|Disorder|false|false||sepsis
null|Septicemia|Disorder|false|false||sepsisnull|Sepsis <Sepsidae>|Entity|false|false||sepsisnull|Blood Circulation|Finding|false|false||bloodstreamnull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Respiratory attachment|Finding|false|false||respiratory
null|respiratory|Finding|false|false||respiratory
null|null|Finding|false|false||respiratory
null|Respiratory specimen|Finding|false|false||respiratorynull|Respiratory rate|Attribute|false|false||respiratorynull|Failure (biologic function)|Finding|false|false||failure
null|Failure|Finding|false|false||failure
null|Personal failure|Finding|false|false||failurenull|Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE|Drug|false|false||antibiotics
null|Antibiotics|Drug|false|false||antibiotics
null|Antibiotics, ophthalmologic|Drug|false|false||antibiotics
null|Antibiotics, Gynecological|Drug|false|false||antibiotics
null|antibiotics, intestinal|Drug|false|false||antibiotics
null|Antibiotic throat preparations|Drug|false|false||antibiotics
null|Antibiotics, Antitubercular|Drug|false|false||antibiotics
null|Antibiotics for systemic use|Drug|false|false||antibiotics
null|Antifungal Antibiotics, Topical|Drug|false|false||antibioticsnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Rehabilitation therapy|Procedure|false|false||rehabnull|Diagnostic Service Section ID - Physical Therapy|Finding|false|false||physical therapynull|Physical therapy|Procedure|false|false||physical therapynull|Physical therapy (field)|Title|false|false||physical therapynull|physical examination (physical finding)|Finding|false|false||physical
null|Physical|Finding|false|false||physicalnull|Physical Examination|Procedure|false|false||physicalnull|Therapy Object (animal model)|Finding|false|false||therapy
null|therapeutic aspects|Finding|false|false||therapynull|Therapeutic procedure|Procedure|false|false||therapynull|Nutrition (function)|Finding|false|false||nutrition
null|Nutritional status|Finding|false|false||nutrition
null|Nutrition outcomes|Finding|false|false||nutritionnull|Feeding and dietary regimes|Procedure|false|false||nutrition
null|Nutritional Study|Procedure|false|false||nutritionnull|Science of nutrition|Title|false|false||nutritionnull|Help document|Finding|false|false||helpnull|Assisted (qualifier value)|Modifier|false|false||helpnull|Strength (attribute)|Finding|false|false||strengthnull|Pharmaceutical Strength|LabModifier|false|false||strength
null|Physical Strength|LabModifier|false|false||strengthnull|Rehabilitation therapy|Procedure|false|false||rehabnull|Primary care provider|Subject|false|false||primary care doctornull|Location Service Code - Primary Care|Finding|false|false||primary carenull|Primary Health Care|Procedure|false|false||primary carenull|True primary (qualifier value)|Time|false|false||primarynull|Primary|Modifier|false|false||primarynull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Doctor - Title|Finding|false|false||doctornull|Physicians|Subject|false|false||doctornull|Following|Time|false|false||following
null|Status post|Time|false|false||followingnull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|famotidine|Drug|false|false||famotidine
null|famotidine|Drug|false|false||famotidinenull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Twice a day|Time|false|false||twice dailynull|Daily|Time|false|false||dailynull|Gastroesophageal reflux disease|Disorder|false|false||heartburnnull|Heartburn|Finding|false|false||heartburnnull|triamcinolone acetonide|Drug|false|false||triamcinolone acetonide
null|triamcinolone acetonide|Drug|false|false||triamcinolone acetonidenull|triamcinolone|Drug|false|false||triamcinolone
null|triamcinolone|Drug|false|false||triamcinolonenull|Emollient Cream|Drug|false|false||cream
null|Cream|Drug|false|false||cream
null|Dairy Cream|Drug|false|false||creamnull|Thrice|LabModifier|false|false||three timesnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Daily|Time|false|false||dailynull|Eruption of skin (disorder)|Disorder|false|false||rashnull|Skin rash|Finding|false|false||rash
null|Eruptions|Finding|false|false||rash
null|Exanthema|Finding|false|false||rashnull|lisinopril|Drug|false|false||lisinopril
null|lisinopril|Drug|false|false||lisinoprilnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Daily|Time|false|false||dailynull|Message Waiting Priority - High|Finding|false|false||high
null|high - ActExposureLevelCode|Finding|false|false||high
null|IPSS Risk Category High|Finding|false|false||high
null|IPSS-R Risk Category High|Finding|false|false||high
null|High (finding)|Finding|false|false||highnull|Observation Value - High|Modifier|false|false||high
null|High|Modifier|false|false||high
null|Abnormally high|Modifier|false|false||highnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|Congestive heart failure|Disorder|false|false||heart failure
null|Heart failure|Disorder|false|false||heart failurenull|Malignant neoplasm of heart|Disorder|false|false||heart
null|benign neoplasm of heart|Disorder|false|false||heartnull|HEART PROBLEM|Finding|false|false||heartnull|Chest>Heart|Anatomy|false|false||heart
null|Heart|Anatomy|false|false||heartnull|Failure (biologic function)|Finding|false|false||failure
null|Failure|Finding|false|false||failure
null|Personal failure|Finding|false|false||failurenull|Started|Modifier|false|false||STARTEDnull|docusate|Drug|false|false||docusate
null|docusate|Drug|false|false||docusatenull|Colace|Drug|false|false||Colace
null|Colace|Drug|false|false||Colacenull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Twice a day|Time|false|false||twice dailynull|Daily|Time|false|false||dailynull|Constipation|Finding|false|false||constipationnull|Continuous|Finding|false|false||CONTINUEDnull|null|Drug|false|false||vancomycin oralnull|vancomycin|Drug|false|false||vancomycin
null|vancomycin|Drug|false|false||vancomycinnull|Vancomycin measurement|Procedure|false|false||vancomycinnull|Oral Liquid Product|Drug|false|false||oral liquidnull|Oral Dosage Form|Drug|false|false||oralnull|Oral Route of Administration|Finding|false|false||oral
null|Oral (intended site)|Finding|false|false||oralnull|Oral cavity|Anatomy|false|false||oralnull|Oral|Modifier|false|false||oralnull|Liquid Dosage Form|Drug|false|false||liquid
null|Liquid substance|Drug|false|false||liquidnull|Liquid (finding)|Finding|false|false||liquidnull|Liquid diet|Procedure|false|false||liquidnull|Liquid (state of matter)|Modifier|false|false||liquidnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|6 Hours|Time|false|false||6 hoursnull|Hour|Time|false|false||hoursnull|Last|Modifier|false|false||lastnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Start brand of breakfast cereal|Drug|false|false||STARTnull|start - HtmlLinkType|Finding|false|false||STARTnull|Collagen Tile Brachytherapy|Procedure|false|false||STARTnull|Beginning|Time|false|false||STARTnull|Daily|Time|false|false||dailynull|CIAO3 gene|Finding|false|false||prnnull|As required|Time|false|false||prn
null|Pro Re Nata|Time|false|false||prnnull|Hypervolemia (finding)|Finding|false|false||volume overloadnull|Volume (publication)|Finding|false|false||volumenull|Volume|LabModifier|false|false||volumenull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions