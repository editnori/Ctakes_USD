CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|true|false||Unit
null|Unit device|Device|true|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|true|false||Unit
null|Unit of Measure|LabModifier|true|false||Unit
null|Unit|LabModifier|true|false||Unit
null|Enzyme Unit|LabModifier|true|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Pharmaceutical Preparations|Drug|false|false||MEDICINEnull|Medicine|Title|false|false||MEDICINEnull|codeine|Drug|false|false||Codeine
null|codeine|Drug|false|false||Codeinenull|Augmentin|Drug|false|false||Augmentin
null|Augmentin|Drug|false|false||Augmentinnull|Topamax|Drug|false|false||Topamax
null|Topamax|Drug|false|false||Topamaxnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Dyspnea|Finding|false|false||Shortness of Breathnull|null|Attribute|false|false||Shortness of Breathnull|Breath|Finding|false|false||Breathnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|History of cerebral aneurysm|Finding|false|false||history of cerebral aneurysmnull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Cerebral Aneurysm|Disorder|false|false||cerebral aneurysmnull|Cerebral hemisphere structure (body structure)|Anatomy|false|false||cerebral
null|Brain|Anatomy|false|false||cerebralnull|Aneurysm|Finding|false|false||aneurysmnull|Dyspnea|Finding|false|false||shortness of breathnull|null|Attribute|false|false||shortness of breathnull|Breath|Finding|false|false||breathnull|Further|Modifier|false|false||furthernull|Disease Management|Procedure|false|false||managementnull|Management Occupations|Subject|false|false||managementnull|Management procedure|Event|false|false||management
null|Administration occupational activities|Event|false|false||managementnull|Early|Time|false|false||Earliernull|Transaction counts and value totals - month|Finding|false|false||month
null|Precision - month|Finding|false|false||monthnull|month|Time|false|false||month
null|Monthly (qualifier value)|Time|false|false||monthnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|Physiologic warmth|Finding|false|false||warmth
null|Social warmth|Finding|false|false||warmthnull|Erythema|Disorder|false|false||erythemanull|Consistent with|Finding|false|false||consistent withnull|Compatible|Modifier|false|false||consistent withnull|Consistent with|Finding|false|false||consistentnull|Cellulitis|Disorder|false|false||cellulitisnull|cellulitis on exam (physical finding)|Finding|false|false||cellulitisnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|true|false||time
null|Time (foundation metadata concept)|Finding|true|false||time
null|Value type - Time|Finding|true|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|true|false||time
null|Data types - Time|Finding|true|false||time
null|null|Finding|true|false||timenull|Time|Time|true|false||timenull|Deep thrombophlebitis|Disorder|true|false||DVT
null|Deep Vein Thrombosis|Disorder|true|false||DVTnull|area DVT|Anatomy|true|false||DVTnull|null|Attribute|true|false||DVTnull|Course|Time|false|false||coursenull|cephalexin|Drug|false|false||cephalexin
null|cephalexin|Drug|false|false||cephalexinnull|Improvement|Finding|false|false||improvementnull|Erythema|Disorder|false|false||erythemanull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|2 days ago|Time|false|false||2 days agonull|2 Days|Time|false|false||2 daysnull|day|Time|false|false||daysnull|FBXW7 wt Allele|Finding|false|false||ago
null|FBXW7 gene|Finding|false|false||agonull|Dyspnea on exertion|Finding|false|false||dyspnea on exertionnull|null|Finding|false|false||dyspnea
null|Dyspnea|Finding|false|false||dyspneanull|Exertion|Finding|false|false||exertionnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|true|false||pain
null|Pain|Finding|true|false||painnull|null|Attribute|true|false||painnull|Upper Respiratory Infections|Disorder|true|false||URInull|Uniform Resource Identifier|Finding|true|false||URI
null|URI1 gene|Finding|true|false||URI
null|URI1 wt Allele|Finding|true|false||URInull|Symptoms aspect|Finding|true|false||symptoms
null|Symptoms|Finding|true|false||symptomsnull|null|Time|true|false||priornull|Deep thrombophlebitis|Disorder|true|false||DVT
null|Deep Vein Thrombosis|Disorder|true|false||DVTnull|area DVT|Anatomy|true|false||DVTnull|null|Attribute|true|false||DVTnull|Relationship modifier - Patient|Finding|true|false||patient
null|Specimen Type - Patient|Finding|true|false||patient
null|Mail Claim Party - Patient|Finding|true|false||patient
null|Report source - Patient|Finding|true|false||patient
null|null|Finding|true|false||patient
null|Disabled Person Code - Patient|Finding|true|false||patientnull|Patients|Subject|true|false||patientnull|Veterinary Patient|Entity|true|false||patientnull|Fever symptoms (finding)|Finding|true|false||fever
null|Fever|Finding|true|false||fevernull|Chills|Finding|true|false||chillsnull|Abdominal Pain|Finding|true|false||abdominal painnull|Abdomen|Anatomy|true|false||abdominalnull|Abdominal (qualifier value)|Modifier|true|false||abdominalnull|Administration Method - Pain|Finding|true|false||pain
null|Pain|Finding|true|false||painnull|null|Attribute|true|false||painnull|Intestines|Anatomy|false|false||bowelnull|Neoplasm of uncertain or unknown behavior of bladder|Disorder|false|false||bladder
null|Benign neoplasm of bladder|Disorder|false|false||bladder
null|Carcinoma in situ of bladder|Disorder|false|false||bladdernull|Procedures on bladder|Procedure|false|false||bladdernull|Urinary Bladder|Anatomy|false|false||bladdernull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|Glycation End Products, Advanced|Drug|false|false||age
null|Glycation End Products, Advanced|Drug|false|false||agenull|null|Attribute|false|false||agenull|Age|Subject|false|false||agenull|Appropriate|Modifier|false|false||appropriatenull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Screening - procedure intent|Finding|false|false||screening
null|Special screening finding|Finding|false|false||screening
null|Aspects of disease screening|Finding|false|false||screeningnull|research subject screening|Procedure|false|false||screening
null|Disease Screening|Procedure|false|false||screening
null|Screening|Procedure|false|false||screening
null|Screening for cancer|Procedure|false|false||screening
null|Screening procedure|Procedure|false|false||screeningnull|Recent|Time|true|false||recentnull|Weight Loss|Finding|true|false||weight loss
null|Losing Weight (question)|Finding|true|false||weight lossnull|Measured weight loss (observable entity)|LabModifier|true|false||weight lossnull|infant weight for previous delivery (history)|Finding|true|false||weight
null|Weight symptom (finding)|Finding|true|false||weightnull|Weighing patient|Procedure|true|false||weightnull|null|Attribute|true|false||weightnull|Body Weight|Subject|true|false||weightnull|Importance Weight|Modifier|true|false||weightnull|Weight|LabModifier|true|false||weightnull|Loss (adaptation)|Finding|true|false||lossnull|Loss (quantitative)|LabModifier|true|false||lossnull|Has patient|Finding|false|false||patient hasnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Known|Modifier|false|false||knownnull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Brain Aneurysm|Disorder|false|false||brain aneurysmnull|Brain Diseases|Disorder|false|false||brainnull|Head>Brain|Anatomy|false|false||brain
null|Brain|Anatomy|false|false||brainnull|Aneurysm|Finding|false|false||aneurysmnull|Referral category - Inpatient|Finding|false|false||inpatient
null|Patient Class - Inpatient|Finding|false|false||inpatientnull|inpatient encounter|Procedure|false|false||inpatientnull|inpatient|Subject|false|false||inpatientnull|Team|Subject|false|false||teamnull|Clinical Study Case|Finding|false|false||case
null|Case - situation|Finding|false|false||casenull|True Case Status|Modifier|false|false||casenull|Case unit dose|LabModifier|false|false||casenull|Fibrinolytic Agents|Drug|false|false||thrombolyticsnull|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparinnull|null|Time|false|false||prior tonull|null|Time|false|false||priornull|Transfer - product ownership|Finding|false|false||transfer
null|Transfer Technique|Finding|false|false||transfer
null|ActClass - transfer|Finding|false|false||transfer
null|null|Finding|false|false||transfernull|Transfer (immobility management)|Procedure|false|false||transfernull|Initial (abbreviation)|Finding|false|false||initialnull|Initially|Time|false|false||initialnull|Firstly|Modifier|false|false||initialnull|Taking vital signs|Procedure|false|false||vital signsnull|null|Attribute|false|false||vital signs
null|Vital signs|Attribute|false|false||vital signsnull|Vital High Nitrogen Enteral Nutrition|Drug|false|false||vitalnull|Vital (qualifier value)|Modifier|false|false||vitalnull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|null|Modifier|false|false||unremarkablenull|ECHO protocol|Procedure|true|false||echo
null|Extension for Community Healthcare Outcomes|Procedure|true|false||echonull|Echo <Calopterygidae>|Entity|true|false||echonull|Obvious|Modifier|true|false||obviousnull|Aspects of signs|Finding|true|false||signs
null|Physical findings|Finding|true|false||signsnull|Manufactured sign|Device|true|false||signsnull|Right side of heart|Anatomy|true|false||right heartnull|Table Cell Horizontal Align - right|Finding|true|false||rightnull|Right sided|Modifier|true|false||right
null|Right|Modifier|true|false||rightnull|Malignant neoplasm of heart|Disorder|true|false||heart
null|benign neoplasm of heart|Disorder|true|false||heartnull|HEART PROBLEM|Finding|true|false||heartnull|Chest>Heart|Anatomy|true|false||heart
null|Heart|Anatomy|true|false||heartnull|Muscle strain|Disorder|true|false||strainnull|Nature of Abnormal Testing - Strain|Finding|true|false||strain
null|Straining (finding)|Finding|true|false||strain
null|strain symptom|Finding|true|false||strain
null|Emotional Strain|Finding|true|false||strainnull|Organism Strain|Entity|true|false||strainnull|Microbiological strain|Modifier|true|false||strainnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparinnull|AML Lab Table|Finding|false|false||lab
null|LAT2 gene|Finding|false|false||lab
null|EWS Lab Table|Finding|false|false||labnull|Laboratory|Device|false|false||labnull|Labrador retriever|Entity|false|false||lab
null|Laboratory|Entity|false|false||labnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Transfer - product ownership|Finding|false|false||Transfer
null|Transfer Technique|Finding|false|false||Transfer
null|ActClass - transfer|Finding|false|false||Transfer
null|null|Finding|false|false||Transfernull|Transfer (immobility management)|Procedure|false|false||Transfernull|Oxygen nasal cannula|Device|false|false||Nasal Cannula
null|Nasal Cannula|Device|false|false||Nasal Cannulanull|Nasal brand of oxymetazoline|Drug|false|false||Nasal
null|Nasal brand of oxymetazoline|Drug|false|false||Nasal
null|Nasal dosage form|Drug|false|false||Nasalnull|Nasal Route of Administration|Finding|false|false||Nasal
null|Nasal (intended site)|Finding|false|false||Nasalnull|null|Anatomy|false|false||Nasalnull|Specimen Type - Cannula|Finding|false|false||Cannula
null|null|Finding|false|false||Cannulanull|Body Parts - Cannula|Anatomy|false|false||Cannulanull|Cannula device|Device|false|false||Cannulanull|Calamus <grasshoppers>|Entity|false|false||Cannulanull|outcomes otolaryngology breathing|Finding|false|false||breathing
null|Inspiration (function)|Finding|false|false||breathing
null|Respiration|Finding|false|false||breathingnull|null|Attribute|false|false||breathingnull|respiratory system process|Phenomenon|false|false||breathingnull|Greatly|Finding|false|false||greatlynull|Admission Level of Care Code - Improved|Finding|false|false||improved
null|Improved - answer to question|Finding|false|false||improved
null|Improved|Finding|false|false||improvednull|Better|Modifier|false|false||improvednull|Chest Pain|Finding|true|false||chest painnull|null|Attribute|true|false||chest painnull|Chest problem|Finding|true|false||chestnull|Chest|Anatomy|true|false||chest
null|Anterior thoracic region|Anatomy|true|false||chestnull|Administration Method - Pain|Finding|true|false||pain
null|Pain|Finding|true|false||painnull|null|Attribute|true|false||painnull|Cerebral Aneurysm|Disorder|false|false||CEREBRAL ANEURYSMnull|Cerebral hemisphere structure (body structure)|Anatomy|false|false||CEREBRAL
null|Brain|Anatomy|false|false||CEREBRALnull|Aneurysm|Finding|false|false||ANEURYSMnull|Incidental Findings|Finding|false|false||incidental findingnull|Incidental|Finding|false|false||incidentalnull|Experimental Finding|Finding|false|false||finding
null|Signs and Symptoms|Finding|false|false||finding
null|Finding|Finding|false|false||findingnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Dizziness|Finding|false|false||dizziness
null|Vertigo|Finding|false|false||dizzinessnull|CAT scan of head|Procedure|false|false||Head CTnull|Problems with head|Disorder|false|false||Headnull|Procedure on head|Procedure|false|false||Headnull|Structure of head of caudate nucleus|Anatomy|false|false||Head
null|Head|Anatomy|false|false||Headnull|Head Device|Device|false|false||Headnull|Infarction, Lacunar|Disorder|false|false||lacunar infarctsnull|Infarction|Finding|false|false||infarctsnull|null|Anatomy|false|false||basal ganglia
null|Basal Ganglia|Anatomy|false|false||basal ganglianull|Basal|Modifier|false|false||basalnull|Ganglia|Anatomy|false|false||ganglianull|Most Recent|Time|false|false||most recentnull|Recent|Time|false|false||recentnull|Contrast Media|Drug|true|false||contrastnull|Contrast|Modifier|true|false||contrastnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Protuberance|Anatomy|false|false||protuberancenull|Structure of genu of corpus callosum|Anatomy|false|false||genu
null|Knee|Anatomy|false|false||genunull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Code System Type - Internal|Modifier|false|false||internal
null|Internal Surface|Modifier|false|false||internal
null|Internal|Modifier|false|false||internalnull|Head+Neck>Carotid artery|Anatomy|false|false||carotid artery
null|Carotid Arteries|Anatomy|false|false||carotid artery
null|Common carotid artery|Anatomy|false|false||carotid artery
null|null|Anatomy|false|false||carotid arterynull|Carotid Arteries|Anatomy|false|false||carotidnull|Arterial system|Anatomy|false|false||artery
null|Arteries|Anatomy|false|false||arterynull|tocilizumab|Drug|false|false||MRA
null|tocilizumab|Drug|false|false||MRA
null|tocilizumab|Drug|false|false||MRAnull|Magnetic Resonance Angiography|Procedure|false|false||MRAnull|MRI-Based Angiogram|Lab|false|false||MRAnull|year|Time|false|false||yearsnull|BRCA1 gene mutation|Disorder|false|false||BRCA1 GENE MUTATIONnull|BRCA1 gene|Finding|false|false||BRCA1 GENEnull|BRCA1 gene (lab test)|Procedure|false|false||BRCA1 GENEnull|BRCA1 protein, human|Drug|false|false||BRCA1
null|BRCA1 protein, human|Drug|false|false||BRCA1null|BRCA1 gene|Finding|false|false||BRCA1null|Gene Mutation|Finding|false|false||GENE MUTATION
null|Gene Mutant|Finding|false|false||GENE MUTATIONnull|Gross Extranodal Extension|Finding|false|false||GENE
null|Genes|Finding|false|false||GENEnull|Mutation Abnormality|Disorder|false|false||MUTATIONnull|Mutation|Finding|false|false||MUTATIONnull|Chronic Obstructive Airway Disease|Disorder|false|false||CHRONIC OBSTRUCTIVE PULMONARY DISEASEnull|Chronic - Admission Level of Care Code|Finding|false|false||CHRONICnull|Provision of recurring care for chronic illness|Procedure|false|false||CHRONICnull|chronic|Time|false|false||CHRONICnull|Lung Diseases, Obstructive|Disorder|false|false||OBSTRUCTIVE PULMONARY DISEASEnull|Obstructed|Finding|false|false||OBSTRUCTIVEnull|Lung diseases|Disorder|false|false||PULMONARY DISEASEnull|History of - respiratory disease|Finding|false|false||PULMONARY DISEASEnull|Pulmonary (intended site)|Finding|false|false||PULMONARYnull|Lung|Anatomy|false|false||PULMONARYnull|null|Attribute|false|false||PULMONARYnull|Pulmonary (qualifier value)|Modifier|false|false||PULMONARYnull|Disease|Disorder|false|false||DISEASEnull|Sleep Apnea Syndromes|Disorder|false|false||SLEEP APNEAnull|SLEEP APNEA (device)|Device|false|false||SLEEP APNEAnull|Sleep brand of diphenhydramine hydrochloride|Drug|false|false||SLEEP
null|Sleep brand of diphenhydramine hydrochloride|Drug|false|false||SLEEPnull|Sleep|Finding|false|false||SLEEPnull|Apnea|Finding|false|false||APNEAnull|Colonic Polyps|Disorder|false|false||COLONIC POLYPSnull|Encounter due to family history of colonic polyps|Finding|false|false||COLONIC POLYPSnull|Colon structure (body structure)|Anatomy|false|false||COLONICnull|polyps|Disorder|false|false||POLYPSnull|null|Finding|false|false||POLYPSnull|Gastroesophageal reflux disease|Disorder|false|false||GASTROESOPHAGEAL REFLUXnull|Infantile Gastroesophageal Reflux|Finding|false|false||GASTROESOPHAGEAL REFLUX
null|Acid reflux|Finding|false|false||GASTROESOPHAGEAL REFLUXnull|gastroesophageal|Anatomy|false|false||GASTROESOPHAGEALnull|Reflux|Finding|false|false||REFLUXnull|Cancer patients and suicide and depression|Disorder|false|false||DEPRESSION
null|Mental Depression|Disorder|false|false||DEPRESSION
null|Depressive disorder|Disorder|false|false||DEPRESSION
null|Depressed mood|Disorder|false|false||DEPRESSIONnull|Depression - motion|Finding|false|false||DEPRESSION
null|null|Finding|false|false||DEPRESSIONnull|Depression - recess|Modifier|false|false||DEPRESSIONnull|Prediabetes syndrome|Disorder|false|false||PRE-DIABETESnull|Hematuria|Disorder|false|false||HEMATURIAnull|Low Back Pain|Finding|false|false||LOW BACK PAINnull|IPSS-R Risk Category Low|Finding|false|false||LOW
null|IPSS Risk Category Low|Finding|false|false||LOW
null|low confidentiality|Finding|false|false||LOWnull|Low - MessageWaitingPriority|Modifier|false|false||LOW
null|low|Modifier|false|false||LOW
null|low exposure|Modifier|false|false||LOWnull|null|LabModifier|false|false||LOWnull|Back Pain|Finding|false|false||BACK PAINnull|Administration Method - Pain|Finding|false|false||PAIN
null|Pain|Finding|false|false||PAINnull|null|Attribute|false|false||PAINnull|Varicosity|Disorder|false|false||VARICOSE VEINSnull|Varicose|Modifier|false|false||VARICOSEnull|Procedure on vein|Procedure|false|false||VEINSnull|Veins|Anatomy|false|false||VEINSnull|Scabies infestation|Disorder|false|false||SCABIESnull|Scabies <Mollusca>|Entity|false|false||SCABIESnull|Hyperlipidemia|Disorder|false|false||HYPERLIPIDEMIA
null|Hyperlipoproteinemias|Disorder|false|false||HYPERLIPIDEMIAnull|Serum lipids high (finding)|Finding|false|false||HYPERLIPIDEMIAnull|Rotator cuff syndrome|Disorder|false|false||ROTATOR CUFF TEARnull|Rotator Cuff Tears|Finding|false|false||ROTATOR CUFF TEARnull|Rotator Cuff|Anatomy|false|false||ROTATOR CUFFnull|null|Device|false|false||ROTATORnull|Cuffing (morphologic abnormality)|Finding|false|false||CUFFnull|Cuff - body part|Anatomy|false|false||CUFFnull|Cuff Device|Device|false|false||CUFFnull|Laceration|Disorder|false|false||TEAR
null|Rupture|Disorder|false|false||TEARnull|Tears (substance)|Finding|false|false||TEARnull|Tear Shape|Modifier|false|false||TEARnull|Syncope|Finding|false|false||syncopenull|Syncope <Gastrophryninae>|Entity|false|false||syncopenull|Transient Cerebral Ischemia|Disorder|true|false||TIA
null|Transient Ischemic Attack|Disorder|true|false||TIAnull|Tacca leontopetaloides|Entity|true|false||TIAnull|Carotid Arteries|Anatomy|true|false||carotidnull|Significant|Finding|true|false||significantnull|Event Seriousness - Significant|Modifier|true|false||significantnull|Stenosis|Finding|true|false||stenosisnull|Stenosis <Pimeliinae>|Entity|true|false||stenosisnull|Stenosis Morphology|Modifier|true|false||stenosisnull|ECHO protocol|Procedure|true|false||ECHO
null|Extension for Community Healthcare Outcomes|Procedure|true|false||ECHOnull|Echo <Calopterygidae>|Entity|true|false||ECHOnull|Total abdominal hysterectomy with bilateral salpingo-oophorectomy|Procedure|false|false||TAH/BSOnull|Total abdominal hysterectomy|Procedure|false|false||TAHnull|Tahitian language|Entity|false|false||TAHnull|Buthionine Sulfoximine|Drug|false|false||BSO
null|Buthionine Sulfoximine|Drug|false|false||BSO
null|Buthionine Sulfoximine|Drug|false|false||BSOnull|Cholecystectomy procedure|Procedure|false|false||CHOLECYSTECTOMYnull|Entity Name Part Type - family|Finding|true|false||family
null|Last Name|Finding|true|false||family
null|Living Arrangement - Family|Finding|true|false||family
null|Family (taxonomic)|Finding|true|false||family
null|Family Collection|Finding|true|false||familynull|Family|Subject|true|false||familynull|Deep thrombophlebitis|Disorder|true|true||DVT
null|Deep Vein Thrombosis|Disorder|true|true||DVTnull|area DVT|Anatomy|true|false||DVTnull|null|Attribute|true|true||DVTnull|Sister|Subject|false|false||sistersnull|Atrial Fibrillation|Disorder|false|true||atrial fibrillationnull|null|Attribute|false|true||atrial fibrillationnull|Atrial Fibrillation by ECG Finding|Lab|false|true||atrial fibrillationnull|Heart Atrium|Anatomy|false|false||atrialnull|Fibrillation|Disorder|false|false||fibrillationnull|On admission|Time|false|false||ON ADMISSIONnull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||GENERALnull|General medical service|Procedure|false|false||GENERALnull|Generalized|Modifier|false|false||GENERALnull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|Obesity|Disorder|false|false||obesenull|HEENT|Anatomy|false|false||HEENTnull|Pupil equal round and reacting to light|Finding|false|false||PERRLnull|Anicteric|Finding|false|false||anictericnull|Scleral Diseases|Disorder|false|false||scleranull|examination of sclera|Procedure|false|false||scleranull|Sclera|Anatomy|false|false||scleranull|Pink color|Modifier|false|false||pinknull|Malignant neoplasm of conjunctiva|Disorder|false|false||conjunctiva
null|Benign neoplasm of conjunctiva|Disorder|false|false||conjunctiva
null|Conjunctival Diseases|Disorder|false|false||conjunctivanull|Specimen Type - Conjunctiva|Finding|false|false||conjunctiva
null|null|Finding|false|false||conjunctivanull|examination of conjunctiva|Procedure|false|false||conjunctiva
null|Procedure on conjunctiva|Procedure|false|false||conjunctivanull|Structure of palpebral conjunctiva|Anatomy|false|false||conjunctiva
null|conjunctiva|Anatomy|false|false||conjunctivanull|Myelofibrosis|Disorder|false|false||MMMnull|Medial part of medial mammillary nucleus|Anatomy|false|false||MMMnull|Language Ability Proficiency - Good|Finding|false|false||good
null|Language Proficiency - Good|Finding|false|false||goodnull|Specimen Quality - Good|Modifier|false|false||good
null|Good|Modifier|false|false||goodnull|Dentition|Anatomy|false|false||dentition
null|Tooth structure|Anatomy|false|false||dentitionnull|Passive joint movement of neck (finding)|Finding|false|false||NECK
null|Neck problem|Finding|false|false||NECKnull|dendritic spine neck|Anatomy|false|false||NECK
null|Neck|Anatomy|false|false||NECKnull|Supple neck|Finding|true|false||supple necknull|Supple|Finding|true|false||supplenull|Passive joint movement of neck (finding)|Finding|true|false||neck
null|Neck problem|Finding|true|false||necknull|dendritic spine neck|Anatomy|true|false||neck
null|Neck|Anatomy|true|false||necknull|Leukocyte adhesion deficiency type 1|Disorder|true|false||LAD
null|Leukocyte adhesion deficiency|Disorder|true|false||LADnull|ITGB2 wt Allele|Finding|true|false||LAD
null|DLD gene|Finding|true|false||LADnull|Anterior descending branch of left coronary artery|Anatomy|true|false||LADnull|Ladino Language|Entity|true|false||LADnull|Jugular venous engorgement|Finding|true|false||JVDnull|Cardiac attachment|Finding|true|false||CARDIACnull|Heart|Anatomy|true|false||CARDIACnull|Cardiac - anatomy qualifier|Modifier|true|false||CARDIACnull|Heart murmur|Finding|true|false||murmursnull|Pericardial friction rub|Finding|true|false||rubsnull|Lung diseases|Disorder|false|false||LUNGnull|Lung Problem|Finding|false|false||LUNGnull|Chest>Lung|Anatomy|false|false||LUNG
null|Lung|Anatomy|false|false||LUNGnull|cetrimonium bromide|Drug|true|false||CTABnull|Wheezing|Finding|true|false||wheezesnull|Basilar Rales|Finding|true|false||rales
null|Rales|Finding|true|false||ralesnull|Rhonchi|Finding|true|false||rhonchinull|Use of accessory muscles|Finding|true|false||use of accessory musclesnull|Use of|Finding|true|false||use ofnull|Use - dosing instruction imperative|Finding|true|false||use
null|utilization qualifier|Finding|true|false||use
null|Usage|Finding|true|false||usenull|Accessory skeletal muscle|Disorder|true|false||accessory musclesnull|Accessory|Device|true|false||accessorynull|Set of muscles|Anatomy|true|false||muscles
null|Muscle (organ)|Anatomy|true|false||muscles
null|Muscle Tissue|Anatomy|true|false||musclesnull|Malignant neoplasm of abdomen|Disorder|true|false||ABDOMENnull|Abdomen problem|Finding|true|false||ABDOMENnull|Abdomen|Anatomy|true|false||ABDOMEN
null|Abdominal Cavity|Anatomy|true|false||ABDOMENnull|Protective muscle spasm|Finding|true|false||guardingnull|Hepatosplenomegaly|Finding|true|false||hepatosplenomegalynull|All extremities|Anatomy|true|false||EXTREMITIES
null|Limb structure|Anatomy|true|false||EXTREMITIESnull|Body Site Modifier - Lower|Anatomy|true|false||lowernull|Lower (action)|Event|true|false||lowernull|Lower - spatial qualifier|Modifier|true|false||lowernull|Exam|Finding|true|false||examnull|Medical Examination|Procedure|true|false||examnull|Swelling|Finding|true|false||swelling
null|Edema|Finding|true|false||swellingnull|Posterior part of right leg|Anatomy|true|false||R calfnull|Structure of calf of leg|Anatomy|true|false||calf
null|null|Anatomy|true|false||calfnull|Cattle calf (organism)|Entity|true|false||calfnull|Tender|Modifier|false|false||tendernull|Palpation|Procedure|false|false||palpationnull|null|Drug|false|false||PULSESnull|Physiologic pulse|Finding|false|false||PULSESnull|Pulse taking|Procedure|false|false||PULSESnull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false||pulsesnull|Neurology speciality|Title|false|false||NEUROnull|Neurologic (qualifier value)|Modifier|false|false||NEUROnull|Gender Status - Intact|Finding|true|false||intactnull|Intact|Modifier|true|false||intactnull|Focal|Modifier|true|false||focalnull|Deficit|Modifier|true|false||deficitsnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|true|false||SKIN
null|Skin and subcutaneous tissue disorders|Disorder|true|false||SKINnull|Skin Specimen Source Code|Finding|true|false||SKIN
null|Skin Specimen|Finding|true|false||SKINnull|Skin, Human|Anatomy|true|false||SKIN
null|Skin|Anatomy|true|false||SKINnull|Feels warm|Finding|true|false||warmnull|warming process|Phenomenon|true|false||warmnull|Well (answer to question)|Finding|true|false||wellnull|Well (container)|Device|true|false||wellnull|Microplate Well|Modifier|true|false||well
null|Good|Modifier|true|false||well
null|Healthy|Modifier|true|false||wellnull|Excoriation|Disorder|true|false||excoriationsnull|Lesion|Finding|true|false||lesionsnull|Skin rash|Finding|true|false||rashes
null|Exanthema|Finding|true|false||rashesnull|On discharge|Time|true|false||ON DISCHARGEnull|Body Substance Discharge|Finding|true|false||DISCHARGE
null|Discharge Body Fluid|Finding|true|false||DISCHARGE
null|Body Fluid Discharge|Finding|true|false||DISCHARGE
null|null|Finding|true|false||DISCHARGEnull|Patient Discharge|Procedure|true|false||DISCHARGEnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||GENERALnull|General medical service|Procedure|false|false||GENERALnull|Generalized|Modifier|false|false||GENERALnull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|Obesity|Disorder|false|false||obesenull|HEENT|Anatomy|false|false||HEENTnull|Pupil equal round and reacting to light|Finding|false|false||PERRLnull|Anicteric|Finding|false|false||anictericnull|Scleral Diseases|Disorder|false|false||scleranull|examination of sclera|Procedure|false|false||scleranull|Sclera|Anatomy|false|false||scleranull|Pink color|Modifier|false|false||pinknull|Malignant neoplasm of conjunctiva|Disorder|false|false||conjunctiva
null|Benign neoplasm of conjunctiva|Disorder|false|false||conjunctiva
null|Conjunctival Diseases|Disorder|false|false||conjunctivanull|Specimen Type - Conjunctiva|Finding|false|false||conjunctiva
null|null|Finding|false|false||conjunctivanull|examination of conjunctiva|Procedure|false|false||conjunctiva
null|Procedure on conjunctiva|Procedure|false|false||conjunctivanull|Structure of palpebral conjunctiva|Anatomy|false|false||conjunctiva
null|conjunctiva|Anatomy|false|false||conjunctivanull|Myelofibrosis|Disorder|false|false||MMMnull|Medial part of medial mammillary nucleus|Anatomy|false|false||MMMnull|Language Ability Proficiency - Good|Finding|false|false||good
null|Language Proficiency - Good|Finding|false|false||goodnull|Specimen Quality - Good|Modifier|false|false||good
null|Good|Modifier|false|false||goodnull|Dentition|Anatomy|false|false||dentition
null|Tooth structure|Anatomy|false|false||dentitionnull|Passive joint movement of neck (finding)|Finding|false|false||NECK
null|Neck problem|Finding|false|false||NECKnull|dendritic spine neck|Anatomy|false|false||NECK
null|Neck|Anatomy|false|false||NECKnull|Supple neck|Finding|true|false||supple necknull|Supple|Finding|true|false||supplenull|Passive joint movement of neck (finding)|Finding|true|false||neck
null|Neck problem|Finding|true|false||necknull|dendritic spine neck|Anatomy|true|false||neck
null|Neck|Anatomy|true|false||necknull|Leukocyte adhesion deficiency type 1|Disorder|true|false||LAD
null|Leukocyte adhesion deficiency|Disorder|true|false||LADnull|ITGB2 wt Allele|Finding|true|false||LAD
null|DLD gene|Finding|true|false||LADnull|Anterior descending branch of left coronary artery|Anatomy|true|false||LADnull|Ladino Language|Entity|true|false||LADnull|Jugular venous engorgement|Finding|true|false||JVDnull|Cardiac attachment|Finding|true|false||CARDIACnull|Heart|Anatomy|true|false||CARDIACnull|Cardiac - anatomy qualifier|Modifier|true|false||CARDIACnull|Heart murmur|Finding|true|false||murmursnull|Pericardial friction rub|Finding|true|false||rubsnull|Lung diseases|Disorder|false|false||LUNGnull|Lung Problem|Finding|false|false||LUNGnull|Chest>Lung|Anatomy|false|false||LUNG
null|Lung|Anatomy|false|false||LUNGnull|cetrimonium bromide|Drug|true|false||CTABnull|Wheezing|Finding|true|false||wheezesnull|Basilar Rales|Finding|true|false||rales
null|Rales|Finding|true|false||ralesnull|Rhonchi|Finding|true|false||rhonchinull|Use of accessory muscles|Finding|true|false||use of accessory musclesnull|Use of|Finding|true|false||use ofnull|Use - dosing instruction imperative|Finding|true|false||use
null|utilization qualifier|Finding|true|false||use
null|Usage|Finding|true|false||usenull|Accessory skeletal muscle|Disorder|true|false||accessory musclesnull|Accessory|Device|true|false||accessorynull|Set of muscles|Anatomy|true|false||muscles
null|Muscle (organ)|Anatomy|true|false||muscles
null|Muscle Tissue|Anatomy|true|false||musclesnull|Malignant neoplasm of abdomen|Disorder|true|false||ABDOMENnull|Abdomen problem|Finding|true|false||ABDOMENnull|Abdomen|Anatomy|true|false||ABDOMEN
null|Abdominal Cavity|Anatomy|true|false||ABDOMENnull|Protective muscle spasm|Finding|true|false||guardingnull|Hepatosplenomegaly|Finding|true|false||hepatosplenomegalynull|All extremities|Anatomy|true|false||EXTREMITIES
null|Limb structure|Anatomy|true|false||EXTREMITIESnull|Body Site Modifier - Lower|Anatomy|true|false||lowernull|Lower (action)|Event|true|false||lowernull|Lower - spatial qualifier|Modifier|true|false||lowernull|Exam|Finding|true|false||examnull|Medical Examination|Procedure|true|false||examnull|Swelling|Finding|true|false||swelling
null|Edema|Finding|true|false||swellingnull|Posterior part of right leg|Anatomy|true|false||R calfnull|Structure of calf of leg|Anatomy|true|false||calf
null|null|Anatomy|true|false||calfnull|Cattle calf (organism)|Entity|true|false||calfnull|Tender|Modifier|false|false||tendernull|Palpation|Procedure|false|false||palpationnull|null|Drug|false|false||PULSESnull|Physiologic pulse|Finding|false|false||PULSESnull|Pulse taking|Procedure|false|false||PULSESnull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false||pulsesnull|Neurology speciality|Title|false|false||NEUROnull|Neurologic (qualifier value)|Modifier|false|false||NEUROnull|Gender Status - Intact|Finding|true|false||intactnull|Intact|Modifier|true|false||intactnull|Focal|Modifier|true|false||focalnull|Deficit|Modifier|true|false||deficitsnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|true|false||SKIN
null|Skin and subcutaneous tissue disorders|Disorder|true|false||SKINnull|Skin Specimen Source Code|Finding|true|false||SKIN
null|Skin Specimen|Finding|true|false||SKINnull|Skin, Human|Anatomy|true|false||SKIN
null|Skin|Anatomy|true|false||SKINnull|Feels warm|Finding|true|false||warmnull|warming process|Phenomenon|true|false||warmnull|Well (answer to question)|Finding|true|false||wellnull|Well (container)|Device|true|false||wellnull|Microplate Well|Modifier|true|false||well
null|Good|Modifier|true|false||well
null|Healthy|Modifier|true|false||wellnull|Excoriation|Disorder|true|false||excoriationsnull|Lesion|Finding|true|false||lesionsnull|Skin rash|Finding|true|false||rashes
null|Exanthema|Finding|true|false||rashesnull|On discharge|Time|true|false||ON DISCHARGEnull|Body Substance Discharge|Finding|true|false||DISCHARGE
null|Discharge Body Fluid|Finding|true|false||DISCHARGE
null|Body Fluid Discharge|Finding|true|false||DISCHARGE
null|null|Finding|true|false||DISCHARGEnull|Patient Discharge|Procedure|true|false||DISCHARGEnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Primed lymphocyte test|Procedure|false|false||PLTnull|Count Dosing Unit|LabModifier|false|false||COUNT
null|Count|LabModifier|false|false||COUNTnull|Monos|Drug|false|false||MONOS
null|Mono-S|Drug|false|false||MONOS
null|Monos|Drug|false|false||MONOSnull|SARCOIDOSIS, EARLY-ONSET|Disorder|false|false||EOS
null|Familial eosinophilia|Disorder|false|false||EOSnull|PRSS33 gene|Finding|false|false||EOS
null|IKZF4 gene|Finding|false|false||EOSnull|Eos <Loriini>|Entity|false|false||EOSnull|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSEnull|Glucose measurement|Procedure|false|false||GLUCOSEnull|Glucose^1.5H post dose glucagon|Lab|false|false||GLUCOSEnull|urea|Drug|false|false||UREA
null|urea|Drug|false|false||UREA
null|urea|Drug|false|false||UREAnull|Urea measurement|Procedure|false|false||UREAnull|Sodium supplements|Drug|false|false||SODIUM
null|sodium|Drug|false|false||SODIUM
null|sodium|Drug|false|false||SODIUM
null|Sodium Drug Class|Drug|false|false||SODIUMnull|Sodium metabolic function|Finding|false|false||SODIUMnull|Sodium measurement|Procedure|false|false||SODIUMnull|Potassium Drug Class|Drug|false|false||POTASSIUM
null|Dietary Potassium|Drug|false|false||POTASSIUM
null|potassium|Drug|false|false||POTASSIUM
null|potassium|Drug|false|false||POTASSIUM
null|potassium|Drug|false|false||POTASSIUM
null|Potassium supplement|Drug|false|false||POTASSIUM
null|Potassium supplement|Drug|false|false||POTASSIUMnull|Potassium metabolic function|Finding|false|false||POTASSIUMnull|Potassium measurement|Procedure|false|false||POTASSIUMnull|chloride ion|Drug|false|false||CHLORIDE
null|Chlorides|Drug|false|false||CHLORIDEnull|Chloride metabolic function|Finding|false|false||CHLORIDEnull|Chloride measurement|Procedure|false|false||CHLORIDEnull|Total|Modifier|false|false||TOTALnull|carbon dioxide|Drug|false|false||CO2
null|carbon dioxide|Drug|false|false||CO2null|MT-CO2 gene|Finding|false|false||CO2
null|null|Finding|false|false||CO2
null|C2 wt Allele|Finding|false|false||CO2null|blood anion gap (lab test)|Procedure|false|false||ANION GAP
null|Anion gap measurement|Procedure|false|false||ANION GAPnull|Anion Gap|Attribute|false|false||ANION GAPnull|Anion gap result|Lab|false|false||ANION GAPnull|Anions|Drug|false|false||ANIONnull|Ras GTPase-Activating Protein 1, Human|Drug|false|false||GAP
null|Ras GTPase-Activating Protein 1, Human|Drug|false|false||GAP
null|GTPase-Activating Proteins|Drug|false|false||GAP
null|GTPase-Activating Proteins|Drug|false|false||GAPnull|RASA1 wt Allele|Finding|false|false||GAP
null|RASA1 gene|Finding|false|false||GAPnull|Gap (space)|Modifier|false|false||GAPnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|History of cerebral aneurysm|Finding|false|false||history of cerebral aneurysmnull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Cerebral Aneurysm|Disorder|false|false||cerebral aneurysmnull|Cerebral hemisphere structure (body structure)|Anatomy|false|false||cerebral
null|Brain|Anatomy|false|false||cerebralnull|Aneurysm|Finding|false|false||aneurysmnull|Recent|Time|false|false||recentnull|Biomaterial Treatment|Finding|false|false||treatment
null|Treating|Finding|false|false||treatment
null|therapeutic aspects|Finding|false|false||treatmentnull|treatment - ActInformationManagementReason|Procedure|false|false||treatment
null|Administration (procedure)|Procedure|false|false||treatment
null|Therapeutic procedure|Procedure|false|false||treatmentnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|Erythema|Disorder|false|false||erythemanull|Keflex|Drug|false|false||keflex
null|Keflex|Drug|false|false||keflexnull|5 Days|Time|false|false||5 daysnull|day|Time|false|false||daysnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Dyspnea|Finding|false|false||shortness of breathnull|null|Attribute|false|false||shortness of breathnull|Breath|Finding|false|false||breathnull|Pulmonary Embolism|Finding|false|false||Pulmonary embolismnull|Pulmonary (intended site)|Finding|false|false||Pulmonarynull|Lung|Anatomy|false|false||Pulmonarynull|null|Attribute|false|false||Pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||Pulmonarynull|Embolism|Finding|false|false||embolism
null|Embolus|Finding|false|false||embolismnull|Lovenox|Drug|false|false||lovenox
null|Lovenox|Drug|false|false||lovenoxnull|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarinnull|At discharge|Time|false|false||at dischargenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Dyspnea|Finding|false|false||Shortness of breathnull|null|Attribute|false|false||Shortness of breathnull|Breath|Finding|false|false||breathnull|Patient need for (contextual qualifier)|Finding|true|false||need fornull|Patient need for (contextual qualifier)|Finding|true|false||neednull|Needs|Modifier|true|false||neednull|Supplement|Finding|true|false||supplementalnull|oxygen|Drug|true|false||oxygen
null|oxygen|Drug|true|false||oxygen
null|oxygen|Drug|true|false||oxygennull|Oxygen Therapy Care|Procedure|true|false||oxygennull|Oxygen Equipment Location|Modifier|true|false||oxygennull|History of cerebral aneurysm|Finding|false|false||History of cerebral aneurysmnull|Medical History|Finding|false|false||History ofnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Cerebral Aneurysm|Disorder|false|false||cerebral aneurysmnull|Cerebral hemisphere structure (body structure)|Anatomy|false|false||cerebral
null|Brain|Anatomy|false|false||cerebralnull|Aneurysm|Finding|false|false||aneurysmnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Aneurysm|Finding|false|false||aneurysmnull|Follow - dosing instruction imperative|Finding|false|false||follow
null|Follow|Finding|false|false||follownull|Followed by|Time|false|false||follownull|CYREN gene|Finding|false|false||MRInull|Magnetic resonance imaging service|Procedure|false|false||MRI
null|Magnetic Resonance Imaging|Procedure|false|false||MRInull|Maori Language|Entity|false|false||MRInull|Last|Modifier|false|false||lastnull|size|Modifier|false|false||sizenull|size - solid dosage form|LabModifier|false|false||sizenull|Aneurysm|Finding|false|false||aneurysmnull|Consideration|Finding|false|false||considerationnull|aspirin|Drug|false|false||aspirin
null|aspirin|Drug|false|false||aspirinnull|Aneurysm|Finding|false|false||aneurysmnull|Anti-coagulant [EPC]|Drug|false|false||anti-coagulantnull|TNFSF14 protein, human|Drug|false|false||light
null|TNFSF14 protein, human|Drug|false|false||lightnull|Light - subjective measurement|Finding|false|false||light
null|TNFSF14 wt Allele|Finding|false|false||light
null|TNFSF14 gene|Finding|false|false||light
null|Light color|Finding|false|false||lightnull|Phototherapy|Procedure|false|false||lightnull|Light|Phenomenon|false|false||lightnull|Light (qualifier)|Modifier|false|false||lightnull|Aneurysm|Finding|false|false||aneurysmnull|Risk|Finding|false|false||risk ofnull|Risk|Finding|false|false||risknull|Hemorrhage|Finding|false|false||bleedingnull|Discussion (communication)|Finding|false|false||discussionnull|Discussion (procedure)|Procedure|false|false||discussionnull|Decision|Finding|false|false||decisionnull|Fixation of dental bridge|Procedure|false|false||bridgenull|Type of bridge device|Device|false|false||bridgenull|Coumadin|Drug|false|false||Coumadin
null|Coumadin|Drug|false|false||Coumadinnull|Lovenox|Drug|false|false||lovenox
null|Lovenox|Drug|false|false||lovenoxnull|Hold - dosing instruction fragment|Finding|false|false||hold
null|hold - Data Operation|Finding|false|false||holdnull|Hold (action)|Event|false|false||holdnull|aspirin|Drug|false|false||aspirin
null|aspirin|Drug|false|false||aspirinnull|tocilizumab|Drug|false|false||MRA
null|tocilizumab|Drug|false|false||MRA
null|tocilizumab|Drug|false|false||MRAnull|Magnetic Resonance Angiography|Procedure|false|false||MRAnull|MRI-Based Angiogram|Lab|false|false||MRAnull|size|Modifier|false|false||sizenull|size - solid dosage form|LabModifier|false|false||sizenull|Aneurysm|Finding|false|false||aneurysmnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|size|Modifier|false|false||sizenull|size - solid dosage form|LabModifier|false|false||sizenull|Aneurysm|Finding|false|false||aneurysmnull|Changing|Finding|true|false||changenull|Change - procedure|Procedure|true|false||changenull|Delta (difference)|LabModifier|true|false||change
null|Changed status|LabModifier|true|false||changenull|Hyperlipidemia|Disorder|false|false||Hyperlipidemia
null|Hyperlipoproteinemias|Disorder|false|false||Hyperlipidemianull|Serum lipids high (finding)|Finding|false|false||Hyperlipidemianull|atorvastatin|Drug|false|false||atorvastatin
null|atorvastatin|Drug|false|false||atorvastatinnull|Cancer patients and suicide and depression|Disorder|false|false||Depression
null|Mental Depression|Disorder|false|false||Depression
null|Depressive disorder|Disorder|false|false||Depression
null|Depressed mood|Disorder|false|false||Depressionnull|Depression - motion|Finding|false|false||Depression
null|null|Finding|false|false||Depressionnull|Depression - recess|Modifier|false|false||Depressionnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Gastroesophageal reflux disease|Disorder|false|false||GERDnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|omeprazole|Drug|false|false||omeprazole
null|omeprazole|Drug|false|false||omeprazolenull|Asthma|Disorder|false|false||Asthmanull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Reactive airway disease|Disorder|true|false||reactive airway disease
null|Chronic obstructive pulmonary disease of horses|Disorder|true|false||reactive airway diseasenull|Reactive Therapy|Procedure|true|false||reactivenull|Reactive|Modifier|true|false||reactivenull|airway disease|Disorder|true|false||airway diseasenull|Airway structure|Anatomy|true|false||airway
null|Chest>Airway|Anatomy|true|false||airwaynull|Artificial Airways|Device|true|false||airwaynull|Disease|Disorder|true|false||diseasenull|Exam|Finding|true|false||examnull|Medical Examination|Procedure|true|false||examnull|albuterol|Drug|false|false||albuterol
null|albuterol|Drug|false|false||albuterolnull|Inhaler (unit of presentation)|Finding|false|false||inhalernull|Inhaler|Device|false|false||inhalernull|Inhaler Dosing Unit|LabModifier|false|false||inhalernull|Marketing basis - Transitional|Finding|false|false||Transitionalnull|Transitional cell morphology|Modifier|false|false||Transitionalnull|Decreased Coagulation Activity [PE]|Finding|false|false||Anti-coagulationnull|Outpatient Physical Therapy Improvement in Movement and Assessment Log (OPTIMAL) Survey|Finding|false|false||optimalnull|Optimum|Modifier|false|false||optimalnull|Length|LabModifier|false|false||lengthnull|Biomaterial Treatment|Finding|false|false||treatment
null|Treating|Finding|false|false||treatment
null|therapeutic aspects|Finding|false|false||treatmentnull|treatment - ActInformationManagementReason|Procedure|false|false||treatment
null|Administration (procedure)|Procedure|false|false||treatment
null|Therapeutic procedure|Procedure|false|false||treatmentnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Cigarette smoke (substance)|Drug|false|false||Cigarette smokingnull|Cigarette smoking behavior|Finding|false|false||Cigarette smokingnull|Cigarette Dosage Form|Drug|false|false||Cigarettenull|Cigarette|Device|false|false||Cigarettenull|Location characteristic ID - Smoking|Finding|false|false||smoking
null|Smoking|Finding|false|false||smoking
null|Tobacco smoking behavior|Finding|false|false||smokingnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|On admission|Time|false|false||on admissionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|encouragement|Finding|false|false||encouragementnull|Resources|Finding|false|false||resourcesnull|Cessation of smoking|Finding|false|false||smoking cessationnull|Smoking cessation therapy|Procedure|false|false||smoking cessationnull|Location characteristic ID - Smoking|Finding|false|false||smoking
null|Smoking|Finding|false|false||smoking
null|Tobacco smoking behavior|Finding|false|false||smokingnull|Cessation|Event|false|false||cessationnull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|MEDICATION LIST|Finding|false|false||Medication listnull|Pharmaceutical Preparations|Drug|false|false||Medicationnull|medication - HL7 publishing domain|Finding|false|false||Medication
null|Medications|Finding|false|false||Medicationnull|List|Finding|false|false||list
null|Sequence Data Type|Finding|false|false||listnull|Accurate (qualifier value)|Modifier|false|false||accuratenull|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||completenull|Completion Status for valid values - Complete|Finding|false|false||complete
null|Data operation - complete|Finding|false|false||complete
null|Finish - dosing instruction imperative|Finding|false|false||completenull|Complete|Modifier|false|false||completenull|lovastatin|Drug|false|false||Lovastatin
null|lovastatin|Drug|false|false||Lovastatinnull|Oral Dosage Form|Drug|false|false||oralnull|Oral Route of Administration|Finding|false|false||oral
null|Oral (intended site)|Finding|false|false||oralnull|Oral cavity|Anatomy|false|false||oralnull|Oral|Modifier|false|false||oralnull|Daily|Time|false|false||dailynull|sertraline|Drug|false|false||Sertraline
null|sertraline|Drug|false|false||Sertralinenull|Daily|Time|false|false||DAILYnull|aspirin|Drug|false|false||Aspirin
null|aspirin|Drug|false|false||Aspirinnull|Daily|Time|false|false||DAILYnull|omeprazole|Drug|false|false||Omeprazole
null|omeprazole|Drug|false|false||Omeprazolenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|albuterol sulfate|Drug|false|false||albuterol sulfate
null|albuterol sulfate|Drug|false|false||albuterol sulfatenull|albuterol|Drug|false|false||albuterol
null|albuterol|Drug|false|false||albuterolnull|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||sulfate
null|Sulfates, Inorganic|Drug|false|false||sulfate
null|sulfate ion|Drug|false|false||sulfate
null|sulfate ion|Drug|false|false||sulfate
null|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||sulfatenull|mcg/actuation|LabModifier|false|false||mcg/actuationnull|microgram|LabModifier|false|false||mcgnull|Actuation (unit of presentation)|LabModifier|false|false||actuationnull|Inhalation Route of Administration|Finding|false|false||inhalation
null|Inspiration (function)|Finding|false|false||inhalationnull|Inhalation Dosing Unit|LabModifier|false|false||inhalationnull|CIAO3 gene|Finding|false|false||prnnull|As required|Time|false|false||prn
null|Pro Re Nata|Time|false|false||prnnull|Wheezing|Finding|false|false||wheezingnull|Vitamin D Drug Class|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|D Vitamin|Drug|false|false||Vitamin D
null|Vitamin D [EPC]|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|Vitamin D Drug Class|Drug|false|false||Vitamin Dnull|Vitamin D measurement|Procedure|false|false||Vitamin Dnull|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitaminnull|Storage Unit|Device|false|false||UNIT
null|Unit device|Device|false|false||UNITnull|Unit - NCI Thesaurus Property|LabModifier|false|false||UNIT
null|Unit of Measure|LabModifier|false|false||UNIT
null|Unit|LabModifier|false|false||UNIT
null|Enzyme Unit|LabModifier|false|false||UNITnull|Daily|Time|false|false||DAILYnull|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin Drug Class|Drug|false|false||Multivitamins
null|Multivitamin Drug Class|Drug|false|false||Multivitaminsnull|Minerals|Drug|false|false||mineralsnull|Tablet Dosage Form|Drug|false|false||TABnull|Tablet Dosing Unit|LabModifier|false|false||TABnull|Daily|Time|false|false||DAILYnull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|lovastatin|Drug|false|false||Lovastatin
null|lovastatin|Drug|false|false||Lovastatinnull|Oral Dosage Form|Drug|false|false||oralnull|Oral Route of Administration|Finding|false|false||oral
null|Oral (intended site)|Finding|false|false||oralnull|Oral cavity|Anatomy|false|false||oralnull|Oral|Modifier|false|false||oralnull|Daily|Time|false|false||dailynull|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin Drug Class|Drug|false|false||Multivitamins
null|Multivitamin Drug Class|Drug|false|false||Multivitaminsnull|Minerals|Drug|false|false||mineralsnull|Tablet Dosage Form|Drug|false|false||TABnull|Tablet Dosing Unit|LabModifier|false|false||TABnull|Daily|Time|false|false||DAILYnull|omeprazole|Drug|false|false||Omeprazole
null|omeprazole|Drug|false|false||Omeprazolenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|sertraline|Drug|false|false||Sertraline
null|sertraline|Drug|false|false||Sertralinenull|Daily|Time|false|false||DAILYnull|Vitamin D Drug Class|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|D Vitamin|Drug|false|false||Vitamin D
null|Vitamin D [EPC]|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|Vitamin D Drug Class|Drug|false|false||Vitamin Dnull|Vitamin D measurement|Procedure|false|false||Vitamin Dnull|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitaminnull|Storage Unit|Device|false|false||UNIT
null|Unit device|Device|false|false||UNITnull|Unit - NCI Thesaurus Property|LabModifier|false|false||UNIT
null|Unit of Measure|LabModifier|false|false||UNIT
null|Unit|LabModifier|false|false||UNIT
null|Enzyme Unit|LabModifier|false|false||UNITnull|Daily|Time|false|false||DAILYnull|enoxaparin sodium|Drug|false|false||Enoxaparin Sodium
null|enoxaparin sodium|Drug|false|false||Enoxaparin Sodiumnull|enoxaparin|Drug|false|false||Enoxaparin
null|enoxaparin|Drug|false|false||Enoxaparinnull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|Every twelve hours|Time|false|false||Q12Hnull|Firstly|Modifier|false|false||Firstnull|First (number)|LabModifier|false|false||Firstnull|Unit dose|LabModifier|false|false||Dose
null|Dosage|LabModifier|false|false||Dosenull|next - HtmlLinkType|Finding|false|false||Nextnull|Following|Time|false|false||Next
null|Then|Time|false|false||Nextnull|Adjacent|Modifier|false|false||Nextnull|Extended Priority Codes - Routine|Finding|false|false||Routine
null|Report priority - Routine|Finding|false|false||Routine
null|Admission Type - Routine|Finding|false|false||Routine
null|Level of Care - Routine|Finding|false|false||Routine
null|Processing priority - Routine|Finding|false|false||Routine
null|Referral priority - Routine|Finding|false|false||Routinenull|Routine coag|Procedure|false|false||Routinenull|Priority - Routine|Time|false|false||Routinenull|Routine|Modifier|false|false||Routinenull|Administration (procedure)|Procedure|false|false||Administrationnull|Administration occupational activities|Event|false|false||Administrationnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||Time
null|Time (foundation metadata concept)|Finding|false|false||Time
null|Value type - Time|Finding|false|false||Time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||Time
null|Data types - Time|Finding|false|false||Time
null|null|Finding|false|false||Timenull|Time|Time|false|false||Timenull|enoxaparin|Drug|false|false||enoxaparin
null|enoxaparin|Drug|false|false||enoxaparinnull|Hour|Time|false|false||hoursnull|Syringes|Device|false|false||Syringenull|Syringe (unit of presentation)|LabModifier|false|false||Syringe
null|Syringe Dosing Unit|LabModifier|false|false||Syringenull|refill|Finding|false|false||Refillsnull|Nicotine Transdermal Patch|Drug|false|false||Nicotine Patchnull|nicotine|Drug|false|false||Nicotine
null|nicotine|Drug|false|false||Nicotinenull|Patch - Extended Release Film|Drug|false|false||Patch
null|Human patch material|Drug|false|false||Patch
null|Body tissue patch material|Drug|false|false||Patchnull|Plaque (lesion)|Finding|false|false||Patchnull|Patch Dosage Form|Device|false|false||Patch
null|Surgical patch|Device|false|false||Patchnull|Patch (unit of presentation)|LabModifier|false|false||Patch
null|Patch Dosing Unit|LabModifier|false|false||Patchnull|Daily|Time|false|false||DAILYnull|nicotine|Drug|false|false||nicotine
null|nicotine|Drug|false|false||nicotinenull|Nicoderm C-Q|Drug|false|false||Nicoderm CQ
null|Nicoderm C-Q|Drug|false|false||Nicoderm CQnull|Nicoderm|Drug|false|false||Nicoderm
null|Nicoderm|Drug|false|false||Nicodermnull|Hour|Time|false|false||hournull|Apply (administration method)|Finding|false|false||Apply
null|Apply (instruction)|Finding|false|false||Apply
null|null|Finding|false|false||Apply
null|Apply|Finding|false|false||Applynull|Patch - Extended Release Film|Drug|false|false||patch
null|Human patch material|Drug|false|false||patch
null|Body tissue patch material|Drug|false|false||patchnull|Plaque (lesion)|Finding|false|false||patchnull|Patch Dosage Form|Device|false|false||patch
null|Surgical patch|Device|false|false||patchnull|Patch (unit of presentation)|LabModifier|false|false||patch
null|Patch Dosing Unit|LabModifier|false|false||patchnull|Daily|Time|false|false||dailynull|Patch - Extended Release Film|Drug|false|false||Patch
null|Human patch material|Drug|false|false||Patch
null|Body tissue patch material|Drug|false|false||Patchnull|Plaque (lesion)|Finding|false|false||Patchnull|Patch Dosage Form|Device|false|false||Patch
null|Surgical patch|Device|false|false||Patchnull|Patch (unit of presentation)|LabModifier|false|false||Patch
null|Patch Dosing Unit|LabModifier|false|false||Patchnull|refill|Finding|false|false||Refillsnull|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarinnull|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarinnull|Coumadin|Drug|false|false||Coumadin
null|Coumadin|Drug|false|false||Coumadinnull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|PRSS30P gene|Finding|false|false||Dispnull|Dispense (activity)|Event|false|false||Dispnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|albuterol sulfate|Drug|false|false||albuterol sulfate
null|albuterol sulfate|Drug|false|false||albuterol sulfatenull|albuterol|Drug|false|false||albuterol
null|albuterol|Drug|false|false||albuterolnull|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||sulfate
null|Sulfates, Inorganic|Drug|false|false||sulfate
null|sulfate ion|Drug|false|false||sulfate
null|sulfate ion|Drug|false|false||sulfate
null|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||sulfatenull|mcg/actuation|LabModifier|false|false||mcg/actuationnull|microgram|LabModifier|false|false||mcgnull|Actuation (unit of presentation)|LabModifier|false|false||actuationnull|Inhalation Route of Administration|Finding|false|false||inhalation
null|Inspiration (function)|Finding|false|false||inhalationnull|Inhalation Dosing Unit|LabModifier|false|false||inhalationnull|CIAO3 gene|Finding|false|false||prnnull|As required|Time|false|false||prn
null|Pro Re Nata|Time|false|false||prnnull|Wheezing|Finding|false|false||wheezingnull|Referral category - Outpatient|Finding|false|false||Outpatient
null|Patient Class - Outpatient|Finding|false|false||Outpatientnull|Outpatients|Subject|false|false||Outpatientnull|AML Lab Table|Finding|false|false||Lab
null|LAT2 gene|Finding|false|false||Lab
null|EWS Lab Table|Finding|false|false||Labnull|Laboratory|Device|false|false||Labnull|Labrador retriever|Entity|false|false||Lab
null|Laboratory|Entity|false|false||Labnull|Work|Event|false|false||Worknull|Integrated Neuromusculoskeletal Release|Procedure|false|false||INR
null|International Normalized Ratio|Procedure|false|false||INRnull|Coagulation tissue factor induced.INR|Attribute|false|false||INRnull|ICD-9|Finding|false|false||ICD-9
null|International Classification of Diseases, Ninth Revision|Finding|false|false||ICD-9null|Disruptive, Impulse Control, and Conduct Disorders|Disorder|false|false||ICD
null|Type II Mucolipidosis|Disorder|false|false||ICDnull|International Classification of Diseases|Finding|false|false||ICD
null|GNPTAB wt Allele|Finding|false|false||ICDnull|Icd Regimen|Procedure|false|false||ICDnull|between lunch and dinner|Time|false|false||ICDnull|What subject filter - Result|Finding|false|false||result
null|Result|Finding|false|false||result
null|Experimental Result|Finding|false|false||resultnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|null|Attribute|false|false||Primary Diagnosisnull|Principal diagnosis|Modifier|false|false||Primary Diagnosisnull|True primary (qualifier value)|Time|false|false||Primarynull|Primary|Modifier|false|false||Primarynull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Pulmonary Embolism|Finding|false|false||Pulmonary embolismnull|Pulmonary (intended site)|Finding|false|false||Pulmonarynull|Lung|Anatomy|false|false||Pulmonarynull|null|Attribute|false|false||Pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||Pulmonarynull|Embolism|Finding|false|false||embolism
null|Embolus|Finding|false|false||embolismnull|Secondary diagnosis|Finding|false|false||Secondary Diagnosisnull|null|Attribute|false|false||Secondary Diagnosisnull|Neoplasm Metastasis|Disorder|false|false||Secondarynull|metastatic qualifier|Finding|false|false||Secondarynull|Secondary to|Modifier|false|false||Secondarynull|second (number)|LabModifier|false|false||Secondarynull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Superficial Thrombophlebitis|Disorder|false|false||Superficial thrombophlebitisnull|Superficial|Modifier|false|false||Superficialnull|Thrombophlebitis|Finding|false|false||thrombophlebitisnull|null|Attribute|false|false||Primary Diagnosisnull|Principal diagnosis|Modifier|false|false||Primary Diagnosisnull|True primary (qualifier value)|Time|false|false||Primarynull|Primary|Modifier|false|false||Primarynull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Pulmonary Embolism|Finding|false|false||Pulmonary embolismnull|Pulmonary (intended site)|Finding|false|false||Pulmonarynull|Lung|Anatomy|false|false||Pulmonarynull|null|Attribute|false|false||Pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||Pulmonarynull|Embolism|Finding|false|false||embolism
null|Embolus|Finding|false|false||embolismnull|Secondary diagnosis|Finding|false|false||Secondary Diagnosisnull|null|Attribute|false|false||Secondary Diagnosisnull|Neoplasm Metastasis|Disorder|false|false||Secondarynull|metastatic qualifier|Finding|false|false||Secondarynull|Secondary to|Modifier|false|false||Secondarynull|second (number)|LabModifier|false|false||Secondarynull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Superficial Thrombophlebitis|Disorder|false|false||Superficial thrombophlebitisnull|Superficial|Modifier|false|false||Superficialnull|Thrombophlebitis|Finding|false|false||thrombophlebitisnull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Coordination of Benefits - Independent|Finding|false|false||Independent
null|Religious Affiliation - Independent|Finding|false|false||Independent
null|Independence|Finding|false|false||Independent
null|Independently able|Finding|false|false||Independentnull|FBXW7-AS1 gene|Finding|false|false||Dearnull|Production Class Code - Pleasure|Finding|false|false||pleasure
null|pleasurable emotion|Finding|false|false||pleasurenull|Pleasure - Animals raised for recreation|Entity|false|false||pleasurenull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Embolism|Finding|false|false||embolism
null|Embolus|Finding|false|false||embolismnull|Blood Clot|Finding|false|false||blood clot
null|Thrombus|Finding|false|false||blood clotnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|In Blood|Finding|false|false||blood
null|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||bloodnull|clotrimazole|Drug|false|false||clot
null|clotrimazole|Drug|false|false||clotnull|Blood Clot|Finding|false|false||clotnull|Lung|Anatomy|false|false||lungsnull|Blood Clot|Finding|false|false||blood clot
null|Thrombus|Finding|false|false||blood clotnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|clotrimazole|Drug|false|false||clot
null|clotrimazole|Drug|false|false||clotnull|Blood Clot|Finding|false|false||clotnull|Pharmaceutical Preparations|Drug|false|false||medicinenull|Medicine|Title|false|false||medicinenull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Primary care provider|Subject|false|false||primary care doctornull|Location Service Code - Primary Care|Finding|false|false||primary carenull|Primary Health Care|Procedure|false|false||primary carenull|True primary (qualifier value)|Time|false|false||primarynull|Primary|Modifier|false|false||primarynull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Doctor - Title|Finding|false|false||doctornull|Physicians|Subject|false|false||doctornull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|month|Time|false|false||monthsnull|Neurosurgeon|Subject|false|false||neurosurgeonnull|Aneurysm|Finding|false|false||aneurysmnull|Repeat Object|Finding|false|false||repeat
null|Repeat|Finding|false|false||repeatnull|Repeat Pattern|Time|false|false||repeatnull|CYREN gene|Finding|false|false||MRInull|Magnetic resonance imaging service|Procedure|false|false||MRI
null|Magnetic Resonance Imaging|Procedure|false|false||MRInull|Maori Language|Entity|false|false||MRInull|Brain Diseases|Disorder|false|false||brainnull|Head>Brain|Anatomy|false|false||brain
null|Brain|Anatomy|false|false||brainnull|CYREN gene|Finding|true|false||MRInull|Magnetic resonance imaging service|Procedure|true|false||MRI
null|Magnetic Resonance Imaging|Procedure|true|false||MRInull|Maori Language|Entity|true|false||MRInull|size|Modifier|true|false||sizenull|size - solid dosage form|LabModifier|true|false||sizenull|Still|Disorder|false|false||stillnull|size|Modifier|false|false||sizenull|size - solid dosage form|LabModifier|false|false||sizenull|Continuous|Finding|false|false||continuednull|Recovery - healing process|Finding|false|false||recoverynull|null|Event|false|false||recoverynull|recovery - adjustment|LabModifier|false|false||recoverynull|Team|Subject|false|false||Teamnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions