 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|25,29
No|30,32
:|32,33
_|36,37
_|37,38
_|38,39
<EOL>|39,40
<EOL>|41,42
Admission|42,51
Date|52,56
:|56,57
_|59,60
_|60,61
_|61,62
Discharge|76,85
Date|86,90
:|90,91
_|94,95
_|95,96
_|96,97
<EOL>|97,98
<EOL>|99,100
Date|100,104
of|105,107
Birth|108,113
:|113,114
_|116,117
_|117,118
_|118,119
Sex|132,135
:|135,136
F|139,140
<EOL>|140,141
<EOL>|142,143
Service|143,150
:|150,151
MEDICINE|152,160
<EOL>|160,161
<EOL>|162,163
No|175,177
Known|178,183
Allergies|184,193
/|194,195
Adverse|196,203
Drug|204,208
Reactions|209,218
<EOL>|218,219
<EOL>|220,221
Attending|221,230
:|230,231
_|232,233
_|233,234
_|234,235
.|235,236
<EOL>|236,237
<EOL>|238,239
s|256,257
/|257,258
p|258,259
tachyarrhythmia|260,275
<EOL>|275,276
<EOL>|277,278
Major|278,283
Surgical|284,292
or|293,295
Invasive|296,304
Procedure|305,314
:|314,315
<EOL>|315,316
None|316,320
<EOL>|320,321
<EOL>|321,322
<EOL>|323,324
_|352,353
_|353,354
_|354,355
yo|356,358
F|359,360
smoker|361,367
with|368,372
PMH|373,376
of|377,379
asthma|380,386
/|386,387
COPD|387,391
on|392,394
theophylline|395,407
,|407,408
CAD|409,412
,|412,413
<EOL>|414,415
HTN|415,418
,|418,419
hyperlipidemia|420,434
,|434,435
and|436,439
atypical|440,448
chest|449,454
pain|455,459
presenting|460,470
with|471,475
<EOL>|476,477
malaise|477,484
and|485,488
SOB|489,492
during|493,499
an|500,502
episode|503,510
of|511,513
tachyarrythmia|514,528
at|529,531
home|532,536
<EOL>|537,538
which|538,543
has|544,547
since|548,553
resolved|554,562
.|562,563
Pt|565,567
recalls|568,575
that|576,580
she|581,584
took|585,589
her|590,593
VS|594,596
on|597,599
<EOL>|600,601
the|601,604
telehealth|605,615
monitor|616,623
,|623,624
then|625,629
nurse|630,635
called|636,642
and|643,646
asked|647,652
her|653,656
to|657,659
<EOL>|660,661
recheck|661,668
them|669,673
.|673,674
_|676,677
_|677,678
_|678,679
services|680,688
came|689,693
and|694,697
measured|698,706
HR|707,709
at|710,712
110s|713,717
,|717,718
but|719,722
pt|723,725
<EOL>|726,727
was|727,730
without|731,738
CP|739,741
,|741,742
SOB|743,746
,|746,747
visual|748,754
sx|755,757
,|757,758
HA|759,761
,|761,762
palps|763,768
.|768,769
Also|771,775
denies|776,782
F|783,784
/|784,785
C|785,786
,|786,787
<EOL>|788,789
N|789,790
/|790,791
V|791,792
,|792,793
abd|794,797
pain|798,802
,|802,803
change|804,810
in|811,813
bowel|814,819
or|820,822
bladder|823,830
.|830,831
Per|833,836
her|837,840
PCP|841,844
,|844,845
_|846,847
_|847,848
_|848,849
<EOL>|850,851
_|851,852
_|852,853
_|853,854
,|854,855
the|856,859
patient|860,867
does|868,872
have|873,877
a|878,879
history|880,887
of|888,890
tachyarrythmias|891,906
even|907,911
<EOL>|912,913
though|913,919
the|920,923
patient|924,931
denies|932,938
this|939,943
history|944,951
.|951,952
She|954,957
also|958,962
took|963,967
<EOL>|968,969
theophylline|969,981
for|982,985
some|986,990
time|991,995
,|995,996
although|997,1005
it|1006,1008
is|1009,1011
not|1012,1015
on|1016,1018
her|1019,1022
med|1023,1026
list|1027,1031
<EOL>|1032,1033
and|1033,1036
she|1037,1040
states|1041,1047
she|1048,1051
has|1052,1055
n't|1055,1058
taken|1059,1064
it|1065,1067
since|1068,1073
_|1074,1075
_|1075,1076
_|1076,1077
.|1077,1078
However|1080,1087
,|1087,1088
PCP|1089,1092
<EOL>|1093,1094
concern|1094,1101
is|1102,1104
that|1105,1109
the|1110,1113
theophylline|1114,1126
may|1127,1130
be|1131,1133
contributing|1134,1146
.|1146,1147
Recent|1149,1155
<EOL>|1156,1157
stress|1157,1163
test|1164,1168
with|1169,1173
reversible|1174,1184
lesion|1185,1191
being|1192,1197
treated|1198,1205
conservatively|1206,1220
.|1220,1221
<EOL>|1222,1223
<EOL>|1226,1227
.|1227,1228
<EOL>|1228,1229
In|1229,1231
ED|1232,1234
VS|1235,1237
were|1238,1242
98.8|1243,1247
78|1248,1250
154|1251,1254
/|1254,1255
82|1255,1257
20|1258,1260
95|1261,1263
%|1263,1264
.|1264,1265
Has|1267,1270
CXR|1271,1274
in|1275,1277
ED|1278,1280
which|1281,1286
was|1287,1290
<EOL>|1291,1292
unremarkable|1292,1304
.|1304,1305
Transfer|1307,1315
VS|1316,1318
were|1319,1323
HR|1324,1326
=|1326,1327
60|1327,1329
,|1329,1330
BP|1331,1333
=|1333,1334
126|1334,1337
/|1337,1338
75|1338,1340
,|1340,1341
RR|1342,1344
=|1344,1345
18|1345,1347
,|1347,1348
POx|1349,1352
=|1352,1353
94|1353,1355
%|1355,1356
<EOL>|1357,1358
RA|1358,1360
<EOL>|1360,1361
.|1361,1362
<EOL>|1362,1363
On|1363,1365
the|1366,1369
floor|1370,1375
,|1375,1376
pt|1377,1379
asymptomatic|1380,1392
and|1393,1396
feels|1397,1402
well|1403,1407
.|1407,1408
Only|1410,1414
upset|1415,1420
<EOL>|1421,1422
because|1422,1429
she|1430,1433
's|1433,1435
been|1436,1440
in|1441,1443
the|1444,1447
hospital|1448,1456
every|1457,1462
month|1463,1468
so|1469,1471
far|1472,1475
this|1476,1480
year|1481,1485
.|1485,1486
<EOL>|1486,1487
<EOL>|1487,1488
<EOL>|1489,1490
-|1512,1513
ASTHMA|1513,1519
<EOL>|1522,1523
-|1523,1524
HYPERTENSION|1524,1536
<EOL>|1539,1540
-|1540,1541
HYPERLIPIDEMIA|1541,1555
<EOL>|1558,1559
-|1559,1560
HEADACHE|1560,1568
<EOL>|1571,1572
-|1572,1573
OSTEOARTHRITIS|1573,1587
<EOL>|1590,1591
-|1591,1592
ATYPICAL|1592,1600
CHEST|1601,1606
PAIN|1607,1611
<EOL>|1614,1615
-|1615,1616
TOBACCO|1616,1623
ABUSE|1624,1629
<EOL>|1632,1633
-|1633,1634
ABNORMAL|1634,1642
CHEST|1643,1648
XRAY|1649,1653
<EOL>|1656,1657
-|1657,1658
COPD|1658,1662
<EOL>|1664,1665
<EOL>|1665,1666
<EOL>|1667,1668
:|1682,1683
<EOL>|1683,1684
_|1684,1685
_|1685,1686
_|1686,1687
<EOL>|1687,1688
:|1702,1703
<EOL>|1703,1704
Mother|1704,1710
:|1710,1711
_|1712,1713
_|1713,1714
_|1714,1715
,|1715,1716
HTN|1717,1720
<EOL>|1722,1723
Father|1723,1729
:|1729,1730
_|1731,1732
_|1732,1733
_|1733,1734
CA|1735,1737
<EOL>|1739,1740
Brother|1740,1747
:|1747,1748
CA|1749,1751
?|1751,1752
<EOL>|1754,1755
Brother|1755,1762
:|1762,1763
_|1764,1765
_|1765,1766
_|1766,1767
<EOL>|1768,1769
<EOL>|1769,1770
<EOL>|1771,1772
Physical|1772,1780
_|1781,1782
_|1782,1783
_|1783,1784
:|1784,1785
<EOL>|1785,1786
ADMISSION|1786,1795
PEx|1796,1799
:|1799,1800
<EOL>|1800,1801
VS|1801,1803
:|1803,1804
97.9|1805,1809
,|1809,1810
155|1811,1814
/|1814,1815
90|1815,1817
,|1817,1818
64|1819,1821
,|1821,1822
16|1823,1825
@|1825,1826
94|1826,1828
%|1828,1829
(|1829,1830
RA|1830,1832
)|1832,1833
<EOL>|1833,1834
GA|1834,1836
:|1836,1837
AOx3|1838,1842
,|1842,1843
NAD|1844,1847
<EOL>|1847,1848
HEENT|1848,1853
:|1853,1854
PERRLA|1856,1862
.|1862,1863
MMM|1864,1867
.|1867,1868
no|1869,1871
LAD|1872,1875
.|1875,1876
no|1877,1879
JVD|1880,1883
.|1883,1884
neck|1885,1889
supple|1890,1896
.|1896,1897
<EOL>|1898,1899
Cards|1899,1904
:|1904,1905
PMI|1906,1909
palpable|1910,1918
at|1919,1921
_|1922,1923
_|1923,1924
_|1924,1925
IC|1926,1928
space|1929,1934
.|1934,1935
No|1936,1938
RVH|1939,1942
.|1942,1943
RRR|1944,1947
S1|1948,1950
/|1950,1951
S2|1951,1953
heard|1954,1959
.|1959,1960
<EOL>|1961,1962
no|1962,1964
murmurs|1965,1972
/|1972,1973
gallops|1973,1980
/|1980,1981
rubs|1981,1985
.|1985,1986
<EOL>|1986,1987
Pulm|1987,1991
:|1991,1992
scattered|1993,2002
exp|2003,2006
wheezing|2007,2015
with|2016,2020
minimal|2021,2028
air|2029,2032
movment|2033,2040
<EOL>|2040,2041
Abd|2041,2044
:|2044,2045
soft|2046,2050
,|2050,2051
NT|2052,2054
,|2054,2055
+|2056,2057
BS|2057,2059
.|2059,2060
no|2061,2063
g|2064,2065
/|2065,2066
rt|2066,2068
.|2068,2069
<EOL>|2069,2070
Extremities|2070,2081
:|2081,2082
wwp|2083,2086
,|2086,2087
no|2088,2090
edema|2091,2096
.|2096,2097
DPs|2098,2101
,|2101,2102
PTs|2103,2106
2|2107,2108
+|2108,2109
.|2109,2110
<EOL>|2110,2111
Skin|2111,2115
:|2115,2116
no|2117,2119
rashes|2120,2126
,|2126,2127
eccymoses|2128,2137
,|2137,2138
lesions|2139,2146
<EOL>|2147,2148
Neuro|2148,2153
/|2153,2154
Psych|2154,2159
:|2159,2160
CNs|2161,2164
II|2165,2167
-|2167,2168
XII|2168,2171
intact|2172,2178
.|2178,2179
_|2180,2181
_|2181,2182
_|2182,2183
strength|2184,2192
in|2193,2195
muscle|2196,2202
groups|2203,2209
<EOL>|2210,2211
tested|2211,2217
,|2217,2218
sensation|2219,2228
symmetric|2229,2238
.|2238,2239
<EOL>|2240,2241
<EOL>|2241,2242
DISCHARGE|2242,2251
PEx|2252,2255
:|2255,2256
<EOL>|2256,2257
<EOL>|2257,2258
<EOL>|2259,2260
Pertinent|2260,2269
Results|2270,2277
:|2277,2278
<EOL>|2278,2279
Relevant|2279,2287
and|2288,2291
representative|2292,2306
labs|2307,2311
:|2311,2312
<EOL>|2312,2313
CBC|2313,2316
and|2317,2320
coags|2321,2326
:|2326,2327
<EOL>|2327,2328
-|2328,2329
_|2329,2330
_|2330,2331
_|2331,2332
03|2333,2335
:|2335,2336
30PM|2336,2340
BLOOD|2341,2346
WBC|2347,2350
-|2350,2351
6.7|2351,2354
RBC|2355,2358
-|2358,2359
4|2359,2360
.|2360,2361
40|2361,2363
Hgb|2364,2367
-|2367,2368
13.2|2368,2372
Hct|2373,2376
-|2376,2377
38.9|2377,2381
<EOL>|2382,2383
MCV|2383,2386
-|2386,2387
88|2387,2389
MCH|2390,2393
-|2393,2394
29.9|2394,2398
MCHC|2399,2403
-|2403,2404
33.9|2404,2408
RDW|2409,2412
-|2412,2413
15|2413,2415
.|2415,2416
7|2416,2417
*|2417,2418
Plt|2419,2422
_|2423,2424
_|2424,2425
_|2425,2426
<EOL>|2426,2427
-|2427,2428
_|2428,2429
_|2429,2430
_|2430,2431
05|2432,2434
:|2434,2435
55AM|2435,2439
BLOOD|2440,2445
WBC|2446,2449
-|2449,2450
5.9|2450,2453
RBC|2454,2457
-|2457,2458
4|2458,2459
.|2459,2460
32|2460,2462
Hgb|2463,2466
-|2466,2467
12.8|2467,2471
Hct|2472,2475
-|2475,2476
38.4|2476,2480
<EOL>|2481,2482
MCV|2482,2485
-|2485,2486
89|2486,2488
MCH|2489,2492
-|2492,2493
29.6|2493,2497
MCHC|2498,2502
-|2502,2503
33.2|2503,2507
RDW|2508,2511
-|2511,2512
15|2512,2514
.|2514,2515
6|2515,2516
*|2516,2517
Plt|2518,2521
_|2522,2523
_|2523,2524
_|2524,2525
<EOL>|2525,2526
-|2526,2527
_|2527,2528
_|2528,2529
_|2529,2530
03|2531,2533
:|2533,2534
30PM|2534,2538
BLOOD|2539,2544
_|2545,2546
_|2546,2547
_|2547,2548
PTT|2549,2552
-|2552,2553
26.2|2553,2557
_|2558,2559
_|2559,2560
_|2560,2561
<EOL>|2561,2562
<EOL>|2562,2563
Chem|2563,2567
:|2567,2568
<EOL>|2568,2569
-|2569,2570
_|2570,2571
_|2571,2572
_|2572,2573
03|2574,2576
:|2576,2577
30PM|2577,2581
BLOOD|2582,2587
Glucose|2588,2595
-|2595,2596
105|2596,2599
*|2599,2600
UreaN|2601,2606
-|2606,2607
18|2607,2609
Creat|2610,2615
-|2615,2616
0.9|2616,2619
Na|2620,2622
-|2622,2623
139|2623,2626
<EOL>|2627,2628
K|2628,2629
-|2629,2630
3.5|2630,2633
Cl|2634,2636
-|2636,2637
101|2637,2640
HCO3|2641,2645
-|2645,2646
31|2646,2648
<EOL>|2649,2650
-|2650,2651
_|2651,2652
_|2652,2653
_|2653,2654
05|2655,2657
:|2657,2658
55AM|2658,2662
BLOOD|2663,2668
Glucose|2669,2676
-|2676,2677
101|2677,2680
*|2680,2681
UreaN|2682,2687
-|2687,2688
20|2688,2690
Creat|2691,2696
-|2696,2697
0.9|2697,2700
Na|2701,2703
-|2703,2704
139|2704,2707
<EOL>|2708,2709
K|2709,2710
-|2710,2711
4.2|2711,2714
Cl|2715,2717
-|2717,2718
99|2718,2720
HCO3|2721,2725
-|2725,2726
32|2726,2728
<EOL>|2728,2729
<EOL>|2729,2730
CEs|2730,2733
:|2733,2734
<EOL>|2734,2735
-|2735,2736
_|2736,2737
_|2737,2738
_|2738,2739
03|2740,2742
:|2742,2743
30PM|2743,2747
BLOOD|2748,2753
cTropnT|2754,2761
-|2761,2762
<|2762,2763
0|2763,2764
.|2764,2765
01|2765,2767
<EOL>|2767,2768
-|2768,2769
_|2769,2770
_|2770,2771
_|2771,2772
09|2773,2775
:|2775,2776
10PM|2776,2780
BLOOD|2781,2786
CK|2787,2789
-|2789,2790
MB|2790,2792
-|2792,2793
4|2793,2794
cTropnT|2795,2802
-|2802,2803
<|2803,2804
0|2804,2805
.|2805,2806
01|2806,2808
<EOL>|2808,2809
-|2809,2810
_|2810,2811
_|2811,2812
_|2812,2813
05|2814,2816
:|2816,2817
55AM|2817,2821
BLOOD|2822,2827
CK|2828,2830
-|2830,2831
MB|2831,2833
-|2833,2834
3|2834,2835
cTropnT|2836,2843
-|2843,2844
<|2844,2845
0|2845,2846
.|2846,2847
01|2847,2849
<EOL>|2849,2850
<EOL>|2850,2851
Misc|2851,2855
:|2855,2856
<EOL>|2856,2857
-|2857,2858
_|2858,2859
_|2859,2860
_|2860,2861
05|2862,2864
:|2864,2865
55AM|2865,2869
BLOOD|2870,2875
Triglyc|2876,2883
-|2883,2884
96|2884,2886
HDL|2887,2890
-|2890,2891
50|2891,2893
CHOL|2894,2898
/|2898,2899
HD|2899,2901
-|2901,2902
3.2|2902,2905
LDLcalc|2906,2913
-|2913,2914
90|2914,2916
<EOL>|2917,2918
Cholest|2918,2925
-|2925,2926
159|2926,2929
<EOL>|2929,2930
<EOL>|2931,2932
To|2955,2957
Do|2958,2960
:|2960,2961
<EOL>|2961,2962
1|2962,2963
)|2963,2964
follow|2965,2971
-|2971,2972
up|2972,2974
theophylline|2975,2987
level|2988,2993
<EOL>|2993,2994
_|2994,2995
_|2995,2996
_|2996,2997
yo|2998,3000
F|3001,3002
smoker|3003,3009
with|3010,3014
PMH|3015,3018
of|3019,3021
asthma|3022,3028
/|3028,3029
COPD|3029,3033
managed|3034,3041
with|3042,3046
theophylline|3047,3059
<EOL>|3060,3061
until|3061,3066
_|3067,3068
_|3068,3069
_|3069,3070
when|3071,3075
theophylline|3076,3088
was|3089,3092
discontinued|3093,3105
because|3106,3113
of|3114,3116
<EOL>|3117,3118
tachycardia|3118,3129
,|3129,3130
CAD|3131,3134
,|3134,3135
HTN|3136,3139
,|3139,3140
and|3141,3144
hyperlipidemia|3145,3159
who|3160,3163
presented|3164,3173
from|3174,3178
<EOL>|3179,3180
home|3180,3184
with|3185,3189
asymptomatic|3190,3202
tachyarrythmia|3203,3217
.|3217,3218
<EOL>|3218,3219
.|3219,3220
<EOL>|3222,3223
ACTIVE|3223,3229
ISSUES|3230,3236
:|3236,3237
<EOL>|3237,3238
.|3238,3239
<EOL>|3239,3240
#|3240,3241
Tachycarrhymia|3242,3256
in|3257,3259
context|3260,3267
of|3268,3270
recent|3271,3277
inducible|3278,3287
ischemia|3288,3296
seen|3297,3301
on|3302,3304
<EOL>|3305,3306
ECHO|3306,3310
stress|3311,3317
test|3318,3322
(|3323,3324
_|3324,3325
_|3325,3326
_|3326,3327
)|3327,3328
:|3328,3329
At|3331,3333
the|3334,3337
time|3338,3342
of|3343,3345
admission|3346,3355
,|3355,3356
her|3357,3360
<EOL>|3361,3362
symptoms|3362,3370
had|3371,3374
resolved|3375,3383
,|3383,3384
no|3385,3387
abnormalities|3388,3401
were|3402,3406
seen|3407,3411
on|3412,3414
imaging|3415,3422
or|3423,3425
<EOL>|3426,3427
labs|3427,3431
,|3431,3432
and|3433,3436
her|3437,3440
VS|3441,3443
and|3444,3447
PEx|3448,3451
were|3452,3456
remarkable|3457,3467
only|3468,3472
for|3473,3476
non-acute|3477,3486
lung|3487,3491
<EOL>|3492,3493
.|3501,3502
MI|3504,3506
was|3507,3510
ruled|3511,3516
out|3517,3520
by|3521,3523
trop|3524,3528
negative|3529,3537
x3|3538,3540
,|3540,3541
no|3542,3544
EKG|3545,3548
changes|3549,3556
.|3556,3557
<EOL>|3558,3559
Cardiology|3560,3570
was|3571,3574
consulted|3575,3584
to|3585,3587
evaluate|3588,3596
need|3597,3601
for|3602,3605
catheterization|3606,3621
<EOL>|3622,3623
vs|3623,3625
other|3626,3631
intervention|3632,3644
,|3644,3645
but|3646,3649
did|3650,3653
not|3654,3657
feel|3658,3662
that|3663,3667
any|3668,3671
urgent|3672,3678
<EOL>|3679,3680
inpatient|3680,3689
work|3690,3694
-|3694,3695
up|3695,3697
was|3698,3701
necessary|3702,3711
,|3711,3712
especially|3713,3723
in|3724,3726
the|3727,3730
context|3731,3738
of|3739,3741
<EOL>|3742,3743
asymptomatic|3743,3755
tachycardia|3756,3767
.|3767,3768
She|3770,3773
had|3774,3777
already|3778,3785
had|3786,3789
Holter|3790,3796
and|3797,3800
ECHO|3801,3805
<EOL>|3806,3807
prior|3807,3812
to|3813,3815
this|3816,3820
admission|3821,3830
.|3830,3831
Cardiology|3833,3843
recommended|3844,3855
restarting|3856,3866
<EOL>|3867,3868
theophylline|3868,3880
if|3881,3883
,|3883,3884
in|3885,3887
fact|3888,3892
,|3892,3893
she|3894,3897
received|3898,3906
such|3907,3911
benefit|3912,3919
from|3920,3924
<EOL>|3925,3926
pulmonary|3926,3935
point|3936,3941
of|3942,3944
view|3945,3949
.|3949,3950
She|3952,3955
was|3956,3959
restarted|3960,3969
on|3970,3972
theophylline|3973,3985
<EOL>|3986,3987
200mg|3987,3992
TID|3993,3996
,|3996,3997
which|3998,4003
was|4004,4007
her|4008,4011
dose|4012,4016
prior|4017,4022
to|4023,4025
discontinuation|4026,4041
.|4041,4042
She|4044,4047
<EOL>|4048,4049
received|4049,4057
tobacco|4058,4065
cessation|4066,4075
education|4076,4085
,|4085,4086
was|4087,4090
continued|4091,4100
on|4101,4103
home|4104,4108
<EOL>|4109,4110
diltiazem|4110,4119
and|4120,4123
aspirin|4124,4131
(|4132,4133
dose|4133,4137
was|4138,4141
temporarily|4142,4153
increased|4154,4163
to|4164,4166
325mg|4167,4172
<EOL>|4173,4174
prior|4174,4179
to|4180,4182
ruling|4183,4189
out|4190,4193
MI|4194,4196
)|4196,4197
.|4197,4198
Admission|4200,4209
theopylline|4210,4221
level|4222,4227
was|4228,4231
<EOL>|4232,4233
pending|4233,4240
at|4241,4243
the|4244,4247
time|4248,4252
of|4253,4255
discharge|4256,4265
.|4265,4266
<EOL>|4266,4267
.|4267,4268
<EOL>|4270,4271
#|4271,4272
Asthma|4273,4279
and|4280,4283
COPD|4284,4288
:|4288,4289
patient|4290,4297
was|4298,4301
given|4302,4307
Albuterol|4308,4317
and|4318,4321
ipratropium|4322,4333
<EOL>|4334,4335
nebs|4335,4339
,|4339,4340
and|4341,4344
she|4345,4348
was|4349,4352
continued|4353,4362
on|4363,4365
her|4366,4369
home|4370,4374
doses|4375,4380
of|4381,4383
fluticasone|4384,4395
,|4395,4396
<EOL>|4397,4398
montelukast|4398,4409
,|4409,4410
fluticasone|4411,4422
-|4422,4423
salmetrol|4423,4432
.|4432,4433
She|4435,4438
was|4439,4442
given|4443,4448
O2|4449,4451
PRN|4452,4455
.|4455,4456
<EOL>|4458,4459
After|4459,4464
cardiology|4465,4475
consult|4476,4483
,|4483,4484
she|4485,4488
was|4489,4492
restarted|4493,4502
on|4503,4505
her|4506,4509
theophylline|4510,4522
<EOL>|4523,4524
at|4524,4526
200mg|4527,4532
TID|4533,4536
,|4536,4537
with|4538,4542
pulm|4543,4547
and|4548,4551
cardiology|4552,4562
follow|4563,4569
-|4569,4570
up|4570,4572
.|4572,4573
<EOL>|4573,4574
.|4574,4575
<EOL>|4577,4578
#|4578,4579
Tobacco|4580,4587
abuse|4588,4593
:|4593,4594
she|4595,4598
declined|4599,4607
nicotine|4608,4616
patch|4617,4622
,|4622,4623
and|4624,4627
education|4628,4637
was|4638,4641
<EOL>|4642,4643
given|4643,4648
regarding|4649,4658
the|4659,4662
health|4663,4669
hazards|4670,4677
of|4678,4680
smoking|4681,4688
.|4688,4689
<EOL>|4689,4690
.|4690,4691
<EOL>|4693,4694
#|4694,4695
HL|4696,4698
:|4698,4699
patient|4700,4707
was|4708,4711
continued|4712,4721
oh|4722,4724
her|4725,4728
simvastatin|4729,4740
,|4740,4741
but|4742,4745
because|4746,4753
her|4754,4757
<EOL>|4758,4759
LDL|4759,4762
was|4763,4766
not|4767,4770
at|4771,4773
goal|4774,4778
(|4779,4780
<|4780,4781
70|4781,4783
)|4783,4784
,|4784,4785
her|4786,4789
dose|4790,4794
was|4795,4798
increased|4799,4808
to|4809,4811
40mg|4812,4816
daily|4817,4822
.|4822,4823
<EOL>|4823,4824
.|4824,4825
<EOL>|4825,4826
INACTIVE|4826,4834
ISSUES|4835,4841
:|4841,4842
<EOL>|4842,4843
.|4843,4844
<EOL>|4844,4845
#|4845,4846
HTN|4847,4850
:|4850,4851
continued|4852,4861
isosorbide|4862,4872
and|4873,4876
hydrochlorothiazide|4877,4896
at|4897,4899
home|4900,4904
<EOL>|4905,4906
doses|4906,4911
.|4911,4912
<EOL>|4912,4913
.|4913,4914
<EOL>|4914,4915
#|4915,4916
Code|4917,4921
:|4921,4922
Full|4923,4927
<EOL>|4927,4928
<EOL>|4929,4930
Medications|4930,4941
on|4942,4944
Admission|4945,4954
:|4954,4955
<EOL>|4955,4956
-|4956,4957
acetaminophen|4957,4970
325|4971,4974
mg|4975,4977
Tablet|4978,4984
Sig|4985,4988
:|4988,4989
One|4990,4993
(|4994,4995
1|4995,4996
)|4996,4997
Tablet|4998,5004
PO|5005,5007
every|5008,5013
four|5014,5018
<EOL>|5019,5020
(|5020,5021
4|5021,5022
)|5022,5023
hours|5024,5029
as|5030,5032
needed|5033,5039
for|5040,5043
pain|5044,5048
.|5048,5049
<EOL>|5051,5052
-|5052,5053
albuterol|5053,5062
sulfate|5063,5070
90|5071,5073
mcg|5074,5077
/|5077,5078
Actuation|5078,5087
HFA|5088,5091
Aerosol|5092,5099
Inhaler|5100,5107
Sig|5108,5111
:|5111,5112
<EOL>|5113,5114
Two|5114,5117
(|5118,5119
2|5119,5120
)|5120,5121
Inhalation|5123,5133
every|5134,5139
_|5140,5141
_|5141,5142
_|5142,5143
hours|5144,5149
.|5149,5150
<EOL>|5152,5153
-|5153,5154
diltiazem|5154,5163
HCl|5164,5167
180|5168,5171
mg|5172,5174
Capsule|5175,5182
,|5182,5183
Extended|5184,5192
Release|5193,5200
Sig|5201,5204
:|5204,5205
Two|5206,5209
(|5210,5211
2|5211,5212
)|5212,5213
<EOL>|5214,5215
Capsule|5215,5222
,|5222,5223
Extended|5224,5232
Release|5233,5240
PO|5241,5243
DAILY|5244,5249
(|5250,5251
Daily|5251,5256
)|5256,5257
.|5257,5258
<EOL>|5260,5261
-|5261,5262
fluticasone|5262,5273
50|5274,5276
mcg|5277,5280
/|5280,5281
Actuation|5281,5290
Spray|5291,5296
,|5296,5297
Suspension|5298,5308
Sig|5309,5312
:|5312,5313
One|5314,5317
(|5318,5319
1|5319,5320
)|5320,5321
<EOL>|5322,5323
Spray|5323,5328
Nasal|5329,5334
DAILY|5335,5340
(|5341,5342
Daily|5342,5347
)|5347,5348
.|5348,5349
<EOL>|5351,5352
-|5352,5353
fluticasone|5353,5364
-|5364,5365
salmeterol|5365,5375
500|5376,5379
-|5379,5380
50|5380,5382
mcg|5383,5386
/|5386,5387
dose|5387,5391
Disk|5392,5396
with|5397,5401
Device|5402,5408
Sig|5409,5412
:|5412,5413
<EOL>|5414,5415
One|5415,5418
(|5419,5420
1|5420,5421
)|5421,5422
Disk|5423,5427
with|5428,5432
Device|5433,5439
Inhalation|5440,5450
BID|5451,5454
(|5455,5456
2|5456,5457
times|5458,5463
a|5464,5465
day|5466,5469
)|5469,5470
.|5470,5471
<EOL>|5473,5474
-|5474,5475
hydrochlorothiazide|5475,5494
12.5|5495,5499
mg|5500,5502
Capsule|5503,5510
Sig|5511,5514
:|5514,5515
One|5516,5519
(|5520,5521
1|5521,5522
)|5522,5523
Capsule|5524,5531
PO|5532,5534
<EOL>|5535,5536
DAILY|5536,5541
(|5542,5543
Daily|5543,5548
)|5548,5549
.|5549,5550
<EOL>|5552,5553
-|5553,5554
isosorbide|5554,5564
mononitrate|5565,5576
60|5577,5579
mg|5580,5582
Tablet|5583,5589
Extended|5590,5598
Release|5599,5606
24|5607,5609
hr|5610,5612
<EOL>|5613,5614
Sig|5614,5617
:|5617,5618
One|5619,5622
(|5623,5624
1|5624,5625
)|5625,5626
Tablet|5627,5633
Extended|5634,5642
Release|5643,5650
24|5651,5653
hr|5654,5656
PO|5657,5659
DAILY|5660,5665
(|5666,5667
Daily|5667,5672
)|5672,5673
.|5673,5674
<EOL>|5676,5677
-|5677,5678
montelukast|5678,5689
10|5690,5692
mg|5693,5695
Tablet|5696,5702
Sig|5703,5706
:|5706,5707
One|5708,5711
(|5712,5713
1|5713,5714
)|5714,5715
Tablet|5716,5722
PO|5723,5725
DAILY|5726,5731
<EOL>|5732,5733
(|5733,5734
Daily|5734,5739
)|5739,5740
.|5740,5741
<EOL>|5743,5744
-|5744,5745
omeprazole|5745,5755
20|5756,5758
mg|5759,5761
Capsule|5762,5769
,|5769,5770
Delayed|5771,5778
Release|5779,5786
(|5786,5787
E.C|5787,5790
.|5790,5791
)|5791,5792
Sig|5793,5796
:|5796,5797
One|5798,5801
(|5802,5803
1|5803,5804
)|5804,5805
<EOL>|5806,5807
Capsule|5807,5814
,|5814,5815
Delayed|5816,5823
Release|5824,5831
(|5831,5832
E.C|5832,5835
.|5835,5836
)|5836,5837
PO|5838,5840
DAILY|5841,5846
(|5847,5848
Daily|5848,5853
)|5853,5854
.|5854,5855
<EOL>|5857,5858
-|5858,5859
tiotropium|5859,5869
bromide|5870,5877
18|5878,5880
mcg|5881,5884
Capsule|5885,5892
,|5892,5893
w|5894,5895
/|5895,5896
Inhalation|5896,5906
Device|5907,5913
Sig|5914,5917
:|5917,5918
<EOL>|5919,5920
One|5920,5923
(|5924,5925
1|5925,5926
)|5926,5927
Cap|5928,5931
Inhalation|5932,5942
DAILY|5943,5948
(|5949,5950
Daily|5950,5955
)|5955,5956
.|5956,5957
<EOL>|5959,5960
-|5960,5961
calcium|5961,5968
carbonate|5969,5978
200|5979,5982
mg|5983,5985
(|5986,5987
500|5987,5990
mg|5991,5993
)|5993,5994
Tablet|5995,6001
,|6001,6002
Chewable|6003,6011
Sig|6012,6015
:|6015,6016
One|6017,6020
<EOL>|6021,6022
(|6022,6023
1|6023,6024
)|6024,6025
Tablet|6026,6032
,|6032,6033
Chewable|6034,6042
PO|6043,6045
DAILY|6046,6051
(|6052,6053
Daily|6053,6058
)|6058,6059
.|6059,6060
<EOL>|6062,6063
-|6063,6064
multivitamin|6064,6076
Tablet|6081,6087
Sig|6088,6091
:|6091,6092
One|6093,6096
(|6097,6098
1|6098,6099
)|6099,6100
Tablet|6101,6107
PO|6108,6110
DAILY|6111,6116
<EOL>|6117,6118
(|6118,6119
Daily|6119,6124
)|6124,6125
.|6125,6126
<EOL>|6128,6129
-|6129,6130
aspirin|6130,6137
81|6138,6140
mg|6141,6143
Tablet|6144,6150
Sig|6151,6154
:|6154,6155
One|6156,6159
(|6160,6161
1|6161,6162
)|6162,6163
Tablet|6164,6170
PO|6171,6173
once|6174,6178
a|6179,6180
day|6181,6184
.|6184,6185
<EOL>|6187,6188
-|6188,6189
simvastatin|6189,6200
20mg|6201,6205
qday|6206,6210
<EOL>|6210,6211
<EOL>|6212,6213
Discharge|6213,6222
Medications|6223,6234
:|6234,6235
<EOL>|6235,6236
1.|6236,6238
simvastatin|6239,6250
40|6251,6253
mg|6254,6256
Tablet|6257,6263
Sig|6264,6267
:|6267,6268
One|6269,6272
(|6273,6274
1|6274,6275
)|6275,6276
Tablet|6277,6283
PO|6284,6286
DAILY|6287,6292
<EOL>|6293,6294
(|6294,6295
Daily|6295,6300
)|6300,6301
.|6301,6302
<EOL>|6302,6303
Disp|6303,6307
:|6307,6308
*|6308,6309
30|6309,6311
Tablet|6312,6318
(|6318,6319
s|6319,6320
)|6320,6321
*|6321,6322
Refills|6323,6330
:|6330,6331
*|6331,6332
0|6332,6333
*|6333,6334
<EOL>|6334,6335
2.|6335,6337
hydrochlorothiazide|6338,6357
12.5|6358,6362
mg|6363,6365
Capsule|6366,6373
Sig|6374,6377
:|6377,6378
One|6379,6382
(|6383,6384
1|6384,6385
)|6385,6386
Capsule|6387,6394
PO|6395,6397
<EOL>|6398,6399
DAILY|6399,6404
(|6405,6406
Daily|6406,6411
)|6411,6412
.|6412,6413
<EOL>|6415,6416
3.|6416,6418
fluticasone|6419,6430
50|6431,6433
mcg|6434,6437
/|6437,6438
Actuation|6438,6447
Spray|6448,6453
,|6453,6454
Suspension|6455,6465
Sig|6466,6469
:|6469,6470
_|6471,6472
_|6472,6473
_|6473,6474
<EOL>|6475,6476
Sprays|6476,6482
Nasal|6483,6488
DAILY|6489,6494
(|6495,6496
Daily|6496,6501
)|6501,6502
as|6503,6505
needed|6506,6512
for|6513,6516
congestion|6517,6527
.|6527,6528
<EOL>|6530,6531
4.|6531,6533
isosorbide|6534,6544
mononitrate|6545,6556
60|6557,6559
mg|6560,6562
Tablet|6563,6569
Extended|6570,6578
Release|6579,6586
24|6587,6589
hr|6590,6592
<EOL>|6593,6594
Sig|6594,6597
:|6597,6598
One|6599,6602
(|6603,6604
1|6604,6605
)|6605,6606
Tablet|6607,6613
Extended|6614,6622
Release|6623,6630
24|6631,6633
hr|6634,6636
PO|6637,6639
DAILY|6640,6645
(|6646,6647
Daily|6647,6652
)|6652,6653
.|6653,6654
<EOL>|6656,6657
5.|6657,6659
montelukast|6660,6671
10|6672,6674
mg|6675,6677
Tablet|6678,6684
Sig|6685,6688
:|6688,6689
One|6690,6693
(|6694,6695
1|6695,6696
)|6696,6697
Tablet|6698,6704
PO|6705,6707
DAILY|6708,6713
<EOL>|6714,6715
(|6715,6716
Daily|6716,6721
)|6721,6722
.|6722,6723
<EOL>|6725,6726
6.|6726,6728
fluticasone|6729,6740
-|6740,6741
salmeterol|6741,6751
500|6752,6755
-|6755,6756
50|6756,6758
mcg|6759,6762
/|6762,6763
dose|6763,6767
Disk|6768,6772
with|6773,6777
Device|6778,6784
Sig|6785,6788
:|6788,6789
<EOL>|6790,6791
One|6791,6794
(|6795,6796
1|6796,6797
)|6797,6798
Disk|6799,6803
with|6804,6808
Device|6809,6815
Inhalation|6816,6826
BID|6827,6830
(|6831,6832
2|6832,6833
times|6834,6839
a|6840,6841
day|6842,6845
)|6845,6846
.|6846,6847
<EOL>|6849,6850
7.|6850,6852
acetaminophen|6853,6866
-|6866,6867
codeine|6867,6874
300|6875,6878
-|6878,6879
30|6879,6881
mg|6882,6884
Tablet|6885,6891
Sig|6892,6895
:|6895,6896
One|6897,6900
(|6901,6902
1|6902,6903
)|6903,6904
Tablet|6905,6911
PO|6912,6914
<EOL>|6915,6916
every|6916,6921
four|6922,6926
(|6927,6928
4|6928,6929
)|6929,6930
hours|6931,6936
as|6937,6939
needed|6940,6946
for|6947,6950
pain|6951,6955
.|6955,6956
<EOL>|6958,6959
8.|6959,6961
albuterol|6962,6971
sulfate|6972,6979
90|6980,6982
mcg|6983,6986
/|6986,6987
Actuation|6987,6996
HFA|6997,7000
Aerosol|7001,7008
Inhaler|7009,7016
Sig|7017,7020
:|7020,7021
<EOL>|7022,7023
Two|7023,7026
(|7027,7028
2|7028,7029
)|7029,7030
puffs|7031,7036
Inhalation|7037,7047
every|7048,7053
_|7054,7055
_|7055,7056
_|7056,7057
hours|7058,7063
as|7064,7066
needed|7067,7073
for|7074,7077
shortness|7078,7087
<EOL>|7088,7089
of|7089,7091
breath|7092,7098
or|7099,7101
wheezing|7102,7110
.|7110,7111
<EOL>|7113,7114
9.|7114,7116
omeprazole|7117,7127
20|7128,7130
mg|7131,7133
Capsule|7134,7141
,|7141,7142
Delayed|7143,7150
Release|7151,7158
(|7158,7159
E.C|7159,7162
.|7162,7163
)|7163,7164
Sig|7165,7168
:|7168,7169
One|7170,7173
(|7174,7175
1|7175,7176
)|7176,7177
<EOL>|7178,7179
Capsule|7179,7186
,|7186,7187
Delayed|7188,7195
Release|7196,7203
(|7203,7204
E.C|7204,7207
.|7207,7208
)|7208,7209
PO|7210,7212
DAILY|7213,7218
(|7219,7220
Daily|7220,7225
)|7225,7226
.|7226,7227
<EOL>|7229,7230
10.|7230,7233
Spiriva|7234,7241
with|7242,7246
HandiHaler|7247,7257
18|7258,7260
mcg|7261,7264
Capsule|7265,7272
,|7272,7273
w|7274,7275
/|7275,7276
Inhalation|7276,7286
Device|7287,7293
<EOL>|7294,7295
Sig|7295,7298
:|7298,7299
One|7300,7303
(|7304,7305
1|7305,7306
)|7306,7307
capsule|7308,7315
Inhalation|7316,7326
once|7327,7331
a|7332,7333
day|7334,7337
.|7337,7338
<EOL>|7340,7341
11.|7341,7344
aspirin|7345,7352
81|7353,7355
mg|7356,7358
Tablet|7359,7365
Sig|7366,7369
:|7369,7370
One|7371,7374
(|7375,7376
1|7376,7377
)|7377,7378
Tablet|7379,7385
PO|7386,7388
once|7389,7393
a|7394,7395
day|7396,7399
.|7399,7400
<EOL>|7402,7403
12.|7403,7406
calcium|7407,7414
carbonate|7415,7424
200|7425,7428
mg|7429,7431
(|7432,7433
500|7433,7436
mg|7437,7439
)|7439,7440
Tablet|7441,7447
,|7447,7448
Chewable|7449,7457
Sig|7458,7461
:|7461,7462
One|7463,7466
<EOL>|7467,7468
(|7468,7469
1|7469,7470
)|7470,7471
Tablet|7472,7478
,|7478,7479
Chewable|7480,7488
PO|7489,7491
DAILY|7492,7497
(|7498,7499
Daily|7499,7504
)|7504,7505
.|7505,7506
<EOL>|7508,7509
13.|7509,7512
diltiazem|7513,7522
HCl|7523,7526
180|7527,7530
mg|7531,7533
Capsule|7534,7541
,|7541,7542
Extended|7543,7551
Release|7552,7559
Sig|7560,7563
:|7563,7564
Two|7565,7568
(|7569,7570
2|7570,7571
)|7571,7572
<EOL>|7573,7574
Capsule|7574,7581
,|7581,7582
Extended|7583,7591
Release|7592,7599
PO|7600,7602
DAILY|7603,7608
(|7609,7610
Daily|7610,7615
)|7615,7616
.|7616,7617
<EOL>|7619,7620
14.|7620,7623
multivitamin|7624,7636
Tablet|7641,7647
Sig|7648,7651
:|7651,7652
One|7653,7656
(|7657,7658
1|7658,7659
)|7659,7660
Tablet|7661,7667
PO|7668,7670
DAILY|7671,7676
<EOL>|7677,7678
(|7678,7679
Daily|7679,7684
)|7684,7685
.|7685,7686
<EOL>|7688,7689
15.|7689,7692
theophylline|7693,7705
200|7706,7709
mg|7710,7712
Capsule|7713,7720
,|7720,7721
Ext|7722,7725
Release|7726,7733
24|7734,7736
hr|7737,7739
Sig|7740,7743
:|7743,7744
One|7745,7748
(|7749,7750
1|7750,7751
)|7751,7752
<EOL>|7753,7754
Capsule|7754,7761
,|7761,7762
Ext|7763,7766
Release|7767,7774
24|7775,7777
hr|7778,7780
PO|7781,7783
three|7784,7789
times|7790,7795
a|7796,7797
day|7798,7801
.|7801,7802
<EOL>|7802,7803
Disp|7803,7807
:|7807,7808
*|7808,7809
90|7809,7811
Capsule|7812,7819
,|7819,7820
Ext|7821,7824
Release|7825,7832
24|7833,7835
hr|7836,7838
(|7838,7839
s|7839,7840
)|7840,7841
*|7841,7842
Refills|7843,7850
:|7850,7851
*|7851,7852
0|7852,7853
*|7853,7854
<EOL>|7854,7855
16.|7855,7858
albuterol|7859,7868
sulfate|7869,7876
0.63|7877,7881
mg|7882,7884
/|7884,7885
3|7885,7886
mL|7887,7889
Solution|7890,7898
for|7899,7902
Nebulization|7903,7915
<EOL>|7916,7917
Sig|7917,7920
:|7920,7921
One|7922,7925
(|7926,7927
1|7927,7928
)|7928,7929
treatment|7930,7939
Inhalation|7940,7950
every|7951,7956
_|7957,7958
_|7958,7959
_|7959,7960
hours|7961,7966
as|7967,7969
needed|7970,7976
for|7977,7980
<EOL>|7981,7982
shortness|7982,7991
of|7992,7994
breath|7995,8001
or|8002,8004
wheezing|8005,8013
for|8014,8017
15|8018,8020
doses|8021,8026
.|8026,8027
<EOL>|8027,8028
Disp|8028,8032
:|8032,8033
*|8033,8034
15|8034,8036
ampules|8037,8044
*|8044,8045
Refills|8046,8053
:|8053,8054
*|8054,8055
0|8055,8056
*|8056,8057
<EOL>|8057,8058
<EOL>|8058,8059
<EOL>|8060,8061
Discharge|8061,8070
Disposition|8071,8082
:|8082,8083
<EOL>|8083,8084
Home|8084,8088
With|8089,8093
Service|8094,8101
<EOL>|8101,8102
<EOL>|8103,8104
Facility|8104,8112
:|8112,8113
<EOL>|8113,8114
_|8114,8115
_|8115,8116
_|8116,8117
<EOL>|8117,8118
<EOL>|8119,8120
Discharge|8120,8129
Diagnosis|8130,8139
:|8139,8140
<EOL>|8140,8141
Primary|8141,8148
:|8148,8149
<EOL>|8149,8150
-|8150,8151
Tachyarrhythmia|8151,8166
<EOL>|8166,8167
-|8167,8168
Hyperlipidemia|8168,8182
<EOL>|8182,8183
-|8183,8184
Asthma|8184,8190
,|8190,8191
COPD|8192,8196
<EOL>|8196,8197
<EOL>|8197,8198
Secondary|8198,8207
:|8207,8208
<EOL>|8208,8209
-|8209,8210
Hypertension|8210,8222
<EOL>|8223,8224
-|8224,8225
Tobacco|8225,8232
Use|8233,8236
<EOL>|8238,8239
<EOL>|8239,8240
<EOL>|8241,8242
Mental|8263,8269
Status|8270,8276
:|8276,8277
Clear|8278,8283
and|8284,8287
coherent|8288,8296
.|8296,8297
<EOL>|8297,8298
Level|8298,8303
of|8304,8306
Consciousness|8307,8320
:|8320,8321
Alert|8322,8327
and|8328,8331
interactive|8332,8343
.|8343,8344
<EOL>|8344,8345
Activity|8345,8353
Status|8354,8360
:|8360,8361
Ambulatory|8362,8372
-|8373,8374
Independent|8375,8386
.|8386,8387
<EOL>|8387,8388
<EOL>|8388,8389
<EOL>|8390,8391
Mrs.|8415,8419
_|8420,8421
_|8421,8422
_|8422,8423
,|8423,8424
<EOL>|8424,8425
<EOL>|8425,8426
_|8426,8427
_|8427,8428
_|8428,8429
were|8430,8434
hospitalized|8435,8447
because|8448,8455
the|8456,8459
visiting|8460,8468
nurses|8469,8475
were|8476,8480
concerned|8481,8490
<EOL>|8491,8492
about|8492,8497
an|8498,8500
elevated|8501,8509
heart|8510,8515
rate|8516,8520
,|8520,8521
but|8522,8525
by|8526,8528
the|8529,8532
time|8533,8537
_|8538,8539
_|8539,8540
_|8540,8541
came|8542,8546
to|8547,8549
the|8550,8553
<EOL>|8554,8555
hospital|8555,8563
,|8563,8564
your|8565,8569
elevated|8570,8578
heart|8579,8584
rate|8585,8589
had|8590,8593
resolved|8594,8602
.|8602,8603
Nevertheless|8605,8617
,|8617,8618
<EOL>|8619,8620
_|8620,8621
_|8621,8622
_|8622,8623
were|8624,8628
admitted|8629,8637
to|8638,8640
ensure|8641,8647
that|8648,8652
your|8653,8657
heart|8658,8663
had|8664,8667
n't|8667,8670
suffered|8671,8679
any|8680,8683
<EOL>|8684,8685
damage|8685,8691
,|8691,8692
and|8693,8696
to|8697,8699
see|8700,8703
the|8704,8707
inpatient|8708,8717
cardiologist|8718,8730
.|8730,8731
Your|8733,8737
labs|8738,8742
were|8743,8747
<EOL>|8748,8749
unremarkable|8749,8761
from|8762,8766
a|8767,8768
cardiac|8769,8776
standpoint|8777,8787
,|8787,8788
and|8789,8792
_|8793,8794
_|8794,8795
_|8795,8796
saw|8797,8800
the|8801,8804
<EOL>|8805,8806
cardiologist|8806,8818
(|8819,8820
who|8820,8823
recommend|8824,8833
no|8834,8836
intervention|8837,8849
at|8850,8852
this|8853,8857
time|8858,8862
)|8862,8863
.|8863,8864
_|8866,8867
_|8867,8868
_|8868,8869
<EOL>|8870,8871
should|8871,8877
follow|8878,8884
-|8884,8885
up|8885,8887
with|8888,8892
your|8893,8897
pulmonologist|8898,8911
as|8912,8914
an|8915,8917
outpatient|8918,8928
for|8929,8932
<EOL>|8933,8934
your|8934,8938
breathing|8939,8948
issues|8949,8955
.|8955,8956
The|8958,8961
best|8962,8966
thing|8967,8972
_|8973,8974
_|8974,8975
_|8975,8976
can|8977,8980
do|8981,8983
for|8984,8987
your|8988,8992
lung|8993,8997
<EOL>|8998,8999
health|8999,9005
is|9006,9008
to|9009,9011
quit|9012,9016
smoking|9017,9024
,|9024,9025
and|9026,9029
we|9030,9032
encourage|9033,9042
_|9043,9044
_|9044,9045
_|9045,9046
to|9047,9049
do|9050,9052
so|9053,9055
.|9055,9056
<EOL>|9056,9057
<EOL>|9057,9058
The|9058,9061
following|9062,9071
changes|9072,9079
were|9080,9084
made|9085,9089
to|9090,9092
your|9093,9097
medications|9098,9109
:|9109,9110
<EOL>|9110,9111
-|9111,9112
INCREASE|9112,9120
your|9121,9125
simvastatin|9126,9137
to|9138,9140
40mg|9141,9145
daily|9146,9151
in|9152,9154
order|9155,9160
to|9161,9163
lower|9164,9169
your|9170,9174
<EOL>|9175,9176
cholesterol|9176,9187
to|9188,9190
goal|9191,9195
(|9196,9197
as|9197,9199
recommended|9200,9211
by|9212,9214
the|9215,9218
cardiologist|9219,9231
)|9231,9232
<EOL>|9232,9233
-|9233,9234
RESTART|9234,9241
theophylline|9242,9254
200mg|9255,9260
three|9261,9266
times|9267,9272
a|9273,9274
day|9275,9278
<EOL>|9278,9279
-|9279,9280
We|9280,9282
will|9283,9287
also|9288,9292
be|9293,9295
giving|9296,9302
_|9303,9304
_|9304,9305
_|9305,9306
a|9307,9308
prescription|9309,9321
for|9322,9325
albuterol|9326,9335
<EOL>|9336,9337
nebulizers|9337,9347
to|9348,9350
use|9351,9354
instead|9355,9362
of|9363,9365
your|9366,9370
inhaler|9371,9378
(|9379,9380
when|9380,9384
needed|9385,9391
)|9391,9392
,|9392,9393
but|9394,9397
<EOL>|9398,9399
refills|9399,9406
will|9407,9411
have|9412,9416
to|9417,9419
be|9420,9422
through|9423,9430
your|9431,9435
primary|9436,9443
physician|9444,9453
or|9454,9456
<EOL>|9457,9458
pulmonologist|9458,9471
<EOL>|9471,9472
<EOL>|9472,9473
_|9473,9474
_|9474,9475
_|9475,9476
discuss|9477,9484
your|9485,9489
theophylline|9490,9502
dose|9503,9507
and|9508,9511
breathing|9512,9521
status|9522,9528
with|9529,9533
<EOL>|9534,9535
your|9535,9539
primary|9540,9547
provider|9548,9556
(|9557,9558
Dr|9558,9560
.|9560,9561
_|9562,9563
_|9563,9564
_|9564,9565
and|9566,9569
your|9570,9574
pulmonologist|9575,9588
(|9589,9590
Dr|9590,9592
.|9592,9593
<EOL>|9594,9595
_|9595,9596
_|9596,9597
_|9597,9598
.|9598,9599
<EOL>|9601,9602
<EOL>|9603,9604
Followup|9604,9612
Instructions|9613,9625
:|9625,9626
<EOL>|9626,9627
_|9627,9628
_|9628,9629
_|9629,9630
<EOL>|9630,9631

