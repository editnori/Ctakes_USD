 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|42,51|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|42,51|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|42,56|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|76,85|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|76,85|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|76,85|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|76,85|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|76,85|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|76,90|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|108,113|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|108,113|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|108,113|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|132,135|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|143,150|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|143,150|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|152,160|true|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|Allergies|184,193|true|false|false|C1717415||Allergies
Event|Event|Allergies|184,193|true|false|false|||Allergies
Finding|Pathologic Function|Allergies|184,193|true|false|false|C0020517|Hypersensitivity|Allergies
Finding|Pathologic Function|Allergies|196,218|true|false|false|C0041755|Adverse reaction to drug|Adverse Drug Reactions
Drug|Pharmacologic Substance|Allergies|204,208|true|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|Drug
Finding|Finding|Allergies|204,208|true|false|false|C0740721|Drug problem|Drug
Finding|Pathologic Function|Allergies|204,218|true|false|false|C0041755|Adverse reaction to drug|Drug Reactions
Event|Event|Allergies|209,218|true|false|false|||Reactions
Event|Event|Allergies|221,230|false|false|false|||Attending
Finding|Functional Concept|Allergies|221,230|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|Chief Complaint|256,264|false|false|false|C0741302|atypia morphology|Atypical
Finding|Sign or Symptom|Chief Complaint|256,275|false|false|false|C0262384|Atypical chest pain|Atypical chest pain
Anatomy|Body Location or Region|Chief Complaint|265,270|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Chief Complaint|265,270|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Chief Complaint|265,275|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|Chief Complaint|265,275|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Chief Complaint|271,275|false|true|false|C2598155||pain
Event|Event|Chief Complaint|271,275|false|false|false|||pain
Finding|Functional Concept|Chief Complaint|271,275|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Chief Complaint|271,275|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Classification|Chief Complaint|278,283|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|284,292|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|284,292|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|296,314|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|305,314|false|false|false|C0945766||Procedure
Event|Event|Chief Complaint|305,314|false|false|false|||Procedure
Event|Occupational Activity|Chief Complaint|305,314|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|305,314|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|305,314|false|false|false|C0184661|Interventional procedure|Procedure
Procedure|Health Care Activity|Chief Complaint|322,326|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|Echo
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|322,326|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|Echo
Anatomy|Body Location or Region|History of Present Illness|390,395|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|390,395|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|History of Present Illness|390,400|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|History of Present Illness|390,400|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|History of Present Illness|396,400|false|false|false|C2598155||pain
Event|Event|History of Present Illness|396,400|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|396,400|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|396,400|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|History of Present Illness|423,427|false|false|false|C2598155||Pain
Event|Event|History of Present Illness|423,427|false|false|false|||Pain
Finding|Functional Concept|History of Present Illness|423,427|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|History of Present Illness|423,427|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Functional Concept|History of Present Illness|442,446|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Disorder|Disease or Syndrome|History of Present Illness|447,456|false|false|false|C0751438|Posterior pituitary disease|posterior
Anatomy|Body Location or Region|History of Present Illness|457,465|false|false|false|C0037004;C4299050|Shoulder;Upper extremity>Shoulder|shoulder
Procedure|Diagnostic Procedure|History of Present Illness|457,465|false|false|false|C0221590;C0869975|Examination of shoulder(s);Procedures on Shoulder|shoulder
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|457,465|false|false|false|C0221590;C0869975|Examination of shoulder(s);Procedures on Shoulder|shoulder
Event|Event|History of Present Illness|470,478|false|false|false|||radiates
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|484,487|false|false|false|C0446516;C1140618;C1269078|Upper Extremity;Upper arm|arm
Disorder|Anatomical Abnormality|History of Present Illness|484,487|false|false|false|C3495676|Anorectal Malformations|arm
Event|Event|History of Present Illness|484,487|false|false|false|||arm
Finding|Gene or Genome|History of Present Illness|484,487|false|false|false|C1824218;C3715044|AKR1A1 wt Allele;ARMC9 gene|arm
Procedure|Diagnostic Procedure|History of Present Illness|484,487|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Research Activity|History of Present Illness|484,487|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|484,487|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|492,499|false|false|false|C0016129|Fingers|fingers
Event|Event|History of Present Illness|509,514|false|false|false|||turns
Finding|Gene or Genome|History of Present Illness|521,525|false|false|false|C1428865|GPSM2 gene|pins
Event|Event|History of Present Illness|528,535|false|false|false|||needles
Attribute|Clinical Attribute|History of Present Illness|537,544|false|false|false|C3854129||symptom
Event|Event|History of Present Illness|537,544|false|false|false|||symptom
Finding|Sign or Symptom|History of Present Illness|537,544|false|false|false|C1457887|Symptoms|symptom
Event|Event|History of Present Illness|550,553|true|false|false|||SOB
Finding|Sign or Symptom|History of Present Illness|550,553|true|false|false|C0013404|Dyspnea|SOB
Finding|Body Substance|History of Present Illness|559,566|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|559,566|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|559,566|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|History of Present Illness|572,579|false|false|false|||endorse
Event|Event|History of Present Illness|593,604|false|false|false|||diaphoresis
Finding|Finding|History of Present Illness|593,604|false|true|false|C0700590|Increased sweating|diaphoresis
Disorder|Disease or Syndrome|History of Present Illness|609,613|false|false|false|C0017168|Gastroesophageal reflux disease|gerd
Event|Event|History of Present Illness|609,613|false|false|false|||gerd
Event|Event|History of Present Illness|620,628|false|false|false|||symptoms
Finding|Functional Concept|History of Present Illness|620,628|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|History of Present Illness|620,628|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|History of Present Illness|629,641|false|false|false|||accompanying
Attribute|Clinical Attribute|History of Present Illness|646,650|false|false|false|C2598155||Pain
Event|Event|History of Present Illness|646,650|false|false|false|||Pain
Finding|Functional Concept|History of Present Illness|646,650|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|History of Present Illness|646,650|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Event|Event|History of Present Illness|660,670|false|false|false|||controlled
Drug|Organic Chemical|History of Present Illness|677,684|false|false|false|C0699142|Tylenol|tylenol
Drug|Pharmacologic Substance|History of Present Illness|677,684|false|false|false|C0699142|Tylenol|tylenol
Event|Event|History of Present Illness|677,684|false|false|false|||tylenol
Disorder|Disease or Syndrome|Past Medical History|714,717|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|Past Medical History|714,717|false|false|false|||HTN
Disorder|Disease or Syndrome|Past Medical History|720,726|false|false|false|C0004096|Asthma|Asthma
Event|Event|Past Medical History|720,726|false|false|false|||Asthma
Disorder|Disease or Syndrome|Past Medical History|729,743|false|false|false|C0012813|Diverticulitis|Diverticulitis
Event|Event|Past Medical History|729,743|false|false|false|||Diverticulitis
Finding|Gene or Genome|Past Medical History|758,761|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Anatomy|Body Location or Region|Past Medical History|764,769|false|false|false|C0524470|Right hip region structure|R hip
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|766,769|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|hip
Drug|Amino Acid, Peptide, or Protein|Past Medical History|766,769|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Biologically Active Substance|Past Medical History|766,769|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Pharmacologic Substance|Past Medical History|766,769|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Finding|Gene or Genome|Past Medical History|766,769|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|hip
Procedure|Therapeutic or Preventive Procedure|Past Medical History|766,769|false|false|false|C1292890|Procedure on hip|hip
Procedure|Therapeutic or Preventive Procedure|Past Medical History|766,781|false|false|false|C0392806|Prosthetic arthroplasty of hip (procedure)|hip replacement
Event|Event|Past Medical History|770,781|false|false|false|||replacement
Finding|Functional Concept|Past Medical History|770,781|false|false|false|C0559956|Replacement|replacement
Procedure|Health Care Activity|Past Medical History|770,781|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|replacement
Procedure|Therapeutic or Preventive Procedure|Past Medical History|770,781|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|replacement
Finding|Idea or Concept|Family Medical History|830,836|false|false|false|C1546508|Relationship - Mother|Mother
Disorder|Disease or Syndrome|Family Medical History|843,846|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|Family Medical History|843,846|false|false|false|||HTN
Finding|Conceptual Entity|Family Medical History|849,855|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Idea or Concept|Family Medical History|849,855|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Event|Event|Family Medical History|866,873|false|false|false|||Brother
Finding|Conceptual Entity|Family Medical History|866,873|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Finding|Idea or Concept|Family Medical History|866,873|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Event|Event|Family Medical History|881,888|false|false|false|||Brother
Finding|Conceptual Entity|Family Medical History|881,888|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Finding|Idea or Concept|Family Medical History|881,888|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Event|Event|Family Medical History|899,907|false|false|false|||Physical
Finding|Finding|Family Medical History|899,907|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|Family Medical History|899,907|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|Family Medical History|899,907|false|false|false|C0031809|Physical Examination|Physical
Event|Event|Family Medical History|964,971|false|false|false|||General
Finding|Classification|Family Medical History|964,971|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|Family Medical History|964,971|false|false|false|C3812897|General medical service|General
Attribute|Clinical Attribute|Family Medical History|973,978|true|false|false|C5890168||Alert
Drug|Organic Chemical|Family Medical History|973,978|true|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Family Medical History|973,978|true|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|Family Medical History|973,978|true|false|false|||Alert
Finding|Finding|Family Medical History|973,978|true|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Family Medical History|973,978|true|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Family Medical History|973,978|true|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|Family Medical History|980,988|true|false|false|||oriented
Finding|Intellectual Product|Family Medical History|993,998|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|Family Medical History|999,1007|true|false|false|||distress
Finding|Finding|Family Medical History|999,1007|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|Family Medical History|999,1007|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Anatomy|Body Location or Region|Family Medical History|1010,1015|true|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1017,1023|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|Family Medical History|1017,1023|false|false|false|C0036412|Scleral Diseases|Sclera
Event|Event|Family Medical History|1017,1023|false|false|false|||Sclera
Procedure|Health Care Activity|Family Medical History|1017,1023|false|false|false|C2228481|examination of sclera|Sclera
Event|Event|Family Medical History|1024,1033|false|false|false|||anicteric
Finding|Finding|Family Medical History|1024,1033|false|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1035,1038|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|Family Medical History|1035,1038|false|false|false|C0026987|Myelofibrosis|MMM
Anatomy|Body Location or Region|Family Medical History|1040,1050|false|false|false|C0521367|Oropharyngeal|oropharynx
Event|Event|Family Medical History|1051,1056|false|false|false|||clear
Finding|Idea or Concept|Family Medical History|1051,1056|false|false|false|C1550016|Remote control command - Clear|clear
Anatomy|Body Location or Region|Family Medical History|1059,1063|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Anatomy|Cell Component|Family Medical History|1059,1063|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Finding|Finding|Family Medical History|1059,1063|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|Neck
Event|Event|Family Medical History|1065,1071|true|false|false|||supple
Finding|Functional Concept|Family Medical History|1065,1071|true|false|false|C0332254|Supple|supple
Event|Event|Family Medical History|1073,1076|true|false|false|||JVP
Finding|Finding|Family Medical History|1073,1076|true|false|false|C0428897|Jugular venous pressure|JVP
Event|Event|Family Medical History|1081,1089|true|false|false|||elevated
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1094,1097|true|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|Family Medical History|1094,1097|true|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|Family Medical History|1094,1097|true|false|false|||LAD
Finding|Gene or Genome|Family Medical History|1094,1097|true|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1100,1105|true|false|false|C0024109|Lung|Lungs
Event|Event|Family Medical History|1107,1112|true|false|false|||Clear
Finding|Idea or Concept|Family Medical History|1107,1112|true|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|Family Medical History|1116,1128|true|false|false|||auscultation
Procedure|Diagnostic Procedure|Family Medical History|1116,1128|true|false|false|C0004339|Auscultation|auscultation
Event|Event|Family Medical History|1145,1152|true|false|false|||wheezes
Finding|Sign or Symptom|Family Medical History|1145,1152|true|false|false|C0043144|Wheezing|wheezes
Event|Event|Family Medical History|1154,1159|true|false|false|||rales
Finding|Finding|Family Medical History|1154,1159|true|false|false|C0034642;C0240859|Basilar Rales;Rales|rales
Event|Activity|Family Medical History|1183,1187|false|false|false|C0871208|Rating (action)|rate
Event|Event|Family Medical History|1183,1187|false|false|false|||rate
Finding|Idea or Concept|Family Medical History|1183,1187|false|false|false|C1549480|Amount type - Rate|rate
Event|Event|Family Medical History|1192,1198|true|false|false|||rhythm
Finding|Finding|Family Medical History|1192,1198|true|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|Family Medical History|1192,1198|true|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Event|Event|Family Medical History|1219,1226|true|false|false|||murmurs
Finding|Finding|Family Medical History|1219,1226|true|false|false|C0018808|Heart murmur|murmurs
Event|Event|Family Medical History|1228,1232|true|false|false|||rubs
Finding|Finding|Family Medical History|1228,1232|true|false|false|C0232267|Pericardial friction rub|rubs
Event|Event|Family Medical History|1235,1242|true|false|false|||gallops
Anatomy|Body Location or Region|Family Medical History|1245,1252|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|Family Medical History|1245,1252|false|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Event|Event|Family Medical History|1245,1252|false|false|false|||Abdomen
Finding|Finding|Family Medical History|1245,1252|false|false|false|C0941288|Abdomen problem|Abdomen
Disorder|Disease or Syndrome|Family Medical History|1254,1258|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|Family Medical History|1254,1258|false|false|false|||soft
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1287,1292|true|false|false|C0021853|Intestines|bowel
Finding|Finding|Family Medical History|1287,1299|true|false|false|C0232693|Bowel sounds|bowel sounds
Event|Event|Family Medical History|1293,1299|true|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|Family Medical History|1293,1299|true|false|false|C0037709||sounds
Finding|Finding|Family Medical History|1300,1307|true|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|Family Medical History|1300,1307|true|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Sign or Symptom|Family Medical History|1313,1331|true|false|false|C0234246|Rebound tenderness|rebound tenderness
Event|Event|Family Medical History|1321,1331|true|false|false|||tenderness
Finding|Mental Process|Family Medical History|1321,1331|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|Family Medical History|1321,1331|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Event|Event|Family Medical History|1335,1343|true|false|false|||guarding
Finding|Finding|Family Medical History|1335,1343|true|false|false|C0427198|Protective muscle spasm|guarding
Event|Event|Family Medical History|1348,1360|true|false|false|||organomegaly
Finding|Finding|Family Medical History|1348,1360|true|false|false|C4054315|Organomegaly|organomegaly
Disorder|Congenital Abnormality|Family Medical History|1363,1366|true|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Event|Event|Family Medical History|1363,1366|true|false|false|||Ext
Finding|Gene or Genome|Family Medical History|1363,1366|true|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Event|Event|Family Medical History|1368,1372|false|false|false|||Warm
Finding|Finding|Family Medical History|1368,1372|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|Family Medical History|1368,1372|false|false|false|C0687712|warming process|Warm
Finding|Finding|Family Medical History|1374,1378|true|false|false|C5575035|Well (answer to question)|well
Event|Event|Family Medical History|1379,1387|true|false|false|||perfused
Drug|Food|Family Medical History|1392,1398|true|false|false|C5890763||pulses
Event|Event|Family Medical History|1392,1398|true|false|false|||pulses
Finding|Physiologic Function|Family Medical History|1392,1398|true|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|Family Medical History|1392,1398|true|false|false|C0034107|Pulse taking|pulses
Disorder|Anatomical Abnormality|Family Medical History|1403,1411|true|false|false|C0149651|Clubbing|clubbing
Event|Event|Family Medical History|1403,1411|true|false|false|||clubbing
Event|Event|Family Medical History|1413,1421|true|false|false|||cyanosis
Finding|Sign or Symptom|Family Medical History|1413,1421|true|false|false|C0010520|Cyanosis|cyanosis
Attribute|Clinical Attribute|Family Medical History|1426,1431|true|false|false|C1717255||edema
Event|Event|Family Medical History|1426,1431|true|false|false|||edema
Finding|Pathologic Function|Family Medical History|1426,1431|true|false|false|C0013604|Edema|edema
Disorder|Disease or Syndrome|Family Medical History|1468,1473|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|1468,1473|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|1468,1473|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|Family Medical History|1474,1477|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|Family Medical History|1482,1485|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|Family Medical History|1482,1485|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|Family Medical History|1482,1485|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|Family Medical History|1491,1494|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|Family Medical History|1491,1494|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|Family Medical History|1491,1494|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|Family Medical History|1491,1494|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|Family Medical History|1500,1503|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|Family Medical History|1500,1503|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|Family Medical History|1509,1512|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|Family Medical History|1509,1512|false|false|false|||MCV
Lab|Laboratory or Test Result|Family Medical History|1509,1512|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|Family Medical History|1509,1512|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|Family Medical History|1509,1512|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|Family Medical History|1517,1520|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|Family Medical History|1517,1520|false|false|false|C0600370|methacholine|MCH
Event|Event|Family Medical History|1517,1520|false|false|false|||MCH
Finding|Gene or Genome|Family Medical History|1517,1520|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|Family Medical History|1517,1520|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|Family Medical History|1517,1520|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|Family Medical History|1526,1530|false|false|false|||MCHC
Procedure|Laboratory Procedure|Family Medical History|1526,1530|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|Family Medical History|1545,1548|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|Family Medical History|1565,1570|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|1565,1570|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|1565,1570|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|Family Medical History|1571,1574|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|Family Medical History|1579,1582|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|Family Medical History|1579,1582|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|Family Medical History|1579,1582|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|Family Medical History|1588,1591|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|Family Medical History|1588,1591|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|Family Medical History|1588,1591|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|Family Medical History|1588,1591|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|Family Medical History|1597,1600|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|Family Medical History|1597,1600|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|Family Medical History|1606,1609|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|Family Medical History|1606,1609|false|false|false|||MCV
Lab|Laboratory or Test Result|Family Medical History|1606,1609|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|Family Medical History|1606,1609|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|Family Medical History|1606,1609|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|Family Medical History|1614,1617|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|Family Medical History|1614,1617|false|false|false|C0600370|methacholine|MCH
Event|Event|Family Medical History|1614,1617|false|false|false|||MCH
Finding|Gene or Genome|Family Medical History|1614,1617|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|Family Medical History|1614,1617|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|Family Medical History|1614,1617|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|Family Medical History|1623,1627|false|false|false|||MCHC
Procedure|Laboratory Procedure|Family Medical History|1623,1627|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|Family Medical History|1642,1645|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|Family Medical History|1662,1667|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|1662,1667|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|1662,1667|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|Family Medical History|1668,1671|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|Family Medical History|1676,1679|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|Family Medical History|1676,1679|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|Family Medical History|1676,1679|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|Family Medical History|1685,1688|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|Family Medical History|1685,1688|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|Family Medical History|1685,1688|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|Family Medical History|1685,1688|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|Family Medical History|1694,1697|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|Family Medical History|1694,1697|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|Family Medical History|1703,1706|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|Family Medical History|1703,1706|false|false|false|||MCV
Lab|Laboratory or Test Result|Family Medical History|1703,1706|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|Family Medical History|1703,1706|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|Family Medical History|1703,1706|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|Family Medical History|1711,1714|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|Family Medical History|1711,1714|false|false|false|C0600370|methacholine|MCH
Event|Event|Family Medical History|1711,1714|false|false|false|||MCH
Finding|Gene or Genome|Family Medical History|1711,1714|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|Family Medical History|1711,1714|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|Family Medical History|1711,1714|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|Family Medical History|1720,1724|false|false|false|||MCHC
Procedure|Laboratory Procedure|Family Medical History|1720,1724|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|Family Medical History|1739,1742|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|Family Medical History|1759,1764|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|1759,1764|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|1759,1764|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|Family Medical History|1759,1772|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|Family Medical History|1759,1772|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|Family Medical History|1759,1772|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|Family Medical History|1765,1772|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|Family Medical History|1765,1772|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|Family Medical History|1765,1772|false|false|false|C0017725|glucose|Glucose
Event|Event|Family Medical History|1765,1772|false|false|false|||Glucose
Lab|Laboratory or Test Result|Family Medical History|1765,1772|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|Family Medical History|1765,1772|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|Family Medical History|1817,1821|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|Family Medical History|1817,1821|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|Family Medical History|1817,1821|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|Family Medical History|1846,1851|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|1846,1851|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|1846,1851|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|Family Medical History|1846,1859|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|Family Medical History|1846,1859|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|Family Medical History|1846,1859|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|Family Medical History|1852,1859|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|Family Medical History|1852,1859|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|Family Medical History|1852,1859|false|false|false|C0017725|glucose|Glucose
Event|Event|Family Medical History|1852,1859|false|false|false|||Glucose
Lab|Laboratory or Test Result|Family Medical History|1852,1859|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|Family Medical History|1852,1859|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|Family Medical History|1904,1908|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|Family Medical History|1904,1908|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|Family Medical History|1904,1908|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|Family Medical History|1933,1938|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|1933,1938|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|1933,1938|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|Family Medical History|1933,1946|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|Family Medical History|1933,1946|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|Family Medical History|1933,1946|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|Family Medical History|1939,1946|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|Family Medical History|1939,1946|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|Family Medical History|1939,1946|false|false|false|C0017725|glucose|Glucose
Event|Event|Family Medical History|1939,1946|false|false|false|||Glucose
Lab|Laboratory or Test Result|Family Medical History|1939,1946|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|Family Medical History|1939,1946|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|Family Medical History|1990,1994|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|Family Medical History|1990,1994|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|Family Medical History|1990,1994|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|Family Medical History|2019,2024|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|2019,2024|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|2019,2024|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|Family Medical History|2051,2056|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|2051,2056|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|2051,2056|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|Family Medical History|2057,2062|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|Family Medical History|2057,2062|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|Family Medical History|2057,2062|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|Family Medical History|2057,2062|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Drug|Organic Chemical|Family Medical History|2060,2064|false|false|false|C0602254|MB 3|MB-3
Disorder|Disease or Syndrome|Family Medical History|2091,2096|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|2091,2096|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|2091,2096|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|Family Medical History|2097,2102|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|Family Medical History|2097,2102|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|Family Medical History|2097,2102|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|Family Medical History|2097,2102|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Anatomy|Body System|Family Medical History|2144,2154|false|false|false|C0007226|Cardiovascular system|Cardiology
Attribute|Clinical Attribute|Family Medical History|2155,2161|false|false|false|C4255046||Report
Event|Event|Family Medical History|2155,2161|false|false|false|||Report
Finding|Intellectual Product|Family Medical History|2155,2161|false|false|false|C0684224|Report (document)|Report
Procedure|Health Care Activity|Family Medical History|2155,2161|false|false|false|C0700287|Reporting|Report
Attribute|Clinical Attribute|Family Medical History|2162,2168|false|false|false|C1718621|W stress|Stress
Drug|Organic Chemical|Family Medical History|2162,2168|false|false|false|C0723460|Stress bismuth subsalicylate|Stress
Drug|Pharmacologic Substance|Family Medical History|2162,2168|false|false|false|C0723460|Stress bismuth subsalicylate|Stress
Finding|Finding|Family Medical History|2162,2168|false|false|false|C0038435|Stress|Stress
Procedure|Diagnostic Procedure|Family Medical History|2162,2174|false|false|false|C0809864|stress study|Stress Study
Event|Event|Family Medical History|2169,2174|false|false|false|||Study
Finding|Intellectual Product|Family Medical History|2169,2174|false|false|false|C1705923|Study Object|Study
Procedure|Research Activity|Family Medical History|2169,2174|false|false|false|C0008972;C0947630;C2603343|Clinical Research;Scientific Study;Study|Study
Finding|Daily or Recreational Activity|Family Medical History|2195,2203|false|false|false|C0015259|Exercise|EXERCISE
Procedure|Therapeutic or Preventive Procedure|Family Medical History|2195,2203|false|false|false|C1522704|Exercise Pain Management|EXERCISE
Event|Event|Family Medical History|2204,2211|false|false|false|||RESULTS
Finding|Daily or Recreational Activity|Family Medical History|2219,2226|false|false|false|C0035253|Rest|RESTING
Event|Event|Family Medical History|2227,2231|false|false|false|||DATA
Finding|Idea or Concept|Family Medical History|2227,2231|false|false|false|C1511726|Data|DATA
Event|Event|Family Medical History|2233,2236|false|false|false|||EKG
Finding|Intellectual Product|Family Medical History|2233,2236|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|Family Medical History|2233,2236|false|false|false|C1623258|Electrocardiography|EKG
Anatomy|Body Space or Junction|Family Medical History|2239,2244|false|false|false|C0030471;C1305231|Nasal sinus;Sinus - general anatomical term|SINUS
Disorder|Anatomical Abnormality|Family Medical History|2239,2244|false|false|false|C0016169|pathologic fistula|SINUS
Drug|Organic Chemical|Family Medical History|2239,2244|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|SINUS
Drug|Pharmacologic Substance|Family Medical History|2239,2244|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|SINUS
Event|Event|Family Medical History|2239,2244|false|false|false|||SINUS
Event|Event|Family Medical History|2250,2253|false|false|false|||AEA
Finding|Finding|Family Medical History|2250,2253|false|false|false|C5676667|Anti-enterocyte antibody positivity|AEA
Disorder|Disease or Syndrome|Family Medical History|2255,2259|false|false|false|C0023211|Left Bundle-Branch Block|LBBB
Event|Event|Family Medical History|2255,2259|false|false|false|||LBBB
Lab|Laboratory or Test Result|Family Medical History|2255,2259|false|false|false|C0344420||LBBB
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2263,2268|false|false|false|C0018787;C4037974|Chest>Heart;Heart|HEART
Disorder|Neoplastic Process|Family Medical History|2263,2268|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|HEART
Finding|Sign or Symptom|Family Medical History|2263,2268|false|false|false|C0795691|HEART PROBLEM|HEART
Attribute|Clinical Attribute|Family Medical History|2263,2273|false|false|false|C0018810;C0488794|heart rate|HEART RATE
Finding|Finding|Family Medical History|2263,2273|false|false|false|C2041121||HEART RATE
Procedure|Health Care Activity|Family Medical History|2263,2273|false|false|false|C2197023|examination of heart rate|HEART RATE
Event|Activity|Family Medical History|2269,2273|false|false|false|C0871208|Rating (action)|RATE
Event|Event|Family Medical History|2269,2273|false|false|false|||RATE
Finding|Idea or Concept|Family Medical History|2269,2273|false|false|false|C1549480|Amount type - Rate|RATE
Disorder|Disease or Syndrome|Family Medical History|2279,2284|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|2279,2284|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|2279,2284|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Finding|Finding|Family Medical History|2279,2293|false|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|BLOOD PRESSURE
Finding|Organism Function|Family Medical History|2279,2293|false|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|BLOOD PRESSURE
Procedure|Health Care Activity|Family Medical History|2279,2293|false|false|false|C0005824|Blood pressure determination|BLOOD PRESSURE
Event|Event|Family Medical History|2285,2293|false|false|false|||PRESSURE
Finding|Finding|Family Medical History|2285,2293|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|PRESSURE
Finding|Functional Concept|Family Medical History|2285,2293|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|PRESSURE
Finding|Organ or Tissue Function|Family Medical History|2285,2293|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|PRESSURE
Phenomenon|Phenomenon or Process|Family Medical History|2285,2293|false|false|false|C0033095||PRESSURE
Finding|Finding|Family Medical History|2307,2315|false|false|false|C0442711;C1507394;C1522729;C2348563;C3715209|Clinical trial protocol document;Library Protocol;Protocol - answer to question;Protocols documentation;Study Protocol|PROTOCOL
Finding|Intellectual Product|Family Medical History|2307,2315|false|false|false|C0442711;C1507394;C1522729;C2348563;C3715209|Clinical trial protocol document;Library Protocol;Protocol - answer to question;Protocols documentation;Study Protocol|PROTOCOL
Event|Event|Family Medical History|2316,2324|false|false|false|||MODIFIED
Attribute|Clinical Attribute|Family Medical History|2341,2346|false|false|false|C1300072|Tumor stage|STAGE
Event|Event|Family Medical History|2347,2351|false|false|false|||TIME
Finding|Finding|Family Medical History|2347,2351|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|TIME
Finding|Idea or Concept|Family Medical History|2347,2351|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|TIME
Finding|Intellectual Product|Family Medical History|2347,2351|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|TIME
Drug|Hazardous or Poisonous Substance|Family Medical History|2352,2357|false|false|false|C0002658;C0025611|amphetamine;methamphetamine|SPEED
Drug|Organic Chemical|Family Medical History|2352,2357|false|false|false|C0002658;C0025611|amphetamine;methamphetamine|SPEED
Drug|Pharmacologic Substance|Family Medical History|2352,2357|false|false|false|C0002658;C0025611|amphetamine;methamphetamine|SPEED
Procedure|Therapeutic or Preventive Procedure|Family Medical History|2358,2367|false|false|false|C0439775|Elevation procedure|ELEVATION
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2368,2373|false|false|false|C0018787;C4037974|Chest>Heart;Heart|HEART
Disorder|Neoplastic Process|Family Medical History|2368,2373|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|HEART
Finding|Sign or Symptom|Family Medical History|2368,2373|false|false|false|C0795691|HEART PROBLEM|HEART
Disorder|Disease or Syndrome|Family Medical History|2374,2379|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|2374,2379|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|2374,2379|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Event|Event|Family Medical History|2380,2383|false|false|false|||RPP
Drug|Organic Chemical|Family Medical History|2394,2397|false|false|false|C0025810;C0048853|5,10-dihydro-5-methylphenazine;methylphenidate|MPH
Drug|Pharmacologic Substance|Family Medical History|2394,2397|false|false|false|C0025810;C0048853|5,10-dihydro-5-methylphenazine;methylphenidate|MPH
Event|Event|Family Medical History|2394,2397|false|false|false|||MPH
Finding|Intellectual Product|Family Medical History|2394,2397|false|false|false|C1513008|Master of Public Health|MPH
Event|Activity|Family Medical History|2403,2407|false|false|false|C0871208|Rating (action)|RATE
Finding|Idea or Concept|Family Medical History|2403,2407|false|false|false|C1549480|Amount type - Rate|RATE
Event|Event|Family Medical History|2408,2416|false|false|false|||PRESSURE
Finding|Finding|Family Medical History|2408,2416|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|PRESSURE
Finding|Functional Concept|Family Medical History|2408,2416|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|PRESSURE
Finding|Organ or Tissue Function|Family Medical History|2408,2416|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|PRESSURE
Phenomenon|Phenomenon or Process|Family Medical History|2408,2416|false|false|false|C0033095||PRESSURE
Event|Event|Family Medical History|2508,2516|false|false|false|||EXERCISE
Finding|Daily or Recreational Activity|Family Medical History|2508,2516|false|false|false|C0015259|Exercise|EXERCISE
Procedure|Therapeutic or Preventive Procedure|Family Medical History|2508,2516|false|false|false|C1522704|Exercise Pain Management|EXERCISE
Event|Event|Family Medical History|2517,2521|false|false|false|||TIME
Finding|Finding|Family Medical History|2517,2521|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|TIME
Finding|Idea or Concept|Family Medical History|2517,2521|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|TIME
Finding|Intellectual Product|Family Medical History|2517,2521|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|TIME
Drug|Amino Acid, Peptide, or Protein|Family Medical History|2528,2531|false|false|false|C1506708|MAX protein, human|MAX
Drug|Biologically Active Substance|Family Medical History|2528,2531|false|false|false|C1506708|MAX protein, human|MAX
Finding|Finding|Family Medical History|2528,2531|false|false|false|C0919516;C0919551;C4760036|MAX gene;Max (cigarettes);Oncogene MAX|MAX
Finding|Gene or Genome|Family Medical History|2528,2531|false|false|false|C0919516;C0919551;C4760036|MAX gene;Max (cigarettes);Oncogene MAX|MAX
Attribute|Clinical Attribute|Family Medical History|2532,2535|false|false|false|C5848651;C5848652||HRT
Event|Event|Family Medical History|2532,2535|false|false|false|||HRT
Procedure|Therapeutic or Preventive Procedure|Family Medical History|2532,2535|false|false|false|C0282402|Hormone replacement therapy|HRT
Event|Activity|Family Medical History|2536,2540|false|false|false|C0871208|Rating (action)|RATE
Event|Event|Family Medical History|2536,2540|false|false|false|||RATE
Finding|Idea or Concept|Family Medical History|2536,2540|false|false|false|C1549480|Amount type - Rate|RATE
Finding|Finding|Family Medical History|2541,2549|false|false|false|C5453128|Achieved|ACHIEVED
Event|Event|Family Medical History|2558,2566|false|false|false|||SYMPTOMS
Finding|Functional Concept|Family Medical History|2558,2566|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|SYMPTOMS
Finding|Sign or Symptom|Family Medical History|2558,2566|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|SYMPTOMS
Finding|Finding|Family Medical History|2568,2576|false|false|false|C0741302|atypia morphology|ATYPICAL
Attribute|Clinical Attribute|Family Medical History|2603,2617|false|false|false|C3173575||INTERPRETATION
Event|Event|Family Medical History|2603,2617|false|false|false|||INTERPRETATION
Finding|Intellectual Product|Family Medical History|2603,2617|false|false|false|C0459471|Interpretation Process|INTERPRETATION
Event|Event|Family Medical History|2636,2644|false|false|false|||referred
Event|Event|Family Medical History|2648,2656|false|false|false|||evaluate
Event|Event|Family Medical History|2660,2668|false|false|false|||atypical
Finding|Finding|Family Medical History|2660,2668|false|false|false|C0741302|atypia morphology|atypical
Anatomy|Body Location or Region|Family Medical History|2671,2676|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Family Medical History|2671,2676|false|false|false|C0741025|Chest problem|chest
Finding|Sign or Symptom|Family Medical History|2671,2687|false|false|false|C0235710|Chest discomfort|chest discomfort
Event|Event|Family Medical History|2677,2687|false|false|false|||discomfort
Finding|Sign or Symptom|Family Medical History|2677,2687|false|false|false|C2364135|Discomfort|discomfort
Finding|Body Substance|Family Medical History|2693,2700|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Family Medical History|2693,2700|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Family Medical History|2693,2700|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Family Medical History|2701,2710|false|false|false|||completed
Event|Event|Family Medical History|2735,2743|false|false|false|||protocol
Finding|Finding|Family Medical History|2735,2743|false|false|false|C0442711;C1507394;C1522729;C2348563;C3715209|Clinical trial protocol document;Library Protocol;Protocol - answer to question;Protocols documentation;Study Protocol|protocol
Finding|Intellectual Product|Family Medical History|2735,2743|false|false|false|C0442711;C1507394;C1522729;C2348563;C3715209|Clinical trial protocol document;Library Protocol;Protocol - answer to question;Protocols documentation;Study Protocol|protocol
Event|Event|Family Medical History|2745,2757|false|false|false|||representing
Event|Event|Family Medical History|2765,2773|false|false|false|||exercise
Finding|Daily or Recreational Activity|Family Medical History|2765,2773|false|false|false|C0015259|Exercise|exercise
Procedure|Therapeutic or Preventive Procedure|Family Medical History|2765,2773|false|false|false|C1522704|Exercise Pain Management|exercise
Attribute|Clinical Attribute|Family Medical History|2765,2783|false|false|false|C0162521;C2709256|Exercise Tolerance|exercise tolerance
Finding|Finding|Family Medical History|2765,2783|false|false|false|C2024889||exercise tolerance
Event|Event|Family Medical History|2774,2783|false|false|false|||tolerance
Finding|Finding|Family Medical History|2774,2783|false|false|false|C0013220;C0020963;C0220929;C0231197|Drug Tolerance;Immune Tolerance;Mental tolerance;Physiologic tolerance|tolerance
Finding|Mental Process|Family Medical History|2774,2783|false|false|false|C0013220;C0020963;C0220929;C0231197|Drug Tolerance;Immune Tolerance;Mental tolerance;Physiologic tolerance|tolerance
Finding|Pathologic Function|Family Medical History|2774,2783|false|false|false|C0013220;C0020963;C0220929;C0231197|Drug Tolerance;Immune Tolerance;Mental tolerance;Physiologic tolerance|tolerance
Finding|Physiologic Function|Family Medical History|2774,2783|false|false|false|C0013220;C0020963;C0220929;C0231197|Drug Tolerance;Immune Tolerance;Mental tolerance;Physiologic tolerance|tolerance
Attribute|Clinical Attribute|Family Medical History|2792,2795|false|true|false|C1114365||age
Drug|Biologically Active Substance|Family Medical History|2792,2795|false|true|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|Family Medical History|2792,2795|false|true|false|C0162574|Glycation End Products, Advanced|age
Event|Event|Family Medical History|2792,2795|false|false|false|||age
Event|Event|Family Medical History|2803,2807|false|false|false|||METS
Finding|Gene or Genome|Family Medical History|2803,2807|false|false|false|C0812270;C1705694|ETV3 gene;ETV3 wt Allele|METS
Event|Event|Family Medical History|2815,2823|false|false|false|||exercise
Finding|Daily or Recreational Activity|Family Medical History|2815,2823|false|false|false|C0015259|Exercise|exercise
Procedure|Therapeutic or Preventive Procedure|Family Medical History|2815,2823|false|false|false|C1522704|Exercise Pain Management|exercise
Procedure|Diagnostic Procedure|Family Medical History|2815,2828|false|false|false|C0015260|Exercise stress test|exercise test
Anatomy|Body Location or Region|Family Medical History|2824,2828|false|false|false|C4318744|Test - temporal region|test
Event|Event|Family Medical History|2824,2828|false|false|false|||test
Finding|Functional Concept|Family Medical History|2824,2828|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Finding|Intellectual Product|Family Medical History|2824,2828|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Lab|Laboratory or Test Result|Family Medical History|2824,2828|false|false|false|C0456984|Test Result|test
Procedure|Laboratory Procedure|Family Medical History|2824,2828|false|false|false|C0022885|Laboratory Procedures|test
Event|Event|Family Medical History|2833,2840|false|false|false|||stopped
Finding|Body Substance|Family Medical History|2848,2855|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Family Medical History|2848,2855|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Family Medical History|2848,2855|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Activity|Family Medical History|2858,2865|false|false|false|C1272683||request
Event|Event|Family Medical History|2858,2865|false|false|false|||request
Finding|Idea or Concept|Family Medical History|2858,2865|false|false|false|C1522634;C1553397;C1553888|Question (inquiry);Request - ActReason;request - ActMood|request
Finding|Intellectual Product|Family Medical History|2858,2865|false|false|false|C1522634;C1553397;C1553888|Question (inquiry);Request - ActReason;request - ActMood|request
Disorder|Neoplastic Process|Family Medical History|2866,2875|false|false|false|C0027627|Neoplasm Metastasis|secondary
Event|Event|Family Medical History|2866,2875|false|false|false|||secondary
Finding|Functional Concept|Family Medical History|2866,2875|false|false|false|C1522484|metastatic qualifier|secondary
Event|Event|Family Medical History|2880,2887|false|false|false|||fatigue
Finding|Sign or Symptom|Family Medical History|2880,2887|false|false|false|C0015672|Fatigue|fatigue
Event|Event|Family Medical History|2897,2905|false|false|false|||exercise
Finding|Daily or Recreational Activity|Family Medical History|2897,2905|false|false|false|C0015259|Exercise|exercise
Procedure|Therapeutic or Preventive Procedure|Family Medical History|2897,2905|false|false|false|C1522704|Exercise Pain Management|exercise
Finding|Body Substance|Family Medical History|2911,2918|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Family Medical History|2911,2918|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Family Medical History|2911,2918|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Family Medical History|2919,2927|false|false|false|||reported
Finding|Functional Concept|Family Medical History|2948,2956|false|false|false|C0205409;C1548221|Bed Status - Isolated;Isolated|isolated
Finding|Idea or Concept|Family Medical History|2948,2956|false|false|false|C0205409;C1548221|Bed Status - Isolated;Isolated|isolated
Finding|Functional Concept|Family Medical History|2964,2968|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|Family Medical History|2975,2980|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Family Medical History|2975,2980|false|false|false|C0741025|Chest problem|chest
Finding|Sign or Symptom|Family Medical History|2975,2991|false|false|false|C0235710|Chest discomfort|chest discomfort
Event|Event|Family Medical History|2981,2991|false|false|false|||discomfort
Finding|Sign or Symptom|Family Medical History|2981,2991|false|false|false|C2364135|Discomfort|discomfort
Event|Governmental or Regulatory Activity|Family Medical History|3002,3006|false|false|false|C1510751|Academic Research Enhancement Awards|area
Event|Event|Family Medical History|3010,3020|false|false|false|||discomfort
Finding|Sign or Symptom|Family Medical History|3010,3020|false|false|false|C2364135|Discomfort|discomfort
Event|Event|Family Medical History|3038,3044|false|false|false|||tender
Event|Event|Family Medical History|3048,3057|false|false|false|||palpation
Procedure|Diagnostic Procedure|Family Medical History|3048,3057|false|false|false|C0030247|Palpation|palpation
Event|Event|Family Medical History|3064,3074|true|false|false|||discomfort
Finding|Sign or Symptom|Family Medical History|3064,3074|true|false|false|C2364135|Discomfort|discomfort
Event|Event|Family Medical History|3075,3083|true|false|false|||resolved
Drug|Amino Acid, Peptide, or Protein|Family Medical History|3089,3093|true|false|false|C1742913|REST protein, human|rest
Drug|Biologically Active Substance|Family Medical History|3089,3093|true|false|false|C1742913|REST protein, human|rest
Event|Event|Family Medical History|3089,3093|true|false|false|||rest
Finding|Daily or Recreational Activity|Family Medical History|3089,3093|true|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Gene or Genome|Family Medical History|3089,3093|true|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Molecular Function|Family Medical History|3089,3093|true|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Functional Concept|Family Medical History|3103,3109|false|false|false|C0332197|Absent|absent
Lab|Laboratory or Test Result|Family Medical History|3103,3109|false|false|false|C5237010|Expression Negative|absent
Event|Event|Family Medical History|3145,3153|false|false|false|||presence
Procedure|Therapeutic or Preventive Procedure|Family Medical History|3145,3153|false|false|false|C0392148|Providing presence (regime/therapy)|presence
Finding|Finding|Family Medical History|3145,3156|false|false|false|C0150312|Present|presence of
Disorder|Disease or Syndrome|Family Medical History|3161,3165|false|false|false|C0023211|Left Bundle-Branch Block|LBBB
Event|Event|Family Medical History|3161,3165|false|false|false|||LBBB
Lab|Laboratory or Test Result|Family Medical History|3161,3165|false|false|false|C0344420||LBBB
Event|Event|Family Medical History|3189,3204|false|false|false|||uninterpretable
Event|Event|Family Medical History|3209,3217|false|false|false|||ischemia
Finding|Pathologic Function|Family Medical History|3209,3217|false|false|false|C0022116|Ischemia|ischemia
Procedure|Therapeutic or Preventive Procedure|Family Medical History|3209,3217|false|false|false|C4321499|Ischemia Procedure|ischemia
Event|Event|Family Medical History|3223,3229|false|false|false|||rhythm
Finding|Finding|Family Medical History|3223,3229|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|Family Medical History|3223,3229|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Anatomy|Body Space or Junction|Family Medical History|3234,3239|false|false|false|C0030471;C1305231|Nasal sinus;Sinus - general anatomical term|sinus
Disorder|Anatomical Abnormality|Family Medical History|3234,3239|false|false|false|C0016169|pathologic fistula|sinus
Drug|Organic Chemical|Family Medical History|3234,3239|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Drug|Pharmacologic Substance|Family Medical History|3234,3239|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Event|Event|Family Medical History|3234,3239|false|false|false|||sinus
Finding|Functional Concept|Family Medical History|3256,3264|false|false|false|C0205409;C1548221|Bed Status - Isolated;Isolated|isolated
Finding|Idea or Concept|Family Medical History|3256,3264|false|false|false|C0205409;C1548221|Bed Status - Isolated;Isolated|isolated
Disorder|Disease or Syndrome|Family Medical History|3265,3269|false|false|false|C3714976|ACTIVATED PI3K-DELTA SYNDROME|APDs
Drug|Organic Chemical|Family Medical History|3265,3269|false|false|false|C0043603|pamidronate|APDs
Drug|Pharmacologic Substance|Family Medical History|3265,3269|false|false|false|C0043603|pamidronate|APDs
Event|Event|Family Medical History|3265,3269|false|false|false|||APDs
Finding|Gene or Genome|Family Medical History|3265,3269|false|false|false|C3714973|PIK3CD wt Allele|APDs
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|3285,3291|false|false|false|C0018792|Heart Atrium|atrial
Event|Event|Family Medical History|3292,3300|false|false|false|||couplets
Finding|Finding|Family Medical History|3292,3300|false|false|false|C0429001|Paired ventricular premature complexes|couplets
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|3305,3311|false|false|false|C0018792|Heart Atrium|atrial
Event|Event|Family Medical History|3313,3321|false|false|false|||triplets
Finding|Daily or Recreational Activity|Family Medical History|3324,3331|false|false|false|C0035253|Rest|Resting
Finding|Intellectual Product|Family Medical History|3332,3336|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Organ or Tissue Function|Family Medical History|3337,3345|false|false|false|C0039155|Systole|systolic
Disorder|Disease or Syndrome|Family Medical History|3337,3358|false|false|false|C0221155|Systolic Hypertension|systolic hypertension
Disorder|Disease or Syndrome|Family Medical History|3346,3358|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|Family Medical History|3346,3358|false|false|false|||hypertension
Disorder|Disease or Syndrome|Family Medical History|3371,3376|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Family Medical History|3371,3376|false|false|false|||blood
Finding|Body Substance|Family Medical History|3371,3376|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Finding|Family Medical History|3371,3385|false|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|blood pressure
Finding|Organism Function|Family Medical History|3371,3385|false|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|blood pressure
Procedure|Health Care Activity|Family Medical History|3371,3385|false|false|false|C0005824|Blood pressure determination|blood pressure
Event|Event|Family Medical History|3377,3385|false|false|false|||pressure
Finding|Finding|Family Medical History|3377,3385|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|Family Medical History|3377,3385|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|Family Medical History|3377,3385|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|Family Medical History|3377,3385|false|false|false|C0033095||pressure
Event|Event|Family Medical History|3387,3395|false|false|false|||response
Finding|Finding|Family Medical History|3387,3395|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Intellectual Product|Family Medical History|3387,3395|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Mental Process|Family Medical History|3387,3395|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Event|Event|Family Medical History|3400,3408|false|false|false|||exercise
Finding|Daily or Recreational Activity|Family Medical History|3400,3408|false|false|false|C0015259|Exercise|exercise
Procedure|Therapeutic or Preventive Procedure|Family Medical History|3400,3408|false|false|false|C1522704|Exercise Pain Management|exercise
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|3414,3419|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Family Medical History|3414,3419|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Family Medical History|3414,3419|false|false|false|C0795691|HEART PROBLEM|heart
Attribute|Clinical Attribute|Family Medical History|3414,3424|false|false|false|C0018810;C0488794|heart rate|heart rate
Finding|Finding|Family Medical History|3414,3424|false|false|false|C2041121||heart rate
Procedure|Health Care Activity|Family Medical History|3414,3424|false|false|false|C2197023|examination of heart rate|heart rate
Attribute|Clinical Attribute|Family Medical History|3414,3433|false|false|false|C1997754|Heart rate response (observable entity)|heart rate response
Event|Activity|Family Medical History|3420,3424|false|false|false|C0871208|Rating (action)|rate
Event|Event|Family Medical History|3420,3424|false|false|false|||rate
Finding|Idea or Concept|Family Medical History|3420,3424|false|false|false|C1549480|Amount type - Rate|rate
Event|Event|Family Medical History|3425,3433|false|false|false|||response
Finding|Finding|Family Medical History|3425,3433|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Intellectual Product|Family Medical History|3425,3433|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Mental Process|Family Medical History|3425,3433|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Organism Function|Family Medical History|3425,3445|false|false|false|C2265833|response to exercise|response to exercise
Event|Event|Family Medical History|3437,3445|false|false|false|||exercise
Finding|Daily or Recreational Activity|Family Medical History|3437,3445|false|false|false|C0015259|Exercise|exercise
Procedure|Therapeutic or Preventive Procedure|Family Medical History|3437,3445|false|false|false|C1522704|Exercise Pain Management|exercise
Event|Event|Family Medical History|3458,3465|false|false|false|||blunted
Event|Event|Family Medical History|3471,3481|false|false|false|||IMPRESSION
Finding|Intellectual Product|Family Medical History|3471,3481|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|Family Medical History|3471,3481|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Event|Event|Family Medical History|3488,3496|false|false|false|||exercise
Finding|Daily or Recreational Activity|Family Medical History|3488,3496|false|false|false|C0015259|Exercise|exercise
Procedure|Therapeutic or Preventive Procedure|Family Medical History|3488,3496|false|false|false|C1522704|Exercise Pain Management|exercise
Attribute|Clinical Attribute|Family Medical History|3488,3506|false|false|false|C0162521;C2709256|Exercise Tolerance|exercise tolerance
Finding|Finding|Family Medical History|3488,3506|false|false|false|C2024889||exercise tolerance
Event|Event|Family Medical History|3497,3506|false|false|false|||tolerance
Finding|Finding|Family Medical History|3497,3506|false|false|false|C0013220;C0020963;C0220929;C0231197|Drug Tolerance;Immune Tolerance;Mental tolerance;Physiologic tolerance|tolerance
Finding|Mental Process|Family Medical History|3497,3506|false|false|false|C0013220;C0020963;C0220929;C0231197|Drug Tolerance;Immune Tolerance;Mental tolerance;Physiologic tolerance|tolerance
Finding|Pathologic Function|Family Medical History|3497,3506|false|false|false|C0013220;C0020963;C0220929;C0231197|Drug Tolerance;Immune Tolerance;Mental tolerance;Physiologic tolerance|tolerance
Finding|Physiologic Function|Family Medical History|3497,3506|false|false|false|C0013220;C0020963;C0220929;C0231197|Drug Tolerance;Immune Tolerance;Mental tolerance;Physiologic tolerance|tolerance
Event|Event|Family Medical History|3519,3527|true|false|false|||symptoms
Finding|Functional Concept|Family Medical History|3519,3527|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Family Medical History|3519,3527|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Drug|Amino Acid, Peptide, or Protein|Family Medical History|3550,3553|true|false|false|C0018064|Equine Gonadotropins|ECG
Drug|Hormone|Family Medical History|3550,3553|true|false|false|C0018064|Equine Gonadotropins|ECG
Drug|Pharmacologic Substance|Family Medical History|3550,3553|true|false|false|C0018064|Equine Gonadotropins|ECG
Event|Event|Family Medical History|3550,3553|true|false|false|||ECG
Finding|Intellectual Product|Family Medical History|3550,3553|true|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|ECG
Procedure|Diagnostic Procedure|Family Medical History|3550,3553|true|false|false|C1623258|Electrocardiography|ECG
Event|Event|Family Medical History|3557,3565|false|false|false|||achieved
Event|Event|Family Medical History|3566,3574|false|false|false|||workload
Finding|Daily or Recreational Activity|Family Medical History|3576,3583|false|false|false|C0035253|Rest|Resting
Finding|Intellectual Product|Family Medical History|3584,3588|false|false|false|C1547225|Mild Severity of Illness Code|mild
Event|Event|Family Medical History|3589,3597|false|false|false|||systolic
Finding|Organ or Tissue Function|Family Medical History|3589,3597|false|false|false|C0039155|Systole|systolic
Disorder|Disease or Syndrome|Family Medical History|3599,3611|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|Family Medical History|3599,3611|false|false|false|||hypertension
Disorder|Disease or Syndrome|Family Medical History|3629,3634|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Family Medical History|3629,3634|false|false|false|||blood
Finding|Body Substance|Family Medical History|3629,3634|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Finding|Family Medical History|3629,3643|false|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|blood pressure
Finding|Organism Function|Family Medical History|3629,3643|false|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|blood pressure
Procedure|Health Care Activity|Family Medical History|3629,3643|false|false|false|C0005824|Blood pressure determination|blood pressure
Attribute|Clinical Attribute|Family Medical History|3629,3652|false|false|false|C1997183|Speed of blood pressure response|blood pressure response
Event|Event|Family Medical History|3635,3643|false|false|false|||pressure
Finding|Finding|Family Medical History|3635,3643|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|Family Medical History|3635,3643|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|Family Medical History|3635,3643|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|Family Medical History|3635,3643|false|false|false|C0033095||pressure
Event|Event|Family Medical History|3644,3652|false|false|false|||response
Finding|Finding|Family Medical History|3644,3652|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Intellectual Product|Family Medical History|3644,3652|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Mental Process|Family Medical History|3644,3652|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Event|Event|Family Medical History|3657,3665|false|false|false|||exercise
Finding|Daily or Recreational Activity|Family Medical History|3657,3665|false|false|false|C0015259|Exercise|exercise
Procedure|Therapeutic or Preventive Procedure|Family Medical History|3657,3665|false|false|false|C1522704|Exercise Pain Management|exercise
Event|Event|Family Medical History|3679,3684|true|false|false|||study
Finding|Intellectual Product|Family Medical History|3679,3684|true|false|false|C1705923|Study Object|study
Procedure|Research Activity|Family Medical History|3679,3684|true|false|false|C0008972;C0947630;C2603343|Clinical Research;Scientific Study;Study|study
Event|Event|Family Medical History|3687,3693|true|false|false|||target
Finding|Functional Concept|Family Medical History|3687,3693|true|false|false|C1521840|Target|target
Procedure|Research Activity|Family Medical History|3687,3693|true|false|false|C5575831|Therapeutically Applicable Research to Generate Effective Treatments|target
Procedure|Therapeutic or Preventive Procedure|Family Medical History|3687,3704|true|false|false|C0744682|Target heart rate|target heart rate
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|3694,3699|true|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Family Medical History|3694,3699|true|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Family Medical History|3694,3699|true|false|false|C0795691|HEART PROBLEM|heart
Attribute|Clinical Attribute|Family Medical History|3694,3704|true|false|false|C0018810;C0488794|heart rate|heart rate
Finding|Finding|Family Medical History|3694,3704|true|false|false|C2041121||heart rate
Procedure|Health Care Activity|Family Medical History|3694,3704|true|false|false|C2197023|examination of heart rate|heart rate
Event|Activity|Family Medical History|3700,3704|true|false|false|C0871208|Rating (action)|rate
Event|Event|Family Medical History|3700,3704|true|false|false|||rate
Finding|Idea or Concept|Family Medical History|3700,3704|true|false|false|C1549480|Amount type - Rate|rate
Event|Event|Family Medical History|3709,3717|true|false|false|||achieved
Event|Event|Family Medical History|3722,3728|false|false|false|||SIGNED
Finding|Idea or Concept|Hospital Course|3785,3790|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Intellectual Product|Hospital Course|3785,3790|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Event|Event|Hospital Course|3791,3798|false|false|false|||history
Finding|Conceptual Entity|Hospital Course|3791,3798|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|3791,3798|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Hospital Course|3791,3798|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|3791,3801|false|false|false|C0262926|Medical History|history of
Finding|Functional Concept|Hospital Course|3802,3806|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|3813,3816|false|false|false|C0446516;C1140618;C1269078|Upper Extremity;Upper arm|arm
Disorder|Anatomical Abnormality|Hospital Course|3813,3816|false|false|false|C3495676|Anorectal Malformations|arm
Event|Event|Hospital Course|3813,3816|false|false|false|||arm
Finding|Gene or Genome|Hospital Course|3813,3816|false|false|false|C1824218;C3715044|AKR1A1 wt Allele;ARMC9 gene|arm
Procedure|Diagnostic Procedure|Hospital Course|3813,3816|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Research Activity|Hospital Course|3813,3816|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3813,3816|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Anatomy|Body Location or Region|Hospital Course|3821,3826|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Hospital Course|3821,3826|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Hospital Course|3833,3837|false|true|false|C2598155||pain
Event|Event|Hospital Course|3833,3837|false|false|false|||pain
Finding|Functional Concept|Hospital Course|3833,3837|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|3833,3837|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Mental Process|Hospital Course|3845,3852|false|false|false|C0542559|contextual factors|setting
Disorder|Disease or Syndrome|Hospital Course|3856,3860|false|false|false|C0023211|Left Bundle-Branch Block|LBBB
Event|Event|Hospital Course|3856,3860|false|false|false|||LBBB
Lab|Laboratory or Test Result|Hospital Course|3856,3860|false|false|false|C0344420||LBBB
Event|Event|Hospital Course|3861,3871|false|false|false|||presenting
Anatomy|Body Location or Region|Hospital Course|3893,3898|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|Hospital Course|3893,3898|false|false|false|C0741025|Chest problem|Chest
Attribute|Clinical Attribute|Hospital Course|3893,3903|false|false|false|C2926613||Chest Pain
Finding|Sign or Symptom|Hospital Course|3893,3903|false|false|false|C0008031|Chest Pain|Chest Pain
Attribute|Clinical Attribute|Hospital Course|3899,3903|false|false|false|C2598155||Pain
Event|Event|Hospital Course|3899,3903|false|false|false|||Pain
Finding|Functional Concept|Hospital Course|3899,3903|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|Hospital Course|3899,3903|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Body Substance|Hospital Course|3908,3915|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|3908,3915|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|3908,3915|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|3918,3926|true|false|false|||symptoms
Finding|Functional Concept|Hospital Course|3918,3926|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Hospital Course|3918,3926|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|Hospital Course|3946,3953|true|false|false|||anginal
Finding|Functional Concept|Hospital Course|3958,3964|true|false|false|C0349590;C1262865|Nature;Natures|nature
Finding|Idea or Concept|Hospital Course|3958,3964|true|false|false|C0349590;C1262865|Nature;Natures|nature
Event|Event|Hospital Course|3968,3975|true|false|false|||suggest
Anatomy|Body Space or Junction|Hospital Course|3976,3979|false|false|false|C0262187|anterior calcarine sulcus (human only)|ACS
Disorder|Disease or Syndrome|Hospital Course|3976,3979|false|false|false|C0742343;C0796147|Acrocallosal Syndrome;Acute Chest Syndrome|ACS
Drug|Amino Acid, Peptide, or Protein|Hospital Course|3976,3979|false|false|false|C4042561|ACSS2 protein, human|ACS
Drug|Enzyme|Hospital Course|3976,3979|false|false|false|C4042561|ACSS2 protein, human|ACS
Event|Event|Hospital Course|3976,3979|false|false|false|||ACS
Finding|Gene or Genome|Hospital Course|3976,3979|false|false|false|C1150760;C1424787;C1825842;C1842089;C2266615;C4318612;C5400867;C5551036|ACCS gene;ACS - Activity Card Sort;ACSS2 gene;ACSS2 wt Allele;American Community Survey;CO-methylating acetyl-CoA synthase activity;PLA2G15 gene;acetate-CoA ligase activity|ACS
Finding|Intellectual Product|Hospital Course|3976,3979|false|false|false|C1150760;C1424787;C1825842;C1842089;C2266615;C4318612;C5400867;C5551036|ACCS gene;ACS - Activity Card Sort;ACSS2 gene;ACSS2 wt Allele;American Community Survey;CO-methylating acetyl-CoA synthase activity;PLA2G15 gene;acetate-CoA ligase activity|ACS
Finding|Molecular Function|Hospital Course|3976,3979|false|false|false|C1150760;C1424787;C1825842;C1842089;C2266615;C4318612;C5400867;C5551036|ACCS gene;ACS - Activity Card Sort;ACSS2 gene;ACSS2 wt Allele;American Community Survey;CO-methylating acetyl-CoA synthase activity;PLA2G15 gene;acetate-CoA ligase activity|ACS
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4011,4018|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|Hospital Course|4011,4018|false|true|false|C1314974|Cardiac attachment|cardiac
Finding|Idea or Concept|Hospital Course|4020,4024|false|false|false|C0035647|Risk|risk
Attribute|Clinical Attribute|Hospital Course|4020,4032|false|false|false|C1830376||risk factors
Finding|Finding|Hospital Course|4020,4032|false|false|false|C0035648;C0455624;C1553898|History of - risk factor;risk factors;risk factors - observation list|risk factors
Finding|Intellectual Product|Hospital Course|4020,4032|false|false|false|C0035648;C0455624;C1553898|History of - risk factor;risk factors;risk factors - observation list|risk factors
Event|Event|Hospital Course|4025,4032|false|false|false|||factors
Disorder|Disease or Syndrome|Hospital Course|4039,4043|true|false|false|C0023211|Left Bundle-Branch Block|LBBB
Event|Event|Hospital Course|4039,4043|true|false|false|||LBBB
Lab|Laboratory or Test Result|Hospital Course|4039,4043|true|false|false|C0344420||LBBB
Event|Event|Hospital Course|4049,4059|true|false|false|||physicians
Event|Event|Hospital Course|4071,4072|true|false|false|||r
Event|Event|Hospital Course|4073,4076|true|false|false|||oMI
Finding|Gene or Genome|Hospital Course|4073,4076|true|true|false|C1825553|HTRA2 gene|oMI
Event|Event|Hospital Course|4083,4086|true|false|false|||EKG
Finding|Intellectual Product|Hospital Course|4083,4086|true|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|Hospital Course|4083,4086|true|false|false|C1623258|Electrocardiography|EKG
Finding|Finding|Hospital Course|4087,4092|true|false|false|C0439044|Living Alone|alone
Event|Event|Hospital Course|4094,4098|false|false|false|||Trop
Event|Event|Hospital Course|4100,4107|false|false|false|||results
Event|Event|Hospital Course|4113,4121|false|false|false|||negative
Finding|Classification|Hospital Course|4113,4121|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|4113,4121|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|4113,4121|false|false|false|C5237010|Expression Negative|negative
Attribute|Clinical Attribute|Hospital Course|4126,4132|false|false|false|C1718621|W stress|Stress
Drug|Organic Chemical|Hospital Course|4126,4132|false|false|false|C0723460|Stress bismuth subsalicylate|Stress
Drug|Pharmacologic Substance|Hospital Course|4126,4132|false|false|false|C0723460|Stress bismuth subsalicylate|Stress
Event|Event|Hospital Course|4126,4132|false|false|false|||Stress
Finding|Finding|Hospital Course|4126,4132|false|false|false|C0038435|Stress|Stress
Procedure|Diagnostic Procedure|Hospital Course|4126,4137|false|false|false|C0920208|Echocardiography, Stress|Stress Echo
Event|Event|Hospital Course|4133,4137|false|false|false|||Echo
Procedure|Health Care Activity|Hospital Course|4133,4137|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|Echo
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4133,4137|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|Echo
Event|Event|Hospital Course|4138,4146|false|false|false|||revealed
Finding|Finding|Hospital Course|4148,4151|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Hospital Course|4148,4151|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Disorder|Disease or Syndrome|Hospital Course|4161,4172|false|false|false|C3887505|DYSFUNCTION - SKIN DISORDERS|dysfunction
Event|Event|Hospital Course|4161,4172|false|false|false|||dysfunction
Finding|Conceptual Entity|Hospital Course|4161,4172|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Functional Concept|Hospital Course|4161,4172|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Pathologic Function|Hospital Course|4161,4172|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Event|Event|Hospital Course|4178,4189|false|false|false|||hypokinesis
Finding|Finding|Hospital Course|4178,4189|false|false|false|C0086439|Hypokinesia|hypokinesis
Event|Event|Hospital Course|4197,4205|false|false|false|||inferior
Finding|Social Behavior|Hospital Course|4197,4205|false|false|false|C0678975|inferiority|inferior
Event|Event|Hospital Course|4231,4241|false|false|false|||consistent
Finding|Idea or Concept|Hospital Course|4231,4241|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|Hospital Course|4231,4246|false|false|false|C0332290|Consistent with|consistent with
Finding|Finding|Hospital Course|4247,4253|false|false|false|C0087136;C1549113|Marital Status - Single;Unmarried|single
Disorder|Disease or Syndrome|Hospital Course|4247,4268|false|false|false|C0856737|Single vessel disease|single vessel disease
Anatomy|Body Location or Region|Hospital Course|4254,4260|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4254,4260|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Disorder|Disease or Syndrome|Hospital Course|4261,4268|false|true|false|C0012634|Disease|disease
Event|Event|Hospital Course|4261,4268|false|false|false|||disease
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4277,4280|false|false|false|C0226047|Posterior interventricular branch of right coronary artery|PDA
Disorder|Congenital Abnormality|Hospital Course|4277,4280|false|false|false|C0013274;C1335302;C4282128|PATENT DUCTUS ARTERIOSUS 1;Pancreatic Ductal Adenocarcinoma;Patent ductus arteriosus|PDA
Disorder|Neoplastic Process|Hospital Course|4277,4280|false|false|false|C0013274;C1335302;C4282128|PATENT DUCTUS ARTERIOSUS 1;Pancreatic Ductal Adenocarcinoma;Patent ductus arteriosus|PDA
Event|Event|Hospital Course|4281,4293|false|false|false|||distribution
Finding|Cell Function|Hospital Course|4281,4293|false|false|false|C1704711;C5779816|Distribution;Distribution [PK]|distribution
Finding|Functional Concept|Hospital Course|4281,4293|false|false|false|C1704711;C5779816|Distribution;Distribution [PK]|distribution
Anatomy|Body System|Hospital Course|4297,4307|false|false|false|C0007226|Cardiovascular system|cardiology
Event|Event|Hospital Course|4308,4315|false|false|false|||consult
Procedure|Health Care Activity|Hospital Course|4308,4315|false|false|false|C0009818|Consultation|consult
Event|Event|Hospital Course|4320,4328|false|false|false|||obtained
Event|Event|Hospital Course|4333,4337|false|false|false|||they
Event|Event|Hospital Course|4339,4343|false|false|false|||felt
Event|Event|Hospital Course|4357,4364|false|false|false|||managed
Finding|Body Substance|Hospital Course|4376,4383|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|4376,4383|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|4376,4383|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Organic Chemical|Hospital Course|4403,4410|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|Hospital Course|4403,4410|false|false|false|C0004057|aspirin|aspirin
Event|Event|Hospital Course|4403,4410|false|false|false|||aspirin
Drug|Organic Chemical|Hospital Course|4418,4424|false|false|false|C0360714|Hydroxymethylglutaryl-CoA Reductase Inhibitors|statin
Drug|Pharmacologic Substance|Hospital Course|4418,4424|false|false|false|C0360714|Hydroxymethylglutaryl-CoA Reductase Inhibitors|statin
Event|Event|Hospital Course|4418,4424|false|false|false|||statin
Finding|Gene or Genome|Hospital Course|4418,4424|false|false|false|C1414273|EEF1A2 gene|statin
Event|Event|Hospital Course|4432,4439|false|false|false|||history
Finding|Conceptual Entity|Hospital Course|4432,4439|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|4432,4439|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Hospital Course|4432,4439|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Event|Event|Hospital Course|4443,4450|false|false|false|||suggest
Disorder|Disease or Syndrome|Hospital Course|4451,4457|false|false|false|C0004096|Asthma|asthma
Event|Event|Hospital Course|4451,4457|false|false|false|||asthma
Event|Event|Hospital Course|4460,4467|false|false|false|||blocker
Event|Event|Hospital Course|4473,4488|false|false|false|||contraindicated
Event|Event|Hospital Course|4498,4508|false|false|false|||discharged
Event|Event|Hospital Course|4519,4527|false|false|false|||extended
Event|Event|Hospital Course|4529,4536|false|false|false|||release
Finding|Functional Concept|Hospital Course|4529,4536|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|release
Procedure|Health Care Activity|Hospital Course|4529,4536|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4529,4536|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|release
Drug|Organic Chemical|Hospital Course|4537,4546|false|false|false|C0012373|diltiazem|diltiazem
Drug|Pharmacologic Substance|Hospital Course|4537,4546|false|false|false|C0012373|diltiazem|diltiazem
Event|Event|Hospital Course|4537,4546|false|false|false|||diltiazem
Attribute|Clinical Attribute|Hospital Course|4552,4564|false|false|false|C3263700||instructions
Event|Event|Hospital Course|4552,4564|false|false|false|||instructions
Finding|Intellectual Product|Hospital Course|4552,4564|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|instructions
Event|Event|Hospital Course|4568,4574|false|false|false|||follow
Anatomy|Body System|Hospital Course|4581,4591|false|false|false|C0007226|Cardiovascular system|cardiology
Disorder|Disease or Syndrome|Hospital Course|4606,4609|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|Hospital Course|4606,4609|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|Hospital Course|4606,4609|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|Hospital Course|4606,4609|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|Hospital Course|4606,4609|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|Hospital Course|4606,4609|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|Hospital Course|4606,4609|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|Hospital Course|4606,4609|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|Hospital Course|4606,4609|false|false|false|||PCP
Finding|Gene or Genome|Hospital Course|4606,4609|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|Hospital Course|4606,4609|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Disorder|Disease or Syndrome|Hospital Course|4616,4644|false|false|false|C0039240|Supraventricular tachycardia|Supraventricular tachycardia
Finding|Finding|Hospital Course|4616,4644|false|false|false|C3815188|Supraventricular Tachycardia by ECG Finding|Supraventricular tachycardia
Event|Event|Hospital Course|4633,4644|false|false|false|||tachycardia
Finding|Finding|Hospital Course|4633,4644|false|false|false|C0039231;C3827868|Tachycardia;Tachycardia by ECG Finding|tachycardia
Finding|Body Substance|Hospital Course|4650,4657|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|4650,4657|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|4650,4657|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|4671,4675|false|false|false|||runs
Finding|Finding|Hospital Course|4671,4675|false|false|false|C0600140|Does run (finding)|runs
Disorder|Disease or Syndrome|Hospital Course|4680,4683|false|false|false|C0039240|Supraventricular tachycardia|SVT
Event|Event|Hospital Course|4680,4683|false|false|false|||SVT
Finding|Finding|Hospital Course|4680,4683|false|false|false|C3815188|Supraventricular Tachycardia by ECG Finding|SVT
Event|Event|Hospital Course|4700,4703|false|false|false|||MAT
Finding|Finding|Hospital Course|4700,4703|false|false|false|C0221158;C1151970;C1412111;C1417038;C3714902;C5780814;C5890859|ACAT1 gene;ACAT1 wt Allele;MAT1A gene;MAT1A wt Allele;Multifocal atrial tachycardia;Multinational Association of Supportive Care in Cancer Antiemesis Tool;[acyl-carrier-protein] S-malonyltransferase activity|MAT
Finding|Gene or Genome|Hospital Course|4700,4703|false|false|false|C0221158;C1151970;C1412111;C1417038;C3714902;C5780814;C5890859|ACAT1 gene;ACAT1 wt Allele;MAT1A gene;MAT1A wt Allele;Multifocal atrial tachycardia;Multinational Association of Supportive Care in Cancer Antiemesis Tool;[acyl-carrier-protein] S-malonyltransferase activity|MAT
Finding|Intellectual Product|Hospital Course|4700,4703|false|false|false|C0221158;C1151970;C1412111;C1417038;C3714902;C5780814;C5890859|ACAT1 gene;ACAT1 wt Allele;MAT1A gene;MAT1A wt Allele;Multifocal atrial tachycardia;Multinational Association of Supportive Care in Cancer Antiemesis Tool;[acyl-carrier-protein] S-malonyltransferase activity|MAT
Finding|Molecular Function|Hospital Course|4700,4703|false|false|false|C0221158;C1151970;C1412111;C1417038;C3714902;C5780814;C5890859|ACAT1 gene;ACAT1 wt Allele;MAT1A gene;MAT1A wt Allele;Multifocal atrial tachycardia;Multinational Association of Supportive Care in Cancer Antiemesis Tool;[acyl-carrier-protein] S-malonyltransferase activity|MAT
Finding|Mental Process|Hospital Course|4711,4718|false|false|false|C0542559|contextual factors|setting
Finding|Finding|Hospital Course|4722,4728|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|Hospital Course|4722,4728|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Event|Event|Hospital Course|4729,4740|false|false|false|||obstructive
Finding|Functional Concept|Hospital Course|4729,4740|false|false|false|C0549186|Obstructed|obstructive
Anatomy|Body Location or Region|Hospital Course|4742,4746|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4742,4746|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Hospital Course|4742,4746|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Hospital Course|4742,4746|false|false|false|C0740941|Lung Problem|lung
Disorder|Disease or Syndrome|Hospital Course|4742,4754|false|false|false|C0024115|Lung diseases|lung disease
Disorder|Disease or Syndrome|Hospital Course|4747,4754|false|false|false|C0012634|Disease|disease
Event|Event|Hospital Course|4747,4754|false|false|false|||disease
Finding|Intellectual Product|Hospital Course|4759,4766|false|true|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|Hospital Course|4759,4766|false|true|false|C1555457|Provision of recurring care for chronic illness|chronic
Drug|Organic Chemical|Hospital Course|4767,4779|false|false|false|C0039771|theophylline|theophylline
Drug|Pharmacologic Substance|Hospital Course|4767,4779|false|false|false|C0039771|theophylline|theophylline
Event|Event|Hospital Course|4767,4779|false|false|false|||theophylline
Procedure|Laboratory Procedure|Hospital Course|4767,4779|false|false|false|C0039773|Assay of theophylline|theophylline
Finding|Finding|Hospital Course|4767,4783|false|false|false|C0241361|theophylline use|theophylline use
Event|Event|Hospital Course|4780,4783|false|false|false|||use
Finding|Functional Concept|Hospital Course|4780,4783|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|Hospital Course|4780,4783|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Anatomy|Body System|Hospital Course|4785,4795|false|false|false|C0007226|Cardiovascular system|Cardiology
Event|Event|Hospital Course|4797,4808|false|false|false|||reccomended
Event|Event|Hospital Course|4817,4828|false|false|false|||discontinue
Drug|Organic Chemical|Hospital Course|4833,4845|false|false|false|C0039771|theophylline|theophylline
Drug|Pharmacologic Substance|Hospital Course|4833,4845|false|false|false|C0039771|theophylline|theophylline
Event|Event|Hospital Course|4833,4845|false|false|false|||theophylline
Procedure|Laboratory Procedure|Hospital Course|4833,4845|false|false|false|C0039773|Assay of theophylline|theophylline
Event|Event|Hospital Course|4850,4855|false|false|false|||spoke
Event|Event|Hospital Course|4884,4890|false|false|false|||agreed
Disorder|Disease or Syndrome|Hospital Course|4909,4913|false|true|false|C0339510|Vitelliform Macular Dystrophy|best
Finding|Gene or Genome|Hospital Course|4909,4913|false|true|false|C1826421;C5781213|BEST1 gene;BEST1 wt Allele|best
Event|Event|Hospital Course|4914,4920|false|false|false|||course
Event|Activity|Hospital Course|4925,4931|false|false|false|C3266814|Action|action
Event|Event|Hospital Course|4925,4931|false|false|false|||action
Finding|Functional Concept|Hospital Course|4925,4931|false|false|false|C0441472;C1552007|Clinical action|action
Finding|Idea or Concept|Hospital Course|4925,4931|false|false|false|C0441472;C1552007|Clinical action|action
Event|Event|Hospital Course|4949,4959|false|false|false|||discharged
Attribute|Clinical Attribute|Hospital Course|4965,4977|false|false|false|C3263700||instructions
Event|Event|Hospital Course|4965,4977|false|false|false|||instructions
Finding|Intellectual Product|Hospital Course|4965,4977|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|instructions
Event|Event|Hospital Course|4994,4997|false|false|false|||use
Finding|Functional Concept|Hospital Course|4994,4997|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|Hospital Course|4994,4997|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Functional Concept|Hospital Course|4994,5000|false|false|false|C1524063|Use of|use of
Drug|Organic Chemical|Hospital Course|5001,5013|false|false|false|C0039771|theophylline|theophylline
Drug|Pharmacologic Substance|Hospital Course|5001,5013|false|false|false|C0039771|theophylline|theophylline
Event|Event|Hospital Course|5001,5013|false|false|false|||theophylline
Procedure|Laboratory Procedure|Hospital Course|5001,5013|false|false|false|C0039773|Assay of theophylline|theophylline
Event|Event|Hospital Course|5018,5024|false|false|false|||follow
Event|Event|Hospital Course|5038,5051|false|false|false|||pulmonologist
Anatomy|Body System|Hospital Course|5056,5066|false|false|false|C0007226|Cardiovascular system|cardiology
Attribute|Clinical Attribute|Hospital Course|5071,5082|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|5071,5082|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|5071,5082|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|5071,5082|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|5071,5095|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|Hospital Course|5086,5095|false|false|false|||Admission
Procedure|Health Care Activity|Hospital Course|5086,5095|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Organic Chemical|Hospital Course|5097,5104|false|false|false|C0699142|Tylenol|Tylenol
Drug|Pharmacologic Substance|Hospital Course|5097,5104|false|false|false|C0699142|Tylenol|Tylenol
Finding|Gene or Genome|Hospital Course|5113,5116|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|5117,5121|false|false|false|C2598155||pain
Event|Event|Hospital Course|5117,5121|false|false|false|||pain
Finding|Functional Concept|Hospital Course|5117,5121|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|5117,5121|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|Hospital Course|5124,5133|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|Hospital Course|5124,5133|false|false|false|C0001927|albuterol|Albuterol
Drug|Organic Chemical|Hospital Course|5124,5141|false|false|false|C0543495|albuterol sulfate|Albuterol Sulfate
Drug|Pharmacologic Substance|Hospital Course|5124,5141|false|false|false|C0543495|albuterol sulfate|Albuterol Sulfate
Drug|Element, Ion, or Isotope|Hospital Course|5134,5141|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Inorganic Chemical|Hospital Course|5134,5141|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Pharmacologic Substance|Hospital Course|5134,5141|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Finding|Gene or Genome|Hospital Course|5156,5159|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|Hospital Course|5160,5163|false|false|false|||SOB
Finding|Sign or Symptom|Hospital Course|5160,5163|false|false|false|C0013404|Dyspnea|SOB
Drug|Organic Chemical|Hospital Course|5166,5177|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Hospital Course|5166,5177|false|false|false|C0082607|fluticasone|Fluticasone
Event|Event|Hospital Course|5166,5177|false|false|false|||Fluticasone
Drug|Biomedical or Dental Material|Hospital Course|5185,5190|false|false|false|C1154182|Spray Dosage Form|spray
Event|Activity|Hospital Course|5185,5190|false|false|false|C2003858|Spray (action)|spray
Event|Event|Hospital Course|5185,5190|false|false|false|||spray
Finding|Functional Concept|Hospital Course|5185,5190|false|false|false|C4521772|Spray (administration method)|spray
Drug|Biomedical or Dental Material|Hospital Course|5191,5201|false|false|false|C0038960;C1382107|Suspension substance;Suspensions|suspension
Drug|Substance|Hospital Course|5191,5201|false|false|false|C0038960;C1382107|Suspension substance;Suspensions|suspension
Event|Event|Hospital Course|5191,5201|false|false|false|||suspension
Finding|Functional Concept|Hospital Course|5191,5201|false|false|false|C1705537|Suspension (action)|suspension
Finding|Gene or Genome|Hospital Course|5211,5214|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|5215,5224|false|false|false|C1717415||allergies
Event|Event|Hospital Course|5215,5224|false|false|false|||allergies
Finding|Pathologic Function|Hospital Course|5215,5224|false|false|false|C0020517|Hypersensitivity|allergies
Drug|Biomedical or Dental Material|Hospital Course|5243,5246|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Organic Chemical|Hospital Course|5243,5246|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Pharmacologic Substance|Hospital Course|5243,5246|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Event|Event|Hospital Course|5243,5246|false|false|false|||INH
Finding|Functional Concept|Hospital Course|5243,5246|false|false|false|C0205535|Inhalation Route of Administration|INH
Disorder|Mental or Behavioral Dysfunction|Hospital Course|5247,5250|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5247,5250|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|5247,5250|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|5247,5250|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|5247,5250|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|5253,5257|false|false|false|C0020261|hydrochlorothiazide|HCTZ
Drug|Pharmacologic Substance|Hospital Course|5253,5257|false|false|false|C0020261|hydrochlorothiazide|HCTZ
Drug|Biomedical or Dental Material|Hospital Course|5293,5299|false|false|false|C0039225|Tablet Dosage Form|tablet
Event|Event|Hospital Course|5293,5299|false|false|false|||tablet
Drug|Organic Chemical|Hospital Course|5312,5322|false|false|false|C0028978|omeprazole|omeprazole
Drug|Pharmacologic Substance|Hospital Course|5312,5322|false|false|false|C0028978|omeprazole|omeprazole
Event|Event|Hospital Course|5312,5322|false|false|false|||omeprazole
Drug|Organic Chemical|Hospital Course|5338,5349|false|false|false|C0074554|simvastatin|simvastatin
Drug|Pharmacologic Substance|Hospital Course|5338,5349|false|false|false|C0074554|simvastatin|simvastatin
Event|Event|Hospital Course|5338,5349|false|false|false|||simvastatin
Drug|Organic Chemical|Hospital Course|5365,5377|false|false|false|C0039771|theophylline|theophylline
Drug|Pharmacologic Substance|Hospital Course|5365,5377|false|false|false|C0039771|theophylline|theophylline
Event|Event|Hospital Course|5365,5377|false|false|false|||theophylline
Procedure|Laboratory Procedure|Hospital Course|5365,5377|false|false|false|C0039773|Assay of theophylline|theophylline
Finding|Functional Concept|Hospital Course|5384,5393|false|false|false|C0443318|Sustained|sustained
Drug|Biomedical or Dental Material|Hospital Course|5384,5401|false|false|false|C1710261|Sustained Release Dosage Form|sustained release
Event|Event|Hospital Course|5394,5401|false|false|false|||release
Finding|Functional Concept|Hospital Course|5394,5401|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|release
Procedure|Health Care Activity|Hospital Course|5394,5401|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5394,5401|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|release
Event|Event|Hospital Course|5409,5412|false|false|false|||TID
Drug|Organic Chemical|Hospital Course|5415,5422|false|false|false|C0905678|Spiriva|spiriva
Drug|Pharmacologic Substance|Hospital Course|5415,5422|false|false|false|C0905678|Spiriva|spiriva
Event|Event|Hospital Course|5415,5422|false|false|false|||spiriva
Event|Event|Hospital Course|5426,5429|false|false|false|||mcg
Event|Event|Hospital Course|5433,5443|false|false|false|||inhalation
Finding|Functional Concept|Hospital Course|5433,5443|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Finding|Organism Function|Hospital Course|5433,5443|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5446,5449|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Enzyme|Hospital Course|5446,5449|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Organic Chemical|Hospital Course|5446,5449|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Pharmacologic Substance|Hospital Course|5446,5449|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Event|Event|Hospital Course|5446,5449|false|false|false|||ASA
Finding|Gene or Genome|Hospital Course|5446,5449|false|false|false|C1412553|ARSA gene|ASA
Drug|Biologically Active Substance|Hospital Course|5457,5464|false|true|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|Hospital Course|5457,5464|false|true|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|Hospital Course|5457,5464|false|true|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|Hospital Course|5457,5464|false|true|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|Hospital Course|5457,5464|false|true|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|Hospital Course|5457,5464|false|false|false|||Calcium
Finding|Physiologic Function|Hospital Course|5457,5464|false|true|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|Hospital Course|5457,5464|false|true|false|C0201925|Calcium measurement|Calcium
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5465,5468|false|false|false|C0262329|Short insular gyrus|sig
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5465,5468|false|false|false|C0034789|Receptors, Antigen, B-Cell|sig
Drug|Immunologic Factor|Hospital Course|5465,5468|false|false|false|C0034789|Receptors, Antigen, B-Cell|sig
Finding|Receptor|Hospital Course|5465,5468|false|false|false|C0034789|Receptors, Antigen, B-Cell|sig
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5469,5476|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Immunologic Factor|Hospital Course|5469,5476|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Pharmacologic Substance|Hospital Course|5469,5476|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Event|Event|Hospital Course|5469,5476|false|false|false|||unknown
Finding|Finding|Hospital Course|5469,5476|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Functional Concept|Hospital Course|5469,5476|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Idea or Concept|Hospital Course|5469,5476|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Intellectual Product|Hospital Course|5469,5476|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5479,5482|false|false|false|C0056632;C0459207;C2702357;C3488428|Cyclophosphamide/Dacarbazine/Vincristine;cod, unspecified preparation;codfish allergenic extract|Cod
Drug|Food|Hospital Course|5479,5482|false|false|false|C0056632;C0459207;C2702357;C3488428|Cyclophosphamide/Dacarbazine/Vincristine;cod, unspecified preparation;codfish allergenic extract|Cod
Drug|Immunologic Factor|Hospital Course|5479,5482|false|false|false|C0056632;C0459207;C2702357;C3488428|Cyclophosphamide/Dacarbazine/Vincristine;cod, unspecified preparation;codfish allergenic extract|Cod
Drug|Pharmacologic Substance|Hospital Course|5479,5482|false|false|false|C0056632;C0459207;C2702357;C3488428|Cyclophosphamide/Dacarbazine/Vincristine;cod, unspecified preparation;codfish allergenic extract|Cod
Event|Event|Hospital Course|5479,5482|false|false|false|||Cod
Finding|Finding|Hospital Course|5479,5482|false|false|false|C0007465;C0457523;C1420285;C5444130|Cancerization of Pancreatic Ducts;Cause of Death;Cemento-osseous dysplasia;SNRPB gene|Cod
Finding|Gene or Genome|Hospital Course|5479,5482|false|false|false|C0007465;C0457523;C1420285;C5444130|Cancerization of Pancreatic Ducts;Cause of Death;Cemento-osseous dysplasia;SNRPB gene|Cod
Finding|Pathologic Function|Hospital Course|5479,5482|false|false|false|C0007465;C0457523;C1420285;C5444130|Cancerization of Pancreatic Ducts;Cause of Death;Cemento-osseous dysplasia;SNRPB gene|Cod
Drug|Food|Hospital Course|5479,5492|false|false|false|C0009213|cod liver oil|Cod liver oil
Drug|Organic Chemical|Hospital Course|5479,5492|false|false|false|C0009213|cod liver oil|Cod liver oil
Drug|Pharmacologic Substance|Hospital Course|5479,5492|false|false|false|C0009213|cod liver oil|Cod liver oil
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5483,5488|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|Hospital Course|5483,5488|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|Hospital Course|5483,5488|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|Hospital Course|5483,5488|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|Hospital Course|5483,5488|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|Hospital Course|5483,5488|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|Hospital Course|5483,5488|false|false|false|||liver
Finding|Finding|Hospital Course|5483,5488|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|Hospital Course|5483,5488|false|false|false|C0872387|Procedures on liver|liver
Drug|Biomedical or Dental Material|Hospital Course|5489,5492|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|oil
Drug|Food|Hospital Course|5489,5492|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|oil
Drug|Organic Chemical|Hospital Course|5489,5492|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|oil
Drug|Pharmacologic Substance|Hospital Course|5489,5492|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|oil
Event|Event|Hospital Course|5489,5492|false|false|false|||oil
Event|Event|Hospital Course|5493,5496|false|false|false|||Sig
Finding|Gene or Genome|Hospital Course|5497,5500|false|false|false|C1823916|UNK gene|unk
Drug|Organic Chemical|Hospital Course|5503,5515|false|false|false|C0301532|Multivitamin preparation|Multivitamin
Drug|Pharmacologic Substance|Hospital Course|5503,5515|false|false|false|C0301532|Multivitamin preparation|Multivitamin
Drug|Vitamin|Hospital Course|5503,5515|false|false|false|C0301532|Multivitamin preparation|Multivitamin
Event|Event|Hospital Course|5521,5530|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|5521,5530|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|5521,5530|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|5521,5530|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|5521,5530|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|5521,5542|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|5531,5542|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|5531,5542|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|5531,5542|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|5531,5542|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Hospital Course|5547,5560|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Drug|Pharmacologic Substance|Hospital Course|5547,5560|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Event|Event|Hospital Course|5547,5560|false|false|false|||acetaminophen
Procedure|Laboratory Procedure|Hospital Course|5547,5560|false|false|false|C0373527|Acetaminophen measurement|acetaminophen
Drug|Biomedical or Dental Material|Hospital Course|5568,5574|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|5588,5594|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|5588,5594|false|false|false|||Tablet
Event|Event|Hospital Course|5598,5601|false|false|false|||Q4H
Event|Event|Hospital Course|5603,5608|false|false|false|||every
Finding|Intellectual Product|Hospital Course|5603,5608|false|false|false|C1720374|Every - dosing instruction fragment|every
Event|Event|Hospital Course|5622,5628|false|false|false|||needed
Attribute|Clinical Attribute|Hospital Course|5633,5637|false|false|false|C2598155||pain
Event|Event|Hospital Course|5633,5637|false|false|false|||pain
Finding|Functional Concept|Hospital Course|5633,5637|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|5633,5637|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|Hospital Course|5644,5653|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|Hospital Course|5644,5653|false|false|false|C0001927|albuterol|albuterol
Event|Event|Hospital Course|5644,5653|false|false|false|||albuterol
Drug|Organic Chemical|Hospital Course|5644,5661|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Pharmacologic Substance|Hospital Course|5644,5661|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Element, Ion, or Isotope|Hospital Course|5654,5661|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Inorganic Chemical|Hospital Course|5654,5661|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Pharmacologic Substance|Hospital Course|5654,5661|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Event|Event|Hospital Course|5654,5661|false|false|false|||sulfate
Disorder|Disease or Syndrome|Hospital Course|5679,5682|false|false|false|C0015458|Facial Hemiatrophy|HFA
Event|Event|Hospital Course|5679,5682|false|false|false|||HFA
Procedure|Diagnostic Procedure|Hospital Course|5679,5682|false|false|false|C0430649|High frequency audiometry|HFA
Drug|Biomedical or Dental Material|Hospital Course|5683,5690|false|false|false|C1112870|Aerosol Dose Form|Aerosol
Event|Event|Hospital Course|5691,5698|false|false|false|||Inhaler
Finding|Functional Concept|Hospital Course|5691,5698|false|false|false|C4319647|Inhaler (unit of presentation)|Inhaler
Finding|Functional Concept|Hospital Course|5718,5728|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Finding|Organism Function|Hospital Course|5718,5728|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Event|Event|Hospital Course|5752,5758|false|false|false|||needed
Event|Event|Hospital Course|5763,5766|false|false|false|||SOB
Finding|Sign or Symptom|Hospital Course|5763,5766|false|false|false|C0013404|Dyspnea|SOB
Event|Event|Hospital Course|5768,5774|false|false|false|||wheeze
Finding|Sign or Symptom|Hospital Course|5768,5774|false|false|false|C0043144|Wheezing|wheeze
Drug|Organic Chemical|Hospital Course|5781,5792|false|false|false|C0082607|fluticasone|fluticasone
Drug|Pharmacologic Substance|Hospital Course|5781,5792|false|false|false|C0082607|fluticasone|fluticasone
Event|Event|Hospital Course|5781,5792|false|false|false|||fluticasone
Drug|Pharmacologic Substance|Hospital Course|5781,5803|false|false|false|C0939232|fluticasone / salmeterol|fluticasone-salmeterol
Drug|Organic Chemical|Hospital Course|5793,5803|false|false|false|C0073992|salmeterol|salmeterol
Drug|Pharmacologic Substance|Hospital Course|5793,5803|false|false|false|C0073992|salmeterol|salmeterol
Event|Event|Hospital Course|5793,5803|false|false|false|||salmeterol
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5820,5824|false|false|false|C1556138|Disc - Body Part|Disk
Drug|Biomedical or Dental Material|Hospital Course|5820,5824|false|false|false|C0993608|Disk Drug Form|Disk
Finding|Functional Concept|Hospital Course|5830,5836|false|false|false|C1550509|Participation Type - device|Device
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5837,5840|false|false|false|C0262329|Short insular gyrus|Sig
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5837,5840|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Drug|Immunologic Factor|Hospital Course|5837,5840|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Finding|Receptor|Hospital Course|5837,5840|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5851,5855|false|false|false|C1556138|Disc - Body Part|Disk
Drug|Biomedical or Dental Material|Hospital Course|5851,5855|false|false|false|C0993608|Disk Drug Form|Disk
Finding|Functional Concept|Hospital Course|5861,5867|false|false|false|C1550509|Participation Type - device|Device
Event|Event|Hospital Course|5868,5878|false|false|false|||Inhalation
Finding|Functional Concept|Hospital Course|5868,5878|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Finding|Organism Function|Hospital Course|5868,5878|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Disorder|Mental or Behavioral Dysfunction|Hospital Course|5879,5882|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5879,5882|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|5879,5882|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|5879,5882|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|5879,5882|false|false|false|C1332410|BID gene|BID
Finding|Finding|Hospital Course|5884,5891|false|false|false|C4035627|2 times|2 times
Disorder|Disease or Syndrome|Hospital Course|5886,5891|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|Hospital Course|5894,5897|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|5894,5897|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|Hospital Course|5905,5916|false|false|false|C0082607|fluticasone|fluticasone
Drug|Pharmacologic Substance|Hospital Course|5905,5916|false|false|false|C0082607|fluticasone|fluticasone
Event|Event|Hospital Course|5905,5916|false|false|false|||fluticasone
Drug|Biomedical or Dental Material|Hospital Course|5934,5939|false|false|false|C1154182|Spray Dosage Form|Spray
Event|Activity|Hospital Course|5934,5939|false|false|false|C2003858|Spray (action)|Spray
Event|Event|Hospital Course|5934,5939|false|false|false|||Spray
Finding|Functional Concept|Hospital Course|5934,5939|false|false|false|C4521772|Spray (administration method)|Spray
Drug|Biomedical or Dental Material|Hospital Course|5934,5951|false|false|false|C1710170|SPRAY, SUSPENSION|Spray, Suspension
Drug|Biomedical or Dental Material|Hospital Course|5941,5951|false|false|false|C0038960;C1382107|Suspension substance;Suspensions|Suspension
Drug|Substance|Hospital Course|5941,5951|false|false|false|C0038960;C1382107|Suspension substance;Suspensions|Suspension
Event|Event|Hospital Course|5941,5951|false|false|false|||Suspension
Finding|Functional Concept|Hospital Course|5941,5951|false|false|false|C1705537|Suspension (action)|Suspension
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5963,5968|false|false|false|C0028429||Nasal
Drug|Biomedical or Dental Material|Hospital Course|5963,5968|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Organic Chemical|Hospital Course|5963,5968|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Pharmacologic Substance|Hospital Course|5963,5968|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Finding|Finding|Hospital Course|5963,5968|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Finding|Functional Concept|Hospital Course|5963,5968|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Finding|Intellectual Product|Hospital Course|5969,5973|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|Hospital Course|5969,5979|false|false|false|C3537736|Once A Day|once a day
Finding|Idea or Concept|Hospital Course|5976,5979|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|5976,5979|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Hospital Course|5983,5989|false|false|false|||needed
Finding|Finding|Hospital Course|5994,6001|false|false|false|C0020517;C0489531;C1314973;C1527304;C1547542;C3539909|Allergic Reaction;Allergic disposition;Allergy - Charge Type Reason;History of allergies;Hypersensitivity;Response to antigens|allergy
Finding|Idea or Concept|Hospital Course|5994,6001|false|false|false|C0020517;C0489531;C1314973;C1527304;C1547542;C3539909|Allergic Reaction;Allergic disposition;Allergy - Charge Type Reason;History of allergies;Hypersensitivity;Response to antigens|allergy
Finding|Pathologic Function|Hospital Course|5994,6001|false|false|false|C0020517;C0489531;C1314973;C1527304;C1547542;C3539909|Allergic Reaction;Allergic disposition;Allergy - Charge Type Reason;History of allergies;Hypersensitivity;Response to antigens|allergy
Finding|Physiologic Function|Hospital Course|5994,6001|false|false|false|C0020517;C0489531;C1314973;C1527304;C1547542;C3539909|Allergic Reaction;Allergic disposition;Allergy - Charge Type Reason;History of allergies;Hypersensitivity;Response to antigens|allergy
Event|Event|Hospital Course|6002,6010|false|false|false|||symptoms
Finding|Functional Concept|Hospital Course|6002,6010|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Hospital Course|6002,6010|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Drug|Organic Chemical|Hospital Course|6017,6036|false|false|false|C0020261|hydrochlorothiazide|hydrochlorothiazide
Drug|Pharmacologic Substance|Hospital Course|6017,6036|false|false|false|C0020261|hydrochlorothiazide|hydrochlorothiazide
Drug|Biomedical or Dental Material|Hospital Course|6043,6049|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|6063,6069|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Intellectual Product|Hospital Course|6073,6077|false|false|false|C1720092|Once - dosing instruction fragment|once
Finding|Idea or Concept|Hospital Course|6081,6084|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|6081,6084|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|Hospital Course|6091,6101|false|false|false|C0028978|omeprazole|omeprazole
Drug|Pharmacologic Substance|Hospital Course|6091,6101|false|false|false|C0028978|omeprazole|omeprazole
Event|Event|Hospital Course|6091,6101|false|false|false|||omeprazole
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6108,6115|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|6108,6115|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|6108,6115|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Attribute|Clinical Attribute|Hospital Course|6117,6124|false|false|false|C1545665|Views delayed|Delayed
Drug|Biomedical or Dental Material|Hospital Course|6117,6132|false|false|false|C1707664|Delayed Release Dosage Form|Delayed Release
Event|Event|Hospital Course|6125,6132|false|false|false|||Release
Finding|Functional Concept|Hospital Course|6125,6132|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|6125,6132|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6125,6132|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Event|Event|Hospital Course|6139,6142|false|false|false|||Sig
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6153,6160|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|6153,6160|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|6153,6160|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Attribute|Clinical Attribute|Hospital Course|6162,6169|false|false|false|C1545665|Views delayed|Delayed
Drug|Biomedical or Dental Material|Hospital Course|6162,6177|false|false|false|C1707664|Delayed Release Dosage Form|Delayed Release
Event|Event|Hospital Course|6170,6177|false|false|false|||Release
Finding|Functional Concept|Hospital Course|6170,6177|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|6170,6177|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6170,6177|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|Hospital Course|6207,6218|false|false|false|C0074554|simvastatin|simvastatin
Drug|Pharmacologic Substance|Hospital Course|6207,6218|false|false|false|C0074554|simvastatin|simvastatin
Event|Event|Hospital Course|6207,6218|false|false|false|||simvastatin
Drug|Biomedical or Dental Material|Hospital Course|6225,6231|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|6245,6251|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|6245,6251|false|false|false|||Tablet
Event|Event|Hospital Course|6252,6254|false|false|false|||PO
Finding|Intellectual Product|Hospital Course|6255,6259|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|Hospital Course|6255,6265|false|false|false|C3537736|Once A Day|once a day
Finding|Idea or Concept|Hospital Course|6262,6265|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|6262,6265|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|Hospital Course|6272,6282|false|false|false|C0213771|tiotropium|tiotropium
Drug|Pharmacologic Substance|Hospital Course|6272,6282|false|false|false|C0213771|tiotropium|tiotropium
Event|Event|Hospital Course|6272,6282|false|false|false|||tiotropium
Drug|Organic Chemical|Hospital Course|6272,6290|false|false|false|C1306772|tiotropium bromide|tiotropium bromide
Drug|Pharmacologic Substance|Hospital Course|6272,6290|false|false|false|C1306772|tiotropium bromide|tiotropium bromide
Drug|Inorganic Chemical|Hospital Course|6283,6290|false|false|false|C0006222|Bromides|bromide
Event|Event|Hospital Course|6283,6290|false|false|false|||bromide
Procedure|Laboratory Procedure|Hospital Course|6283,6290|false|false|false|C0202341|Bromides measurement|bromide
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6298,6305|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|6298,6305|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|6298,6305|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Finding|Functional Concept|Hospital Course|6309,6319|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Finding|Organism Function|Hospital Course|6309,6319|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Finding|Functional Concept|Hospital Course|6320,6326|false|false|false|C1550509|Participation Type - device|Device
Disorder|Congenital Abnormality|Hospital Course|6341,6344|false|false|false|C1855179|CATARACT, ANTERIOR POLAR|Cap
Drug|Biomedical or Dental Material|Hospital Course|6341,6344|false|false|false|C0006935|capsule (pharmacologic)|Cap
Event|Event|Hospital Course|6341,6344|false|false|false|||Cap
Finding|Gene or Genome|Hospital Course|6341,6344|false|false|false|C1416891;C1418551;C1419093;C1422073;C1422760;C2985259;C4522312|BRD4 gene;BRD4 wt Allele;CAP1 gene;HACD1 gene;LNPEP gene;SERPINB6 gene;SORBS1 gene|Cap
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6341,6344|false|false|false|C0278651;C0280547;C1879916|CAP Regimen;cisplatin/cyclophosphamide/doxorubicin protocol;cyclophosphamide/doxorubicin/prednisone protocol|Cap
Finding|Functional Concept|Hospital Course|6345,6355|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Finding|Organism Function|Hospital Course|6345,6355|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Event|Event|Hospital Course|6356,6361|false|false|false|||DAILY
Drug|Organic Chemical|Hospital Course|6376,6383|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|Hospital Course|6376,6383|false|false|false|C0004057|aspirin|aspirin
Event|Event|Hospital Course|6376,6383|false|false|false|||aspirin
Drug|Biomedical or Dental Material|Hospital Course|6390,6396|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|6397,6400|false|false|false|||Sig
Drug|Biomedical or Dental Material|Hospital Course|6410,6416|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|6410,6416|false|false|false|||Tablet
Event|Event|Hospital Course|6417,6419|false|false|false|||PO
Finding|Intellectual Product|Hospital Course|6420,6424|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|Hospital Course|6420,6430|false|false|false|C3537736|Once A Day|once a day
Finding|Idea or Concept|Hospital Course|6427,6430|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|6427,6430|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|Hospital Course|6438,6450|false|false|false|C0301532|Multivitamin preparation|multivitamin
Drug|Pharmacologic Substance|Hospital Course|6438,6450|false|false|false|C0301532|Multivitamin preparation|multivitamin
Drug|Vitamin|Hospital Course|6438,6450|false|false|false|C0301532|Multivitamin preparation|multivitamin
Drug|Pharmacologic Substance|Hospital Course|6438,6461|false|false|false|C0978787|Multivitamin tablet|multivitamin     Tablet
Drug|Biomedical or Dental Material|Hospital Course|6455,6461|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|6455,6461|false|false|false|||Tablet
Drug|Biomedical or Dental Material|Hospital Course|6475,6481|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|6475,6481|false|false|false|||Tablet
Drug|Organic Chemical|Hospital Course|6507,6516|false|false|false|C0012373|diltiazem|diltiazem
Drug|Pharmacologic Substance|Hospital Course|6507,6516|false|false|false|C0012373|diltiazem|diltiazem
Event|Event|Hospital Course|6507,6516|false|false|false|||diltiazem
Drug|Organic Chemical|Hospital Course|6507,6520|false|false|false|C0700579|diltiazem hydrochloride|diltiazem HCl
Drug|Pharmacologic Substance|Hospital Course|6507,6520|false|false|false|C0700579|diltiazem hydrochloride|diltiazem HCl
Disorder|Neoplastic Process|Hospital Course|6517,6520|false|false|false|C0023443|Hairy Cell Leukemia|HCl
Drug|Immunologic Factor|Hospital Course|6517,6520|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Inorganic Chemical|Hospital Course|6517,6520|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Pharmacologic Substance|Hospital Course|6517,6520|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Event|Event|Hospital Course|6517,6520|false|false|false|||HCl
Drug|Biomedical or Dental Material|Hospital Course|6528,6534|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|6545,6552|false|false|false|||Release
Finding|Functional Concept|Hospital Course|6545,6552|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|6545,6552|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6545,6552|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Biomedical or Dental Material|Hospital Course|6573,6579|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|6573,6579|false|false|false|||Tablet
Event|Event|Hospital Course|6590,6597|false|false|false|||Release
Finding|Functional Concept|Hospital Course|6590,6597|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|6590,6597|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6590,6597|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Finding|Intellectual Product|Hospital Course|6607,6611|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|Hospital Course|6607,6617|false|false|false|C3537736|Once A Day|once a day
Finding|Idea or Concept|Hospital Course|6614,6617|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|6614,6617|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Biomedical or Dental Material|Hospital Course|6628,6634|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|6645,6652|false|false|false|||Release
Finding|Functional Concept|Hospital Course|6645,6652|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|6645,6652|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6645,6652|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Finding|Idea or Concept|Hospital Course|6663,6670|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|6679,6692|false|false|false|C0017887|nitroglycerin|nitroglycerin
Drug|Pharmacologic Substance|Hospital Course|6679,6692|false|false|false|C0017887|nitroglycerin|nitroglycerin
Event|Event|Hospital Course|6679,6692|false|false|false|||nitroglycerin
Drug|Biomedical or Dental Material|Hospital Course|6700,6706|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|6700,6706|false|false|false|||Tablet
Drug|Biomedical or Dental Material|Hospital Course|6700,6718|false|false|false|C0991582|Sublingual Tablet|Tablet, Sublingual
Finding|Finding|Hospital Course|6708,6718|false|false|false|C0001565;C4521982|Sublingual (intended site);Sublingual Route of Administration|Sublingual
Finding|Functional Concept|Hospital Course|6708,6718|false|false|false|C0001565;C4521982|Sublingual (intended site);Sublingual Route of Administration|Sublingual
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6719,6722|false|false|false|C0262329|Short insular gyrus|Sig
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6719,6722|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Drug|Immunologic Factor|Hospital Course|6719,6722|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Finding|Receptor|Hospital Course|6719,6722|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Finding|Finding|Hospital Course|6734,6744|false|false|false|C0001565;C4521982|Sublingual (intended site);Sublingual Route of Administration|Sublingual
Finding|Functional Concept|Hospital Course|6734,6744|false|false|false|C0001565;C4521982|Sublingual (intended site);Sublingual Route of Administration|Sublingual
Event|Event|Hospital Course|6760,6766|false|false|false|||needed
Anatomy|Body Location or Region|Hospital Course|6771,6776|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Hospital Course|6771,6776|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Hospital Course|6771,6781|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|Hospital Course|6771,6781|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Hospital Course|6777,6781|false|false|false|C2598155||pain
Event|Event|Hospital Course|6777,6781|false|false|false|||pain
Finding|Functional Concept|Hospital Course|6777,6781|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|6777,6781|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|6783,6787|false|false|false|||take
Event|Event|Hospital Course|6796,6801|false|false|false|||onset
Anatomy|Body Location or Region|Hospital Course|6805,6810|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Hospital Course|6805,6810|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Hospital Course|6805,6815|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|Hospital Course|6805,6815|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Hospital Course|6811,6815|false|true|false|C2598155||pain
Event|Event|Hospital Course|6811,6815|false|false|false|||pain
Finding|Functional Concept|Hospital Course|6811,6815|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|6811,6815|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|6821,6827|false|false|false|||repeat
Finding|Functional Concept|Hospital Course|6821,6827|false|false|false|C0205341;C1705914|Repeat;Repeat Object|repeat
Event|Event|Hospital Course|6848,6857|false|false|false|||continued
Finding|Idea or Concept|Hospital Course|6848,6857|false|false|false|C0549178|Continuous|continued
Anatomy|Body Location or Region|Hospital Course|6859,6864|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Hospital Course|6859,6864|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Hospital Course|6859,6869|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|Hospital Course|6859,6869|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Hospital Course|6865,6869|false|false|false|C2598155||pain
Event|Event|Hospital Course|6865,6869|false|false|false|||pain
Finding|Functional Concept|Hospital Course|6865,6869|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|6865,6869|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Disorder|Disease or Syndrome|Hospital Course|6876,6879|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|Hospital Course|6876,6879|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|Hospital Course|6876,6879|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6876,6879|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|Hospital Course|6876,6879|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|Hospital Course|6876,6879|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|Hospital Course|6876,6879|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|Hospital Course|6876,6879|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|Hospital Course|6876,6879|false|false|false|||PCP
Finding|Gene or Genome|Hospital Course|6876,6879|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|Hospital Course|6876,6879|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Anatomy|Body Location or Region|Hospital Course|6883,6888|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Hospital Course|6883,6888|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Hospital Course|6883,6893|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|Hospital Course|6883,6893|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Hospital Course|6889,6893|false|false|false|C2598155||pain
Event|Event|Hospital Course|6889,6893|false|false|false|||pain
Finding|Functional Concept|Hospital Course|6889,6893|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|6889,6893|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|6894,6902|false|false|false|||persists
Finding|Idea or Concept|Hospital Course|6919,6926|false|false|false|C0807726|refill|Refills
Event|Event|Hospital Course|6934,6943|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|6934,6943|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|6934,6943|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|6934,6943|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|6934,6943|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|6934,6955|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|6934,6955|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|6944,6955|false|false|false|C2926604||Disposition
Event|Event|Hospital Course|6944,6955|false|false|false|||Disposition
Procedure|Health Care Activity|Hospital Course|6944,6955|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|Hospital Course|6957,6961|false|false|false|||Home
Finding|Idea or Concept|Hospital Course|6957,6961|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|6957,6961|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|6957,6961|false|false|false|C1553498|home health encounter|Home
Event|Event|Hospital Course|6964,6973|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|6964,6973|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|6964,6973|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|6964,6973|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|6964,6973|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|6964,6983|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|6974,6983|false|false|false|C0945731||Diagnosis
Event|Event|Hospital Course|6974,6983|false|false|false|||Diagnosis
Finding|Classification|Hospital Course|6974,6983|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|6974,6983|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|6974,6983|false|false|false|C0011900|Diagnosis|Diagnosis
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6985,6993|false|false|false|C0018787|Heart|Coronary
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6985,7000|false|false|false|C0205042|Coronary artery|Coronary Artery
Disorder|Disease or Syndrome|Hospital Course|6985,7008|false|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|Coronary Artery Disease
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6994,7000|false|false|false|C0003842;C0226004|Arterial system;Arteries|Artery
Anatomy|Body System|Hospital Course|6994,7000|false|false|false|C0003842;C0226004|Arterial system;Arteries|Artery
Disorder|Disease or Syndrome|Hospital Course|6994,7008|false|false|false|C0852949|Arteriopathic disease|Artery Disease
Disorder|Disease or Syndrome|Hospital Course|7001,7008|false|false|false|C0012634|Disease|Disease
Event|Event|Hospital Course|7001,7008|false|false|false|||Disease
Finding|Mental Process|Discharge Condition|7033,7039|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|7033,7046|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|7033,7046|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|7040,7046|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|7040,7046|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|7048,7053|false|false|false|||Clear
Finding|Idea or Concept|Discharge Condition|7048,7053|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|Discharge Condition|7058,7066|false|false|false|||coherent
Finding|Finding|Discharge Condition|7058,7066|false|false|false|C4068804|Coherent|coherent
Event|Event|Discharge Condition|7068,7073|false|false|false|||Level
Attribute|Clinical Attribute|Discharge Condition|7068,7090|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|7068,7090|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|Discharge Condition|7077,7090|false|false|false|||Consciousness
Finding|Finding|Discharge Condition|7077,7090|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|7077,7090|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|7092,7097|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|7092,7097|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|7092,7097|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|Discharge Condition|7092,7097|false|false|false|||Alert
Finding|Finding|Discharge Condition|7092,7097|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|7092,7097|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|7092,7097|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|Discharge Condition|7102,7113|false|false|false|||interactive
Finding|Functional Concept|Discharge Condition|7102,7113|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|7115,7123|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|7115,7123|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|7115,7123|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|7124,7130|false|false|false|C5889824||Status
Event|Event|Discharge Condition|7124,7130|false|false|false|||Status
Finding|Idea or Concept|Discharge Condition|7124,7130|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|7132,7142|false|false|false|||Ambulatory
Finding|Functional Concept|Discharge Condition|7132,7142|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|Discharge Condition|7132,7142|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|Discharge Condition|7132,7142|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|Discharge Condition|7132,7142|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|Discharge Condition|7145,7156|false|false|false|||Independent
Finding|Finding|Discharge Condition|7145,7156|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|Discharge Condition|7145,7156|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Event|Event|Discharge Instructions|7194,7202|false|false|false|||admitted
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|7235,7238|false|false|false|C0446516;C1140618;C1269078|Upper Extremity;Upper arm|arm
Disorder|Anatomical Abnormality|Discharge Instructions|7235,7238|false|false|false|C3495676|Anorectal Malformations|arm
Finding|Gene or Genome|Discharge Instructions|7235,7238|false|false|false|C1824218;C3715044|AKR1A1 wt Allele;ARMC9 gene|arm
Procedure|Diagnostic Procedure|Discharge Instructions|7235,7238|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Research Activity|Discharge Instructions|7235,7238|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|7235,7238|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Finding|Sign or Symptom|Discharge Instructions|7235,7243|false|false|false|C0239377|Arm Pain|arm pain
Attribute|Clinical Attribute|Discharge Instructions|7239,7243|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|7239,7243|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|7239,7243|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|7239,7243|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Discharge Instructions|7254,7263|false|false|false|||worrisome
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|7268,7273|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Discharge Instructions|7268,7273|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Discharge Instructions|7268,7273|false|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|Discharge Instructions|7268,7281|false|false|false|C0018799|Heart Diseases|heart disease
Disorder|Disease or Syndrome|Discharge Instructions|7274,7281|false|false|false|C0012634|Disease|disease
Event|Event|Discharge Instructions|7274,7281|false|false|false|||disease
Anatomy|Body Location or Region|Discharge Instructions|7292,7296|false|false|false|C4318744|Test - temporal region|test
Event|Event|Discharge Instructions|7292,7296|false|false|false|||test
Finding|Functional Concept|Discharge Instructions|7292,7296|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Finding|Intellectual Product|Discharge Instructions|7292,7296|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Lab|Laboratory or Test Result|Discharge Instructions|7292,7296|false|false|false|C0456984|Test Result|test
Procedure|Laboratory Procedure|Discharge Instructions|7292,7296|false|false|false|C0022885|Laboratory Procedures|test
Event|Event|Discharge Instructions|7297,7302|false|false|false|||found
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|7318,7326|false|false|false|C0018787|Heart|coronary
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|7318,7333|false|false|false|C0205042|Coronary artery|coronary artery
Disorder|Disease or Syndrome|Discharge Instructions|7318,7341|false|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|coronary artery disease
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|7327,7333|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|Discharge Instructions|7327,7333|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Disorder|Disease or Syndrome|Discharge Instructions|7327,7341|false|false|false|C0852949|Arteriopathic disease|artery disease
Disorder|Disease or Syndrome|Discharge Instructions|7334,7341|false|false|false|C0012634|Disease|disease
Event|Event|Discharge Instructions|7334,7341|false|false|false|||disease
Event|Event|Discharge Instructions|7352,7359|false|false|false|||started
Event|Event|Discharge Instructions|7365,7368|false|false|false|||new
Finding|Finding|Discharge Instructions|7365,7368|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Discharge Instructions|7365,7368|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Disorder|Disease or Syndrome|Discharge Instructions|7370,7375|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Discharge Instructions|7370,7375|false|false|false|||blood
Finding|Body Substance|Discharge Instructions|7370,7375|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Finding|Discharge Instructions|7370,7384|false|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|blood pressure
Finding|Organism Function|Discharge Instructions|7370,7384|false|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|blood pressure
Procedure|Health Care Activity|Discharge Instructions|7370,7384|false|false|false|C0005824|Blood pressure determination|blood pressure
Event|Event|Discharge Instructions|7376,7384|false|false|false|||pressure
Finding|Finding|Discharge Instructions|7376,7384|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|Discharge Instructions|7376,7384|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|Discharge Instructions|7376,7384|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|Discharge Instructions|7376,7384|false|false|false|C0033095||pressure
Drug|Pharmacologic Substance|Discharge Instructions|7385,7395|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Discharge Instructions|7385,7395|false|false|false|||medication
Finding|Intellectual Product|Discharge Instructions|7385,7395|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|Discharge Instructions|7400,7409|false|false|false|||tolerated
Finding|Finding|Discharge Instructions|7415,7419|false|false|false|C5575035|Well (answer to question)|well
Event|Event|Discharge Instructions|7433,7437|false|false|false|||keep
Event|Event|Discharge Instructions|7449,7455|false|false|false|||follow
Event|Activity|Discharge Instructions|7459,7471|false|false|false|C0003629|Appointments|appointments
Event|Event|Discharge Instructions|7459,7471|false|false|false|||appointments
Event|Event|Discharge Instructions|7475,7481|false|false|false|||listed
Event|Event|Discharge Instructions|7534,7541|false|false|false|||changes
Finding|Functional Concept|Discharge Instructions|7534,7541|false|false|false|C0392747|Changing|changes
Event|Event|Medications|7569,7576|false|false|false|||STARTED
Drug|Organic Chemical|Medications|7584,7593|false|false|false|C0012373|diltiazem|Diltiazem
Drug|Pharmacologic Substance|Medications|7584,7593|false|false|false|C0012373|diltiazem|Diltiazem
Finding|Intellectual Product|Medications|7600,7604|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|Medications|7600,7610|false|false|false|C3537736|Once A Day|once a day
Event|Event|Medications|7607,7610|false|false|false|||day
Finding|Idea or Concept|Medications|7607,7610|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Medications|7607,7610|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|Medications|7628,7640|false|false|false|C0039771|theophylline|theophylline
Drug|Pharmacologic Substance|Medications|7628,7640|false|false|false|C0039771|theophylline|theophylline
Event|Event|Medications|7628,7640|false|false|false|||theophylline
Procedure|Laboratory Procedure|Medications|7628,7640|false|false|false|C0039773|Assay of theophylline|theophylline
Drug|Organic Chemical|Medications|7654,7668|false|false|false|C0017887|nitroglycerin|nitroglycerine
Drug|Pharmacologic Substance|Medications|7654,7668|false|false|false|C0017887|nitroglycerin|nitroglycerine
Event|Event|Medications|7654,7668|false|false|false|||nitroglycerine
Event|Event|Medications|7672,7676|false|false|false|||take
Finding|Intellectual Product|Medications|7686,7701|false|false|false|C4054856|Have Chest Pain|have chest pain
Anatomy|Body Location or Region|Medications|7691,7696|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Medications|7691,7696|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Medications|7691,7701|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|Medications|7691,7701|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Medications|7697,7701|false|false|false|C2598155||pain
Event|Event|Medications|7697,7701|false|false|false|||pain
Finding|Functional Concept|Medications|7697,7701|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Medications|7697,7701|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Medications|7708,7712|false|false|false|||NEED
Drug|Inorganic Chemical|Medications|7716,7720|false|false|false|C0723457|Stop brand of fluoride|STOP
Drug|Pharmacologic Substance|Medications|7716,7720|false|false|false|C0723457|Stop brand of fluoride|STOP
Event|Activity|Medications|7716,7720|false|false|false|C1947925|Stop (Instruction Imperative)|STOP
Event|Event|Medications|7716,7720|false|false|false|||STOP
Finding|Gene or Genome|Medications|7716,7720|false|false|false|C1417022|MAP6 gene|STOP
Event|Event|Medications|7721,7728|false|false|false|||SMOKING
Finding|Individual Behavior|Medications|7721,7728|false|false|false|C0037369;C0453996;C1548578|Location characteristic ID - Smoking;Smoking;Tobacco smoking behavior|SMOKING
Finding|Intellectual Product|Medications|7721,7728|false|false|false|C0037369;C0453996;C1548578|Location characteristic ID - Smoking;Smoking;Tobacco smoking behavior|SMOKING
Event|Event|Medications|7730,7732|false|false|false|||IT
Event|Event|Medications|7738,7742|false|false|false|||KILL
Finding|Functional Concept|Medications|7738,7742|false|false|false|C0162388;C0681205;C1550555|Killing;Sacrifice;kill - ActRelationshipJoin|KILL
Finding|Idea or Concept|Medications|7738,7742|false|false|false|C0162388;C0681205;C1550555|Killing;Sacrifice;kill - ActRelationshipJoin|KILL
Finding|Social Behavior|Medications|7738,7742|false|false|false|C0162388;C0681205;C1550555|Killing;Sacrifice;kill - ActRelationshipJoin|KILL
Event|Event|Medications|7743,7746|false|false|false|||YOU
Procedure|Health Care Activity|Medications|7750,7758|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Medications|7759,7771|false|false|false|C3263700||Instructions
Event|Event|Medications|7759,7771|false|false|false|||Instructions
Finding|Intellectual Product|Medications|7759,7771|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

