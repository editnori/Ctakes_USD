 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|46,55|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|46,55|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|46,60|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|80,89|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|80,89|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|80,94|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|136,139|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|147,154|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|147,154|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|156,164|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|SIMPLE_SEGMENT|167,176|false|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|167,176|false|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|167,176|false|false|false|C0020517|Hypersensitivity|Allergies
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|179,189|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|179,189|false|false|false|C0065374|lisinopril|lisinopril
Event|Event|SIMPLE_SEGMENT|179,189|false|false|false|||lisinopril
Event|Event|SIMPLE_SEGMENT|192,201|false|false|false|||Attending
Finding|Functional Concept|SIMPLE_SEGMENT|192,201|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|SIMPLE_SEGMENT|210,225|false|false|false|C0277786|Chief complaint (finding)|Chief Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|216,225|false|false|false|C3864418||Complaint
Event|Event|SIMPLE_SEGMENT|216,225|false|false|false|||Complaint
Finding|Finding|SIMPLE_SEGMENT|216,225|false|false|false|C5441521|Complaint (finding)|Complaint
Finding|Sign or Symptom|SIMPLE_SEGMENT|227,236|false|true|false|C0004604|Back Pain|Back Pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|232,236|false|false|false|C2598155||Pain
Event|Event|SIMPLE_SEGMENT|232,236|false|false|false|||Pain
Finding|Functional Concept|SIMPLE_SEGMENT|232,236|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|232,236|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Classification|SIMPLE_SEGMENT|239,244|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|SIMPLE_SEGMENT|245,253|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|245,253|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|257,275|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|266,275|false|false|false|C0945766||Procedure
Event|Event|SIMPLE_SEGMENT|266,275|false|false|false|||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|266,275|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|266,275|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|266,275|false|false|false|C0184661|Interventional procedure|Procedure
Event|Event|SIMPLE_SEGMENT|285,292|true|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|285,292|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|285,292|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|285,292|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|285,295|true|false|false|C0262926|Medical History|History of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|285,311|true|false|false|C0488508||History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|285,311|true|false|false|C0262512|History of present illness (finding)|History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|296,303|true|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Idea or Concept|SIMPLE_SEGMENT|296,303|true|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Finding|SIMPLE_SEGMENT|296,311|true|false|false|C4264312|Present illness|Present Illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|304,311|true|false|false|C0221423|Illness (finding)|Illness
Finding|Body Substance|SIMPLE_SEGMENT|317,324|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|317,324|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|317,324|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|350,361|false|false|false|||significant
Finding|Idea or Concept|SIMPLE_SEGMENT|350,361|false|false|false|C0750502|Significant|significant
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|366,369|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|SIMPLE_SEGMENT|366,369|false|false|false|||HTN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|371,375|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Event|Event|SIMPLE_SEGMENT|371,375|false|false|false|||GERD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|378,381|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|378,381|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|378,381|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|378,381|false|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|378,381|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|378,381|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|378,381|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|378,381|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Event|Event|SIMPLE_SEGMENT|386,390|false|false|false|||CABG
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|386,390|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Event|Event|SIMPLE_SEGMENT|395,403|false|false|false|||stenting
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|395,403|false|false|false|C2348535|Stenting|stenting
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|405,409|false|false|false|C0011854|Diabetes Mellitus, Insulin-Dependent|IDDM
Event|Event|SIMPLE_SEGMENT|405,409|false|false|false|||IDDM
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|425,435|false|false|false|C0442874|Neuropathy|neuropathy
Event|Event|SIMPLE_SEGMENT|425,435|false|false|false|||neuropathy
Event|Event|SIMPLE_SEGMENT|441,449|false|false|false|||presents
Anatomy|Body Location or Region|SIMPLE_SEGMENT|457,462|false|false|false|C0230171|Flank (surface region)|flank
Finding|Sign or Symptom|SIMPLE_SEGMENT|457,467|false|false|false|C0016199|Flank Pain|flank pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|463,467|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|463,467|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|463,467|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|463,467|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Body Substance|SIMPLE_SEGMENT|475,482|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|475,482|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|475,482|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Attribute|Clinical Attribute|SIMPLE_SEGMENT|489,493|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|489,493|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|489,493|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|489,493|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|542,550|false|false|false|||worsened
Event|Event|SIMPLE_SEGMENT|579,587|false|false|false|||worsened
Event|Event|SIMPLE_SEGMENT|594,602|false|false|false|||coughing
Finding|Sign or Symptom|SIMPLE_SEGMENT|594,602|false|false|false|C0010200|Coughing|coughing
Event|Event|SIMPLE_SEGMENT|607,613|false|false|false|||moving
Finding|Organism Function|SIMPLE_SEGMENT|607,613|false|false|false|C0560560|Moving|moving
Event|Event|SIMPLE_SEGMENT|629,635|true|false|false|||denies
Event|Event|SIMPLE_SEGMENT|640,647|true|false|false|||dysuria
Finding|Sign or Symptom|SIMPLE_SEGMENT|640,647|true|false|false|C0013428|Dysuria|dysuria
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|649,656|true|false|false|C0042027|Urinary tract|urinary
Event|Event|SIMPLE_SEGMENT|658,667|true|false|false|||frequency
Finding|Intellectual Product|SIMPLE_SEGMENT|658,667|true|false|false|C3898838;C4321352|Frequency;How Often|frequency
Anatomy|Body Location or Region|SIMPLE_SEGMENT|669,678|true|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|SIMPLE_SEGMENT|669,683|true|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|679,683|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|679,683|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|679,683|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|679,683|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Anatomy|Body Location or Region|SIMPLE_SEGMENT|690,695|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|690,695|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|690,700|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|690,700|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|696,700|false|true|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|696,700|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|696,700|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|696,700|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|702,711|false|false|false|||shortness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|702,721|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|SIMPLE_SEGMENT|702,721|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|SIMPLE_SEGMENT|715,721|false|false|false|C0225386|Breath|breath
Event|Event|SIMPLE_SEGMENT|726,735|false|false|false|||dizziness
Finding|Sign or Symptom|SIMPLE_SEGMENT|726,735|false|false|false|C0012833;C0042571|Dizziness;Vertigo|dizziness
Event|Event|SIMPLE_SEGMENT|741,749|false|false|false|||endorses
Event|Event|SIMPLE_SEGMENT|752,760|false|false|false|||episodes
Event|Event|SIMPLE_SEGMENT|764,772|false|false|false|||diarrhea
Finding|Finding|SIMPLE_SEGMENT|764,772|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|SIMPLE_SEGMENT|764,772|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Idea or Concept|SIMPLE_SEGMENT|792,799|false|false|false|C1555582|Initial (abbreviation)|initial
Event|Event|SIMPLE_SEGMENT|800,806|false|false|false|||vitals
Event|Event|SIMPLE_SEGMENT|853,860|false|false|false|||trended
Event|Event|SIMPLE_SEGMENT|886,890|false|false|false|||Labs
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|886,890|false|false|false|C0587081|Laboratory test finding|Labs
Finding|Idea or Concept|SIMPLE_SEGMENT|896,907|false|false|false|C0750502|Significant|significant
Event|Event|SIMPLE_SEGMENT|908,911|false|false|false|||for
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|913,921|false|false|false|C4727483|BRAF Gene Rearrangement|positive
Event|Event|SIMPLE_SEGMENT|913,921|false|false|false|||positive
Finding|Classification|SIMPLE_SEGMENT|913,921|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|SIMPLE_SEGMENT|913,921|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Anatomy|Cell|SIMPLE_SEGMENT|926,929|false|false|false|C0023516|Leukocytes|WBC
Drug|Organic Chemical|SIMPLE_SEGMENT|935,942|false|false|false|C0022924;C0376261|Lactates;lactate|lactate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|935,942|false|false|false|C0022924;C0376261|Lactates;lactate|lactate
Event|Event|SIMPLE_SEGMENT|935,942|false|false|false|||lactate
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|935,942|false|false|false|C0202115|Lactic acid measurement|lactate
Anatomy|Cell|SIMPLE_SEGMENT|948,951|false|false|false|C0023516|Leukocytes|WBC
Event|Event|SIMPLE_SEGMENT|962,965|false|false|false|||PMN
Finding|Cell Function|SIMPLE_SEGMENT|962,965|false|false|false|C2612881;C2825189|Premarket Device Notification;piecemeal microautophagy of the nucleus|PMN
Finding|Intellectual Product|SIMPLE_SEGMENT|962,965|false|false|false|C2612881;C2825189|Premarket Device Notification;piecemeal microautophagy of the nucleus|PMN
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|968,971|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|SIMPLE_SEGMENT|968,971|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|968,971|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|SIMPLE_SEGMENT|968,971|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|SIMPLE_SEGMENT|968,971|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|SIMPLE_SEGMENT|968,971|false|false|false|||AST
Finding|Gene or Genome|SIMPLE_SEGMENT|968,971|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Disorder|Neoplastic Process|SIMPLE_SEGMENT|977,980|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|977,980|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|SIMPLE_SEGMENT|977,980|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|SIMPLE_SEGMENT|977,980|false|false|false|||ALT
Finding|Gene or Genome|SIMPLE_SEGMENT|977,980|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|SIMPLE_SEGMENT|977,980|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|SIMPLE_SEGMENT|977,980|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|977,980|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|985,988|false|false|false|C0023759|Lip structure|Lip
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|985,988|false|false|false|C0153932;C0264511|Benign neoplasm of the lip;Lymphoid interstitial pneumonia|Lip
Disorder|Neoplastic Process|SIMPLE_SEGMENT|985,988|false|false|false|C0153932;C0264511|Benign neoplasm of the lip;Lymphoid interstitial pneumonia|Lip
Finding|Gene or Genome|SIMPLE_SEGMENT|985,988|false|false|false|C1846919;C3889123|SMG1 gene;SMG1 wt Allele|Lip
Event|Event|SIMPLE_SEGMENT|1008,1012|false|false|false|||Chem
Finding|Functional Concept|SIMPLE_SEGMENT|1008,1012|false|false|false|C0079107|chemical aspects|Chem
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1008,1012|false|false|false|C0201682|Chemical procedure|Chem
Event|Event|SIMPLE_SEGMENT|1013,1022|false|false|false|||hemolyzed
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|1036,1044|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|SIMPLE_SEGMENT|1036,1044|false|false|false|||baseline
Finding|Idea or Concept|SIMPLE_SEGMENT|1036,1044|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Finding|Functional Concept|SIMPLE_SEGMENT|1057,1063|false|false|false|C0205341;C1705914|Repeat;Repeat Object|repeat
Event|Event|SIMPLE_SEGMENT|1071,1084|false|false|false|||Hyperglycemic
Event|Event|SIMPLE_SEGMENT|1101,1107|false|false|false|||repeat
Finding|Functional Concept|SIMPLE_SEGMENT|1101,1107|false|false|false|C0205341;C1705914|Repeat;Repeat Object|repeat
Event|Event|SIMPLE_SEGMENT|1109,1112|true|false|false|||CXR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1109,1112|true|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|SIMPLE_SEGMENT|1113,1119|true|false|false|||showed
Finding|Intellectual Product|SIMPLE_SEGMENT|1123,1128|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1129,1136|true|false|false|C1184743|bony process|process
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1129,1136|true|false|false|C1951340|Process Pharmacologic Substance|process
Event|Event|SIMPLE_SEGMENT|1129,1136|true|false|false|||process
Finding|Functional Concept|SIMPLE_SEGMENT|1129,1136|true|false|false|C4521054|Process (qualifier value)|process
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|1129,1136|true|false|false|C1522240|Process|process
Finding|Body Substance|SIMPLE_SEGMENT|1138,1145|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1138,1145|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1138,1145|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1167,1170|false|false|false|C0238052|Xanthomatosis, Cerebrotendinous|CTX
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1167,1170|false|false|false|C0010377;C0010583;C5574748|C-Terminal Telopeptide Type 1 Collagen, human;Crotoxin;cyclophosphamide|CTX
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1167,1170|false|false|false|C0010377;C0010583;C5574748|C-Terminal Telopeptide Type 1 Collagen, human;Crotoxin;cyclophosphamide|CTX
Drug|Enzyme|SIMPLE_SEGMENT|1167,1170|false|false|false|C0010377;C0010583;C5574748|C-Terminal Telopeptide Type 1 Collagen, human;Crotoxin;cyclophosphamide|CTX
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|1167,1170|false|false|false|C0010377;C0010583;C5574748|C-Terminal Telopeptide Type 1 Collagen, human;Crotoxin;cyclophosphamide|CTX
Drug|Organic Chemical|SIMPLE_SEGMENT|1167,1170|false|false|false|C0010377;C0010583;C5574748|C-Terminal Telopeptide Type 1 Collagen, human;Crotoxin;cyclophosphamide|CTX
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1167,1170|false|false|false|C0010377;C0010583;C5574748|C-Terminal Telopeptide Type 1 Collagen, human;Crotoxin;cyclophosphamide|CTX
Event|Event|SIMPLE_SEGMENT|1167,1170|false|false|false|||CTX
Finding|Gene or Genome|SIMPLE_SEGMENT|1167,1170|false|false|false|C1413864;C3539598|CYP27A1 gene;CYP27A1 wt Allele|CTX
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1181,1188|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|SIMPLE_SEGMENT|1181,1188|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1181,1188|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|SIMPLE_SEGMENT|1181,1188|false|false|false|||insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|1181,1188|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1181,1188|false|false|false|C0202098|Insulin measurement|insulin
Event|Event|SIMPLE_SEGMENT|1205,1213|false|false|false|||received
Event|Event|SIMPLE_SEGMENT|1218,1222|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|1218,1222|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|1218,1222|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|1218,1222|false|false|false|C1553498|home health encounter|home
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1236,1243|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|SIMPLE_SEGMENT|1236,1243|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1236,1243|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|SIMPLE_SEGMENT|1236,1243|false|false|false|||insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|1236,1243|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1236,1243|false|false|false|C0202098|Insulin measurement|insulin
Event|Event|SIMPLE_SEGMENT|1245,1248|false|false|false|||UCx
Event|Event|SIMPLE_SEGMENT|1264,1268|false|false|false|||sent
Drug|Antibiotic|SIMPLE_SEGMENT|1275,1286|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|SIMPLE_SEGMENT|1275,1286|false|false|false|||antibiotics
Event|Event|SIMPLE_SEGMENT|1315,1323|false|false|false|||transfer
Finding|Functional Concept|SIMPLE_SEGMENT|1315,1323|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|SIMPLE_SEGMENT|1315,1323|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|SIMPLE_SEGMENT|1315,1323|false|false|false|C4706767|Transfer (immobility management)|transfer
Finding|Finding|SIMPLE_SEGMENT|1365,1385|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Event|Event|SIMPLE_SEGMENT|1370,1377|false|false|false|||Medical
Finding|Functional Concept|SIMPLE_SEGMENT|1370,1377|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|1370,1377|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|1370,1377|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|1370,1377|false|false|false|C0199168|Medical service|Medical
Finding|Finding|SIMPLE_SEGMENT|1370,1385|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1378,1385|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1378,1385|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|1378,1385|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1387,1391|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1387,1391|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|SIMPLE_SEGMENT|1387,1391|false|false|false|||COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|1387,1391|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1394,1397|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1394,1397|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|1394,1397|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|1394,1397|false|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|1394,1397|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1394,1397|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|1394,1397|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1394,1397|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Event|Event|SIMPLE_SEGMENT|1402,1406|false|false|false|||CABG
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1402,1406|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Event|Event|SIMPLE_SEGMENT|1411,1419|false|false|false|||stenting
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1411,1419|false|false|false|C2348535|Stenting|stenting
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|1422,1432|false|false|false|C0011570;C0011581;C0344315;C0812393|Cancer patients and suicide and depression;Depressed mood;Depressive disorder;Mental Depression|Depression
Event|Event|SIMPLE_SEGMENT|1422,1432|false|false|false|||Depression
Finding|Functional Concept|SIMPLE_SEGMENT|1422,1432|false|false|false|C0460137;C1579931|Depression - motion|Depression
Finding|Sign or Symptom|SIMPLE_SEGMENT|1422,1432|false|false|false|C0460137;C1579931|Depression - motion|Depression
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1440,1444|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Event|Event|SIMPLE_SEGMENT|1440,1444|false|false|false|||GERD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1447,1450|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|SIMPLE_SEGMENT|1447,1450|false|false|false|||HTN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1453,1462|false|false|false|C0149931|Migraine Disorders|Migraines
Event|Event|SIMPLE_SEGMENT|1453,1462|false|false|false|||Migraines
Finding|Intellectual Product|SIMPLE_SEGMENT|1465,1472|false|false|false|C1547296|Chronic - Admission Level of Care Code|Chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|1465,1472|false|false|false|C1555457|Provision of recurring care for chronic illness|Chronic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1465,1486|false|false|false|C0748678|shoulder pain chronic|Chronic shoulder pain
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1473,1481|false|false|false|C0037004;C4299050|Shoulder;Upper extremity>Shoulder|shoulder
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1473,1481|false|false|false|C0221590;C0869975|Examination of shoulder(s);Procedures on Shoulder|shoulder
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1473,1481|false|false|false|C0221590;C0869975|Examination of shoulder(s);Procedures on Shoulder|shoulder
Finding|Sign or Symptom|SIMPLE_SEGMENT|1473,1486|false|false|false|C0037011|Shoulder Pain|shoulder pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1482,1486|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|1482,1486|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|1482,1486|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1482,1486|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|1490,1499|false|false|false|C0027415|Narcotics|narcotics
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1490,1499|false|false|false|C0027415|Narcotics|narcotics
Event|Event|SIMPLE_SEGMENT|1490,1499|false|false|false|||narcotics
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1502,1505|false|false|false|C0520679|Sleep Apnea, Obstructive|OSA
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1502,1505|false|false|false|C0764906|OSA protein, Drosophila|OSA
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1502,1505|false|false|false|C0764906|OSA protein, Drosophila|OSA
Event|Event|SIMPLE_SEGMENT|1502,1505|false|false|false|||OSA
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1508,1529|false|false|false|C0031117;C4721453|Peripheral Nervous System Diseases;Peripheral Neuropathy|Peripheral neuropathy
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1519,1529|false|false|false|C0442874|Neuropathy|neuropathy
Event|Event|SIMPLE_SEGMENT|1519,1529|false|false|false|||neuropathy
Finding|Sign or Symptom|SIMPLE_SEGMENT|1532,1540|false|false|false|C0085631;C3887611|Agitation;Restlessness|Restless
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1532,1544|false|false|false|C0035258|Restless Legs Syndrome|Restless leg
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1541,1544|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Finding|Functional Concept|SIMPLE_SEGMENT|1550,1556|false|false|false|C0728831|Social|Social
Finding|Finding|SIMPLE_SEGMENT|1550,1564|false|false|false|C0424945;C3714536|Social History;Social and personal history|Social History
Event|Event|SIMPLE_SEGMENT|1557,1564|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1557,1564|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1557,1564|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|1557,1564|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Classification|SIMPLE_SEGMENT|1570,1576|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|SIMPLE_SEGMENT|1570,1576|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|SIMPLE_SEGMENT|1570,1576|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|SIMPLE_SEGMENT|1570,1576|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Finding|SIMPLE_SEGMENT|1570,1584|false|false|false|C0241889|Family Medical History|Family History
Event|Event|SIMPLE_SEGMENT|1577,1584|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1577,1584|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1577,1584|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|1577,1584|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Event|Event|SIMPLE_SEGMENT|1586,1592|false|false|false|||Mother
Finding|Idea or Concept|SIMPLE_SEGMENT|1586,1592|false|false|false|C1546508|Relationship - Mother|Mother
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1593,1600|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|Unknown
Drug|Immunologic Factor|SIMPLE_SEGMENT|1593,1600|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|Unknown
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1593,1600|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|Unknown
Finding|Finding|SIMPLE_SEGMENT|1593,1600|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|Unknown
Finding|Functional Concept|SIMPLE_SEGMENT|1593,1600|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|Unknown
Finding|Idea or Concept|SIMPLE_SEGMENT|1593,1600|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|Unknown
Finding|Intellectual Product|SIMPLE_SEGMENT|1593,1600|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|Unknown
Drug|Organic Chemical|SIMPLE_SEGMENT|1601,1608|false|false|false|C0001962;C0001975|Alcohols;ethanol|ALCOHOL
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1601,1608|false|false|false|C0001962;C0001975|Alcohols;ethanol|ALCOHOL
Event|Event|SIMPLE_SEGMENT|1601,1608|false|false|false|||ALCOHOL
Finding|Intellectual Product|SIMPLE_SEGMENT|1601,1608|false|false|false|C1547288|Alcohol - Recreational Drug Use Code|ALCOHOL
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|1601,1614|false|false|false|C0085762|Alcohol abuse|ALCOHOL ABUSE
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|1609,1614|false|false|false|C0013146|Drug abuse|ABUSE
Event|Event|SIMPLE_SEGMENT|1609,1614|false|false|false|||ABUSE
Event|Event|SIMPLE_SEGMENT|1609,1614|false|false|false|C1546935|Abuse|ABUSE
Finding|Finding|SIMPLE_SEGMENT|1609,1614|false|false|false|C0562381|Victim of abuse (finding)|ABUSE
Event|Event|SIMPLE_SEGMENT|1622,1626|true|false|false|||ward
Event|Event|SIMPLE_SEGMENT|1630,1635|true|false|false|||state
Finding|Functional Concept|SIMPLE_SEGMENT|1630,1635|true|false|false|C1442792|State|state
Event|Event|SIMPLE_SEGMENT|1645,1649|true|false|false|||know
Event|Event|SIMPLE_SEGMENT|1656,1663|true|false|false|||details
Finding|Finding|SIMPLE_SEGMENT|1656,1673|true|false|false|C0557092|Details of family|details of family
Finding|Classification|SIMPLE_SEGMENT|1667,1673|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|1667,1673|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|1667,1673|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|1667,1673|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|1679,1685|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Idea or Concept|SIMPLE_SEGMENT|1679,1685|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1694,1701|false|false|false|C0019829|Hodgkin Disease|HODGKIN
Event|Event|SIMPLE_SEGMENT|1694,1701|false|false|false|||HODGKIN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1694,1711|false|false|false|C0019829|Hodgkin Disease|HODGKIN'S DISEASE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1704,1711|false|false|false|C0012634|Disease|DISEASE
Event|Event|SIMPLE_SEGMENT|1704,1711|false|false|false|||DISEASE
Event|Event|SIMPLE_SEGMENT|1720,1727|false|false|false|||records
Finding|Idea or Concept|SIMPLE_SEGMENT|1720,1727|false|false|false|C0034869;C1548330|Quantity limited request - Records;Records|records
Finding|Intellectual Product|SIMPLE_SEGMENT|1720,1727|false|false|false|C0034869;C1548330|Quantity limited request - Records;Records|records
Event|Event|SIMPLE_SEGMENT|1733,1741|false|false|false|||Physical
Finding|Finding|SIMPLE_SEGMENT|1733,1741|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|1733,1741|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|1733,1741|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|1733,1746|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|1733,1746|false|false|false|C0031809|Physical Examination|Physical Exam
Event|Event|SIMPLE_SEGMENT|1742,1746|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|1742,1746|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|1742,1746|false|false|false|C0582103|Medical Examination|Exam
Event|Event|SIMPLE_SEGMENT|1748,1757|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|1748,1757|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Finding|Finding|SIMPLE_SEGMENT|1758,1766|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|1758,1766|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|1758,1766|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|1758,1771|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|1758,1771|false|false|false|C0031809|Physical Examination|Physical Exam
Event|Event|SIMPLE_SEGMENT|1767,1771|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|1767,1771|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|1767,1771|false|false|false|C0582103|Medical Examination|Exam
Event|Event|SIMPLE_SEGMENT|1812,1819|false|false|false|||GENERAL
Finding|Classification|SIMPLE_SEGMENT|1812,1819|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|1812,1819|false|false|false|C3812897|General medical service|GENERAL
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1821,1824|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1821,1824|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1821,1824|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|1821,1824|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1821,1824|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|SIMPLE_SEGMENT|1821,1824|false|false|false|||NAD
Finding|Finding|SIMPLE_SEGMENT|1821,1824|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1827,1832|false|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1841,1848|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|SIMPLE_SEGMENT|1841,1848|false|false|false|C1314974|Cardiac attachment|CARDIAC
Event|Event|SIMPLE_SEGMENT|1850,1853|true|false|false|||RRR
Event|Event|SIMPLE_SEGMENT|1865,1872|true|false|false|||murmurs
Finding|Finding|SIMPLE_SEGMENT|1865,1872|true|false|false|C0018808|Heart murmur|murmurs
Event|Event|SIMPLE_SEGMENT|1874,1881|true|false|false|||gallops
Event|Event|SIMPLE_SEGMENT|1886,1890|true|false|false|||rubs
Finding|Finding|SIMPLE_SEGMENT|1886,1890|true|false|false|C0232267|Pericardial friction rub|rubs
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1893,1897|false|false|false|C0024109;C4037972|Chest>Lung;Lung|LUNG
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1893,1897|false|false|false|C0024109;C4037972|Chest>Lung;Lung|LUNG
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1893,1897|false|false|false|C0024115|Lung diseases|LUNG
Event|Event|SIMPLE_SEGMENT|1893,1897|false|false|false|||LUNG
Finding|Finding|SIMPLE_SEGMENT|1893,1897|false|false|false|C0740941|Lung Problem|LUNG
Drug|Organic Chemical|SIMPLE_SEGMENT|1899,1903|true|false|false|C0951233|cetrimonium bromide|CTAB
Event|Event|SIMPLE_SEGMENT|1899,1903|true|false|false|||CTAB
Event|Event|SIMPLE_SEGMENT|1908,1915|true|false|false|||wheezes
Finding|Sign or Symptom|SIMPLE_SEGMENT|1908,1915|true|false|false|C0043144|Wheezing|wheezes
Event|Event|SIMPLE_SEGMENT|1917,1922|true|false|false|||rales
Finding|Finding|SIMPLE_SEGMENT|1917,1922|true|false|false|C0034642;C0240859|Basilar Rales;Rales|rales
Event|Event|SIMPLE_SEGMENT|1924,1931|true|false|false|||rhonchi
Finding|Finding|SIMPLE_SEGMENT|1924,1931|true|false|false|C0035508|Rhonchi|rhonchi
Event|Event|SIMPLE_SEGMENT|1933,1942|true|false|false|||breathing
Event|Event|SIMPLE_SEGMENT|1964,1967|true|false|false|||use
Finding|Functional Concept|SIMPLE_SEGMENT|1964,1967|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|SIMPLE_SEGMENT|1964,1967|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Functional Concept|SIMPLE_SEGMENT|1964,1970|true|false|false|C1524063|Use of|use of
Finding|Finding|SIMPLE_SEGMENT|1964,1988|true|false|false|C1821466|Use of accessory muscles|use of accessory muscles
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|1971,1988|true|false|false|C0158784|Accessory skeletal muscle|accessory muscles
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1981,1988|true|false|false|C0026845;C1995013;C4083049|Muscle (organ);Muscle Tissue;Set of muscles|muscles
Anatomy|Tissue|SIMPLE_SEGMENT|1981,1988|true|false|false|C0026845;C1995013;C4083049|Muscle (organ);Muscle Tissue;Set of muscles|muscles
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1991,1998|true|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1991,1998|true|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Event|Event|SIMPLE_SEGMENT|1991,1998|true|false|false|||ABDOMEN
Finding|Finding|SIMPLE_SEGMENT|1991,1998|true|false|false|C0941288|Abdomen problem|ABDOMEN
Event|Event|SIMPLE_SEGMENT|2015,2017|true|false|false|||BS
Event|Event|SIMPLE_SEGMENT|2019,2028|true|false|false|||nontender
Event|Event|SIMPLE_SEGMENT|2051,2058|true|false|false|||rebound
Event|Event|SIMPLE_SEGMENT|2059,2067|true|false|false|||guarding
Finding|Finding|SIMPLE_SEGMENT|2059,2067|true|false|false|C0427198|Protective muscle spasm|guarding
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2070,2081|true|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Event|Event|SIMPLE_SEGMENT|2086,2094|true|false|false|||cyanosis
Finding|Sign or Symptom|SIMPLE_SEGMENT|2086,2094|true|false|false|C0010520|Cyanosis|cyanosis
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|2096,2104|true|false|false|C0149651|Clubbing|clubbing
Event|Event|SIMPLE_SEGMENT|2096,2104|true|false|false|||clubbing
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2108,2113|true|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|2108,2113|true|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|2108,2113|true|false|false|C0013604|Edema|edema
Event|Event|SIMPLE_SEGMENT|2115,2121|true|false|false|||moving
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2129,2140|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Event|Event|SIMPLE_SEGMENT|2129,2140|false|false|false|||extremities
Drug|Organic Chemical|SIMPLE_SEGMENT|2146,2153|false|false|false|C1995603|PURPOSE (pharmacologic preparation)|purpose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2146,2153|false|false|false|C1995603|PURPOSE (pharmacologic preparation)|purpose
Event|Event|SIMPLE_SEGMENT|2146,2153|false|false|false|||purpose
Finding|Functional Concept|SIMPLE_SEGMENT|2146,2153|false|false|false|C1285529|Purpose|purpose
Event|Event|SIMPLE_SEGMENT|2156,2160|false|false|false|||BACK
Event|Event|SIMPLE_SEGMENT|2165,2175|true|false|false|||tenderness
Finding|Mental Process|SIMPLE_SEGMENT|2165,2175|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|SIMPLE_SEGMENT|2165,2175|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Event|Event|SIMPLE_SEGMENT|2186,2195|true|false|false|||processes
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2200,2204|true|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|2200,2204|true|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|2200,2204|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|2200,2204|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Functional Concept|SIMPLE_SEGMENT|2209,2213|true|false|false|C1552822|Table Cell Horizontal Align - left|left
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2222,2225|false|false|false|C0001365;C0038454|Acute ill-defined cerebrovascular disease;Cerebrovascular accident|CVA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2222,2225|false|false|false|C5779650|Cyclophosphamide/Doxorubicin/Vincristine|CVA
Event|Event|SIMPLE_SEGMENT|2222,2225|false|false|false|||CVA
Finding|Sign or Symptom|SIMPLE_SEGMENT|2222,2236|false|false|false|C0235634|Renal angle tenderness|CVA tenderness
Event|Event|SIMPLE_SEGMENT|2226,2236|false|false|false|||tenderness
Finding|Mental Process|SIMPLE_SEGMENT|2226,2236|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|SIMPLE_SEGMENT|2226,2236|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Event|Event|SIMPLE_SEGMENT|2238,2248|false|false|false|||tenderness
Finding|Mental Process|SIMPLE_SEGMENT|2238,2248|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|SIMPLE_SEGMENT|2238,2248|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Event|Event|SIMPLE_SEGMENT|2252,2261|false|false|false|||palpation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2252,2261|false|false|false|C0030247|Palpation|palpation
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2278,2296|false|false|false|C0448353|Paraspinal Muscles|paraspinal muscles
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2289,2296|false|false|false|C0026845;C1995013;C4083049|Muscle (organ);Muscle Tissue;Set of muscles|muscles
Anatomy|Tissue|SIMPLE_SEGMENT|2289,2296|false|false|false|C0026845;C1995013;C4083049|Muscle (organ);Muscle Tissue;Set of muscles|muscles
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2320,2331|false|false|false|C0037925|Spinal Cord|spinal cord
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2320,2331|false|false|false|C0037928;C0153646;C0154034;C0496938|Benign neoplasm of spinal cord;Malignant neoplasm of spinal cord;Neoplasm of uncertain or unknown behavior of spinal cord;Spinal Cord Diseases|spinal cord
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2320,2331|false|false|false|C0037928;C0153646;C0154034;C0496938|Benign neoplasm of spinal cord;Malignant neoplasm of spinal cord;Neoplasm of uncertain or unknown behavior of spinal cord;Spinal Cord Diseases|spinal cord
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2327,2331|false|false|false|C1550235|Cord - Body Parts|cord
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2327,2331|false|false|false|C3489532|Cone-Rod Dystrophy 2|cord
Event|Event|SIMPLE_SEGMENT|2335,2344|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|2335,2344|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|2335,2344|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|2335,2344|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|2335,2344|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|2345,2353|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|2345,2353|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|2345,2353|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|2345,2358|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2345,2358|false|false|false|C0031809|Physical Examination|Physical Exam
Event|Event|SIMPLE_SEGMENT|2354,2358|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|2354,2358|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2354,2358|false|false|false|C0582103|Medical Examination|Exam
Event|Event|SIMPLE_SEGMENT|2392,2399|false|false|false|||General
Finding|Classification|SIMPLE_SEGMENT|2392,2399|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|SIMPLE_SEGMENT|2392,2399|false|false|false|C3812897|General medical service|General
Event|Event|SIMPLE_SEGMENT|2401,2406|false|false|false|||awake
Finding|Finding|SIMPLE_SEGMENT|2401,2406|false|false|false|C0234422|Awake (finding)|awake
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2408,2413|false|false|false|C5890168||alert
Drug|Organic Chemical|SIMPLE_SEGMENT|2408,2413|false|false|false|C0718338|Alert brand of caffeine|alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2408,2413|false|false|false|C0718338|Alert brand of caffeine|alert
Event|Event|SIMPLE_SEGMENT|2408,2413|false|false|false|||alert
Finding|Finding|SIMPLE_SEGMENT|2408,2413|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Functional Concept|SIMPLE_SEGMENT|2408,2413|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Intellectual Product|SIMPLE_SEGMENT|2408,2413|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2415,2418|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2415,2418|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2415,2418|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|2415,2418|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2415,2418|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|SIMPLE_SEGMENT|2415,2418|false|false|false|||NAD
Finding|Finding|SIMPLE_SEGMENT|2415,2418|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2419,2424|false|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2436,2439|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2436,2439|false|false|false|C0026987|Myelofibrosis|MMM
Event|Event|SIMPLE_SEGMENT|2436,2439|false|false|false|||MMM
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2455,2465|false|false|false|C0521367|Oropharyngeal|oropharynx
Event|Event|SIMPLE_SEGMENT|2470,2473|true|false|false|||RRR
Event|Event|SIMPLE_SEGMENT|2495,2498|true|false|false|||JVD
Finding|Finding|SIMPLE_SEGMENT|2495,2498|true|false|false|C0425687|Jugular venous engorgement|JVD
Event|Event|SIMPLE_SEGMENT|2499,2502|true|false|false|||HJR
Finding|Finding|SIMPLE_SEGMENT|2499,2502|true|false|false|C0239949|Hepatojugular reflux|HJR
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2505,2510|false|false|false|C0024109|Lung|Lungs
Drug|Organic Chemical|SIMPLE_SEGMENT|2512,2516|true|false|false|C0951233|cetrimonium bromide|CTAB
Event|Event|SIMPLE_SEGMENT|2512,2516|true|false|false|||CTAB
Event|Event|SIMPLE_SEGMENT|2524,2525|true|false|false|||r
Event|Event|SIMPLE_SEGMENT|2527,2531|true|false|false|||good
Finding|Idea or Concept|SIMPLE_SEGMENT|2527,2531|true|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Event|Event|SIMPLE_SEGMENT|2532,2540|false|false|false|||movement
Finding|Organism Function|SIMPLE_SEGMENT|2532,2540|false|false|false|C0026649|Movement|movement
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2555,2562|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2555,2562|false|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Event|Event|SIMPLE_SEGMENT|2555,2562|false|false|false|||Abdomen
Finding|Finding|SIMPLE_SEGMENT|2555,2562|false|false|false|C0941288|Abdomen problem|Abdomen
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2564,2569|false|false|false|C0028754|Obesity|obese
Event|Event|SIMPLE_SEGMENT|2564,2569|false|false|false|||obese
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2571,2575|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|SIMPLE_SEGMENT|2594,2596|false|false|false|||BS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2603,2606|false|false|false|C0034155;C1268935|Congenital Thrombotic Thrombocytopenic Purpura;Purpura, Thrombotic Thrombocytopenic|ttp
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2603,2606|false|false|false|C1506603;C4723973|ZFP36 protein, human;thiamine triphosphorate|ttp
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2603,2606|false|false|false|C1506603;C4723973|ZFP36 protein, human;thiamine triphosphorate|ttp
Drug|Organic Chemical|SIMPLE_SEGMENT|2603,2606|false|false|false|C1506603;C4723973|ZFP36 protein, human;thiamine triphosphorate|ttp
Drug|Vitamin|SIMPLE_SEGMENT|2603,2606|false|false|false|C1506603;C4723973|ZFP36 protein, human;thiamine triphosphorate|ttp
Event|Event|SIMPLE_SEGMENT|2603,2606|false|false|false|||ttp
Finding|Gene or Genome|SIMPLE_SEGMENT|2603,2606|false|false|false|C1413036;C1421571;C3539814|ADAMTS13 gene;ZFP36 gene;ZFP36 wt Allele|ttp
Finding|Functional Concept|SIMPLE_SEGMENT|2613,2618|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2619,2636|false|false|false|C5239513|Paraspinal Region|paraspinal region
Drug|Amino Acid Sequence|SIMPLE_SEGMENT|2630,2636|false|false|false|C1514562|Protein Domain|region
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2642,2648|false|false|false|C0036033;C0036037;C3669209;C4299073|Bone structure of sacrum;Pelvis>Sacrum;Sacral Region;Structure of sacrum|sacrum
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2642,2648|false|false|false|C0036033;C0036037;C3669209;C4299073|Bone structure of sacrum;Pelvis>Sacrum;Sacral Region;Structure of sacrum|sacrum
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2652,2660|false|false|false|C0037004;C4299050|Shoulder;Upper extremity>Shoulder|shoulder
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2652,2660|false|false|false|C0221590;C0869975|Examination of shoulder(s);Procedures on Shoulder|shoulder
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2652,2660|false|false|false|C0221590;C0869975|Examination of shoulder(s);Procedures on Shoulder|shoulder
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2665,2668|false|false|false|C0001365;C0038454|Acute ill-defined cerebrovascular disease;Cerebrovascular accident|CVA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2665,2668|false|false|false|C5779650|Cyclophosphamide/Doxorubicin/Vincristine|CVA
Event|Event|SIMPLE_SEGMENT|2665,2668|false|false|false|||CVA
Finding|Sign or Symptom|SIMPLE_SEGMENT|2665,2679|false|false|false|C0235634|Renal angle tenderness|CVA tenderness
Event|Event|SIMPLE_SEGMENT|2669,2679|false|false|false|||tenderness
Finding|Mental Process|SIMPLE_SEGMENT|2669,2679|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|SIMPLE_SEGMENT|2669,2679|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|2681,2684|false|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Event|Event|SIMPLE_SEGMENT|2681,2684|false|false|false|||Ext
Finding|Gene or Genome|SIMPLE_SEGMENT|2681,2684|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Event|Event|SIMPLE_SEGMENT|2694,2697|false|false|false|||WWP
Event|Event|SIMPLE_SEGMENT|2722,2728|false|false|false|||moving
Event|Event|SIMPLE_SEGMENT|2733,2739|false|false|false|||extrem
Drug|Organic Chemical|SIMPLE_SEGMENT|2745,2752|true|false|false|C1995603|PURPOSE (pharmacologic preparation)|purpose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2745,2752|true|false|false|C1995603|PURPOSE (pharmacologic preparation)|purpose
Event|Event|SIMPLE_SEGMENT|2745,2752|true|false|false|||purpose
Finding|Functional Concept|SIMPLE_SEGMENT|2745,2752|true|false|false|C1285529|Purpose|purpose
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2754,2760|true|false|false|C0015450|Face|facial
Event|Event|SIMPLE_SEGMENT|2761,2770|true|false|false|||movements
Finding|Organism Function|SIMPLE_SEGMENT|2761,2770|true|false|false|C0026649|Movement|movements
Event|Event|SIMPLE_SEGMENT|2772,2781|true|false|false|||symmetric
Finding|Conceptual Entity|SIMPLE_SEGMENT|2772,2781|true|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Finding|SIMPLE_SEGMENT|2772,2781|true|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Event|Event|SIMPLE_SEGMENT|2792,2800|true|false|false|||deficits
Anatomy|Body System|SIMPLE_SEGMENT|2802,2806|false|false|false|C1123023;C4520765|Skin;Skin, Human|Skin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2802,2806|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|Skin
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2802,2806|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|Skin
Finding|Body Substance|SIMPLE_SEGMENT|2802,2806|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|Skin
Finding|Intellectual Product|SIMPLE_SEGMENT|2802,2806|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|Skin
Event|Event|SIMPLE_SEGMENT|2811,2817|true|false|false|||rashes
Finding|Sign or Symptom|SIMPLE_SEGMENT|2811,2817|true|false|false|C0015230;C5779628|Exanthema;Skin rash|rashes
Event|Event|SIMPLE_SEGMENT|2819,2826|true|false|false|||lesions
Finding|Finding|SIMPLE_SEGMENT|2819,2826|true|false|false|C0221198|Lesion|lesions
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|2828,2840|true|false|false|C0015256|Excoriation|excoriations
Event|Event|SIMPLE_SEGMENT|2828,2840|true|false|false|||excoriations
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2863,2869|false|false|false|C1644645||CT ABD
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2866,2869|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|ABD
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|2866,2869|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|ABD
Event|Event|SIMPLE_SEGMENT|2866,2869|false|false|false|||ABD
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2870,2876|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|PELVIS
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|2870,2876|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|PELVIS
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2870,2876|false|false|false|C0153663|Malignant neoplasm of pelvis|PELVIS
Finding|Finding|SIMPLE_SEGMENT|2870,2876|false|false|false|C0812455|Pelvis problem|PELVIS
Event|Event|SIMPLE_SEGMENT|2894,2901|false|false|false|||imaging
Finding|Finding|SIMPLE_SEGMENT|2894,2901|false|false|false|C0740845|Imaging problem|imaging
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2894,2901|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|imaging
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2909,2916|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|abdomen
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2909,2916|false|false|false|C0153662|Malignant neoplasm of abdomen|abdomen
Finding|Finding|SIMPLE_SEGMENT|2909,2916|false|false|false|C0941288|Abdomen problem|abdomen
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2909,2920|false|false|false|C0000726|Abdomen|abdomen and
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2909,2927|false|false|false|C1508499|Abdominopelvic structure|abdomen and pelvis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2921,2927|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|2921,2927|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2921,2927|false|false|false|C0153663|Malignant neoplasm of pelvis|pelvis
Finding|Finding|SIMPLE_SEGMENT|2921,2927|false|false|false|C0812455|Pelvis problem|pelvis
Event|Event|SIMPLE_SEGMENT|2928,2940|false|false|false|||demonstrates
Event|Event|SIMPLE_SEGMENT|2969,2977|false|false|false|||calculus
Finding|Body Substance|SIMPLE_SEGMENT|2969,2977|false|false|false|C0006736|Calculi|calculus
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2969,2977|false|false|false|C3668917|Calculus (lab procedure)|calculus
Finding|Functional Concept|SIMPLE_SEGMENT|2985,2990|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|2991,3001|false|false|false|C0424290|Compulsive hoarding|collecting
Event|Event|SIMPLE_SEGMENT|2991,3001|false|false|false|||collecting
Finding|Functional Concept|SIMPLE_SEGMENT|2991,3001|false|false|false|C1516698|Collection (action)|collecting
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3002,3008|false|false|false|C5671121|System (basic dose form)|system
Event|Event|SIMPLE_SEGMENT|3002,3008|false|false|false|||system
Finding|Functional Concept|SIMPLE_SEGMENT|3002,3008|false|false|false|C0449913;C5441654|System;System, LOINC Axis 4|system
Finding|Functional Concept|SIMPLE_SEGMENT|3031,3035|true|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3036,3041|true|false|false|C0022646|Kidney|renal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3036,3041|true|false|false|C0042075|Urologic Diseases|renal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3036,3050|true|false|false|C0392525|Nephrolithiasis|renal calculus
Finding|Body Substance|SIMPLE_SEGMENT|3036,3050|true|false|false|C0022650|Kidney Calculi|renal calculus
Event|Event|SIMPLE_SEGMENT|3042,3050|true|false|false|||calculus
Finding|Body Substance|SIMPLE_SEGMENT|3042,3050|true|false|false|C0006736|Calculi|calculus
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3042,3050|true|false|false|C3668917|Calculus (lab procedure)|calculus
Event|Event|SIMPLE_SEGMENT|3064,3072|true|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|3064,3072|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|3064,3075|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3077,3085|true|false|false|C0041951|Ureter|ureteral
Finding|Functional Concept|SIMPLE_SEGMENT|3077,3085|true|false|false|C1522613|Ureteral Route of Administration|ureteral
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3089,3096|true|false|false|C0042027|Urinary tract|urinary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3089,3104|true|false|false|C0005682;C4037992|Abdomen+Pelvis>Urinary bladder;Urinary Bladder|urinary bladder
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3089,3113|true|false|false|C0005683|Urinary bladder stone (disorder)|urinary bladder calculus
Finding|Body Substance|SIMPLE_SEGMENT|3089,3113|true|false|false|C2712342|Bladder stone (substance)|urinary bladder calculus
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3097,3104|true|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3097,3104|true|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3097,3104|true|false|false|C0872388|Procedures on bladder|bladder
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3097,3113|true|false|false|C0005683|Urinary bladder stone (disorder)|bladder calculus
Finding|Body Substance|SIMPLE_SEGMENT|3097,3113|true|false|false|C2712342|Bladder stone (substance)|bladder calculus
Event|Event|SIMPLE_SEGMENT|3105,3113|false|false|false|||calculus
Finding|Body Substance|SIMPLE_SEGMENT|3105,3113|false|false|false|C0006736|Calculi|calculus
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3105,3113|false|false|false|C3668917|Calculus (lab procedure)|calculus
Finding|Conceptual Entity|SIMPLE_SEGMENT|3124,3133|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Finding|SIMPLE_SEGMENT|3124,3133|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3134,3139|false|false|false|C0022646|Kidney|renal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3134,3139|false|false|false|C0042075|Urologic Diseases|renal
Event|Activity|SIMPLE_SEGMENT|3141,3152|false|false|false|C2349975|Enhance (action)|enhancement
Event|Event|SIMPLE_SEGMENT|3141,3152|false|false|false|||enhancement
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3141,3152|false|false|false|C1627358|Refractive surgery enhancement|enhancement
Event|Event|SIMPLE_SEGMENT|3157,3166|false|false|false|||excretion
Finding|Body Substance|SIMPLE_SEGMENT|3157,3166|false|false|false|C0221102;C0504085|Body Excretions;Excretory function|excretion
Finding|Physiologic Function|SIMPLE_SEGMENT|3157,3166|false|false|false|C0221102;C0504085|Body Excretions;Excretory function|excretion
Finding|Functional Concept|SIMPLE_SEGMENT|3170,3181|false|false|false|C1522726|Intravenous Route of Administration|intravenous
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|3170,3190|false|false|false|C4072741|IV contrast|intravenous contrast
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|3182,3190|false|false|false|C0009924|Contrast Media|contrast
Event|Event|SIMPLE_SEGMENT|3182,3190|false|false|false|||contrast
Event|Event|SIMPLE_SEGMENT|3224,3235|false|false|false|||hypodensity
Finding|Functional Concept|SIMPLE_SEGMENT|3243,3247|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Drug|Amino Acid Sequence|SIMPLE_SEGMENT|3259,3265|false|false|false|C1514562|Protein Domain|region
Event|Event|SIMPLE_SEGMENT|3282,3287|false|false|false|||small
Event|Event|SIMPLE_SEGMENT|3302,3314|false|false|false|||characterize
Finding|Finding|SIMPLE_SEGMENT|3319,3325|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|3319,3325|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|SIMPLE_SEGMENT|3327,3337|false|false|false|||represents
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3338,3343|false|false|false|C0022646|Kidney|renal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3338,3343|false|false|false|C0042075|Urologic Diseases|renal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3338,3348|false|false|false|C0268800;C3887499|Renal cyst;Simple renal cyst|renal cyst
Finding|Finding|SIMPLE_SEGMENT|3338,3348|false|false|false|C2173677||renal cyst
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|3344,3348|false|false|false|C0010709|Cyst|cyst
Event|Event|SIMPLE_SEGMENT|3344,3348|false|false|false|||cyst
Finding|Body Substance|SIMPLE_SEGMENT|3344,3348|false|false|false|C1546594;C1550626|SpecimenType - Cyst|cyst
Finding|Intellectual Product|SIMPLE_SEGMENT|3344,3348|false|false|false|C1546594;C1550626|SpecimenType - Cyst|cyst
Event|Event|SIMPLE_SEGMENT|3362,3370|true|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|3362,3370|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|3362,3373|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|3374,3384|true|false|false|C0424290|Compulsive hoarding|collecting
Event|Event|SIMPLE_SEGMENT|3374,3384|true|false|false|||collecting
Finding|Functional Concept|SIMPLE_SEGMENT|3374,3384|true|false|false|C1516698|Collection (action)|collecting
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3385,3391|true|false|false|C5671121|System (basic dose form)|system
Event|Event|SIMPLE_SEGMENT|3385,3391|true|false|false|||system
Finding|Functional Concept|SIMPLE_SEGMENT|3385,3391|true|false|false|C0449913;C5441654|System;System, LOINC Axis 4|system
Finding|Functional Concept|SIMPLE_SEGMENT|3393,3407|true|false|false|C0332555|Filling defect|filling defect
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3401,3407|true|false|false|C1861101|THYROID HORMONE PLASMA MEMBRANE TRANSPORT DEFECT|defect
Event|Event|SIMPLE_SEGMENT|3401,3407|true|false|false|||defect
Finding|Functional Concept|SIMPLE_SEGMENT|3401,3407|true|false|false|C1457869|Defect|defect
Event|Event|SIMPLE_SEGMENT|3419,3427|false|false|false|||segments
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3442,3448|true|false|false|C4522154|Distal Resection Margin|distal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3449,3456|true|false|false|C0041951|Ureter|ureters
Finding|Finding|SIMPLE_SEGMENT|3466,3470|true|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|3471,3480|true|false|false|||opacified
Finding|Finding|SIMPLE_SEGMENT|3482,3490|true|false|false|C0332149|Possible|possibly
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3491,3500|true|true|false|C0027627|Neoplasm Metastasis|secondary
Event|Event|SIMPLE_SEGMENT|3491,3500|true|false|false|||secondary
Finding|Functional Concept|SIMPLE_SEGMENT|3491,3500|true|true|false|C1522484|metastatic qualifier|secondary
Event|Event|SIMPLE_SEGMENT|3504,3515|true|false|false|||peristalsis
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|3504,3515|true|false|false|C0031133|Peristalsis|peristalsis
Event|Event|SIMPLE_SEGMENT|3538,3546|true|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|3538,3546|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|3538,3549|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Finding|Functional Concept|SIMPLE_SEGMENT|3550,3562|true|false|false|C0333348|Inflammatory|inflammatory
Event|Event|SIMPLE_SEGMENT|3563,3569|true|false|false|||change
Finding|Functional Concept|SIMPLE_SEGMENT|3563,3569|true|false|false|C0392747|Changing|change
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3563,3569|true|false|false|C4319952|Change - procedure|change
Event|Event|SIMPLE_SEGMENT|3573,3577|true|false|false|||mass
Finding|Finding|SIMPLE_SEGMENT|3573,3577|true|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|SIMPLE_SEGMENT|3573,3577|true|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|SIMPLE_SEGMENT|3573,3577|true|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3589,3596|false|false|false|C0041951|Ureter|ureters
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3602,3609|false|false|false|C0001625|Adrenal Glands|adrenal
Finding|Finding|SIMPLE_SEGMENT|3602,3609|false|false|false|C0521428|Adrenal|adrenal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3602,3616|false|false|false|C0001625|Adrenal Glands|adrenal glands
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3610,3616|false|false|false|C1285092|Gland|glands
Event|Event|SIMPLE_SEGMENT|3621,3633|false|false|false|||unremarkable
Finding|Finding|SIMPLE_SEGMENT|3639,3642|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|Low
Finding|Intellectual Product|SIMPLE_SEGMENT|3639,3642|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|Low
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3643,3650|false|false|false|C0205054|Hepatic|hepatic
Event|Activity|SIMPLE_SEGMENT|3651,3662|false|false|false|C0599946|Attenuation|attenuation
Event|Event|SIMPLE_SEGMENT|3651,3662|false|false|false|||attenuation
Event|Event|SIMPLE_SEGMENT|3678,3685|false|false|false|||imaging
Finding|Finding|SIMPLE_SEGMENT|3678,3685|false|false|false|C0740845|Imaging problem|imaging
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3678,3685|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|imaging
Event|Event|SIMPLE_SEGMENT|3689,3699|false|false|false|||consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|3689,3699|false|false|false|C0332290|Consistent with|consistent
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3706,3713|false|false|false|C0205054|Hepatic|hepatic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3715,3724|false|false|false|C2711227|Steatohepatitis|steatosis
Event|Event|SIMPLE_SEGMENT|3715,3724|false|false|false|||steatosis
Finding|Pathologic Function|SIMPLE_SEGMENT|3715,3724|false|false|false|C0152254|Fatty degeneration|steatosis
Event|Event|SIMPLE_SEGMENT|3738,3746|true|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|3738,3746|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|3738,3749|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3756,3763|true|false|false|C0205054|Hepatic|hepatic
Finding|Finding|SIMPLE_SEGMENT|3756,3768|true|false|false|C0240225|Liver mass|hepatic mass
Event|Event|SIMPLE_SEGMENT|3764,3768|true|false|false|||mass
Finding|Finding|SIMPLE_SEGMENT|3764,3768|true|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|SIMPLE_SEGMENT|3764,3768|true|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|SIMPLE_SEGMENT|3764,3768|true|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Event|Event|SIMPLE_SEGMENT|3784,3796|true|false|false|||intrahepatic
Finding|Functional Concept|SIMPLE_SEGMENT|3784,3796|true|false|false|C1512952|Intrahepatic Route of Administration|intrahepatic
Finding|Functional Concept|SIMPLE_SEGMENT|3813,3820|true|false|false|C0521378|Biliary|biliary
Event|Event|SIMPLE_SEGMENT|3828,3838|true|false|false|||dilatation
Finding|Finding|SIMPLE_SEGMENT|3828,3838|true|false|false|C0012359;C0700124|Dilated;Pathological Dilatation|dilatation
Finding|Pathologic Function|SIMPLE_SEGMENT|3828,3838|true|false|false|C0012359;C0700124|Dilated;Pathological Dilatation|dilatation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3828,3838|true|false|false|C1322279|Dilate procedure|dilatation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3860,3870|true|false|false|C0008350;C0947622|Cholecystolithiasis;Cholelithiasis|gallstones
Event|Event|SIMPLE_SEGMENT|3860,3870|true|false|false|||gallstones
Finding|Body Substance|SIMPLE_SEGMENT|3860,3870|true|false|false|C0242216|Biliary calculi|gallstones
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3882,3893|true|false|false|C0016976;C1524055;C4071903|Abdomen>Gallbladder;Gallbladder;Gallbladder (MMHCC)|gallbladder
Anatomy|Tissue|SIMPLE_SEGMENT|3882,3893|true|false|false|C0016976;C1524055;C4071903|Abdomen>Gallbladder;Gallbladder;Gallbladder (MMHCC)|gallbladder
Procedure|Health Care Activity|SIMPLE_SEGMENT|3882,3893|true|false|false|C2032932|examination of gallbladder|gallbladder
Event|Event|SIMPLE_SEGMENT|3902,3910|true|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|3902,3910|true|false|false|C3887511|Evidence|evidence
Finding|Intellectual Product|SIMPLE_SEGMENT|3915,3920|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3915,3934|true|false|false|C0149520|Acute Cholecystitis|acute cholecystitis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3921,3934|true|false|false|C0008325|Cholecystitis|cholecystitis
Event|Event|SIMPLE_SEGMENT|3921,3934|true|false|false|||cholecystitis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3944,3950|true|false|false|C0037993;C4037984|Abdomen>Spleen;Spleen|spleen
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3944,3950|true|false|false|C0153470|Malignant neoplasm of spleen|spleen
Event|Event|SIMPLE_SEGMENT|3944,3950|true|false|false|||spleen
Finding|Finding|SIMPLE_SEGMENT|3944,3950|true|false|false|C0812414|Spleen problem|spleen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3944,3950|true|false|false|C0869677|Procedures on Spleen|spleen
Event|Event|SIMPLE_SEGMENT|3958,3966|true|false|false|||enlarged
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3980,3990|true|false|false|C0030274|Pancreas|pancreatic
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3980,3990|true|false|false|C0030292|Pancreatic Hormones|pancreatic
Drug|Hormone|SIMPLE_SEGMENT|3980,3990|true|false|false|C0030292|Pancreatic Hormones|pancreatic
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3980,3990|true|false|false|C0030292|Pancreatic Hormones|pancreatic
Event|Event|SIMPLE_SEGMENT|3991,3997|true|false|false|||ductal
Event|Event|SIMPLE_SEGMENT|3999,4009|true|false|false|||dilatation
Finding|Finding|SIMPLE_SEGMENT|3999,4009|true|false|false|C0012359;C0700124|Dilated;Pathological Dilatation|dilatation
Finding|Pathologic Function|SIMPLE_SEGMENT|3999,4009|true|false|false|C0012359;C0700124|Dilated;Pathological Dilatation|dilatation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3999,4009|true|false|false|C1322279|Dilate procedure|dilatation
Event|Event|SIMPLE_SEGMENT|4014,4022|true|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|4014,4022|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|4014,4025|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4026,4036|false|false|false|C0030274|Pancreas|pancreatic
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4026,4036|false|false|false|C0030292|Pancreatic Hormones|pancreatic
Drug|Hormone|SIMPLE_SEGMENT|4026,4036|false|false|false|C0030292|Pancreatic Hormones|pancreatic
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4026,4036|false|false|false|C0030292|Pancreatic Hormones|pancreatic
Finding|Finding|SIMPLE_SEGMENT|4026,4041|false|false|false|C0877425|Mass of pancreas|pancreatic mass
Event|Event|SIMPLE_SEGMENT|4037,4041|false|false|false|||mass
Finding|Finding|SIMPLE_SEGMENT|4037,4041|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|SIMPLE_SEGMENT|4037,4041|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|SIMPLE_SEGMENT|4037,4041|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Finding|SIMPLE_SEGMENT|4060,4067|true|false|false|C0700124|Dilated|dilated
Finding|Finding|SIMPLE_SEGMENT|4060,4073|true|false|false|C4697734|Dilated loops|dilated loops
Event|Event|SIMPLE_SEGMENT|4068,4073|true|false|false|||loops
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4077,4082|true|false|false|C0021853|Intestines|bowel
Event|Event|SIMPLE_SEGMENT|4096,4104|true|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|4096,4104|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|4096,4107|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4109,4114|true|false|false|C0021853|Intestines|bowel
Event|Event|SIMPLE_SEGMENT|4121,4131|true|false|false|||thickening
Finding|Finding|SIMPLE_SEGMENT|4121,4131|true|false|false|C0205400|Thickened|thickening
Finding|Finding|SIMPLE_SEGMENT|4145,4160|true|false|false|C1522583;C4760449|Intraperitoneal (intended site);Intraperitoneal Route of Administration|intraperitoneal
Finding|Functional Concept|SIMPLE_SEGMENT|4145,4160|true|false|false|C1522583;C4760449|Intraperitoneal (intended site);Intraperitoneal Route of Administration|intraperitoneal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4145,4169|true|false|false|C0032320|Pneumoperitoneum|intraperitoneal free air
Finding|Functional Concept|SIMPLE_SEGMENT|4161,4165|true|false|false|C0332296|Free of (attribute)|free
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4166,4169|true|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4166,4169|true|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|SIMPLE_SEGMENT|4166,4169|true|false|false|C0001861;C3536832|Air (substance);air|air
Event|Event|SIMPLE_SEGMENT|4166,4169|true|false|false|||air
Finding|Finding|SIMPLE_SEGMENT|4166,4169|true|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|SIMPLE_SEGMENT|4166,4169|true|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|SIMPLE_SEGMENT|4166,4169|true|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Event|Event|SIMPLE_SEGMENT|4173,4177|true|false|false|||free
Finding|Functional Concept|SIMPLE_SEGMENT|4173,4177|true|false|false|C0332296|Free of (attribute)|free
Finding|Pathologic Function|SIMPLE_SEGMENT|4173,4183|true|false|false|C0013687|effusion|free fluid
Drug|Substance|SIMPLE_SEGMENT|4178,4183|true|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|4178,4183|true|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|4178,4183|true|false|false|C1546638|Fluid Specimen Code|fluid
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4202,4210|true|false|false|C1293134|Enlargement procedure|enlarged
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4211,4219|true|false|false|C0018246|Inguinal region|inguinal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4221,4226|true|false|false|C0020889|Bone structure of ilium|iliac
Finding|Idea or Concept|SIMPLE_SEGMENT|4227,4232|true|false|false|C1524075|chain of objects|chain
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4251,4266|false|false|false|C0035359|Retroperitoneal Space|retroperitoneal
Finding|Body Substance|SIMPLE_SEGMENT|4267,4272|false|false|false|C0024202|Lymph|lymph
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4267,4278|false|false|false|C0024204|lymph nodes|lymph nodes
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4267,4278|false|false|false|C0154054|benign neoplasm of lymph nodes|lymph nodes
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4280,4289|false|false|false|C0000726|Abdomen|Abdominal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4280,4295|false|false|false|C0003484;C4037989|Abdomen>Aorta.abdominal;Abdominal aorta structure|Abdominal aorta
Procedure|Health Care Activity|SIMPLE_SEGMENT|4280,4295|false|false|false|C2228415|examination of abdominal aorta|Abdominal aorta
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4290,4295|false|false|false|C0003483;C4037978|Aorta;Chest+Abdomen>Aorta|aorta
Procedure|Health Care Activity|SIMPLE_SEGMENT|4290,4295|false|false|false|C0869784|Procedure on aorta|aorta
Event|Event|SIMPLE_SEGMENT|4309,4315|false|false|false|||course
Event|Event|SIMPLE_SEGMENT|4321,4328|false|false|false|||caliber
Finding|Finding|SIMPLE_SEGMENT|4334,4342|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|SIMPLE_SEGMENT|4334,4342|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Event|Event|SIMPLE_SEGMENT|4343,4358|false|false|false|||atherosclerotic
Finding|Functional Concept|SIMPLE_SEGMENT|4343,4358|false|false|false|C0333482|atherosclerotic|atherosclerotic
Event|Event|SIMPLE_SEGMENT|4359,4372|false|false|false|||calcification
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|4359,4372|false|false|false|C0006660;C0006663;C1533591|Calcification;Calcinosis;Physiologic calcification|calcification
Finding|Pathologic Function|SIMPLE_SEGMENT|4359,4372|false|false|false|C0006660;C0006663;C1533591|Calcification;Calcinosis;Physiologic calcification|calcification
Finding|Functional Concept|SIMPLE_SEGMENT|4384,4399|false|false|false|C0333482|atherosclerotic|atherosclerotic
Event|Event|SIMPLE_SEGMENT|4400,4413|false|false|false|||calcification
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|4400,4413|false|false|false|C0006660;C0006663;C1533591|Calcification;Calcinosis;Physiologic calcification|calcification
Finding|Pathologic Function|SIMPLE_SEGMENT|4400,4413|false|false|false|C0006660;C0006663;C1533591|Calcification;Calcinosis;Physiologic calcification|calcification
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4430,4440|false|false|false|C0025474|Mesentery|mesenteric
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4442,4448|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|SIMPLE_SEGMENT|4442,4448|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Event|Event|SIMPLE_SEGMENT|4449,4455|false|false|false|||origin
Finding|Classification|SIMPLE_SEGMENT|4449,4455|false|false|false|C0079946;C1550512|National origin;Participation Type - origin|origin
Finding|Intellectual Product|SIMPLE_SEGMENT|4449,4455|false|false|false|C0079946;C1550512|National origin;Participation Type - origin|origin
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4480,4487|true|false|false|C0262950;C4520924|Bone Tissue, Human;Skeletal bone|osseous
Anatomy|Tissue|SIMPLE_SEGMENT|4480,4487|true|false|false|C0262950;C4520924|Bone Tissue, Human;Skeletal bone|osseous
Event|Event|SIMPLE_SEGMENT|4488,4494|true|false|false|||lesion
Finding|Finding|SIMPLE_SEGMENT|4488,4494|true|true|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|SIMPLE_SEGMENT|4488,4494|true|true|false|C0221198;C1546698|Lesion|lesion
Event|Event|SIMPLE_SEGMENT|4500,4510|false|false|false|||IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|4500,4510|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|4500,4510|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Functional Concept|SIMPLE_SEGMENT|4536,4541|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|4542,4552|false|false|false|C0424290|Compulsive hoarding|collecting
Event|Event|SIMPLE_SEGMENT|4542,4552|false|false|false|||collecting
Finding|Functional Concept|SIMPLE_SEGMENT|4542,4552|false|false|false|C1516698|Collection (action)|collecting
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4553,4559|false|false|false|C5671121|System (basic dose form)|system
Finding|Functional Concept|SIMPLE_SEGMENT|4553,4559|false|false|false|C0449913;C5441654|System;System, LOINC Axis 4|system
Event|Event|SIMPLE_SEGMENT|4560,4568|false|false|false|||calculus
Finding|Body Substance|SIMPLE_SEGMENT|4560,4568|false|false|false|C0006736|Calculi|calculus
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4560,4568|false|false|false|C3668917|Calculus (lab procedure)|calculus
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4574,4581|false|false|false|C0205054|Hepatic|Hepatic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4574,4591|false|false|false|C0015695;C2711227|Fatty Liver;Steatohepatitis|Hepatic steatosis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4582,4591|false|false|false|C2711227|Steatohepatitis|steatosis
Event|Event|SIMPLE_SEGMENT|4582,4591|false|false|false|||steatosis
Finding|Pathologic Function|SIMPLE_SEGMENT|4582,4591|false|false|false|C0152254|Fatty degeneration|steatosis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4607,4616|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4607,4616|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|4607,4616|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Event|Event|SIMPLE_SEGMENT|4617,4626|false|false|false|||densities
Finding|Functional Concept|SIMPLE_SEGMENT|4634,4638|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Drug|Amino Acid Sequence|SIMPLE_SEGMENT|4647,4653|false|false|false|C1514562|Protein Domain|region
Event|Event|SIMPLE_SEGMENT|4655,4664|false|false|false|||measuring
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4687,4695|false|false|false|C2926606||findings
Event|Event|SIMPLE_SEGMENT|4687,4695|false|false|false|||findings
Finding|Functional Concept|SIMPLE_SEGMENT|4687,4695|false|false|false|C2607943|findings aspects|findings
Event|Event|SIMPLE_SEGMENT|4704,4713|false|false|false|||represent
Event|Event|SIMPLE_SEGMENT|4714,4719|false|false|false|||areas
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4724,4743|false|false|false|C2062952|Round atelectasis|rounded atelectasis
Event|Event|SIMPLE_SEGMENT|4732,4743|false|false|false|||atelectasis
Finding|Pathologic Function|SIMPLE_SEGMENT|4732,4743|false|false|false|C0004144|Atelectasis|atelectasis
Finding|Idea or Concept|SIMPLE_SEGMENT|4759,4763|false|false|false|C0233324;C1705313|Term (lexical);Term Birth|term
Finding|Organism Function|SIMPLE_SEGMENT|4759,4763|false|false|false|C0233324;C1705313|Term (lexical);Term Birth|term
Event|Event|SIMPLE_SEGMENT|4764,4772|false|false|false|||followup
Procedure|Health Care Activity|SIMPLE_SEGMENT|4764,4772|false|false|false|C1522577|follow-up|followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4791,4799|false|false|true|C0881858||CT chest
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4791,4799|false|false|true|C0202823|Chest CT|CT chest
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4794,4799|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Event|Event|SIMPLE_SEGMENT|4794,4799|false|false|false|||chest
Finding|Finding|SIMPLE_SEGMENT|4794,4799|false|false|false|C0741025|Chest problem|chest
Event|Event|SIMPLE_SEGMENT|4803,4814|false|false|false|||recommended
Procedure|Health Care Activity|SIMPLE_SEGMENT|4818,4827|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|SIMPLE_SEGMENT|4828,4832|false|false|false|||LABS
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4828,4832|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4846,4851|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4846,4851|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4846,4851|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|4852,4855|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|4860,4863|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4860,4863|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4860,4863|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4870,4873|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4870,4873|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|4870,4873|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4870,4873|false|false|false|C0019029|Hemoglobin concentration|Hgb
Event|Event|SIMPLE_SEGMENT|4879,4882|false|false|false|||Hct
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4879,4882|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4879,4882|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|4889,4892|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|4889,4892|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4889,4892|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4889,4892|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4889,4892|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|4896,4899|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4896,4899|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|4896,4899|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|4896,4899|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|4896,4899|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4896,4899|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4906,4910|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4926,4929|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4946,4951|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4946,4951|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4946,4951|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Antibiotic|SIMPLE_SEGMENT|4968,4973|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4968,4973|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|SIMPLE_SEGMENT|4968,4973|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4978,4981|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|Eos
Event|Event|SIMPLE_SEGMENT|4978,4981|false|false|false|||Eos
Finding|Gene or Genome|SIMPLE_SEGMENT|4978,4981|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|Eos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5008,5013|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5008,5013|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5008,5013|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|5008,5021|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5008,5021|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5008,5021|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5014,5021|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|5014,5021|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5014,5021|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|5014,5021|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5014,5021|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5014,5021|false|false|false|C0337438|Glucose measurement|Glucose
Event|Event|SIMPLE_SEGMENT|5057,5058|false|false|false|||5
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5068,5072|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5068,5072|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5068,5072|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5099,5104|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5099,5104|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5099,5104|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5105,5108|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5105,5108|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|SIMPLE_SEGMENT|5105,5108|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|SIMPLE_SEGMENT|5105,5108|false|false|false|||ALT
Finding|Gene or Genome|SIMPLE_SEGMENT|5105,5108|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|SIMPLE_SEGMENT|5105,5108|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|SIMPLE_SEGMENT|5105,5108|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5105,5108|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5112,5115|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5112,5115|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5112,5115|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5112,5115|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|SIMPLE_SEGMENT|5112,5115|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|SIMPLE_SEGMENT|5112,5115|false|false|false|||AST
Finding|Gene or Genome|SIMPLE_SEGMENT|5112,5115|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5120,5127|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|SIMPLE_SEGMENT|5120,5127|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5155,5160|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5155,5160|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5155,5160|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5155,5168|false|false|false|C0853248|Blood albumin|BLOOD Albumin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5161,5168|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5161,5168|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5161,5168|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Event|Event|SIMPLE_SEGMENT|5161,5168|false|false|false|||Albumin
Finding|Gene or Genome|SIMPLE_SEGMENT|5161,5168|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Finding|Physiologic Function|SIMPLE_SEGMENT|5161,5168|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5161,5168|false|false|false|C0201838|Albumin measurement|Albumin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5173,5180|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|5173,5180|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5173,5180|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5173,5180|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|5173,5180|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|SIMPLE_SEGMENT|5173,5180|false|false|false|||Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|5173,5180|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5173,5180|false|false|false|C0201925|Calcium measurement|Calcium
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5213,5218|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5213,5218|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5213,5218|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5245,5250|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5245,5250|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5245,5250|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5251,5257|false|false|false|C0023764|lipase|Lipase
Drug|Enzyme|SIMPLE_SEGMENT|5251,5257|false|false|false|C0023764|lipase|Lipase
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5251,5257|false|false|false|C0023764|lipase|Lipase
Event|Event|SIMPLE_SEGMENT|5251,5257|false|false|false|||Lipase
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5251,5257|false|false|false|C0373670|Lipase measurement|Lipase
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5274,5279|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5274,5279|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5274,5279|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Event|Event|SIMPLE_SEGMENT|5284,5287|false|false|false|||pO2
Finding|Classification|SIMPLE_SEGMENT|5284,5287|false|false|false|C0391840;C4521535|Partial pressure of Oxygen;US Military enlisted E5|pO2
Finding|Molecular Function|SIMPLE_SEGMENT|5284,5287|false|false|false|C0391840;C4521535|Partial pressure of Oxygen;US Military enlisted E5|pO2
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5284,5287|false|false|false|C1283004|PO2 measurement|pO2
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5292,5296|false|false|false|C0391839|Carbon dioxide, partial pressure|pCO2
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5292,5296|false|false|false|C0201931|Carbon dioxide measurement, partial pressure|pCO2
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5320,5324|false|false|false|C2987514|Anatomical base|Base
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5320,5324|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|Base
Drug|Chemical Viewed Functionally|SIMPLE_SEGMENT|5320,5324|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|Base
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|5320,5324|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|Base
Finding|Gene or Genome|SIMPLE_SEGMENT|5320,5324|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|Base
Finding|Idea or Concept|SIMPLE_SEGMENT|5320,5324|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|Base
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5342,5347|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5342,5347|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5342,5355|false|false|false|C3824990|lactate in blood (lab test)|BLOOD Lactate
Drug|Organic Chemical|SIMPLE_SEGMENT|5348,5355|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5348,5355|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Event|Event|SIMPLE_SEGMENT|5348,5355|false|false|false|||Lactate
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5348,5355|false|false|false|C0202115|Lactic acid measurement|Lactate
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5379,5384|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5379,5384|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5379,5384|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5388,5391|false|false|false|C2744672|SAT1 protein, human|Sat
Drug|Enzyme|SIMPLE_SEGMENT|5388,5391|false|false|false|C2744672|SAT1 protein, human|Sat
Finding|Gene or Genome|SIMPLE_SEGMENT|5388,5391|false|false|false|C0871290;C1705827;C1822614|College Entrance Examination Board Scholastic Aptitude Test;SAT1 gene;SAT1 wt Allele|Sat
Finding|Intellectual Product|SIMPLE_SEGMENT|5388,5391|false|false|false|C0871290;C1705827;C1822614|College Entrance Examination Board Scholastic Aptitude Test;SAT1 gene;SAT1 wt Allele|Sat
Finding|Body Substance|SIMPLE_SEGMENT|5407,5412|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|5407,5412|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|5407,5412|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5407,5418|false|false|false|C0018965|Hematuria|URINE Blood
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5413,5418|false|false|false|C0851353|Blood and lymphatic system disorders|Blood
Finding|Body Substance|SIMPLE_SEGMENT|5413,5418|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Event|Event|SIMPLE_SEGMENT|5419,5422|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|5419,5422|false|false|false|C5848551|Neg - answer|NEG
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5423,5430|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|Nitrite
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5423,5430|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|Nitrite
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5423,5430|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|Nitrite
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5431,5434|false|false|false|C1744592|Structure of parieto-occipital fissure|POS
Finding|Intellectual Product|SIMPLE_SEGMENT|5431,5434|false|false|false|C5891108|Health Maintenance Organization Point of Service Plan|POS
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5435,5442|false|false|false|C0033684|Proteins|Protein
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5435,5442|false|false|false|C0033684|Proteins|Protein
Event|Event|SIMPLE_SEGMENT|5435,5442|false|false|false|||Protein
Finding|Conceptual Entity|SIMPLE_SEGMENT|5435,5442|false|false|false|C1521746|Protein Info|Protein
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5435,5442|false|false|false|C0202202|Protein measurement|Protein
Event|Event|SIMPLE_SEGMENT|5443,5446|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|5443,5446|false|false|false|C5848551|Neg - answer|NEG
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5448,5455|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|5448,5455|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5448,5455|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|5448,5455|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5448,5455|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5448,5455|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|5461,5467|false|false|false|C0022634|Ketones|Ketone
Finding|Finding|SIMPLE_SEGMENT|5479,5482|false|false|false|C5848551|Neg - answer|NEG
Finding|Finding|SIMPLE_SEGMENT|5491,5494|false|false|false|C5848551|Neg - answer|NEG
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5508,5511|false|false|false|C0011860|Diabetes Mellitus, Non-Insulin-Dependent|MOD
Event|Event|SIMPLE_SEGMENT|5508,5511|false|false|false|||MOD
Finding|Body Substance|SIMPLE_SEGMENT|5524,5529|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|5524,5529|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|5524,5529|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5524,5533|false|false|false|C0221752;C2188659|Red blood cells urine positive|URINE RBC
Anatomy|Cell|SIMPLE_SEGMENT|5530,5533|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5530,5533|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5530,5533|false|false|false|C0014792|Erythrocytes|RBC
Anatomy|Cell|SIMPLE_SEGMENT|5537,5540|false|false|false|C0023516|Leukocytes|WBC
Drug|Food|SIMPLE_SEGMENT|5557,5562|true|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|Yeast
Drug|Immunologic Factor|SIMPLE_SEGMENT|5557,5562|true|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|Yeast
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|5557,5562|true|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|Yeast
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5557,5562|true|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|Yeast
Event|Event|SIMPLE_SEGMENT|5563,5567|false|false|false|||NONE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5569,5572|true|false|false|C0267963|Exocrine pancreatic insufficiency|Epi
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5569,5572|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5569,5572|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Hormone|SIMPLE_SEGMENT|5569,5572|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Organic Chemical|SIMPLE_SEGMENT|5569,5572|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5569,5572|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Event|Event|SIMPLE_SEGMENT|5569,5572|true|false|false|||Epi
Finding|Gene or Genome|SIMPLE_SEGMENT|5569,5572|true|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|Epi
Finding|Intellectual Product|SIMPLE_SEGMENT|5569,5572|true|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|Epi
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5569,5572|true|false|false|C0162734;C3641909|Echo-Planar Imaging;Electronic Portal Imaging|Epi
Finding|Body Substance|SIMPLE_SEGMENT|5597,5602|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|5597,5602|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|5597,5602|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Finding|SIMPLE_SEGMENT|5597,5608|false|false|false|C0278030|Color of urine|URINE Color
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5603,5608|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|Color
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|5603,5608|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|Color
Drug|Organic Chemical|SIMPLE_SEGMENT|5609,5614|false|false|false|C4047917|Cereal plant straw|Straw
Finding|Idea or Concept|SIMPLE_SEGMENT|5622,5627|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|SIMPLE_SEGMENT|5646,5650|false|false|false|||LABS
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5646,5650|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5664,5669|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5664,5669|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5664,5669|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|5670,5673|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|5678,5681|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5678,5681|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5678,5681|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5688,5691|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5688,5691|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|5688,5691|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5688,5691|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5698,5701|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5698,5701|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|5709,5712|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|5709,5712|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5709,5712|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5709,5712|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5709,5712|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|5716,5719|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5716,5719|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|5716,5719|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|5716,5719|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|5716,5719|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5716,5719|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5726,5730|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5746,5749|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5766,5771|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5766,5771|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5766,5771|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Antibiotic|SIMPLE_SEGMENT|5787,5792|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5787,5792|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|SIMPLE_SEGMENT|5787,5792|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5797,5800|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|Eos
Event|Event|SIMPLE_SEGMENT|5797,5800|false|false|false|||Eos
Finding|Gene or Genome|SIMPLE_SEGMENT|5797,5800|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|Eos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5827,5832|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5827,5832|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5827,5832|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|5827,5840|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5827,5840|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5827,5840|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5833,5840|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|5833,5840|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5833,5840|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|5833,5840|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5833,5840|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5833,5840|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5886,5890|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5886,5890|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5886,5890|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5915,5920|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5915,5920|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5915,5920|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5921,5924|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5921,5924|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|SIMPLE_SEGMENT|5921,5924|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|SIMPLE_SEGMENT|5921,5924|false|false|false|||ALT
Finding|Gene or Genome|SIMPLE_SEGMENT|5921,5924|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|SIMPLE_SEGMENT|5921,5924|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|SIMPLE_SEGMENT|5921,5924|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5921,5924|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5928,5931|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5928,5931|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5928,5931|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5928,5931|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|SIMPLE_SEGMENT|5928,5931|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|SIMPLE_SEGMENT|5928,5931|false|false|false|||AST
Finding|Gene or Genome|SIMPLE_SEGMENT|5928,5931|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5935,5942|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|SIMPLE_SEGMENT|5935,5942|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5958,5963|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5958,5963|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5958,5963|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5958,5971|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5964,5971|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|5964,5971|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5964,5971|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5964,5971|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|5964,5971|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|SIMPLE_SEGMENT|5964,5971|false|false|false|||Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|5964,5971|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5964,5971|false|false|false|C0201925|Calcium measurement|Calcium
Finding|Intellectual Product|SIMPLE_SEGMENT|5996,6001|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|Brief
Finding|Idea or Concept|SIMPLE_SEGMENT|6002,6010|false|false|false|C1547192|Organization unit type - Hospital|Hospital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6002,6017|false|false|false|C0488549||Hospital Course
Finding|Finding|SIMPLE_SEGMENT|6002,6017|false|false|false|C0489547|Hospital course|Hospital Course
Event|Event|SIMPLE_SEGMENT|6023,6026|false|false|false|||PMH
Finding|Finding|SIMPLE_SEGMENT|6023,6026|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|PMH
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6032,6035|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|SIMPLE_SEGMENT|6032,6035|false|false|false|||HTN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6037,6041|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Event|Event|SIMPLE_SEGMENT|6037,6041|false|false|false|||GERD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6043,6046|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6043,6046|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|6043,6046|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|6043,6046|false|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|6043,6046|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6043,6046|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|6043,6046|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6043,6046|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Event|Event|SIMPLE_SEGMENT|6051,6055|false|false|false|||CABG
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6051,6055|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Event|Event|SIMPLE_SEGMENT|6060,6068|false|false|false|||stenting
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6060,6068|false|false|false|C2348535|Stenting|stenting
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6070,6074|false|false|false|C0011854|Diabetes Mellitus, Insulin-Dependent|IDDM
Event|Event|SIMPLE_SEGMENT|6070,6074|false|false|false|||IDDM
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6083,6088|false|false|false|C0230171|Flank (surface region)|flank
Finding|Sign or Symptom|SIMPLE_SEGMENT|6083,6093|false|false|false|C0016199|Flank Pain|flank pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6089,6093|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|6089,6093|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|6089,6093|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|6089,6093|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|6094,6102|false|false|false|||presumed
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6106,6121|false|false|false|C2707260||musculoskeletal
Event|Event|SIMPLE_SEGMENT|6106,6121|false|false|false|||musculoskeletal
Finding|Functional Concept|SIMPLE_SEGMENT|6106,6121|false|false|false|C0497254|Musculoskeletal|musculoskeletal
Event|Event|SIMPLE_SEGMENT|6125,6131|false|false|false|||nature
Finding|Functional Concept|SIMPLE_SEGMENT|6125,6131|false|false|false|C0349590;C1262865|Nature;Natures|nature
Finding|Idea or Concept|SIMPLE_SEGMENT|6125,6131|false|false|false|C0349590;C1262865|Nature;Natures|nature
Event|Event|SIMPLE_SEGMENT|6139,6147|false|false|false|||negative
Finding|Classification|SIMPLE_SEGMENT|6139,6147|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|6139,6147|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6139,6147|false|false|false|C5237010|Expression Negative|negative
Event|Event|SIMPLE_SEGMENT|6149,6155|false|false|false|||workup
Finding|Functional Concept|SIMPLE_SEGMENT|6157,6167|false|false|false|C0444507|Incidental|Incidental
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6168,6171|false|false|false|C0042029|Urinary tract infection|UTI
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6168,6171|false|false|false|C0077906|urinastatin|UTI
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6168,6171|false|false|false|C0077906|urinastatin|UTI
Event|Event|SIMPLE_SEGMENT|6168,6171|false|false|false|||UTI
Finding|Gene or Genome|SIMPLE_SEGMENT|6168,6171|false|false|false|C1412376;C5780748|AMBP gene;AMBP wt Allele|UTI
Finding|Finding|SIMPLE_SEGMENT|6174,6186|false|false|false|C0231221;C0332151|Asymptomatic (finding);Asymptomatic diagnosis of|asymptomatic
Event|Event|SIMPLE_SEGMENT|6187,6195|false|false|false|||bacturia
Finding|Intellectual Product|SIMPLE_SEGMENT|6198,6203|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|ACUTE
Event|Event|SIMPLE_SEGMENT|6204,6210|false|false|false|||ISSUES
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6215,6218|false|false|false|C0042029|Urinary tract infection|UTI
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6215,6218|false|false|false|C0077906|urinastatin|UTI
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6215,6218|false|false|false|C0077906|urinastatin|UTI
Event|Event|SIMPLE_SEGMENT|6215,6218|false|false|false|||UTI
Finding|Gene or Genome|SIMPLE_SEGMENT|6215,6218|false|false|false|C1412376;C5780748|AMBP gene;AMBP wt Allele|UTI
Finding|Body Substance|SIMPLE_SEGMENT|6231,6238|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|6231,6238|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|6231,6238|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|6239,6248|true|false|false|||presented
Event|Event|SIMPLE_SEGMENT|6261,6268|true|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|6261,6268|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|6261,6268|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|6261,6268|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|6261,6271|true|false|false|C0262926|Medical History|history of
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6273,6280|true|false|false|C0042027|Urinary tract|urinary
Finding|Functional Concept|SIMPLE_SEGMENT|6284,6292|true|false|false|C0205373;C5849094|Systemic;Systemic Route of Administration|systemic
Finding|Sign or Symptom|SIMPLE_SEGMENT|6284,6301|true|false|false|C2039684|systemic symptoms|systemic symptoms
Event|Event|SIMPLE_SEGMENT|6293,6301|true|false|false|||symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|6293,6301|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|6293,6301|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|SIMPLE_SEGMENT|6311,6318|false|false|false|||started
Drug|Antibiotic|SIMPLE_SEGMENT|6322,6333|false|false|false|C0007561|ceftriaxone|ceftriaxone
Drug|Organic Chemical|SIMPLE_SEGMENT|6322,6333|false|false|false|C0007561|ceftriaxone|ceftriaxone
Event|Event|SIMPLE_SEGMENT|6334,6336|false|false|false|||in
Event|Event|SIMPLE_SEGMENT|6342,6344|false|false|false|||ED
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|6364,6372|false|false|false|C4727483|BRAF Gene Rearrangement|positive
Event|Event|SIMPLE_SEGMENT|6364,6372|false|false|false|||positive
Finding|Classification|SIMPLE_SEGMENT|6364,6372|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|SIMPLE_SEGMENT|6364,6372|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Anatomy|Cell|SIMPLE_SEGMENT|6380,6384|false|false|false|C0023516|Leukocytes|WBCs
Drug|Antibiotic|SIMPLE_SEGMENT|6387,6398|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|Antibiotics
Event|Event|SIMPLE_SEGMENT|6387,6398|false|false|false|||Antibiotics
Event|Event|SIMPLE_SEGMENT|6404,6409|false|false|false|||taken
Event|Event|SIMPLE_SEGMENT|6419,6426|false|false|false|||drawing
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6427,6434|false|false|false|C0042027|Urinary tract|urinary
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6438,6443|true|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|6438,6443|true|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|6438,6443|true|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Event|Event|SIMPLE_SEGMENT|6445,6453|true|false|false|||cultures
Finding|Idea or Concept|SIMPLE_SEGMENT|6445,6453|true|false|false|C0010453|Culture (Anthropological)|cultures
Event|Event|SIMPLE_SEGMENT|6472,6477|true|false|false|||yield
Finding|Body Substance|SIMPLE_SEGMENT|6479,6486|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|6479,6486|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|6479,6486|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|6487,6495|false|false|false|||switched
Drug|Organic Chemical|SIMPLE_SEGMENT|6500,6513|false|false|false|C0008809|ciprofloxacin|ciprofloxacin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6500,6513|false|false|false|C0008809|ciprofloxacin|ciprofloxacin
Event|Event|SIMPLE_SEGMENT|6500,6513|false|false|false|||ciprofloxacin
Event|Event|SIMPLE_SEGMENT|6518,6526|false|false|false|||received
Finding|Idea or Concept|SIMPLE_SEGMENT|6535,6538|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|6535,6538|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Antibiotic|SIMPLE_SEGMENT|6545,6555|false|false|false|C0003232|Antibiotics|antibiotic
Event|Event|SIMPLE_SEGMENT|6556,6562|false|false|false|||course
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6565,6572|true|false|false|C0040405|X-Ray Computed Tomography|CT scan
Event|Event|SIMPLE_SEGMENT|6568,6572|true|false|false|||scan
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6568,6572|true|false|false|C0034606;C0441633|Radionuclide Imaging;Scanning|scan
Event|Event|SIMPLE_SEGMENT|6600,6608|true|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|6600,6608|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|6600,6611|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6612,6626|true|false|false|C0034186|Pyelonephritis|pyelonephritis
Event|Event|SIMPLE_SEGMENT|6612,6626|true|false|false|||pyelonephritis
Drug|Antibiotic|SIMPLE_SEGMENT|6629,6640|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|Antibiotics
Event|Event|SIMPLE_SEGMENT|6629,6640|false|false|false|||Antibiotics
Event|Event|SIMPLE_SEGMENT|6646,6658|false|false|false|||discontinued
Finding|Finding|SIMPLE_SEGMENT|6662,6666|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|6662,6666|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|6662,6666|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|SIMPLE_SEGMENT|6670,6679|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|6670,6679|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|6670,6679|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|6670,6679|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|6670,6679|false|false|false|C0030685|Patient Discharge|discharge
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6684,6689|false|false|false|C0230171|Flank (surface region)|Flank
Finding|Sign or Symptom|SIMPLE_SEGMENT|6684,6694|false|false|false|C0016199|Flank Pain|Flank Pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6690,6694|false|false|false|C2598155||Pain
Event|Event|SIMPLE_SEGMENT|6690,6694|false|false|false|||Pain
Finding|Functional Concept|SIMPLE_SEGMENT|6690,6694|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|6690,6694|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Body Substance|SIMPLE_SEGMENT|6697,6704|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|6697,6704|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|6697,6704|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|6705,6713|false|false|false|||reported
Event|Event|SIMPLE_SEGMENT|6716,6721|false|false|false|||weeks
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6730,6735|false|false|false|C0230171|Flank (surface region)|flank
Finding|Sign or Symptom|SIMPLE_SEGMENT|6730,6740|false|false|false|C0016199|Flank Pain|flank pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6736,6740|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|6736,6740|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|6736,6740|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|6736,6740|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|6742,6750|false|false|false|||constant
Finding|Intellectual Product|SIMPLE_SEGMENT|6742,6750|false|false|false|C1720529|Constant - dosing instruction fragment|constant
Finding|Functional Concept|SIMPLE_SEGMENT|6764,6770|false|false|false|C0349590;C1262865|Nature;Natures|nature
Finding|Idea or Concept|SIMPLE_SEGMENT|6764,6770|false|false|false|C0349590;C1262865|Nature;Natures|nature
Event|Event|SIMPLE_SEGMENT|6775,6783|false|false|false|||worsened
Event|Event|SIMPLE_SEGMENT|6787,6795|false|false|false|||movement
Finding|Organism Function|SIMPLE_SEGMENT|6787,6795|false|false|false|C0026649|Movement|movement
Event|Event|SIMPLE_SEGMENT|6797,6804|false|false|false|||Treated
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6811,6830|false|false|false|C0003209|Anti-Inflammatory Agents|anti-inflammatories
Event|Event|SIMPLE_SEGMENT|6811,6830|false|false|false|||anti-inflammatories
Event|Event|SIMPLE_SEGMENT|6844,6850|false|false|false|||effect
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6852,6859|true|false|false|C0040405|X-Ray Computed Tomography|CT scan
Event|Event|SIMPLE_SEGMENT|6855,6859|true|false|false|||scan
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6855,6859|true|false|false|C0034606;C0441633|Radionuclide Imaging;Scanning|scan
Event|Event|SIMPLE_SEGMENT|6860,6872|true|false|false|||demonstrated
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6877,6892|true|false|false|C0392525|Nephrolithiasis|nephrolithiasis
Event|Event|SIMPLE_SEGMENT|6877,6892|true|false|false|||nephrolithiasis
Event|Event|SIMPLE_SEGMENT|6894,6897|true|false|false|||CXR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6894,6897|true|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|SIMPLE_SEGMENT|6898,6904|true|false|false|||showed
Finding|Functional Concept|SIMPLE_SEGMENT|6908,6912|true|false|false|C0443157|Bony|bony
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|6913,6924|true|false|false|C0000768|Congenital Abnormality|abnormality
Event|Event|SIMPLE_SEGMENT|6913,6924|true|false|false|||abnormality
Finding|Finding|SIMPLE_SEGMENT|6913,6924|true|false|false|C1704258|Abnormality|abnormality
Finding|Finding|SIMPLE_SEGMENT|6941,6948|true|false|false|C4699603|Totally|totally
Event|Event|SIMPLE_SEGMENT|6949,6956|true|false|false|||exclude
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|6957,6979|true|false|false|C0272567|Fracture of multiple ribs|multiple rib fractures
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6966,6969|true|false|false|C0035561|Bone structure of rib|rib
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|6966,6979|true|false|false|C0035522|Rib Fractures|rib fractures
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|6970,6979|true|false|false|C0016658|Fracture|fractures
Event|Event|SIMPLE_SEGMENT|6970,6979|true|false|false|||fractures
Finding|Finding|SIMPLE_SEGMENT|6970,6979|true|false|false|C4554413|Fractured|fractures
Finding|Body Substance|SIMPLE_SEGMENT|6981,6988|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|6981,6988|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|6981,6988|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6991,6995|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|6991,6995|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|6991,6995|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|6991,6995|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|7000,7004|false|false|false|||well
Finding|Finding|SIMPLE_SEGMENT|7000,7004|false|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|7006,7016|false|false|false|||controlled
Event|Event|SIMPLE_SEGMENT|7021,7031|false|false|false|||tolerating
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7035,7046|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7035,7046|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|7035,7046|false|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|7035,7046|false|false|false|C4284232|Medications|medications
Event|Event|SIMPLE_SEGMENT|7059,7069|false|false|false|||discharged
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7076,7079|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|7076,7079|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7076,7079|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7076,7079|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|SIMPLE_SEGMENT|7076,7079|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|7076,7079|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|SIMPLE_SEGMENT|7076,7079|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7076,7079|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|SIMPLE_SEGMENT|7076,7079|false|false|false|||PCP
Finding|Gene or Genome|SIMPLE_SEGMENT|7076,7079|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|SIMPLE_SEGMENT|7076,7079|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Event|SIMPLE_SEGMENT|7080,7089|false|false|false|||following
Event|Event|SIMPLE_SEGMENT|7102,7108|false|false|false|||workup
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7113,7121|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|Diabetes
Event|Event|SIMPLE_SEGMENT|7113,7121|false|false|false|||Diabetes
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7124,7137|false|false|false|C0020456|Hyperglycemia|Hyperglycemia
Event|Event|SIMPLE_SEGMENT|7124,7137|false|false|false|||Hyperglycemia
Finding|Finding|SIMPLE_SEGMENT|7124,7137|false|false|false|C2919432|Glucose in blood specimen above reference range|Hyperglycemia
Finding|Body Substance|SIMPLE_SEGMENT|7139,7146|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|7139,7146|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|7139,7146|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|7151,7163|false|false|false|||persistently
Finding|Idea or Concept|SIMPLE_SEGMENT|7151,7163|false|false|false|C0750508|persistently|persistently
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7168,7172|false|false|false|C0011854|Diabetes Mellitus, Insulin-Dependent|IDDM
Event|Event|SIMPLE_SEGMENT|7168,7172|false|false|false|||IDDM
Event|Event|SIMPLE_SEGMENT|7179,7182|false|false|false|||A1C
Finding|Classification|SIMPLE_SEGMENT|7179,7182|false|false|false|C4521595|United States Military enlisted E3 (qualifier value)|A1C
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7179,7182|false|false|false|C0474680|Hemoglobin A1c measurement|A1C
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|7194,7199|false|false|false|C5575602|Cell Culture Serum|Serum
Finding|Body Substance|SIMPLE_SEGMENT|7194,7199|false|false|false|C0229671;C1546774;C1550100|Serum;Serum specimen|Serum
Finding|Intellectual Product|SIMPLE_SEGMENT|7194,7199|false|false|false|C0229671;C1546774;C1550100|Serum;Serum specimen|Serum
Finding|Finding|SIMPLE_SEGMENT|7194,7207|false|false|false|C3534430|Serum glucose|Serum glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7194,7207|false|false|false|C0202041|Glucose measurement, serum|Serum glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7200,7207|false|false|false|C0017725|glucose|glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|7200,7207|false|false|false|C0017725|glucose|glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7200,7207|false|false|false|C0017725|glucose|glucose
Event|Event|SIMPLE_SEGMENT|7200,7207|false|false|false|||glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|7200,7207|false|false|false|C5781949|Glucose^1.5H post dose glucagon|glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7200,7207|false|false|false|C0337438|Glucose measurement|glucose
Event|Event|SIMPLE_SEGMENT|7235,7239|false|false|false|||Chem
Finding|Functional Concept|SIMPLE_SEGMENT|7235,7239|false|false|false|C0079107|chemical aspects|Chem
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7235,7239|false|false|false|C0201682|Chemical procedure|Chem
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7247,7250|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|gap
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7247,7250|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|gap
Finding|Gene or Genome|SIMPLE_SEGMENT|7247,7250|false|false|false|C1419277;C2984552|RASA1 gene;RASA1 wt Allele|gap
Finding|Finding|SIMPLE_SEGMENT|7270,7276|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|7270,7276|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Drug|Organic Chemical|SIMPLE_SEGMENT|7281,7288|false|false|false|C0022924;C0376261|Lactates;lactate|lactate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7281,7288|false|false|false|C0022924;C0376261|Lactates;lactate|lactate
Event|Event|SIMPLE_SEGMENT|7281,7288|false|false|false|||lactate
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7281,7288|false|false|false|C0202115|Lactic acid measurement|lactate
Event|Event|SIMPLE_SEGMENT|7294,7302|false|false|false|||unlikely
Finding|Finding|SIMPLE_SEGMENT|7294,7302|false|false|false|C0750558|Unlikely|unlikely
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7309,7312|false|false|false|C0011880|Diabetic Ketoacidosis|DKA
Event|Event|SIMPLE_SEGMENT|7309,7312|false|false|false|||DKA
Event|Event|SIMPLE_SEGMENT|7332,7335|false|false|false|||ABG
Finding|Gene or Genome|SIMPLE_SEGMENT|7332,7335|false|false|false|C1412045|A1BG gene|ABG
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7332,7335|false|false|false|C0150411|Analysis of arterial blood gases and pH|ABG
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7340,7347|false|false|false|C0017725|glucose|glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|7340,7347|false|false|false|C0017725|glucose|glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7340,7347|false|false|false|C0017725|glucose|glucose
Event|Event|SIMPLE_SEGMENT|7340,7347|false|false|false|||glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|7340,7347|false|false|false|C5781949|Glucose^1.5H post dose glucagon|glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7340,7347|false|false|false|C0337438|Glucose measurement|glucose
Finding|Idea or Concept|SIMPLE_SEGMENT|7355,7363|false|false|false|C0549178|Continuous|continue
Event|Event|SIMPLE_SEGMENT|7364,7368|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|7364,7368|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|7364,7368|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|7364,7368|false|false|false|C1553498|home health encounter|home
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7374,7380|false|false|false|C0876064|Lantus|lantus
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7374,7380|false|false|false|C0876064|Lantus|lantus
Event|Event|SIMPLE_SEGMENT|7374,7380|false|false|false|||lantus
Event|Event|SIMPLE_SEGMENT|7406,7413|false|false|false|||records
Finding|Idea or Concept|SIMPLE_SEGMENT|7406,7413|false|false|false|C0034869;C1548330|Quantity limited request - Records;Records|records
Finding|Intellectual Product|SIMPLE_SEGMENT|7406,7413|false|false|false|C0034869;C1548330|Quantity limited request - Records;Records|records
Finding|Individual Behavior|SIMPLE_SEGMENT|7428,7438|false|false|false|C0001807;C1547300;C1548760|Aggressive behavior;Precaution Code - Aggressive;Risk Codes - Aggressive|aggressive
Finding|Intellectual Product|SIMPLE_SEGMENT|7428,7438|false|false|false|C0001807;C1547300;C1548760|Aggressive behavior;Precaution Code - Aggressive;Risk Codes - Aggressive|aggressive
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|7439,7442|false|false|false|C1845118|SHORT STATURE, IDIOPATHIC, X-LINKED|ISS
Event|Event|SIMPLE_SEGMENT|7439,7442|false|false|false|||ISS
Event|Event|SIMPLE_SEGMENT|7449,7457|false|false|false|||decrease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7523,7526|false|false|false|C1561643|Chronic Kidney Diseases|CKD
Event|Event|SIMPLE_SEGMENT|7523,7526|false|false|false|||CKD
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7552,7560|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|SIMPLE_SEGMENT|7552,7560|false|false|false|||baseline
Finding|Idea or Concept|SIMPLE_SEGMENT|7552,7560|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Finding|Idea or Concept|SIMPLE_SEGMENT|7566,7577|false|false|false|C0750501|most likely|Most likely
Finding|Finding|SIMPLE_SEGMENT|7571,7577|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|7571,7577|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|SIMPLE_SEGMENT|7579,7588|false|false|false|||pre-renal
Finding|Mental Process|SIMPLE_SEGMENT|7596,7603|false|false|false|C0542559|contextual factors|setting
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7607,7616|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|SIMPLE_SEGMENT|7607,7616|false|false|false|||infection
Finding|Pathologic Function|SIMPLE_SEGMENT|7607,7616|false|false|false|C3714514|Infection|infection
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|7629,7632|false|false|false|C0016520|Structure of interventricular foramen|IVF
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7629,7632|false|false|false|C2751898|Ventricular Fibrillation, Paroxysmal Familial, 1|IVF
Event|Event|SIMPLE_SEGMENT|7629,7632|false|false|false|||IVF
Finding|Gene or Genome|SIMPLE_SEGMENT|7629,7632|false|false|false|C1419864;C4321334|SCN5A gene;SCN5A wt Allele|IVF
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7629,7632|false|false|false|C0015915;C0872104|Assisted Reproductive Technologies;Fertilization in Vitro|IVF
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7648,7658|false|false|false|C0010294|creatinine|creatinine
Drug|Organic Chemical|SIMPLE_SEGMENT|7648,7658|false|false|false|C0010294|creatinine|creatinine
Event|Event|SIMPLE_SEGMENT|7648,7658|false|false|false|||creatinine
Finding|Physiologic Function|SIMPLE_SEGMENT|7648,7658|false|false|false|C4551889|Creatinine metabolic function|creatinine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7648,7658|false|false|false|C0201975|Creatinine measurement|creatinine
Event|Event|SIMPLE_SEGMENT|7663,7672|false|false|false|||corrected
Event|Event|SIMPLE_SEGMENT|7689,7698|false|false|false|||euvolemic
Finding|Finding|SIMPLE_SEGMENT|7700,7705|false|false|false|C3844350|Maybe|maybe
Event|Event|SIMPLE_SEGMENT|7716,7718|false|false|false|||up
Finding|Idea or Concept|SIMPLE_SEGMENT|7723,7731|false|false|false|C0750591|consider|consider
Event|Event|SIMPLE_SEGMENT|7740,7746|false|false|false|||workup
Event|Event|SIMPLE_SEGMENT|7753,7764|true|false|false|||improvement
Finding|Conceptual Entity|SIMPLE_SEGMENT|7753,7764|true|false|false|C2986411|Improvement|improvement
Finding|Body Substance|SIMPLE_SEGMENT|7766,7771|true|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Functional Concept|SIMPLE_SEGMENT|7766,7771|true|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Intellectual Product|SIMPLE_SEGMENT|7766,7771|true|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|7780,7788|true|false|false|C0233591|Twirling|spinning
Event|Event|SIMPLE_SEGMENT|7780,7788|true|false|false|||spinning
Event|Event|SIMPLE_SEGMENT|7789,7794|false|false|false|||urine
Finding|Body Substance|SIMPLE_SEGMENT|7789,7794|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Functional Concept|SIMPLE_SEGMENT|7789,7794|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Intellectual Product|SIMPLE_SEGMENT|7789,7794|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7796,7801|false|false|false|C0022646|Kidney|renal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7796,7801|false|false|false|C0042075|Urologic Diseases|renal
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7824,7835|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7824,7835|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|7824,7835|false|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|7824,7835|false|false|false|C4284232|Medications|medications
Event|Event|SIMPLE_SEGMENT|7847,7854|false|false|false|||CHRONIC
Finding|Intellectual Product|SIMPLE_SEGMENT|7847,7854|false|false|false|C1547296|Chronic - Admission Level of Care Code|CHRONIC
Procedure|Health Care Activity|SIMPLE_SEGMENT|7847,7854|false|false|false|C1555457|Provision of recurring care for chronic illness|CHRONIC
Event|Event|SIMPLE_SEGMENT|7865,7867|false|false|false|||HF
Drug|Antibiotic|SIMPLE_SEGMENT|7873,7876|false|false|false|C0030771|pefloxacin|pEF
Drug|Organic Chemical|SIMPLE_SEGMENT|7873,7876|false|false|false|C0030771|pefloxacin|pEF
Event|Event|SIMPLE_SEGMENT|7873,7876|false|false|false|||pEF
Finding|Finding|SIMPLE_SEGMENT|7873,7876|false|false|false|C1542834|Peak expiratory flow rate|pEF
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7877,7880|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7877,7880|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|7877,7880|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|7877,7880|false|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|7877,7880|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7877,7880|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|7877,7880|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7877,7880|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Event|Event|SIMPLE_SEGMENT|7885,7889|false|false|false|||CABG
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7885,7889|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Event|Event|SIMPLE_SEGMENT|7894,7900|false|false|false|||stents
Event|Activity|SIMPLE_SEGMENT|7920,7925|true|false|false|C5966184|Issue (action)|issue
Event|Event|SIMPLE_SEGMENT|7920,7925|true|false|false|||issue
Finding|Finding|SIMPLE_SEGMENT|7920,7925|true|false|false|C0033213;C1706387|Issue (document);Problem|issue
Finding|Intellectual Product|SIMPLE_SEGMENT|7920,7925|true|false|false|C0033213;C1706387|Issue (document);Problem|issue
Event|Event|SIMPLE_SEGMENT|7932,7941|true|false|false|||inpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|7932,7941|true|false|false|C1548438;C1549404|Patient Class - Inpatient;Referral category - Inpatient|inpatient
Procedure|Health Care Activity|SIMPLE_SEGMENT|7932,7941|true|false|false|C1555324|inpatient encounter|inpatient
Drug|Substance|SIMPLE_SEGMENT|7943,7948|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|Fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|7943,7948|false|false|false|C1546638|Fluid Specimen Code|Fluid
Event|Event|SIMPLE_SEGMENT|7949,7952|false|false|false|||use
Finding|Functional Concept|SIMPLE_SEGMENT|7949,7952|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|SIMPLE_SEGMENT|7949,7952|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Event|Event|SIMPLE_SEGMENT|7957,7966|false|false|false|||judicious
Event|Event|SIMPLE_SEGMENT|7978,7987|false|false|false|||converted
Event|Event|SIMPLE_SEGMENT|7998,8004|false|false|false|||acting
Drug|Organic Chemical|SIMPLE_SEGMENT|8021,8031|false|false|false|C0022251|isosorbide|isosorbide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8021,8031|false|false|false|C0022251|isosorbide|isosorbide
Event|Event|SIMPLE_SEGMENT|8021,8031|false|false|false|||isosorbide
Drug|Organic Chemical|SIMPLE_SEGMENT|8033,8040|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8033,8040|false|false|false|C0004057|aspirin|aspirin
Event|Event|SIMPLE_SEGMENT|8033,8040|false|false|false|||aspirin
Drug|Organic Chemical|SIMPLE_SEGMENT|8046,8058|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8046,8058|false|false|false|C0286651|atorvastatin|atorvastatin
Event|Event|SIMPLE_SEGMENT|8046,8058|false|false|false|||atorvastatin
Event|Event|SIMPLE_SEGMENT|8064,8073|false|false|false|||continued
Drug|Organic Chemical|SIMPLE_SEGMENT|8075,8083|false|false|false|C0126174|losartan|Losartan
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8075,8083|false|false|false|C0126174|losartan|Losartan
Event|Event|SIMPLE_SEGMENT|8084,8088|false|false|false|||held
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8103,8106|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|SIMPLE_SEGMENT|8103,8106|false|false|false|||HTN
Finding|Idea or Concept|SIMPLE_SEGMENT|8108,8112|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|8108,8112|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|8108,8112|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|8113,8123|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8113,8123|false|false|false|C0025859|metoprolol|metoprolol
Event|Event|SIMPLE_SEGMENT|8113,8123|false|false|false|||metoprolol
Drug|Organic Chemical|SIMPLE_SEGMENT|8128,8138|false|false|false|C0022251|isosorbide|isosorbide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8128,8138|false|false|false|C0022251|isosorbide|isosorbide
Event|Event|SIMPLE_SEGMENT|8128,8138|false|false|false|||isosorbide
Event|Event|SIMPLE_SEGMENT|8139,8148|false|false|false|||continued
Drug|Organic Chemical|SIMPLE_SEGMENT|8150,8158|false|false|false|C0126174|losartan|losartan
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8150,8158|false|false|false|C0126174|losartan|losartan
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8159,8163|false|false|false|C0675390|ARID1A protein, human|held
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8159,8163|false|false|false|C0675390|ARID1A protein, human|held
Event|Event|SIMPLE_SEGMENT|8159,8163|false|false|false|||held
Finding|Gene or Genome|SIMPLE_SEGMENT|8159,8163|false|false|false|C1948036;C2985160|ARID1A wt Allele;Held - activity status|held
Finding|Idea or Concept|SIMPLE_SEGMENT|8159,8163|false|false|false|C1948036;C2985160|ARID1A wt Allele;Held - activity status|held
Event|Event|SIMPLE_SEGMENT|8179,8188|false|false|false|||pressures
Finding|Finding|SIMPLE_SEGMENT|8179,8188|false|false|false|C0460139|Pressure (finding)|pressures
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|8179,8188|false|false|false|C0033095||pressures
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8194,8198|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|SIMPLE_SEGMENT|8194,8198|false|false|false|||soft
Event|Event|SIMPLE_SEGMENT|8217,8222|false|false|false|||range
Finding|Intellectual Product|SIMPLE_SEGMENT|8217,8222|false|false|false|C3542016|Concept model range (foundation metadata concept)|range
Event|Event|SIMPLE_SEGMENT|8236,8240|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|8236,8240|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|8236,8240|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|8236,8240|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|8245,8253|false|false|false|C0126174|losartan|losartan
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8245,8253|false|false|false|C0126174|losartan|losartan
Event|Event|SIMPLE_SEGMENT|8245,8253|false|false|false|||losartan
Finding|Sign or Symptom|SIMPLE_SEGMENT|8257,8265|false|false|false|C0085631;C3887611|Agitation;Restlessness|Restless
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8257,8269|false|false|false|C0035258|Restless Legs Syndrome|Restless leg
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8257,8278|false|false|false|C0035258|Restless Legs Syndrome|Restless leg syndrome
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8266,8269|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8270,8278|false|false|false|C0039082|Syndrome|syndrome
Event|Event|SIMPLE_SEGMENT|8270,8278|false|false|false|||syndrome
Finding|Idea or Concept|SIMPLE_SEGMENT|8280,8284|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|8280,8284|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|8280,8284|false|false|false|C1553498|home health encounter|home
Event|Event|SIMPLE_SEGMENT|8285,8295|false|false|false|||ropinarole
Event|Event|SIMPLE_SEGMENT|8296,8305|false|false|false|||continued
Anatomy|Body Location or Region|SIMPLE_SEGMENT|8308,8316|false|false|false|C0037004;C4299050|Shoulder;Upper extremity>Shoulder|Shoulder
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8308,8316|false|false|false|C0221590;C0869975|Examination of shoulder(s);Procedures on Shoulder|Shoulder
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8308,8316|false|false|false|C0221590;C0869975|Examination of shoulder(s);Procedures on Shoulder|Shoulder
Finding|Sign or Symptom|SIMPLE_SEGMENT|8308,8321|false|false|false|C0037011|Shoulder Pain|Shoulder pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8317,8321|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|8317,8321|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|8317,8321|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|8317,8321|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|SIMPLE_SEGMENT|8323,8332|false|false|false|C0030049|oxycodone|oxycodone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8323,8332|false|false|false|C0030049|oxycodone|oxycodone
Event|Event|SIMPLE_SEGMENT|8323,8332|false|false|false|||oxycodone
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8323,8332|false|false|false|C0524222|Oxycodone measurement|oxycodone
Drug|Organic Chemical|SIMPLE_SEGMENT|8337,8344|false|false|false|C0699142|Tylenol|tylenol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8337,8344|false|false|false|C0699142|Tylenol|tylenol
Event|Event|SIMPLE_SEGMENT|8337,8344|false|false|false|||tylenol
Event|Event|SIMPLE_SEGMENT|8356,8360|false|false|false|||dose
Event|Event|SIMPLE_SEGMENT|8368,8377|false|false|false|||inpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|8368,8377|false|false|false|C1548438;C1549404|Patient Class - Inpatient;Referral category - Inpatient|inpatient
Procedure|Health Care Activity|SIMPLE_SEGMENT|8368,8377|false|false|false|C1555324|inpatient encounter|inpatient
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8382,8386|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8382,8386|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|SIMPLE_SEGMENT|8382,8386|false|false|false|||COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|8382,8386|false|false|false|C1412502|ARCN1 gene|COPD
Event|Event|SIMPLE_SEGMENT|8388,8392|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|8388,8392|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|8388,8392|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|8388,8392|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|8393,8399|false|false|false|C0965130|Advair|advair
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8393,8399|false|false|false|C0965130|Advair|advair
Event|Event|SIMPLE_SEGMENT|8393,8399|false|false|false|||advair
Finding|Gene or Genome|SIMPLE_SEGMENT|8404,8407|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Organic Chemical|SIMPLE_SEGMENT|8408,8417|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8408,8417|false|false|false|C0001927|albuterol|albuterol
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8418,8422|false|false|false|C1300458|Nebulizer solution|nebs
Event|Event|SIMPLE_SEGMENT|8418,8422|false|false|false|||nebs
Event|Event|SIMPLE_SEGMENT|8428,8437|false|false|false|||continued
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8442,8446|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Event|Event|SIMPLE_SEGMENT|8442,8446|false|false|false|||GERD
Finding|Idea or Concept|SIMPLE_SEGMENT|8448,8452|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|8448,8452|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|8448,8452|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|8453,8465|false|false|false|C0081876|pantoprazole|pantoprazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8453,8465|false|false|false|C0081876|pantoprazole|pantoprazole
Event|Event|SIMPLE_SEGMENT|8453,8465|false|false|false|||pantoprazole
Event|Event|SIMPLE_SEGMENT|8466,8475|false|false|false|||continued
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8479,8487|false|false|false|C1950154|Insomnia homeopathic medication|Insomnia
Event|Event|SIMPLE_SEGMENT|8479,8487|false|false|false|||Insomnia
Finding|Sign or Symptom|SIMPLE_SEGMENT|8479,8487|false|false|false|C0917801|Sleeplessness|Insomnia
Event|Event|SIMPLE_SEGMENT|8489,8493|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|8489,8493|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|8489,8493|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|8489,8493|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|8494,8503|false|false|false|C0040805|trazodone|trazodone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8494,8503|false|false|false|C0040805|trazodone|trazodone
Event|Event|SIMPLE_SEGMENT|8494,8503|false|false|false|||trazodone
Event|Event|SIMPLE_SEGMENT|8504,8513|false|false|false|||continued
Finding|Idea or Concept|SIMPLE_SEGMENT|8517,8529|false|false|false|C1548597|Marketing basis - Transitional|TRANSITIONAL
Event|Event|SIMPLE_SEGMENT|8530,8536|false|false|false|||ISSUES
Drug|Organic Chemical|SIMPLE_SEGMENT|8540,8548|false|false|false|C0126174|losartan|Losartan
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8540,8548|false|false|false|C0126174|losartan|Losartan
Event|Event|SIMPLE_SEGMENT|8554,8563|false|false|false|||inpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|8554,8563|false|false|false|C1548438;C1549404|Patient Class - Inpatient;Referral category - Inpatient|inpatient
Procedure|Health Care Activity|SIMPLE_SEGMENT|8554,8563|false|false|false|C1555324|inpatient encounter|inpatient
Finding|Body Substance|SIMPLE_SEGMENT|8571,8580|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|8571,8580|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|8571,8580|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|8571,8580|false|false|false|C0030685|Patient Discharge|discharge
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8592,8597|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|8592,8597|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|8592,8597|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Event|Event|SIMPLE_SEGMENT|8599,8608|false|false|false|||pressures
Finding|Finding|SIMPLE_SEGMENT|8599,8608|false|false|false|C0460139|Pressure (finding)|pressures
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|8599,8608|false|false|false|C0033095||pressures
Event|Event|SIMPLE_SEGMENT|8614,8617|false|false|false|||low
Finding|Finding|SIMPLE_SEGMENT|8614,8617|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|SIMPLE_SEGMENT|8614,8617|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Event|Event|SIMPLE_SEGMENT|8618,8624|false|false|false|||normal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8626,8629|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|8626,8629|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|8626,8629|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8626,8629|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|SIMPLE_SEGMENT|8626,8629|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|8626,8629|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|SIMPLE_SEGMENT|8626,8629|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8626,8629|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|SIMPLE_SEGMENT|8626,8629|false|false|false|||PCP
Finding|Gene or Genome|SIMPLE_SEGMENT|8626,8629|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|SIMPLE_SEGMENT|8626,8629|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Event|SIMPLE_SEGMENT|8643,8650|false|false|false|||restart
Finding|Body Substance|SIMPLE_SEGMENT|8654,8661|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|8654,8661|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|8654,8661|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|8665,8671|false|false|false|||follow
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8680,8683|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|8680,8683|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|8680,8683|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8680,8683|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|SIMPLE_SEGMENT|8680,8683|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|8680,8683|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|SIMPLE_SEGMENT|8680,8683|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8680,8683|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|SIMPLE_SEGMENT|8680,8683|false|false|false|||PCP
Finding|Gene or Genome|SIMPLE_SEGMENT|8680,8683|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|SIMPLE_SEGMENT|8680,8683|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Event|SIMPLE_SEGMENT|8688,8698|false|false|false|||resolution
Finding|Conceptual Entity|SIMPLE_SEGMENT|8688,8698|false|false|false|C1514893;C2699488|Resolution;physiologic resolution|resolution
Finding|Pathologic Function|SIMPLE_SEGMENT|8688,8698|false|false|false|C1514893;C2699488|Resolution;physiologic resolution|resolution
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8702,8705|false|false|false|C0042029|Urinary tract infection|UTI
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8702,8705|false|false|false|C0077906|urinastatin|UTI
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8702,8705|false|false|false|C0077906|urinastatin|UTI
Event|Event|SIMPLE_SEGMENT|8702,8705|false|false|false|||UTI
Finding|Gene or Genome|SIMPLE_SEGMENT|8702,8705|false|false|false|C1412376;C5780748|AMBP gene;AMBP wt Allele|UTI
Event|Event|SIMPLE_SEGMENT|8710,8714|false|false|false|||back
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8716,8720|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|8716,8720|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|8716,8720|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|8716,8729|false|false|false|C0030193|Pain|pain symptoms
Event|Event|SIMPLE_SEGMENT|8721,8729|false|false|false|||symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|8721,8729|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|8721,8729|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Body Substance|SIMPLE_SEGMENT|8732,8739|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|8732,8739|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|8732,8739|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8752,8759|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|SIMPLE_SEGMENT|8752,8759|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8752,8759|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|SIMPLE_SEGMENT|8752,8759|false|false|false|||insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|8752,8759|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8752,8759|false|false|false|C0202098|Insulin measurement|insulin
Event|Event|SIMPLE_SEGMENT|8769,8780|true|false|false|||adjustments
Finding|Functional Concept|SIMPLE_SEGMENT|8769,8780|true|false|false|C0456081||adjustments
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8769,8780|true|false|false|C2945673|Clinical adjustment|adjustments
Event|Event|SIMPLE_SEGMENT|8785,8792|true|false|false|||optimal
Finding|Intellectual Product|SIMPLE_SEGMENT|8785,8792|true|false|false|C3260738|Outpatient Physical Therapy Improvement in Movement and Assessment Log (OPTIMAL) Survey|optimal
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8794,8810|true|false|false|C5392125|Glycemic Control|glycemic control
Drug|Organic Chemical|SIMPLE_SEGMENT|8803,8810|true|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8803,8810|true|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Substance|SIMPLE_SEGMENT|8803,8810|true|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Event|Event|SIMPLE_SEGMENT|8803,8810|true|false|false|||control
Finding|Conceptual Entity|SIMPLE_SEGMENT|8803,8810|true|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Functional Concept|SIMPLE_SEGMENT|8803,8810|true|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Idea or Concept|SIMPLE_SEGMENT|8803,8810|true|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Event|Event|SIMPLE_SEGMENT|8816,8823|true|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|8816,8823|true|false|false|C0392747|Changing|changes
Event|Event|SIMPLE_SEGMENT|8827,8834|true|false|false|||regimen
Finding|Intellectual Product|SIMPLE_SEGMENT|8827,8834|true|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8827,8834|true|false|false|C0040808|Treatment Protocols|regimen
Event|Event|SIMPLE_SEGMENT|8840,8844|true|false|false|||made
Event|Event|SIMPLE_SEGMENT|8848,8857|true|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|8848,8857|true|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|8848,8857|true|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|8848,8857|true|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|8848,8857|true|false|false|C0030685|Patient Discharge|discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8861,8872|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8861,8872|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|8861,8872|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|8861,8872|false|false|false|C4284232|Medications|Medications
Finding|Finding|SIMPLE_SEGMENT|8861,8885|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|SIMPLE_SEGMENT|8876,8885|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|8876,8885|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8904,8914|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|8904,8914|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|8904,8919|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|SIMPLE_SEGMENT|8915,8919|false|false|false|||list
Finding|Intellectual Product|SIMPLE_SEGMENT|8915,8919|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|SIMPLE_SEGMENT|8927,8937|false|false|false|||inaccurate
Event|Event|SIMPLE_SEGMENT|8942,8950|false|false|false|||requires
Event|Event|SIMPLE_SEGMENT|8959,8972|false|false|false|||investigation
Finding|Intellectual Product|SIMPLE_SEGMENT|8959,8972|false|false|false|C1552578|Act Class - investigation|investigation
Procedure|Health Care Activity|SIMPLE_SEGMENT|8959,8972|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|investigation
Drug|Organic Chemical|SIMPLE_SEGMENT|8977,8985|false|false|false|C0126174|losartan|Losartan
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8977,8985|false|false|false|C0126174|losartan|Losartan
Event|Event|SIMPLE_SEGMENT|8977,8985|false|false|false|||Losartan
Drug|Organic Chemical|SIMPLE_SEGMENT|8977,8995|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8977,8995|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8986,8995|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|8986,8995|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Food|SIMPLE_SEGMENT|8986,8995|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|8986,8995|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8986,8995|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Event|Event|SIMPLE_SEGMENT|8986,8995|false|false|false|||Potassium
Finding|Physiologic Function|SIMPLE_SEGMENT|8986,8995|false|false|false|C4553027|Potassium metabolic function|Potassium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8986,8995|false|false|false|C0202194|Potassium measurement|Potassium
Drug|Organic Chemical|SIMPLE_SEGMENT|9015,9025|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9015,9025|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Organic Chemical|SIMPLE_SEGMENT|9015,9035|false|false|false|C0724633|metoprolol succinate|Metoprolol Succinate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9015,9035|false|false|false|C0724633|metoprolol succinate|Metoprolol Succinate
Drug|Organic Chemical|SIMPLE_SEGMENT|9026,9035|false|false|false|C0038617;C0220918|Succinates;succinate|Succinate
Event|Event|SIMPLE_SEGMENT|9026,9035|false|false|false|||Succinate
Drug|Organic Chemical|SIMPLE_SEGMENT|9059,9071|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9059,9071|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|SIMPLE_SEGMENT|9088,9098|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9088,9098|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Organic Chemical|SIMPLE_SEGMENT|9088,9110|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9088,9110|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Event|Event|SIMPLE_SEGMENT|9099,9110|false|false|false|||Mononitrate
Finding|Finding|SIMPLE_SEGMENT|9112,9120|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|SIMPLE_SEGMENT|9112,9120|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|SIMPLE_SEGMENT|9121,9128|false|false|false|||Release
Finding|Functional Concept|SIMPLE_SEGMENT|9121,9128|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|9121,9128|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9121,9128|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|SIMPLE_SEGMENT|9150,9163|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9150,9163|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Event|Event|SIMPLE_SEGMENT|9150,9163|false|false|false|||Nitroglycerin
Finding|Gene or Genome|SIMPLE_SEGMENT|9183,9186|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9187,9191|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|9187,9191|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|9187,9191|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|9187,9191|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|SIMPLE_SEGMENT|9196,9206|false|false|false|C0244821|ropinirole|Ropinirole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9196,9206|false|false|false|C0244821|ropinirole|Ropinirole
Event|Event|SIMPLE_SEGMENT|9217,9220|false|false|false|||QPM
Drug|Organic Chemical|SIMPLE_SEGMENT|9225,9234|false|false|false|C0030049|oxycodone|Oxycodone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9225,9234|false|false|false|C0030049|oxycodone|Oxycodone
Event|Event|SIMPLE_SEGMENT|9225,9234|false|false|false|||Oxycodone
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9225,9234|false|false|false|C0524222|Oxycodone measurement|Oxycodone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9225,9248|false|false|false|C0717368|acetaminophen / oxycodone|Oxycodone-Acetaminophen
Drug|Organic Chemical|SIMPLE_SEGMENT|9235,9248|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9235,9248|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|SIMPLE_SEGMENT|9235,9248|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9235,9248|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9263,9266|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|SIMPLE_SEGMENT|9263,9266|false|false|false|||TAB
Event|Event|SIMPLE_SEGMENT|9270,9273|false|false|false|||Q8H
Finding|Gene or Genome|SIMPLE_SEGMENT|9274,9277|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9278,9282|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|9278,9282|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|9278,9282|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|9278,9282|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|SIMPLE_SEGMENT|9287,9298|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9287,9298|false|false|false|C0082607|fluticasone|Fluticasone
Event|Event|SIMPLE_SEGMENT|9287,9298|false|false|false|||Fluticasone
Drug|Organic Chemical|SIMPLE_SEGMENT|9287,9309|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9287,9309|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Organic Chemical|SIMPLE_SEGMENT|9299,9309|false|false|false|C0033474;C0392214|Propionates;propionate|Propionate
Event|Event|SIMPLE_SEGMENT|9319,9323|false|false|false|||PUFF
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|9327,9330|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9327,9330|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9327,9330|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|9327,9330|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|9327,9330|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|9335,9347|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9335,9347|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Organic Chemical|SIMPLE_SEGMENT|9367,9374|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9367,9374|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|SIMPLE_SEGMENT|9396,9405|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9396,9405|false|false|false|C0001927|albuterol|albuterol
Event|Event|SIMPLE_SEGMENT|9396,9405|false|false|false|||albuterol
Drug|Organic Chemical|SIMPLE_SEGMENT|9396,9413|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9396,9413|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|9406,9413|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Inorganic Chemical|SIMPLE_SEGMENT|9406,9413|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9406,9413|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Event|Event|SIMPLE_SEGMENT|9406,9413|false|false|false|||sulfate
Finding|Functional Concept|SIMPLE_SEGMENT|9431,9441|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Finding|Organism Function|SIMPLE_SEGMENT|9431,9441|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Event|Event|SIMPLE_SEGMENT|9442,9447|false|false|false|||q4hrs
Event|Event|SIMPLE_SEGMENT|9448,9456|false|false|false|||wheezing
Finding|Sign or Symptom|SIMPLE_SEGMENT|9448,9456|false|false|false|C0043144|Wheezing|wheezing
Drug|Organic Chemical|SIMPLE_SEGMENT|9463,9472|false|false|false|C0040805|trazodone|TraZODone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9463,9472|false|false|false|C0040805|trazodone|TraZODone
Drug|Organic Chemical|SIMPLE_SEGMENT|9491,9498|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9491,9498|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|SIMPLE_SEGMENT|9491,9498|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|SIMPLE_SEGMENT|9491,9500|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|SIMPLE_SEGMENT|9491,9500|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9491,9500|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|SIMPLE_SEGMENT|9491,9500|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9491,9500|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Event|Event|SIMPLE_SEGMENT|9506,9510|false|false|false|||UNIT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9525,9532|false|false|false|C1314782|Levemir|Levemir
Drug|Hormone|SIMPLE_SEGMENT|9525,9532|false|false|false|C1314782|Levemir|Levemir
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9525,9532|false|false|false|C1314782|Levemir|Levemir
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9542,9549|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|SIMPLE_SEGMENT|9542,9549|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9542,9549|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|SIMPLE_SEGMENT|9542,9549|false|false|false|||insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|9542,9549|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9542,9549|false|false|false|C0202098|Insulin measurement|insulin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9542,9557|false|false|false|C0537270|insulin detemir|insulin detemir
Drug|Hormone|SIMPLE_SEGMENT|9542,9557|false|false|false|C0537270|insulin detemir|insulin detemir
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9542,9557|false|false|false|C0537270|insulin detemir|insulin detemir
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9550,9557|false|false|false|C0537270|insulin detemir|detemir
Drug|Hormone|SIMPLE_SEGMENT|9550,9557|false|false|false|C0537270|insulin detemir|detemir
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9550,9557|false|false|false|C0537270|insulin detemir|detemir
Event|Event|SIMPLE_SEGMENT|9550,9557|false|false|false|||detemir
Finding|Functional Concept|SIMPLE_SEGMENT|9568,9580|false|false|false|C1522438|Subcutaneous Route of Administration|subcutaneous
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9602,9609|false|false|false|C0528249|Humalog|HumaLOG
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9602,9609|false|false|false|C0528249|Humalog|HumaLOG
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9619,9626|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|SIMPLE_SEGMENT|9619,9626|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9619,9626|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|SIMPLE_SEGMENT|9619,9626|false|false|false|||insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|9619,9626|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9619,9626|false|false|false|C0202098|Insulin measurement|insulin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9619,9633|false|false|false|C0293359|insulin lispro|insulin lispro
Drug|Hormone|SIMPLE_SEGMENT|9619,9633|false|false|false|C0293359|insulin lispro|insulin lispro
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9619,9633|false|false|false|C0293359|insulin lispro|insulin lispro
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9627,9633|false|false|false|C0293359|insulin lispro|lispro
Drug|Hormone|SIMPLE_SEGMENT|9627,9633|false|false|false|C0293359|insulin lispro|lispro
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9627,9633|false|false|false|C0293359|insulin lispro|lispro
Event|Event|SIMPLE_SEGMENT|9627,9633|false|false|false|||lispro
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9647,9652|false|false|false|C0222045|Integumentary scale|scale
Event|Activity|SIMPLE_SEGMENT|9647,9652|false|false|false|C1947916|Scaling|scale
Finding|Conceptual Entity|SIMPLE_SEGMENT|9647,9652|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|scale
Finding|Intellectual Product|SIMPLE_SEGMENT|9647,9652|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|scale
Event|Event|SIMPLE_SEGMENT|9655,9667|false|false|false|||subcutaneous
Finding|Functional Concept|SIMPLE_SEGMENT|9655,9667|false|false|false|C1522438|Subcutaneous Route of Administration|subcutaneous
Event|Event|SIMPLE_SEGMENT|9671,9679|false|false|false|||directed
Event|Event|SIMPLE_SEGMENT|9684,9693|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|9684,9693|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|9684,9693|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|9684,9693|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|9684,9693|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|9684,9705|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9694,9705|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9694,9705|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|9694,9705|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|9694,9705|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|SIMPLE_SEGMENT|9710,9719|false|false|false|C0030049|oxycodone|Oxycodone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9710,9719|false|false|false|C0030049|oxycodone|Oxycodone
Event|Event|SIMPLE_SEGMENT|9710,9719|false|false|false|||Oxycodone
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9710,9719|false|false|false|C0524222|Oxycodone measurement|Oxycodone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9710,9733|false|false|false|C0717368|acetaminophen / oxycodone|Oxycodone-Acetaminophen
Drug|Organic Chemical|SIMPLE_SEGMENT|9720,9733|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9720,9733|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|SIMPLE_SEGMENT|9720,9733|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9720,9733|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9748,9751|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|SIMPLE_SEGMENT|9748,9751|false|false|false|||TAB
Event|Event|SIMPLE_SEGMENT|9755,9758|false|false|false|||Q8H
Finding|Gene or Genome|SIMPLE_SEGMENT|9759,9762|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9763,9767|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|9763,9767|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|9763,9767|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|9763,9767|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|SIMPLE_SEGMENT|9772,9785|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9772,9785|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Event|Event|SIMPLE_SEGMENT|9772,9785|false|false|false|||Nitroglycerin
Finding|Gene or Genome|SIMPLE_SEGMENT|9805,9808|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9809,9813|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|9809,9813|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|9809,9813|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|9809,9813|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|SIMPLE_SEGMENT|9818,9828|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9818,9828|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Organic Chemical|SIMPLE_SEGMENT|9818,9838|false|false|false|C0724633|metoprolol succinate|Metoprolol Succinate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9818,9838|false|false|false|C0724633|metoprolol succinate|Metoprolol Succinate
Drug|Organic Chemical|SIMPLE_SEGMENT|9829,9838|false|false|false|C0038617;C0220918|Succinates;succinate|Succinate
Event|Event|SIMPLE_SEGMENT|9829,9838|false|false|false|||Succinate
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9862,9869|false|false|false|C1314782|Levemir|Levemir
Drug|Hormone|SIMPLE_SEGMENT|9862,9869|false|false|false|C1314782|Levemir|Levemir
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9862,9869|false|false|false|C1314782|Levemir|Levemir
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9879,9886|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|SIMPLE_SEGMENT|9879,9886|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9879,9886|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|SIMPLE_SEGMENT|9879,9886|false|false|false|||insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|9879,9886|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9879,9886|false|false|false|C0202098|Insulin measurement|insulin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9879,9894|false|false|false|C0537270|insulin detemir|insulin detemir
Drug|Hormone|SIMPLE_SEGMENT|9879,9894|false|false|false|C0537270|insulin detemir|insulin detemir
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9879,9894|false|false|false|C0537270|insulin detemir|insulin detemir
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9887,9894|false|false|false|C0537270|insulin detemir|detemir
Drug|Hormone|SIMPLE_SEGMENT|9887,9894|false|false|false|C0537270|insulin detemir|detemir
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9887,9894|false|false|false|C0537270|insulin detemir|detemir
Event|Event|SIMPLE_SEGMENT|9887,9894|false|false|false|||detemir
Finding|Functional Concept|SIMPLE_SEGMENT|9905,9917|false|false|false|C1522438|Subcutaneous Route of Administration|subcutaneous
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9938,9945|false|false|false|C0528249|Humalog|HumaLOG
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9938,9945|false|false|false|C0528249|Humalog|HumaLOG
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9955,9962|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|SIMPLE_SEGMENT|9955,9962|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9955,9962|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|SIMPLE_SEGMENT|9955,9962|false|false|false|||insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|9955,9962|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9955,9962|false|false|false|C0202098|Insulin measurement|insulin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9955,9969|false|false|false|C0293359|insulin lispro|insulin lispro
Drug|Hormone|SIMPLE_SEGMENT|9955,9969|false|false|false|C0293359|insulin lispro|insulin lispro
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9955,9969|false|false|false|C0293359|insulin lispro|insulin lispro
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9963,9969|false|false|false|C0293359|insulin lispro|lispro
Drug|Hormone|SIMPLE_SEGMENT|9963,9969|false|false|false|C0293359|insulin lispro|lispro
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9963,9969|false|false|false|C0293359|insulin lispro|lispro
Event|Event|SIMPLE_SEGMENT|9963,9969|false|false|false|||lispro
Event|Event|SIMPLE_SEGMENT|9975,9987|false|false|false|||SUBCUTANEOUS
Finding|Functional Concept|SIMPLE_SEGMENT|9975,9987|false|false|false|C1522438|Subcutaneous Route of Administration|SUBCUTANEOUS
Event|Event|SIMPLE_SEGMENT|9991,9999|false|false|false|||DIRECTED
Drug|Organic Chemical|SIMPLE_SEGMENT|10005,10014|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10005,10014|false|false|false|C0001927|albuterol|albuterol
Event|Event|SIMPLE_SEGMENT|10005,10014|false|false|false|||albuterol
Drug|Organic Chemical|SIMPLE_SEGMENT|10005,10022|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10005,10022|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|10015,10022|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Inorganic Chemical|SIMPLE_SEGMENT|10015,10022|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10015,10022|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Event|Event|SIMPLE_SEGMENT|10015,10022|false|false|false|||sulfate
Finding|Functional Concept|SIMPLE_SEGMENT|10040,10050|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Finding|Organism Function|SIMPLE_SEGMENT|10040,10050|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Event|Event|SIMPLE_SEGMENT|10051,10056|false|false|false|||q4hrs
Event|Event|SIMPLE_SEGMENT|10057,10065|false|false|false|||wheezing
Finding|Sign or Symptom|SIMPLE_SEGMENT|10057,10065|false|false|false|C0043144|Wheezing|wheezing
Drug|Organic Chemical|SIMPLE_SEGMENT|10070,10083|false|false|false|C0008809|ciprofloxacin|Ciprofloxacin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10070,10083|false|false|false|C0008809|ciprofloxacin|Ciprofloxacin
Drug|Antibiotic|SIMPLE_SEGMENT|10070,10087|false|false|false|C0282104|ciprofloxacin hydrochloride|Ciprofloxacin HCl
Drug|Organic Chemical|SIMPLE_SEGMENT|10070,10087|false|false|false|C0282104|ciprofloxacin hydrochloride|Ciprofloxacin HCl
Disorder|Neoplastic Process|SIMPLE_SEGMENT|10084,10087|false|false|false|C0023443|Hairy Cell Leukemia|HCl
Drug|Immunologic Factor|SIMPLE_SEGMENT|10084,10087|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Inorganic Chemical|SIMPLE_SEGMENT|10084,10087|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10084,10087|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Event|Event|SIMPLE_SEGMENT|10084,10087|false|false|false|||HCl
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10103,10111|false|false|false|C0720099|Duration brand of oxymetazoline|Duration
Event|Event|SIMPLE_SEGMENT|10103,10111|false|false|false|||Duration
Event|Event|SIMPLE_SEGMENT|10121,10123|false|false|false|||RX
Drug|Organic Chemical|SIMPLE_SEGMENT|10125,10138|false|false|false|C0008809|ciprofloxacin|ciprofloxacin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10125,10138|false|false|false|C0008809|ciprofloxacin|ciprofloxacin
Drug|Organic Chemical|SIMPLE_SEGMENT|10140,10145|false|false|false|C0701042|Cipro|Cipro
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10140,10145|false|false|false|C0701042|Cipro|Cipro
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10156,10162|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|SIMPLE_SEGMENT|10166,10174|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|10169,10174|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|10169,10174|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Idea or Concept|SIMPLE_SEGMENT|10184,10187|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|10184,10187|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10198,10204|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|10205,10212|false|false|false|||Refills
Finding|Idea or Concept|SIMPLE_SEGMENT|10205,10212|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|10219,10226|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10219,10226|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|SIMPLE_SEGMENT|10219,10226|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|SIMPLE_SEGMENT|10219,10228|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|SIMPLE_SEGMENT|10219,10228|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10219,10228|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|SIMPLE_SEGMENT|10219,10228|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10219,10228|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Event|Event|SIMPLE_SEGMENT|10227,10228|false|false|false|||D
Event|Event|SIMPLE_SEGMENT|10234,10238|false|false|false|||UNIT
Drug|Organic Chemical|SIMPLE_SEGMENT|10252,10261|false|false|false|C0040805|trazodone|TraZODone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10252,10261|false|false|false|C0040805|trazodone|TraZODone
Drug|Organic Chemical|SIMPLE_SEGMENT|10280,10290|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10280,10290|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Organic Chemical|SIMPLE_SEGMENT|10280,10302|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10280,10302|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Event|Event|SIMPLE_SEGMENT|10291,10302|false|false|false|||Mononitrate
Finding|Finding|SIMPLE_SEGMENT|10304,10312|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|SIMPLE_SEGMENT|10304,10312|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|SIMPLE_SEGMENT|10313,10320|false|false|false|||Release
Finding|Functional Concept|SIMPLE_SEGMENT|10313,10320|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|10313,10320|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10313,10320|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|SIMPLE_SEGMENT|10343,10350|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10343,10350|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|SIMPLE_SEGMENT|10372,10384|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10372,10384|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|SIMPLE_SEGMENT|10402,10413|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10402,10413|false|false|false|C0082607|fluticasone|Fluticasone
Event|Event|SIMPLE_SEGMENT|10402,10413|false|false|false|||Fluticasone
Drug|Organic Chemical|SIMPLE_SEGMENT|10402,10424|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10402,10424|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Organic Chemical|SIMPLE_SEGMENT|10414,10424|false|false|false|C0033474;C0392214|Propionates;propionate|Propionate
Event|Event|SIMPLE_SEGMENT|10434,10438|false|false|false|||PUFF
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|10442,10445|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10442,10445|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|10442,10445|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|10442,10445|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|10442,10445|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|10451,10463|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10451,10463|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Organic Chemical|SIMPLE_SEGMENT|10483,10493|false|false|false|C0244821|ropinirole|Ropinirole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10483,10493|false|false|false|C0244821|ropinirole|Ropinirole
Event|Event|SIMPLE_SEGMENT|10504,10507|false|false|false|||QPM
Event|Event|SIMPLE_SEGMENT|10512,10521|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|10512,10521|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|10512,10521|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|10512,10521|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|10512,10521|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10512,10533|false|false|false|C4019243||Discharge Disposition
Finding|Finding|SIMPLE_SEGMENT|10512,10533|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10522,10533|false|false|false|C2926604||Disposition
Event|Event|SIMPLE_SEGMENT|10522,10533|false|false|false|||Disposition
Procedure|Health Care Activity|SIMPLE_SEGMENT|10522,10533|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|SIMPLE_SEGMENT|10535,10539|false|false|false|||Home
Finding|Idea or Concept|SIMPLE_SEGMENT|10535,10539|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|SIMPLE_SEGMENT|10535,10539|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|SIMPLE_SEGMENT|10535,10539|false|false|false|C1553498|home health encounter|Home
Event|Event|SIMPLE_SEGMENT|10542,10551|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|10542,10551|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|10542,10551|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|10542,10551|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|10542,10551|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|10542,10561|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10552,10561|false|false|false|C0945731||Diagnosis
Event|Event|SIMPLE_SEGMENT|10552,10561|false|false|false|||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|10552,10561|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|10552,10561|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10552,10561|false|false|false|C0011900|Diagnosis|Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10563,10580|false|false|false|C0801658||Primary Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10571,10580|false|false|false|C0945731||Diagnosis
Event|Event|SIMPLE_SEGMENT|10571,10580|false|false|false|||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|10571,10580|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|10571,10580|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10571,10580|false|false|false|C0011900|Diagnosis|Diagnosis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10582,10585|false|false|false|C0042029|Urinary tract infection|UTI
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10582,10585|false|false|false|C0077906|urinastatin|UTI
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10582,10585|false|false|false|C0077906|urinastatin|UTI
Event|Event|SIMPLE_SEGMENT|10582,10585|false|false|false|||UTI
Finding|Gene or Genome|SIMPLE_SEGMENT|10582,10585|false|false|false|C1412376;C5780748|AMBP gene;AMBP wt Allele|UTI
Disorder|Neoplastic Process|SIMPLE_SEGMENT|10587,10596|false|false|false|C0027627|Neoplasm Metastasis|Secondary
Event|Event|SIMPLE_SEGMENT|10587,10596|false|false|false|||Secondary
Finding|Functional Concept|SIMPLE_SEGMENT|10587,10596|false|false|false|C1522484|metastatic qualifier|Secondary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10587,10606|false|false|false|C4255018||Secondary Diagnosis
Finding|Finding|SIMPLE_SEGMENT|10587,10606|false|false|false|C0332138|Secondary diagnosis|Secondary Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10597,10606|false|false|false|C0945731||Diagnosis
Event|Event|SIMPLE_SEGMENT|10597,10606|false|false|false|||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|10597,10606|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|10597,10606|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10597,10606|false|false|false|C0011900|Diagnosis|Diagnosis
Finding|Sign or Symptom|SIMPLE_SEGMENT|10608,10617|false|true|false|C0004604|Back Pain|Back Pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10613,10617|false|false|false|C2598155||Pain
Event|Event|SIMPLE_SEGMENT|10613,10617|false|false|false|||Pain
Finding|Functional Concept|SIMPLE_SEGMENT|10613,10617|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|10613,10617|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10618,10626|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|Diabetes
Event|Event|SIMPLE_SEGMENT|10618,10626|false|false|false|||Diabetes
Event|Event|SIMPLE_SEGMENT|10630,10639|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|10630,10639|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|10630,10639|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|10630,10639|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|10630,10639|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10640,10649|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10640,10649|false|false|false|C0012634|Disease|Condition
Event|Event|SIMPLE_SEGMENT|10640,10649|false|false|false|||Condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|10640,10649|false|false|false|C1705253|Logical Condition|Condition
Finding|Mental Process|SIMPLE_SEGMENT|10651,10657|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10651,10664|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|SIMPLE_SEGMENT|10651,10664|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10658,10664|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|10658,10664|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|10666,10671|false|false|false|||Clear
Finding|Idea or Concept|SIMPLE_SEGMENT|10666,10671|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|SIMPLE_SEGMENT|10676,10684|false|false|false|||coherent
Finding|Finding|SIMPLE_SEGMENT|10676,10684|false|false|false|C4068804|Coherent|coherent
Event|Event|SIMPLE_SEGMENT|10686,10691|false|false|false|||Level
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10686,10708|false|false|false|C4050479||Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|10686,10708|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|SIMPLE_SEGMENT|10695,10708|false|false|false|||Consciousness
Finding|Finding|SIMPLE_SEGMENT|10695,10708|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|SIMPLE_SEGMENT|10695,10708|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10710,10715|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|10710,10715|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10710,10715|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|SIMPLE_SEGMENT|10710,10715|false|false|false|||Alert
Finding|Finding|SIMPLE_SEGMENT|10710,10715|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|10710,10715|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|10710,10715|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|SIMPLE_SEGMENT|10720,10731|false|false|false|||interactive
Finding|Functional Concept|SIMPLE_SEGMENT|10720,10731|false|false|false|C1704675|Interaction|interactive
Event|Activity|SIMPLE_SEGMENT|10733,10741|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|10733,10741|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|SIMPLE_SEGMENT|10733,10741|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10742,10748|false|false|false|C5889824||Status
Event|Event|SIMPLE_SEGMENT|10742,10748|false|false|false|||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|10742,10748|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|10750,10760|false|false|false|||Ambulatory
Finding|Functional Concept|SIMPLE_SEGMENT|10750,10760|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|SIMPLE_SEGMENT|10750,10760|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|SIMPLE_SEGMENT|10750,10760|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|SIMPLE_SEGMENT|10750,10760|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|SIMPLE_SEGMENT|10763,10774|false|false|false|||Independent
Finding|Finding|SIMPLE_SEGMENT|10763,10774|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|SIMPLE_SEGMENT|10763,10774|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Event|Event|SIMPLE_SEGMENT|10779,10788|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|10779,10788|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|10779,10788|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|10779,10788|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|10779,10788|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10779,10801|false|false|false|C3669312||Discharge Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|10779,10801|false|false|false|C4282220|Discharge instructions|Discharge Instructions
Procedure|Health Care Activity|SIMPLE_SEGMENT|10779,10801|false|false|false|C2266673|hospital discharge instructions (treatment)|Discharge Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10789,10801|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|10789,10801|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|10789,10801|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Finding|Gene or Genome|SIMPLE_SEGMENT|10803,10807|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Event|Event|SIMPLE_SEGMENT|10823,10827|false|false|false|||seen
Finding|Finding|SIMPLE_SEGMENT|10835,10844|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Idea or Concept|SIMPLE_SEGMENT|10835,10844|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Intellectual Product|SIMPLE_SEGMENT|10835,10844|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Pathologic Function|SIMPLE_SEGMENT|10835,10844|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|10835,10844|false|false|false|C0013956|Emergency Situation|emergency
Procedure|Health Care Activity|SIMPLE_SEGMENT|10835,10844|false|false|false|C1553500|emergency encounter|emergency
Event|Event|SIMPLE_SEGMENT|10845,10855|false|false|false|||department
Finding|Idea or Concept|SIMPLE_SEGMENT|10845,10855|false|false|false|C1547537;C1548283;C1549615|Department - Charge type;Department - No suggested values defined;Organization Unit Type - Department|department
Finding|Sign or Symptom|SIMPLE_SEGMENT|10860,10869|false|true|false|C0004604|Back Pain|back pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10865,10869|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|10865,10869|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|10865,10869|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|10865,10869|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|10881,10889|false|false|false|||admitted
Finding|Idea or Concept|SIMPLE_SEGMENT|10897,10905|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|SIMPLE_SEGMENT|10926,10935|false|false|false|||diagnosed
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10944,10951|false|false|false|C0042027|Urinary tract|urinary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10944,10957|false|false|false|C0042027;C1508753|Urinary system;Urinary tract|urinary tract
Anatomy|Body System|SIMPLE_SEGMENT|10944,10957|false|false|false|C0042027;C1508753|Urinary system;Urinary tract|urinary tract
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10944,10967|false|false|false|C0042029|Urinary tract infection|urinary tract infection
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10952,10957|false|false|false|C1185740|Tract|tract
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10958,10967|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|SIMPLE_SEGMENT|10958,10967|false|false|false|||infection
Finding|Pathologic Function|SIMPLE_SEGMENT|10958,10967|false|false|false|C3714514|Infection|infection
Event|Event|SIMPLE_SEGMENT|10978,10985|false|false|false|||treated
Drug|Antibiotic|SIMPLE_SEGMENT|10991,11002|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|SIMPLE_SEGMENT|10991,11002|false|false|false|||antibiotics
Drug|Substance|SIMPLE_SEGMENT|11008,11014|false|false|false|C0302908|Liquid substance|fluids
Event|Event|SIMPLE_SEGMENT|11008,11014|false|false|false|||fluids
Finding|Body Substance|SIMPLE_SEGMENT|11008,11014|false|false|false|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11008,11014|false|false|false|C0016286|Fluid Therapy|fluids
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11019,11023|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|11019,11023|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|11019,11023|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|11019,11023|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11024,11034|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|11024,11034|false|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|11024,11034|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|SIMPLE_SEGMENT|11047,11054|false|false|false|||concern
Finding|Idea or Concept|SIMPLE_SEGMENT|11047,11054|false|false|false|C2699424|Concern|concern
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11069,11073|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|11069,11073|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|11069,11073|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|11069,11073|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|11077,11084|false|false|false|C0040405|X-Ray Computed Tomography|CT scan
Event|Event|SIMPLE_SEGMENT|11080,11084|false|false|false|||scan
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|11080,11084|false|false|false|C0034606;C0441633|Radionuclide Imaging;Scanning|scan
Event|Event|SIMPLE_SEGMENT|11113,11123|true|false|false|||determined
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11149,11155|true|false|false|C0022646;C0227665|Both kidneys;Kidney|kidney
Disorder|Neoplastic Process|SIMPLE_SEGMENT|11149,11155|true|false|false|C0496892;C0496927|Benign neoplasm of kidney;Neoplasm of uncertain or unknown behavior of kidney|kidney
Finding|Sign or Symptom|SIMPLE_SEGMENT|11149,11155|true|false|false|C0812426|Kidney problem|kidney
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|11149,11155|true|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11149,11155|true|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11149,11161|true|false|false|C0392525|Nephrolithiasis|kidney stone
Finding|Body Substance|SIMPLE_SEGMENT|11149,11161|true|false|false|C0022650|Kidney Calculi|kidney stone
Event|Event|SIMPLE_SEGMENT|11156,11161|true|false|false|||stone
Finding|Body Substance|SIMPLE_SEGMENT|11156,11161|true|false|false|C0006736|Calculi|stone
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11168,11177|true|false|false|C0009450|Communicable Diseases|infection
Event|Event|SIMPLE_SEGMENT|11168,11177|true|false|false|||infection
Finding|Pathologic Function|SIMPLE_SEGMENT|11168,11177|true|false|false|C3714514|Infection|infection
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11184,11192|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|diabetes
Event|Event|SIMPLE_SEGMENT|11184,11192|false|false|false|||diabetes
Event|Event|SIMPLE_SEGMENT|11198,11208|false|false|false|||controlled
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|11217,11224|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|SIMPLE_SEGMENT|11217,11224|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11217,11224|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|SIMPLE_SEGMENT|11217,11224|false|false|false|||insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|11217,11224|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|11217,11224|false|false|false|C0202098|Insulin measurement|insulin
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11225,11230|false|false|false|C0222045|Integumentary scale|scale
Event|Activity|SIMPLE_SEGMENT|11225,11230|false|false|false|C1947916|Scaling|scale
Finding|Conceptual Entity|SIMPLE_SEGMENT|11225,11230|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|scale
Finding|Intellectual Product|SIMPLE_SEGMENT|11225,11230|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|scale
Event|Event|SIMPLE_SEGMENT|11249,11258|false|false|false|||inpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|11249,11258|false|false|false|C1548438;C1549404|Patient Class - Inpatient;Referral category - Inpatient|inpatient
Procedure|Health Care Activity|SIMPLE_SEGMENT|11249,11258|false|false|false|C1555324|inpatient encounter|inpatient
Event|Event|SIMPLE_SEGMENT|11273,11283|false|false|false|||discharged
Event|Event|SIMPLE_SEGMENT|11284,11288|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|11284,11288|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|11284,11288|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|11284,11288|false|false|false|C1553498|home health encounter|home
Drug|Antibiotic|SIMPLE_SEGMENT|11292,11303|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|SIMPLE_SEGMENT|11292,11303|false|false|false|||antibiotics
Event|Event|SIMPLE_SEGMENT|11308,11314|false|false|false|||intent
Finding|Idea or Concept|SIMPLE_SEGMENT|11308,11314|false|false|false|C0162425;C1550453|Act Mood - intent|intent
Finding|Mental Process|SIMPLE_SEGMENT|11308,11314|false|false|false|C0162425;C1550453|Act Mood - intent|intent
Event|Event|SIMPLE_SEGMENT|11318,11324|false|false|false|||follow
Finding|Functional Concept|SIMPLE_SEGMENT|11318,11324|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|SIMPLE_SEGMENT|11318,11324|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|SIMPLE_SEGMENT|11339,11351|false|false|false|C1547426|Location Service Code - Primary Care|primary care
Procedure|Health Care Activity|SIMPLE_SEGMENT|11339,11351|false|false|false|C0033137|Primary Health Care|primary care
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11339,11360|false|false|false|C2735025||primary care provider
Finding|Idea or Concept|SIMPLE_SEGMENT|11339,11360|false|false|false|C1547431|Primary Care Provider - Provider role|primary care provider
Event|Activity|SIMPLE_SEGMENT|11347,11351|false|false|false|C1947933|care activity|care
Finding|Finding|SIMPLE_SEGMENT|11347,11351|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|11347,11351|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Functional Concept|SIMPLE_SEGMENT|11352,11360|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|provider
Finding|Intellectual Product|SIMPLE_SEGMENT|11352,11360|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|provider
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11388,11399|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11388,11399|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|11388,11399|false|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|11388,11399|false|false|false|C4284232|Medications|medications
Event|Event|SIMPLE_SEGMENT|11403,11413|false|false|false|||prescribed
Event|Activity|SIMPLE_SEGMENT|11437,11449|false|false|false|C0003629|Appointments|appointments
Event|Event|SIMPLE_SEGMENT|11437,11449|false|false|false|||appointments
Event|Event|SIMPLE_SEGMENT|11482,11486|false|false|false|||call
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11493,11499|false|false|false|C0944911||weight
Event|Event|SIMPLE_SEGMENT|11493,11499|false|false|false|||weight
Finding|Finding|SIMPLE_SEGMENT|11493,11499|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|SIMPLE_SEGMENT|11493,11499|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|SIMPLE_SEGMENT|11493,11499|false|false|false|C1305866|Weighing patient|weight
Event|Event|SIMPLE_SEGMENT|11500,11504|false|false|false|||goes
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|11521,11524|false|false|false|C3161851|liquid-based cytology (procedure)|lbs
Event|Event|SIMPLE_SEGMENT|11536,11544|false|false|false|||pleasure
Finding|Intellectual Product|SIMPLE_SEGMENT|11536,11544|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|SIMPLE_SEGMENT|11536,11544|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|SIMPLE_SEGMENT|11552,11556|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|11552,11556|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|11552,11556|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|11552,11556|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|11552,11559|false|false|false|C1555558|care of - AddressPartType|care of
Event|Activity|SIMPLE_SEGMENT|11574,11578|false|false|false|C1947933|care activity|Care
Finding|Finding|SIMPLE_SEGMENT|11574,11578|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|SIMPLE_SEGMENT|11574,11578|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11574,11583|false|false|false|C4321316||Care Team
Finding|Finding|SIMPLE_SEGMENT|11574,11583|false|false|false|C4321315|Care team|Care Team
Procedure|Health Care Activity|SIMPLE_SEGMENT|11586,11594|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11595,11607|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|11595,11607|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|11595,11607|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

