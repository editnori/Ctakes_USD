 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|46,55|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|46,55|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|46,60|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|80,89|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|80,89|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|80,94|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|136,139|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|147,154|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|147,154|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|156,164|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|SIMPLE_SEGMENT|167,176|false|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|167,176|false|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|167,176|false|false|false|C0020517|Hypersensitivity|Allergies
Attribute|Clinical Attribute|SIMPLE_SEGMENT|188,197|false|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|188,197|false|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|188,197|false|false|false|C0020517|Hypersensitivity|Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|200,222|true|false|false|C0041755|Adverse reaction to drug|Adverse Drug Reactions
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|208,212|false|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|Drug
Finding|Finding|SIMPLE_SEGMENT|208,212|false|false|false|C0740721|Drug problem|Drug
Finding|Pathologic Function|SIMPLE_SEGMENT|208,222|true|false|false|C0041755|Adverse reaction to drug|Drug Reactions
Event|Event|SIMPLE_SEGMENT|213,222|false|false|false|||Reactions
Event|Event|SIMPLE_SEGMENT|225,234|false|false|false|||Attending
Finding|Functional Concept|SIMPLE_SEGMENT|225,234|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|SIMPLE_SEGMENT|243,258|false|false|false|C0277786|Chief complaint (finding)|Chief Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|249,258|false|false|false|C3864418||Complaint
Event|Event|SIMPLE_SEGMENT|249,258|false|false|false|||Complaint
Finding|Finding|SIMPLE_SEGMENT|249,258|false|false|false|C5441521|Complaint (finding)|Complaint
Anatomy|Body Location or Region|SIMPLE_SEGMENT|260,265|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|SIMPLE_SEGMENT|260,265|false|false|false|C0741025|Chest problem|Chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|260,270|false|false|false|C2926613||Chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|260,270|false|false|false|C0008031|Chest Pain|Chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|266,270|false|true|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|266,270|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|266,270|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|266,270|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Classification|SIMPLE_SEGMENT|275,280|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|SIMPLE_SEGMENT|281,289|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|281,289|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|293,311|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|302,311|false|false|false|C0945766||Procedure
Event|Event|SIMPLE_SEGMENT|302,311|false|false|false|||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|302,311|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|302,311|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|302,311|false|false|false|C0184661|Interventional procedure|Procedure
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|313,320|false|false|false|C0018787|Heart|Cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|313,320|false|false|false|C1314974|Cardiac attachment|Cardiac
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|313,336|false|false|false|C0261588|Cardiac catheterisation as the cause of abnormal reaction of the patient, or of later complication, without mention of misadventure at the time of the procedure|Cardiac catheterization
Finding|Intellectual Product|SIMPLE_SEGMENT|313,336|false|false|false|C1547981|Diagnostic Service Section ID - Cardiac Catheterization|Cardiac catheterization
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|313,336|false|false|false|C0018795;C1548828|Cardiac Catheterization Procedures;Consent Type - Cardiac Catheterization|Cardiac catheterization
Procedure|Health Care Activity|SIMPLE_SEGMENT|313,336|false|false|false|C0018795;C1548828|Cardiac Catheterization Procedures;Consent Type - Cardiac Catheterization|Cardiac catheterization
Event|Event|SIMPLE_SEGMENT|321,336|false|false|false|||catheterization
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|321,336|false|false|false|C0007430|Catheterization|catheterization
Event|Event|SIMPLE_SEGMENT|342,350|false|false|false|||stenting
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|342,350|false|false|false|C2348535|Stenting|stenting
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|356,360|false|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|drug
Finding|Finding|SIMPLE_SEGMENT|356,360|false|false|false|C0740721|Drug problem|drug
Event|Event|SIMPLE_SEGMENT|369,374|false|false|false|||stent
Finding|Functional Concept|SIMPLE_SEGMENT|383,387|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Event|Event|SIMPLE_SEGMENT|402,409|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|402,409|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|402,409|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|402,409|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|402,412|false|false|false|C0262926|Medical History|History of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|402,428|false|false|false|C0488508||History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|402,428|false|false|false|C0262512|History of present illness (finding)|History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|413,420|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Idea or Concept|SIMPLE_SEGMENT|413,420|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Finding|SIMPLE_SEGMENT|413,428|false|false|false|C4264312|Present illness|Present Illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|421,428|false|false|false|C0221423|Illness (finding)|Illness
Finding|Idea or Concept|SIMPLE_SEGMENT|434,438|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|SIMPLE_SEGMENT|434,438|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Event|Event|SIMPLE_SEGMENT|439,442|false|false|false|||old
Attribute|Clinical Attribute|SIMPLE_SEGMENT|454,463|false|false|false|C0012000|Diastole|diastolic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|454,467|false|false|false|C2183328|diastolic congestive heart failure|diastolic CHF
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|464,467|false|false|false|C0262212|Choroidal fissure|CHF
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|464,467|false|false|false|C0018802|Congestive heart failure|CHF
Event|Event|SIMPLE_SEGMENT|464,467|false|false|false|||CHF
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|469,473|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|469,473|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|SIMPLE_SEGMENT|469,473|false|false|false|||COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|469,473|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|479,482|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|SIMPLE_SEGMENT|479,482|false|false|false|||HTN
Event|Event|SIMPLE_SEGMENT|484,487|false|false|false|||HLD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|494,497|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|494,497|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|494,497|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|494,497|false|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|494,497|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|494,497|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|494,497|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|494,497|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|518,521|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|518,521|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|518,521|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Event|Event|SIMPLE_SEGMENT|522,530|false|false|false|||stenting
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|522,530|false|false|false|C2348535|Stenting|stenting
Finding|Functional Concept|SIMPLE_SEGMENT|532,538|false|false|false|C0205341;C1705914|Repeat;Repeat Object|repeat
Event|Event|SIMPLE_SEGMENT|539,547|false|false|false|||stenting
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|539,547|false|false|false|C2348535|Stenting|stenting
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|553,556|false|false|false|C4551552|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|DES
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|553,556|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Biologically Active Substance|SIMPLE_SEGMENT|553,556|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Hormone|SIMPLE_SEGMENT|553,556|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Organic Chemical|SIMPLE_SEGMENT|553,556|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|553,556|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Event|Event|SIMPLE_SEGMENT|553,556|false|false|false|||DES
Finding|Gene or Genome|SIMPLE_SEGMENT|553,556|false|false|false|C1413980|DES gene|DES
Event|Event|SIMPLE_SEGMENT|578,586|false|false|false|||presents
Anatomy|Body Location or Region|SIMPLE_SEGMENT|592,597|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|592,597|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|592,602|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|592,602|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|598,602|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|598,602|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|598,602|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|598,602|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Anatomy|Body Location or Region|SIMPLE_SEGMENT|625,630|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|625,630|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|625,635|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|625,635|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|631,635|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|631,635|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|631,635|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|631,635|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|636,644|false|false|false|||episodes
Event|Event|SIMPLE_SEGMENT|681,688|false|false|false|||located
Anatomy|Body Location or Region|SIMPLE_SEGMENT|704,709|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|704,709|false|false|false|C0741025|Chest problem|chest
Finding|Finding|SIMPLE_SEGMENT|715,722|false|false|false|C3888388|Usually|usually
Event|Event|SIMPLE_SEGMENT|723,729|false|false|false|||occurs
Event|Event|SIMPLE_SEGMENT|736,744|false|false|false|||exertion
Finding|Organism Function|SIMPLE_SEGMENT|736,744|false|false|false|C0015264|Exertion|exertion
Event|Event|SIMPLE_SEGMENT|759,763|false|false|false|||flat
Event|Event|SIMPLE_SEGMENT|792,803|false|false|false|||experienced
Finding|Functional Concept|SIMPLE_SEGMENT|804,811|false|false|false|C0443144|At rest (qualifier value)|at rest
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|807,811|false|false|false|C1742913|REST protein, human|rest
Drug|Biologically Active Substance|SIMPLE_SEGMENT|807,811|false|false|false|C1742913|REST protein, human|rest
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|807,811|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Gene or Genome|SIMPLE_SEGMENT|807,811|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Molecular Function|SIMPLE_SEGMENT|807,811|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Event|Event|SIMPLE_SEGMENT|816,824|false|false|false|||radiates
Finding|Functional Concept|SIMPLE_SEGMENT|832,836|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|832,840|false|false|false|C0230347;C5779993|Left arm;Left upper arm structure|left arm
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|837,840|false|false|false|C0446516;C1140618;C1269078|Upper Extremity;Upper arm|arm
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|837,840|false|false|false|C3495676|Anorectal Malformations|arm
Finding|Gene or Genome|SIMPLE_SEGMENT|837,840|false|false|false|C1824218;C3715044|AKR1A1 wt Allele;ARMC9 gene|arm
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|837,840|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Research Activity|SIMPLE_SEGMENT|837,840|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|837,840|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Event|Event|SIMPLE_SEGMENT|850,858|false|false|false|||relieved
Event|Event|SIMPLE_SEGMENT|864,867|false|false|false|||NTG
Finding|Finding|SIMPLE_SEGMENT|864,867|false|false|false|C1417953;C1847730;C5575300|GLAUCOMA, NORMAL TENSION, SUSCEPTIBILITY TO;OPA1 gene;OPA1 wt Allele|NTG
Finding|Gene or Genome|SIMPLE_SEGMENT|864,867|false|false|false|C1417953;C1847730;C5575300|GLAUCOMA, NORMAL TENSION, SUSCEPTIBILITY TO;OPA1 gene;OPA1 wt Allele|NTG
Event|Event|SIMPLE_SEGMENT|879,888|false|false|false|||pleuritic
Event|Event|SIMPLE_SEGMENT|897,909|false|false|false|||reproducible
Event|Event|SIMPLE_SEGMENT|920,927|false|false|false|||presses
Anatomy|Body Location or Region|SIMPLE_SEGMENT|945,950|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|945,950|false|false|false|C0741025|Chest problem|chest
Finding|Finding|SIMPLE_SEGMENT|952,960|false|false|false|C2984079|Somewhat|Somewhat
Event|Event|SIMPLE_SEGMENT|961,970|false|false|false|||different
Anatomy|Body Location or Region|SIMPLE_SEGMENT|981,986|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|981,986|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|981,991|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|981,991|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|987,991|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|987,991|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|987,991|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|987,991|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|1027,1031|false|false|false|C0228147|Structure of cisterna pontis|PCIs
Event|Event|SIMPLE_SEGMENT|1034,1044|false|false|false|||Associated
Event|Event|SIMPLE_SEGMENT|1050,1058|false|false|false|||dsyspnea
Event|Event|SIMPLE_SEGMENT|1063,1078|false|false|false|||lightheadedness
Finding|Sign or Symptom|SIMPLE_SEGMENT|1063,1078|false|false|false|C0220870|Lightheadedness|lightheadedness
Event|Event|SIMPLE_SEGMENT|1084,1088|false|false|false|||came
Finding|Finding|SIMPLE_SEGMENT|1126,1132|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|SIMPLE_SEGMENT|1126,1132|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Event|Event|SIMPLE_SEGMENT|1141,1150|false|false|false|||yesterday
Finding|Idea or Concept|SIMPLE_SEGMENT|1168,1175|false|false|false|C1555582|Initial (abbreviation)|initial
Event|Event|SIMPLE_SEGMENT|1215,1218|false|false|false|||EKG
Finding|Intellectual Product|SIMPLE_SEGMENT|1215,1218|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1215,1218|false|false|false|C1623258|Electrocardiography|EKG
Event|Event|SIMPLE_SEGMENT|1220,1226|false|false|false|||showed
Event|Event|SIMPLE_SEGMENT|1257,1264|false|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|1257,1264|false|false|false|C0392747|Changing|changes
Event|Event|SIMPLE_SEGMENT|1266,1269|false|false|false|||CXR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1266,1269|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|SIMPLE_SEGMENT|1270,1278|false|false|false|||negative
Finding|Classification|SIMPLE_SEGMENT|1270,1278|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|1270,1278|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1270,1278|false|false|false|C5237010|Expression Negative|negative
Finding|Finding|SIMPLE_SEGMENT|1270,1282|false|false|false|C0205160|Negative|negative for
Finding|Intellectual Product|SIMPLE_SEGMENT|1284,1289|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1290,1297|false|false|false|C1184743|bony process|process
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1290,1297|false|false|false|C1951340|Process Pharmacologic Substance|process
Event|Event|SIMPLE_SEGMENT|1290,1297|false|false|false|||process
Finding|Functional Concept|SIMPLE_SEGMENT|1290,1297|false|false|false|C4521054|Process (qualifier value)|process
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|1290,1297|false|false|false|C1522240|Process|process
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1299,1303|false|false|false|C0587081|Laboratory test finding|Labs
Event|Event|SIMPLE_SEGMENT|1304,1311|false|false|false|||notable
Finding|Finding|SIMPLE_SEGMENT|1312,1324|false|false|false|C0205160|Negative|for negative
Event|Event|SIMPLE_SEGMENT|1316,1324|false|false|false|||negative
Finding|Classification|SIMPLE_SEGMENT|1316,1324|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|1316,1324|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1316,1324|false|false|false|C5237010|Expression Negative|negative
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1325,1333|false|false|false|C0041199|Troponin|troponin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1325,1333|false|false|false|C0041199|Troponin|troponin
Event|Event|SIMPLE_SEGMENT|1325,1333|false|false|false|||troponin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1325,1333|false|false|false|C0523952|Troponin measurement|troponin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1405,1408|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Enzyme|SIMPLE_SEGMENT|1405,1408|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Organic Chemical|SIMPLE_SEGMENT|1405,1408|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1405,1408|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Event|Event|SIMPLE_SEGMENT|1405,1408|false|false|false|||ASA
Finding|Gene or Genome|SIMPLE_SEGMENT|1405,1408|false|false|false|C1412553|ARSA gene|ASA
Event|Event|SIMPLE_SEGMENT|1410,1415|false|false|false|||325mg
Event|Event|SIMPLE_SEGMENT|1429,1437|false|false|false|||transfer
Finding|Functional Concept|SIMPLE_SEGMENT|1429,1437|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|SIMPLE_SEGMENT|1429,1437|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|SIMPLE_SEGMENT|1429,1437|false|false|false|C4706767|Transfer (immobility management)|transfer
Event|Activity|SIMPLE_SEGMENT|1482,1489|false|false|false|C1706079||arrival
Event|Event|SIMPLE_SEGMENT|1482,1489|false|false|false|||arrival
Finding|Functional Concept|SIMPLE_SEGMENT|1482,1489|false|false|false|C1555577|arrival - ActRelationshipType|arrival
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|1497,1502|false|false|false|C3714591|Floor (anatomic)|floor
Finding|Body Substance|SIMPLE_SEGMENT|1504,1511|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1504,1511|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1504,1511|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|1515,1526|false|false|false|||comfortable
Finding|Finding|SIMPLE_SEGMENT|1515,1526|false|false|false|C5546696|Feeling comfortable|comfortable
Event|Event|SIMPLE_SEGMENT|1531,1537|false|false|false|||denies
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1538,1543|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|1538,1543|true|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1545,1549|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|1545,1549|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|1545,1549|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1545,1549|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|1557,1563|false|false|false|||REVIEW
Finding|Idea or Concept|SIMPLE_SEGMENT|1557,1563|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|REVIEW
Finding|Intellectual Product|SIMPLE_SEGMENT|1557,1563|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|REVIEW
Finding|Functional Concept|SIMPLE_SEGMENT|1557,1566|false|false|false|C0699752|Review of|REVIEW OF
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1557,1574|false|false|false|C0488564;C0488565||REVIEW OF SYSTEMS
Procedure|Health Care Activity|SIMPLE_SEGMENT|1557,1574|false|false|false|C0489633|Review of systems (procedure)|REVIEW OF SYSTEMS
Event|Event|SIMPLE_SEGMENT|1567,1574|false|false|false|||SYSTEMS
Finding|Functional Concept|SIMPLE_SEGMENT|1567,1574|false|false|false|C0449913|System|SYSTEMS
Event|Event|SIMPLE_SEGMENT|1579,1584|false|false|false|||noted
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1588,1591|false|false|false|C0268529|Proline dehydrogenase deficiency|HPI
Event|Event|SIMPLE_SEGMENT|1588,1591|false|false|false|||HPI
Finding|Finding|SIMPLE_SEGMENT|1588,1591|false|false|false|C0262512;C1323983|History of present illness (finding);allene oxide synthase activity|HPI
Finding|Molecular Function|SIMPLE_SEGMENT|1588,1591|false|false|false|C0262512;C1323983|History of present illness (finding);allene oxide synthase activity|HPI
Finding|Functional Concept|SIMPLE_SEGMENT|1596,1604|false|false|false|C0332287;C1883712|Add - instruction imperative;In addition to|addition
Event|Event|SIMPLE_SEGMENT|1606,1612|false|false|false|||denies
Event|Event|SIMPLE_SEGMENT|1613,1619|false|false|false|||fevers
Finding|Sign or Symptom|SIMPLE_SEGMENT|1613,1619|true|false|false|C0015967|Fever|fevers
Event|Event|SIMPLE_SEGMENT|1622,1628|false|false|false|||chills
Finding|Sign or Symptom|SIMPLE_SEGMENT|1622,1628|false|false|false|C0085593|Chills|chills
Event|Event|SIMPLE_SEGMENT|1630,1636|false|false|false|||sweats
Finding|Body Substance|SIMPLE_SEGMENT|1630,1636|false|false|false|C0038984;C0038990|Sweat;Sweating|sweats
Finding|Finding|SIMPLE_SEGMENT|1630,1636|false|false|false|C0038984;C0038990|Sweat;Sweating|sweats
Event|Event|SIMPLE_SEGMENT|1638,1648|false|false|false|||presyncope
Finding|Sign or Symptom|SIMPLE_SEGMENT|1638,1648|false|false|false|C0700200|Presyncope|presyncope
Event|Event|SIMPLE_SEGMENT|1650,1657|false|false|false|||syncope
Finding|Sign or Symptom|SIMPLE_SEGMENT|1650,1657|false|false|false|C0039070|Syncope|syncope
Drug|Organic Chemical|SIMPLE_SEGMENT|1659,1664|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1659,1664|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|SIMPLE_SEGMENT|1659,1664|false|false|false|||cough
Finding|Sign or Symptom|SIMPLE_SEGMENT|1659,1664|false|false|false|C0010200|Coughing|cough
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1666,1669|false|false|false|C1956415|Paroxysmal nocturnal dyspnea|PND
Event|Event|SIMPLE_SEGMENT|1666,1669|false|false|false|||PND
Finding|Gene or Genome|SIMPLE_SEGMENT|1666,1669|false|false|false|C1417807;C4552608|NPPA gene;NPPA wt Allele|PND
Event|Event|SIMPLE_SEGMENT|1671,1680|false|false|false|||orthopnea
Finding|Finding|SIMPLE_SEGMENT|1671,1680|false|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|1671,1680|false|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1682,1685|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Event|Event|SIMPLE_SEGMENT|1687,1695|false|false|false|||swelling
Finding|Finding|SIMPLE_SEGMENT|1687,1695|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|SIMPLE_SEGMENT|1687,1695|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1697,1706|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|SIMPLE_SEGMENT|1697,1711|false|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1707,1711|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|1707,1711|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|1707,1711|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1707,1711|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1713,1719|false|false|false|C4255480||nausea
Event|Event|SIMPLE_SEGMENT|1713,1719|false|false|false|||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|1713,1719|false|false|false|C0027497|Nausea|nausea
Event|Event|SIMPLE_SEGMENT|1721,1729|false|false|false|||vomiting
Finding|Sign or Symptom|SIMPLE_SEGMENT|1721,1729|false|false|false|C0042963|Vomiting|vomiting
Event|Event|SIMPLE_SEGMENT|1731,1742|false|false|false|||hematemesis
Finding|Sign or Symptom|SIMPLE_SEGMENT|1731,1742|false|false|false|C0018926|Hematemesis|hematemesis
Event|Event|SIMPLE_SEGMENT|1745,1753|false|false|false|||diarrhea
Finding|Finding|SIMPLE_SEGMENT|1745,1753|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|SIMPLE_SEGMENT|1745,1753|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Event|Event|SIMPLE_SEGMENT|1755,1767|false|false|false|||constipation
Finding|Sign or Symptom|SIMPLE_SEGMENT|1755,1767|false|false|false|C0009806|Constipation|constipation
Finding|Finding|SIMPLE_SEGMENT|1769,1772|false|false|false|C0332575;C1414207;C1416378|DYRK3 gene;IK gene;Redness|red
Finding|Gene or Genome|SIMPLE_SEGMENT|1769,1772|false|false|false|C0332575;C1414207;C1416378|DYRK3 gene;IK gene;Redness|red
Finding|Pathologic Function|SIMPLE_SEGMENT|1776,1788|false|false|false|C0025222;C0474585|Melena|black stools
Finding|Sign or Symptom|SIMPLE_SEGMENT|1776,1788|false|false|false|C0025222;C0474585|Melena|black stools
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1782,1788|false|false|false|C0489144||stools
Event|Event|SIMPLE_SEGMENT|1782,1788|false|false|false|||stools
Finding|Body Substance|SIMPLE_SEGMENT|1782,1788|false|false|false|C0015733|Feces|stools
Event|Event|SIMPLE_SEGMENT|1790,1797|false|false|false|||dysuria
Finding|Sign or Symptom|SIMPLE_SEGMENT|1790,1797|false|false|false|C0013428|Dysuria|dysuria
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1799,1808|false|false|false|C0018965|Hematuria|hematuria
Event|Event|SIMPLE_SEGMENT|1799,1808|false|false|false|||hematuria
Event|Event|SIMPLE_SEGMENT|1811,1819|false|false|false|||myalgias
Finding|Sign or Symptom|SIMPLE_SEGMENT|1811,1819|false|false|false|C0231528|Myalgia|myalgias
Event|Event|SIMPLE_SEGMENT|1821,1832|false|false|false|||arthralgias
Finding|Sign or Symptom|SIMPLE_SEGMENT|1821,1832|false|false|false|C0003862|Arthralgia|arthralgias
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1837,1841|false|false|false|C5779629|Eruption of skin (disorder)|rash
Event|Event|SIMPLE_SEGMENT|1837,1841|false|false|false|||rash
Finding|Pathologic Function|SIMPLE_SEGMENT|1837,1841|false|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Sign or Symptom|SIMPLE_SEGMENT|1837,1841|false|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Event|Event|SIMPLE_SEGMENT|1846,1853|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|1846,1853|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|1846,1853|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|1846,1853|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|1846,1856|true|false|false|C0262926|Medical History|history of
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1857,1860|true|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1857,1860|true|false|false|C2926618||DVT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1857,1860|true|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Event|Event|SIMPLE_SEGMENT|1857,1860|false|false|false|||DVT
Event|Event|SIMPLE_SEGMENT|1864,1866|false|false|false|||PE
Finding|Finding|SIMPLE_SEGMENT|1873,1893|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Event|Event|SIMPLE_SEGMENT|1878,1885|false|false|false|||Medical
Finding|Functional Concept|SIMPLE_SEGMENT|1878,1885|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|1878,1885|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|1878,1885|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|1878,1885|false|false|false|C0199168|Medical service|Medical
Finding|Finding|SIMPLE_SEGMENT|1878,1893|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1886,1893|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1886,1893|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|1886,1893|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1897,1900|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1897,1900|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|1897,1900|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|1897,1900|false|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|1897,1900|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1897,1900|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|1897,1900|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1897,1900|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1917,1920|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1917,1920|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|1917,1920|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Event|Event|SIMPLE_SEGMENT|1921,1929|false|false|false|||stenting
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1921,1929|false|false|false|C2348535|Stenting|stenting
Finding|Functional Concept|SIMPLE_SEGMENT|1931,1937|false|false|false|C0205341;C1705914|Repeat;Repeat Object|repeat
Event|Event|SIMPLE_SEGMENT|1938,1946|false|false|false|||stenting
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1938,1946|false|false|false|C2348535|Stenting|stenting
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1952,1955|false|false|false|C4551552|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|DES
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1952,1955|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1952,1955|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Hormone|SIMPLE_SEGMENT|1952,1955|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Organic Chemical|SIMPLE_SEGMENT|1952,1955|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1952,1955|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Event|Event|SIMPLE_SEGMENT|1952,1955|false|false|false|||DES
Finding|Gene or Genome|SIMPLE_SEGMENT|1952,1955|false|false|false|C1413980|DES gene|DES
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1978,1987|false|false|false|C0012000|Diastole|Diastolic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1978,1991|false|false|false|C2183328|diastolic congestive heart failure|Diastolic CHF
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|1988,1991|false|false|false|C0262212|Choroidal fissure|CHF
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1988,1991|false|false|false|C0018802|Congestive heart failure|CHF
Event|Event|SIMPLE_SEGMENT|1988,1991|false|false|false|||CHF
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2003,2006|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|SIMPLE_SEGMENT|2003,2006|false|false|false|||HTN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2019,2023|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2019,2023|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|SIMPLE_SEGMENT|2019,2023|false|false|false|||COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|2019,2023|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|2028,2038|false|false|false|C0011570;C0011581;C0344315;C0812393|Cancer patients and suicide and depression;Depressed mood;Depressive disorder;Mental Depression|Depression
Event|Event|SIMPLE_SEGMENT|2028,2038|false|false|false|||Depression
Finding|Functional Concept|SIMPLE_SEGMENT|2028,2038|false|false|false|C0460137;C1579931|Depression - motion|Depression
Finding|Sign or Symptom|SIMPLE_SEGMENT|2028,2038|false|false|false|C0460137;C1579931|Depression - motion|Depression
Finding|Functional Concept|SIMPLE_SEGMENT|2043,2048|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2043,2057|false|false|false|C0524468|Structure of right shoulder region|Right shoulder
Finding|Sign or Symptom|SIMPLE_SEGMENT|2043,2062|false|false|false|C0241040;C5700074|Pain of right shoulder region;right shoulder joint pain|Right shoulder pain
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2049,2057|false|false|false|C0037004;C4299050|Shoulder;Upper extremity>Shoulder|shoulder
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2049,2057|false|false|false|C0221590;C0869975|Examination of shoulder(s);Procedures on Shoulder|shoulder
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2049,2057|false|false|false|C0221590;C0869975|Examination of shoulder(s);Procedures on Shoulder|shoulder
Finding|Sign or Symptom|SIMPLE_SEGMENT|2049,2062|false|false|false|C0037011|Shoulder Pain|shoulder pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2058,2062|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|2058,2062|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|2058,2062|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|2058,2062|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2064,2072|false|false|false|C0006444|Bursitis|bursitis
Event|Event|SIMPLE_SEGMENT|2064,2072|false|false|false|||bursitis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2074,2086|false|false|false|C0085515|Rotator Cuff|rotator cuff
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|2074,2093|false|false|false|C0851122|Rotator Cuff Injuries|rotator cuff injury
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2082,2086|false|false|false|C1550244|Cuff - body part|cuff
Finding|Pathologic Function|SIMPLE_SEGMENT|2082,2086|false|false|false|C3668885|Cuffing (morphologic abnormality)|cuff
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|2087,2093|false|false|false|C3263722;C3263723|Traumatic AND/OR non-traumatic injury;Traumatic injury|injury
Event|Event|SIMPLE_SEGMENT|2087,2093|false|false|false|||injury
Finding|Functional Concept|SIMPLE_SEGMENT|2099,2105|false|false|false|C0728831|Social|Social
Finding|Finding|SIMPLE_SEGMENT|2099,2113|false|false|false|C0424945;C3714536|Social History;Social and personal history|Social History
Event|Event|SIMPLE_SEGMENT|2106,2113|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2106,2113|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2106,2113|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2106,2113|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Classification|SIMPLE_SEGMENT|2119,2125|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|SIMPLE_SEGMENT|2119,2125|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|SIMPLE_SEGMENT|2119,2125|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|SIMPLE_SEGMENT|2119,2125|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Finding|SIMPLE_SEGMENT|2119,2133|false|false|false|C0241889|Family Medical History|Family History
Event|Event|SIMPLE_SEGMENT|2126,2133|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2126,2133|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2126,2133|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2126,2133|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Event|Event|SIMPLE_SEGMENT|2174,2178|false|false|false|||know
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2179,2189|false|true|false|C3812393|ErbB Receptors|her family
Drug|Enzyme|SIMPLE_SEGMENT|2179,2189|false|true|false|C3812393|ErbB Receptors|her family
Finding|Receptor|SIMPLE_SEGMENT|2179,2189|false|true|false|C3812393|ErbB Receptors|her family
Event|Event|SIMPLE_SEGMENT|2183,2189|false|false|false|||family
Finding|Classification|SIMPLE_SEGMENT|2183,2189|true|true|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|2183,2189|true|true|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|2183,2189|true|true|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|2183,2189|true|true|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Event|Event|SIMPLE_SEGMENT|2196,2204|false|false|false|||Physical
Finding|Finding|SIMPLE_SEGMENT|2196,2204|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|2196,2204|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|2196,2204|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|2196,2209|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2196,2209|false|false|false|C0031809|Physical Examination|Physical Exam
Event|Event|SIMPLE_SEGMENT|2205,2209|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|2205,2209|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2205,2209|false|false|false|C0582103|Medical Examination|Exam
Event|Event|SIMPLE_SEGMENT|2211,2220|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|2211,2220|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Finding|Finding|SIMPLE_SEGMENT|2221,2229|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Finding|Functional Concept|SIMPLE_SEGMENT|2221,2229|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|2221,2229|false|false|false|C0031809|Physical Examination|physical
Finding|Finding|SIMPLE_SEGMENT|2221,2234|false|false|false|C1509143|physical examination (physical finding)|physical exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2221,2234|false|false|false|C0031809|Physical Examination|physical exam
Event|Event|SIMPLE_SEGMENT|2230,2234|false|false|false|||exam
Finding|Functional Concept|SIMPLE_SEGMENT|2230,2234|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2230,2234|false|false|false|C0582103|Medical Examination|exam
Event|Event|SIMPLE_SEGMENT|2270,2277|false|false|false|||GENERAL
Finding|Classification|SIMPLE_SEGMENT|2270,2277|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|2270,2277|false|false|false|C3812897|General medical service|GENERAL
Event|Event|SIMPLE_SEGMENT|2284,2289|false|false|false|||woman
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2293,2296|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2293,2296|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2293,2296|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|2293,2296|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2293,2296|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|SIMPLE_SEGMENT|2293,2296|false|false|false|||NAD
Finding|Finding|SIMPLE_SEGMENT|2293,2296|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Finding|Finding|SIMPLE_SEGMENT|2298,2306|false|false|false|C1961028|Oriented to place|Oriented
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2311,2315|false|false|false|C2713234||Mood
Event|Event|SIMPLE_SEGMENT|2311,2315|false|false|false|||Mood
Finding|Conceptual Entity|SIMPLE_SEGMENT|2311,2315|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|Mood
Finding|Finding|SIMPLE_SEGMENT|2311,2315|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|Mood
Finding|Mental Process|SIMPLE_SEGMENT|2311,2315|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|Mood
Event|Event|SIMPLE_SEGMENT|2317,2323|false|false|false|||affect
Finding|Mental Process|SIMPLE_SEGMENT|2317,2323|false|false|false|C0001721|Affect (mental function)|affect
Procedure|Health Care Activity|SIMPLE_SEGMENT|2317,2323|false|false|false|C2237113|assessment of affect|affect
Event|Event|SIMPLE_SEGMENT|2325,2336|false|false|false|||appropriate
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2340,2345|false|false|false|C1512338|HEENT|HEENT
Event|Event|SIMPLE_SEGMENT|2347,2351|false|false|false|||NCAT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2353,2359|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2353,2359|false|false|false|C0036412|Scleral Diseases|Sclera
Event|Event|SIMPLE_SEGMENT|2353,2359|false|false|false|||Sclera
Procedure|Health Care Activity|SIMPLE_SEGMENT|2353,2359|false|false|false|C2228481|examination of sclera|Sclera
Event|Event|SIMPLE_SEGMENT|2360,2369|false|false|false|||anicteric
Finding|Finding|SIMPLE_SEGMENT|2360,2369|false|false|false|C0205180|Anicteric|anicteric
Event|Event|SIMPLE_SEGMENT|2371,2376|false|false|false|||PERRL
Finding|Finding|SIMPLE_SEGMENT|2371,2376|false|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Event|Event|SIMPLE_SEGMENT|2378,2382|false|false|false|||EOMI
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2384,2395|false|false|false|C0009758;C0229274|Structure of palpebral conjunctiva;conjunctiva|Conjunctiva
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2384,2395|false|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|Conjunctiva
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2384,2395|false|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|Conjunctiva
Event|Event|SIMPLE_SEGMENT|2384,2395|false|false|false|||Conjunctiva
Finding|Body Substance|SIMPLE_SEGMENT|2384,2395|false|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|Conjunctiva
Finding|Intellectual Product|SIMPLE_SEGMENT|2384,2395|false|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|Conjunctiva
Procedure|Health Care Activity|SIMPLE_SEGMENT|2384,2395|false|false|false|C0872390;C2228431|Procedure on conjunctiva;examination of conjunctiva|Conjunctiva
Event|Event|SIMPLE_SEGMENT|2411,2417|false|false|false|||pallor
Finding|Finding|SIMPLE_SEGMENT|2411,2417|true|false|false|C0241137|Pallor of skin|pallor
Event|Event|SIMPLE_SEGMENT|2421,2429|false|false|false|||cyanosis
Finding|Sign or Symptom|SIMPLE_SEGMENT|2421,2429|true|false|false|C0010520|Cyanosis|cyanosis
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|2437,2441|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|2437,2441|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|2437,2441|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|2437,2441|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2437,2448|false|false|false|C0026639|Oral mucous membrane structure|oral mucosa
Anatomy|Tissue|SIMPLE_SEGMENT|2442,2448|false|false|false|C0026724|Mucous Membrane|mucosa
Finding|Intellectual Product|SIMPLE_SEGMENT|2442,2448|false|false|false|C1561514||mucosa
Event|Event|SIMPLE_SEGMENT|2453,2464|false|false|false|||xanthalesma
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2469,2473|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|SIMPLE_SEGMENT|2469,2473|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|SIMPLE_SEGMENT|2469,2473|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Event|Event|SIMPLE_SEGMENT|2475,2481|false|false|false|||Supple
Finding|Functional Concept|SIMPLE_SEGMENT|2475,2481|false|false|false|C0332254|Supple|Supple
Event|Event|SIMPLE_SEGMENT|2483,2486|false|false|false|||JVP
Finding|Finding|SIMPLE_SEGMENT|2483,2486|false|false|false|C0428897|Jugular venous pressure|JVP
Event|Event|SIMPLE_SEGMENT|2491,2499|false|false|false|||elevated
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2503,2510|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|SIMPLE_SEGMENT|2503,2510|false|false|false|C1314974|Cardiac attachment|CARDIAC
Event|Event|SIMPLE_SEGMENT|2538,2539|false|false|false|||g
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2554,2558|false|false|false|C2598155||Pain
Finding|Functional Concept|SIMPLE_SEGMENT|2554,2558|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|2554,2558|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Event|Event|SIMPLE_SEGMENT|2560,2572|false|false|false|||reproducible
Event|Event|SIMPLE_SEGMENT|2578,2587|false|false|false|||palpation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2578,2587|false|false|false|C0030247|Palpation|palpation
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2597,2602|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|2597,2602|false|false|false|C0741025|Chest problem|chest
Finding|Functional Concept|SIMPLE_SEGMENT|2607,2611|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2613,2619|false|false|false|C0006141|Breast|breast
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2613,2619|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|breast
Event|Event|SIMPLE_SEGMENT|2613,2619|false|false|false|||breast
Finding|Finding|SIMPLE_SEGMENT|2613,2619|false|false|false|C0567499|Breast problem|breast
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2613,2619|false|false|false|C0191838|Procedures on breast|breast
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2623,2628|false|false|false|C0024109|Lung|LUNGS
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2630,2634|false|false|false|C0231832|Respiratory rate|Resp
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2630,2634|false|false|false|C0851355|Respiratory, thoracic and mediastinal disorders|Resp
Event|Event|SIMPLE_SEGMENT|2630,2634|false|false|false|||Resp
Event|Event|SIMPLE_SEGMENT|2635,2644|false|false|false|||unlabored
Finding|Functional Concept|SIMPLE_SEGMENT|2635,2644|false|false|false|C2983702|Unlabored|unlabored
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|2649,2665|true|false|false|C0158784|Accessory skeletal muscle|accessory muscle
Finding|Finding|SIMPLE_SEGMENT|2649,2669|true|false|false|C1821466|Use of accessory muscles|accessory muscle use
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2659,2665|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Anatomy|Tissue|SIMPLE_SEGMENT|2659,2665|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Event|Event|SIMPLE_SEGMENT|2666,2669|false|false|false|||use
Finding|Functional Concept|SIMPLE_SEGMENT|2666,2669|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|SIMPLE_SEGMENT|2666,2669|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Drug|Organic Chemical|SIMPLE_SEGMENT|2671,2675|false|false|false|C0951233|cetrimonium bromide|CTAB
Event|Event|SIMPLE_SEGMENT|2671,2675|false|false|false|||CTAB
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2679,2686|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2679,2686|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Event|Event|SIMPLE_SEGMENT|2679,2686|false|false|false|||ABDOMEN
Finding|Finding|SIMPLE_SEGMENT|2679,2686|false|false|false|C0941288|Abdomen problem|ABDOMEN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2688,2692|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Event|Event|SIMPLE_SEGMENT|2688,2692|false|false|false|||Soft
Event|Event|SIMPLE_SEGMENT|2694,2698|false|false|false|||NTND
Event|Event|SIMPLE_SEGMENT|2703,2706|false|false|false|||HSM
Finding|Gene or Genome|SIMPLE_SEGMENT|2703,2706|true|false|false|C1537594|LRRC4B gene|HSM
Event|Event|SIMPLE_SEGMENT|2710,2720|false|false|false|||tenderness
Finding|Mental Process|SIMPLE_SEGMENT|2710,2720|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|SIMPLE_SEGMENT|2710,2720|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2722,2725|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|Abd
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|2722,2725|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|Abd
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2726,2731|false|false|false|C0003483;C4037978|Aorta;Chest+Abdomen>Aorta|aorta
Procedure|Health Care Activity|SIMPLE_SEGMENT|2726,2731|false|false|false|C0869784|Procedure on aorta|aorta
Event|Event|SIMPLE_SEGMENT|2737,2745|false|false|false|||enlarged
Event|Event|SIMPLE_SEGMENT|2749,2758|false|false|false|||palpation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2749,2758|false|false|false|C0030247|Palpation|palpation
Event|Event|SIMPLE_SEGMENT|2774,2780|false|false|false|||bruits
Finding|Finding|SIMPLE_SEGMENT|2774,2780|true|false|false|C0006318|Bruit|bruits
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2784,2795|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2800,2805|true|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|2800,2805|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|2800,2805|true|false|false|C0013604|Edema|edema
Event|Event|SIMPLE_SEGMENT|2807,2810|false|false|false|||WWP
Anatomy|Body System|SIMPLE_SEGMENT|2814,2818|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2814,2818|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2814,2818|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Event|Event|SIMPLE_SEGMENT|2814,2818|false|false|false|||SKIN
Finding|Body Substance|SIMPLE_SEGMENT|2814,2818|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|SIMPLE_SEGMENT|2814,2818|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Pathologic Function|SIMPLE_SEGMENT|2823,2829|false|false|false|C0333138|Stasis|stasis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2823,2840|true|false|false|C0011620|Stasis dermatitis|stasis dermatitis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2830,2840|true|false|false|C0011603|Dermatitis|dermatitis
Event|Event|SIMPLE_SEGMENT|2830,2840|false|false|false|||dermatitis
Event|Event|SIMPLE_SEGMENT|2842,2848|false|false|false|||ulcers
Finding|Pathologic Function|SIMPLE_SEGMENT|2842,2848|true|false|false|C0041582|Ulcer|ulcers
Event|Event|SIMPLE_SEGMENT|2850,2855|false|false|false|||scars
Finding|Finding|SIMPLE_SEGMENT|2850,2855|true|false|false|C0241158;C2004491|Cicatrix;Scar Tissue|scars
Finding|Pathologic Function|SIMPLE_SEGMENT|2850,2855|true|false|false|C0241158;C2004491|Cicatrix;Scar Tissue|scars
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2860,2869|true|false|false|C0302314|Xanthoma|xanthomas
Event|Event|SIMPLE_SEGMENT|2860,2869|false|false|false|||xanthomas
Drug|Food|SIMPLE_SEGMENT|2873,2879|false|false|false|C5890763||PULSES
Event|Event|SIMPLE_SEGMENT|2873,2879|false|false|false|||PULSES
Finding|Physiologic Function|SIMPLE_SEGMENT|2873,2879|false|false|false|C0391850|Physiologic pulse|PULSES
Procedure|Health Care Activity|SIMPLE_SEGMENT|2873,2879|false|false|false|C0034107|Pulse taking|PULSES
Finding|Functional Concept|SIMPLE_SEGMENT|2883,2888|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2890,2897|false|false|false|C0007272|Carotid Arteries|Carotid
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2901,2908|false|false|false|C0015811|Femur|Femoral
Finding|Functional Concept|SIMPLE_SEGMENT|2927,2931|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2933,2940|false|false|false|C0007272|Carotid Arteries|Carotid
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2944,2951|false|false|false|C0015811|Femur|Femoral
Event|Event|SIMPLE_SEGMENT|2970,2979|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|2970,2979|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|2970,2979|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|2970,2979|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|2970,2979|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|2980,2988|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Finding|Functional Concept|SIMPLE_SEGMENT|2980,2988|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|2980,2988|false|false|false|C0031809|Physical Examination|physical
Finding|Finding|SIMPLE_SEGMENT|2980,2993|false|false|false|C1509143|physical examination (physical finding)|physical exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2980,2993|false|false|false|C0031809|Physical Examination|physical exam
Event|Event|SIMPLE_SEGMENT|2989,2993|false|false|false|||exam
Finding|Functional Concept|SIMPLE_SEGMENT|2989,2993|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2989,2993|false|false|false|C0582103|Medical Examination|exam
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3062,3065|false|false|false|C2744672|SAT1 protein, human|Sat
Drug|Enzyme|SIMPLE_SEGMENT|3062,3065|false|false|false|C2744672|SAT1 protein, human|Sat
Finding|Gene or Genome|SIMPLE_SEGMENT|3062,3065|false|false|false|C0871290;C1705827;C1822614|College Entrance Examination Board Scholastic Aptitude Test;SAT1 gene;SAT1 wt Allele|Sat
Finding|Intellectual Product|SIMPLE_SEGMENT|3062,3065|false|false|false|C0871290;C1705827;C1822614|College Entrance Examination Board Scholastic Aptitude Test;SAT1 gene;SAT1 wt Allele|Sat
Event|Event|SIMPLE_SEGMENT|3074,3081|false|false|false|||General
Finding|Classification|SIMPLE_SEGMENT|3074,3081|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|SIMPLE_SEGMENT|3074,3081|false|false|false|C3812897|General medical service|General
Finding|Body Substance|SIMPLE_SEGMENT|3083,3090|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|3083,3090|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|3083,3090|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|3091,3096|false|false|false|||lying
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3100,3103|false|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Event|Event|SIMPLE_SEGMENT|3100,3103|false|false|false|||bed
Finding|Intellectual Product|SIMPLE_SEGMENT|3100,3103|false|false|false|C2346952|Bachelor of Education|bed
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3107,3110|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3107,3110|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3107,3110|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|3107,3110|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3107,3110|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|SIMPLE_SEGMENT|3107,3110|false|false|false|||NAD
Finding|Finding|SIMPLE_SEGMENT|3107,3110|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3111,3116|false|false|false|C1512338|HEENT|HEENT
Event|Event|SIMPLE_SEGMENT|3118,3122|false|false|false|||EOMI
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3124,3127|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3124,3127|false|false|false|C0026987|Myelofibrosis|MMM
Event|Event|SIMPLE_SEGMENT|3124,3127|false|false|false|||MMM
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3129,3133|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Anatomy|Cell Component|SIMPLE_SEGMENT|3129,3133|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Finding|Finding|SIMPLE_SEGMENT|3129,3133|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|Neck
Event|Event|SIMPLE_SEGMENT|3135,3141|false|false|false|||Supple
Finding|Functional Concept|SIMPLE_SEGMENT|3135,3141|false|false|false|C0332254|Supple|Supple
Event|Event|SIMPLE_SEGMENT|3146,3149|false|false|false|||JVD
Finding|Finding|SIMPLE_SEGMENT|3146,3149|true|false|false|C0425687|Jugular venous engorgement|JVD
Event|Event|SIMPLE_SEGMENT|3150,3161|false|false|false|||appreciated
Event|Event|SIMPLE_SEGMENT|3167,3170|false|false|false|||RRR
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3181,3186|false|false|false|C0024109|Lung|Lungs
Event|Event|SIMPLE_SEGMENT|3188,3193|false|false|false|||Clear
Finding|Idea or Concept|SIMPLE_SEGMENT|3188,3193|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|SIMPLE_SEGMENT|3197,3209|false|false|false|||auscultation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3197,3209|false|false|false|C0004339|Auscultation|auscultation
Event|Event|SIMPLE_SEGMENT|3226,3234|false|false|false|||crackles
Finding|Finding|SIMPLE_SEGMENT|3226,3234|true|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Event|Event|SIMPLE_SEGMENT|3239,3246|false|false|false|||wheezes
Finding|Sign or Symptom|SIMPLE_SEGMENT|3239,3246|false|false|false|C0043144|Wheezing|wheezes
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3248,3251|false|false|false|C0079758|Lymphoma, Mixed-Cell, Follicular|Nml
Finding|Gene or Genome|SIMPLE_SEGMENT|3248,3251|false|false|false|C2680360|RRP8 gene|Nml
Event|Event|SIMPLE_SEGMENT|3252,3256|false|false|false|||work
Event|Occupational Activity|SIMPLE_SEGMENT|3252,3256|false|false|false|C0043227|Work|work
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|3252,3269|false|false|false|C0043229|Work of Breathing|work of breathing
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3260,3269|false|false|false|C5885990||breathing
Event|Event|SIMPLE_SEGMENT|3260,3269|false|false|false|||breathing
Finding|Finding|SIMPLE_SEGMENT|3260,3269|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|SIMPLE_SEGMENT|3260,3269|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|SIMPLE_SEGMENT|3260,3269|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|SIMPLE_SEGMENT|3260,3269|false|false|false|C1160636|respiratory system process|breathing
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3271,3274|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|Abd
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|3271,3274|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|Abd
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3276,3281|false|false|false|C0028754|Obesity|Obese
Event|Event|SIMPLE_SEGMENT|3276,3281|false|false|false|||Obese
Event|Event|SIMPLE_SEGMENT|3283,3287|false|false|false|||NABS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3290,3294|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Event|Event|SIMPLE_SEGMENT|3290,3294|false|false|false|||Soft
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|3303,3306|false|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Event|Event|SIMPLE_SEGMENT|3303,3306|false|false|false|||Ext
Finding|Gene or Genome|SIMPLE_SEGMENT|3303,3306|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Event|Event|SIMPLE_SEGMENT|3308,3311|false|false|false|||WWP
Event|Event|SIMPLE_SEGMENT|3316,3319|false|false|false|||DPs
Finding|Gene or Genome|SIMPLE_SEGMENT|3316,3319|false|false|false|C1843919|PDSS1 gene|DPs
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|3336,3344|true|false|false|C0149651|Clubbing|clubbing
Event|Event|SIMPLE_SEGMENT|3336,3344|false|false|false|||clubbing
Event|Event|SIMPLE_SEGMENT|3346,3354|false|false|false|||cyanosis
Finding|Sign or Symptom|SIMPLE_SEGMENT|3346,3354|true|false|false|C0010520|Cyanosis|cyanosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3359,3364|true|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|3359,3364|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|3359,3364|true|false|false|C0013604|Edema|edema
Procedure|Health Care Activity|SIMPLE_SEGMENT|3387,3396|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3397,3401|false|false|false|C0587081|Laboratory test finding|labs
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3415,3420|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3415,3420|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3415,3420|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|3421,3424|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|3430,3433|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3430,3433|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3430,3433|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3440,3443|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3440,3443|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|3440,3443|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3440,3443|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3449,3452|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3449,3452|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|3459,3462|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|3459,3462|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3459,3462|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3459,3462|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3459,3462|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|3466,3469|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3466,3469|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|3466,3469|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|3466,3469|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|3466,3469|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3466,3469|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3476,3480|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3495,3498|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3515,3520|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3515,3520|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Antibiotic|SIMPLE_SEGMENT|3536,3541|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3536,3541|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|SIMPLE_SEGMENT|3536,3541|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3546,3549|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|Eos
Event|Event|SIMPLE_SEGMENT|3546,3549|false|false|false|||Eos
Finding|Gene or Genome|SIMPLE_SEGMENT|3546,3549|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|Eos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3576,3581|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3576,3581|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3576,3581|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3586,3589|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|SIMPLE_SEGMENT|3586,3589|false|false|false|||PTT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3586,3589|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3611,3616|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3611,3616|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3611,3616|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|3611,3624|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3611,3624|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3611,3624|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3617,3624|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|3617,3624|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3617,3624|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|3617,3624|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3617,3624|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3617,3624|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|SIMPLE_SEGMENT|3672,3676|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3672,3676|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3672,3676|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3702,3707|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3702,3707|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3723,3732|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|3723,3732|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|3723,3732|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|3723,3732|false|false|false|C0030685|Patient Discharge|Discharge
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3733,3737|false|false|false|C0587081|Laboratory test finding|labs
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3751,3756|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3751,3756|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3751,3756|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|3757,3760|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|3766,3769|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3766,3769|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3766,3769|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3776,3779|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3776,3779|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|3776,3779|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3776,3779|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3785,3788|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3785,3788|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|3796,3799|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|3796,3799|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3796,3799|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3796,3799|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3796,3799|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|3803,3806|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3803,3806|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|3803,3806|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|3803,3806|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|3803,3806|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3803,3806|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3813,3817|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3833,3836|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3853,3858|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3853,3858|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3853,3858|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|3853,3866|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3853,3866|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3853,3866|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3859,3866|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|3859,3866|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3859,3866|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|3859,3866|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3859,3866|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3859,3866|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|SIMPLE_SEGMENT|3912,3916|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3912,3916|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3912,3916|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3941,3946|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3941,3946|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3941,3946|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3941,3954|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3947,3954|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|3947,3954|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|3947,3954|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3947,3954|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|3947,3954|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|SIMPLE_SEGMENT|3947,3954|false|false|false|||Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|3947,3954|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3947,3954|false|false|false|C0201925|Calcium measurement|Calcium
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3976,3983|false|false|false|C0018787|Heart|Cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|3976,3983|false|false|false|C1314974|Cardiac attachment|Cardiac
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3976,3991|false|false|false|C2926589||Cardiac enzymes
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3976,3991|false|false|false|C0443763|Cardiac enzymes|Cardiac enzymes
Drug|Enzyme|SIMPLE_SEGMENT|3976,3991|false|false|false|C0443763|Cardiac enzymes|Cardiac enzymes
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3976,3991|false|false|false|C0201934|Cardiac enzymes/isoenzymes measurement|Cardiac enzymes
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3984,3991|false|false|false|C0014442;C3540017;C3540048;C3540772;C3540790;C3541394;C3542456|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS;Enzymes;Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM;Enzymes for ALIMENTARY TRACT AND METABOLISM;Enzymes, antithrombotic;Enzymes, hematological;Enzymes, peripheral vasodilators|enzymes
Drug|Enzyme|SIMPLE_SEGMENT|3984,3991|false|false|false|C0014442;C3540017;C3540048;C3540772;C3540790;C3541394;C3542456|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS;Enzymes;Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM;Enzymes for ALIMENTARY TRACT AND METABOLISM;Enzymes, antithrombotic;Enzymes, hematological;Enzymes, peripheral vasodilators|enzymes
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3984,3991|false|false|false|C0014442;C3540017;C3540048;C3540772;C3540790;C3541394;C3542456|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS;Enzymes;Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM;Enzymes for ALIMENTARY TRACT AND METABOLISM;Enzymes, antithrombotic;Enzymes, hematological;Enzymes, peripheral vasodilators|enzymes
Event|Event|SIMPLE_SEGMENT|3984,3991|false|false|false|||enzymes
Finding|Functional Concept|SIMPLE_SEGMENT|3984,3991|false|false|false|C0014445|enzymology|enzymes
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4005,4010|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4005,4010|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4005,4010|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4014,4017|false|false|false|C0010287|Creatine Kinase|CPK
Drug|Enzyme|SIMPLE_SEGMENT|4014,4017|false|false|false|C0010287|Creatine Kinase|CPK
Event|Event|SIMPLE_SEGMENT|4014,4017|false|false|false|||CPK
Finding|Gene or Genome|SIMPLE_SEGMENT|4014,4017|false|false|false|C1418571|PIK3C2A gene|CPK
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4014,4017|false|false|false|C0201973|Creatine kinase measurement|CPK
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4034,4039|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4034,4039|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4034,4039|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4040,4045|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|SIMPLE_SEGMENT|4040,4045|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|SIMPLE_SEGMENT|4040,4045|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4040,4045|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Drug|Organic Chemical|SIMPLE_SEGMENT|4043,4047|false|false|false|C0602249|MB 2|MB-2
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4074,4079|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4074,4079|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Event|Event|SIMPLE_SEGMENT|4095,4098|false|false|false|||EKG
Finding|Intellectual Product|SIMPLE_SEGMENT|4095,4098|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4095,4098|false|false|false|C1623258|Electrocardiography|EKG
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4100,4105|false|false|false|C0030471;C1305231|Nasal sinus;Sinus - general anatomical term|Sinus
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|4100,4105|false|false|false|C0016169|pathologic fistula|Sinus
Drug|Organic Chemical|SIMPLE_SEGMENT|4100,4105|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|Sinus
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4100,4105|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|Sinus
Finding|Finding|SIMPLE_SEGMENT|4100,4112|false|false|false|C0232201;C2041122|Sinus rhythm|Sinus rhythm
Event|Event|SIMPLE_SEGMENT|4106,4112|false|false|false|||rhythm
Finding|Finding|SIMPLE_SEGMENT|4106,4112|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|SIMPLE_SEGMENT|4106,4112|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Event|Activity|SIMPLE_SEGMENT|4118,4122|false|false|false|C0871208|Rating (action)|rate
Event|Event|SIMPLE_SEGMENT|4118,4122|false|false|false|||rate
Finding|Idea or Concept|SIMPLE_SEGMENT|4118,4122|false|false|false|C1549480|Amount type - Rate|rate
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4137,4141|false|false|false|C0004457|Axis vertebra|axis
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|4137,4141|false|false|false|C0349013|Fracture of second cervical vertebra|axis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4147,4158|false|false|false|C0520877|PR interval feature|PR interval
Finding|Finding|SIMPLE_SEGMENT|4147,4158|false|false|false|C0429087|Finding of electrocardiogram PR interval|PR interval
Event|Event|SIMPLE_SEGMENT|4150,4158|false|false|false|||interval
Finding|Intellectual Product|SIMPLE_SEGMENT|4150,4158|false|false|false|C1552654|Parameterized Data Type - Interval|interval
Event|Event|SIMPLE_SEGMENT|4163,4172|false|false|false|||prolonged
Event|Event|SIMPLE_SEGMENT|4208,4211|false|false|false|||ekg
Finding|Intellectual Product|SIMPLE_SEGMENT|4208,4211|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|ekg
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4208,4211|false|false|false|C1623258|Electrocardiography|ekg
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4214,4220|false|false|false|C1305738|Q wave|Q wave
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4214,4220|false|false|false|C0429089||Q wave
Event|Event|SIMPLE_SEGMENT|4216,4220|false|false|false|||wave
Finding|Gene or Genome|SIMPLE_SEGMENT|4216,4220|false|false|false|C1421479|WASF1 gene|wave
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|4216,4220|false|false|false|C0678544||wave
Event|Event|SIMPLE_SEGMENT|4252,4259|false|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|4252,4259|false|false|false|C0392747|Changing|changes
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4262,4281|false|false|false|C2825165|Nuclear stress test|Nuclear Stress Test
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4270,4276|false|false|false|C1718621|W stress|Stress
Drug|Organic Chemical|SIMPLE_SEGMENT|4270,4276|false|false|false|C0723460|Stress bismuth subsalicylate|Stress
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4270,4276|false|false|false|C0723460|Stress bismuth subsalicylate|Stress
Event|Event|SIMPLE_SEGMENT|4270,4276|false|false|false|||Stress
Finding|Finding|SIMPLE_SEGMENT|4270,4276|false|false|false|C0038435|Stress|Stress
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4270,4281|false|false|false|C0015260;C3494508|Exercise stress test;Stress Test|Stress Test
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4277,4281|false|false|false|C4318744|Test - temporal region|Test
Finding|Functional Concept|SIMPLE_SEGMENT|4277,4281|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|Test
Finding|Intellectual Product|SIMPLE_SEGMENT|4277,4281|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|Test
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4277,4281|false|false|false|C0456984|Test Result|Test
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4277,4281|false|false|false|C0022885|Laboratory Procedures|Test
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4284,4298|false|false|false|C3173575||INTERPRETATION
Event|Event|SIMPLE_SEGMENT|4284,4298|false|false|false|||INTERPRETATION
Finding|Intellectual Product|SIMPLE_SEGMENT|4284,4298|false|false|false|C0459471|Interpretation Process|INTERPRETATION
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4306,4311|false|false|false|C1846009|Intrauterine growth restriction, metaphyseal dysplasia, adrenal hypoplasia congenita, and genital anomaly syndrome|image
Event|Event|SIMPLE_SEGMENT|4306,4311|false|false|false|||image
Finding|Intellectual Product|SIMPLE_SEGMENT|4306,4311|false|false|false|C1696103;C1704254;C1704922;C3542466|Image;Image (foundation metadata concept);Medical Image;image - dosage form|image
Event|Event|SIMPLE_SEGMENT|4323,4331|false|false|false|||adequate
Event|Event|SIMPLE_SEGMENT|4336,4343|false|false|false|||limited
Finding|Functional Concept|SIMPLE_SEGMENT|4336,4343|false|false|false|C0439801;C3542948|Limited (extensiveness);Limited component (foundation metadata concept)|limited
Finding|Intellectual Product|SIMPLE_SEGMENT|4336,4343|false|false|false|C0439801;C3542948|Limited (extensiveness);Limited component (foundation metadata concept)|limited
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4351,4355|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4351,4362|false|false|false|C0225317;C4532079|Neck+Chest>Soft tissue;soft tissue|soft tissue
Anatomy|Tissue|SIMPLE_SEGMENT|4351,4362|false|false|false|C0225317;C4532079|Neck+Chest>Soft tissue;soft tissue|soft tissue
Anatomy|Tissue|SIMPLE_SEGMENT|4356,4362|false|false|false|C0040300|Body tissue|tissue
Finding|Intellectual Product|SIMPLE_SEGMENT|4356,4362|false|false|false|C1547928|Tissue Specimen Code|tissue
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4368,4374|false|false|false|C0006141|Breast|breast
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4368,4374|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|breast
Event|Event|SIMPLE_SEGMENT|4368,4374|false|false|false|||breast
Finding|Finding|SIMPLE_SEGMENT|4368,4374|false|false|false|C0567499|Breast problem|breast
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4368,4374|false|false|false|C0191838|Procedures on breast|breast
Event|Activity|SIMPLE_SEGMENT|4375,4386|false|false|false|C0599946|Attenuation|attenuation
Event|Event|SIMPLE_SEGMENT|4375,4386|false|false|false|||attenuation
Event|Activity|SIMPLE_SEGMENT|4397,4405|false|false|false|C0441655|Activities|activity
Event|Event|SIMPLE_SEGMENT|4397,4405|false|false|false|||activity
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|4397,4405|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|activity
Finding|Finding|SIMPLE_SEGMENT|4397,4405|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|activity
Event|Event|SIMPLE_SEGMENT|4406,4414|false|false|false|||adjacent
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4422,4427|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4422,4427|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|4422,4427|false|false|false|C0795691|HEART PROBLEM|heart
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4436,4440|false|false|false|C1742913|REST protein, human|rest
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4436,4440|false|false|false|C1742913|REST protein, human|rest
Event|Event|SIMPLE_SEGMENT|4436,4440|false|false|false|||rest
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|4436,4440|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Gene or Genome|SIMPLE_SEGMENT|4436,4440|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Molecular Function|SIMPLE_SEGMENT|4436,4440|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4445,4451|false|false|false|C1718621|W stress|stress
Drug|Organic Chemical|SIMPLE_SEGMENT|4445,4451|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4445,4451|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Finding|Finding|SIMPLE_SEGMENT|4445,4451|false|false|false|C0038435|Stress|stress
Event|Event|SIMPLE_SEGMENT|4452,4458|false|false|false|||images
Finding|Functional Concept|SIMPLE_SEGMENT|4461,4465|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4461,4484|false|false|false|C0503990|Cavity of left ventricle|Left ventricular cavity
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4461,4489|false|false|false|C0455830|Left ventricular cavity size|Left ventricular cavity size
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4466,4477|false|false|false|C0018827|Heart Ventricle|ventricular
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4466,4484|false|false|false|C0507083|Cavity of ventricle|ventricular cavity
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4478,4484|false|false|false|C0333343|Body cavities|cavity
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|4478,4484|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4478,4484|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Event|Event|SIMPLE_SEGMENT|4493,4502|false|false|false|||increased
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4505,4509|false|false|false|C1742913|REST protein, human|Rest
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4505,4509|false|false|false|C1742913|REST protein, human|Rest
Event|Event|SIMPLE_SEGMENT|4505,4509|false|false|false|||Rest
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|4505,4509|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|Rest
Finding|Gene or Genome|SIMPLE_SEGMENT|4505,4509|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|Rest
Finding|Molecular Function|SIMPLE_SEGMENT|4505,4509|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|Rest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4514,4520|false|false|false|C1718621|W stress|stress
Drug|Organic Chemical|SIMPLE_SEGMENT|4514,4520|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4514,4520|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Event|Event|SIMPLE_SEGMENT|4514,4520|false|false|false|||stress
Finding|Finding|SIMPLE_SEGMENT|4514,4520|false|false|false|C0038435|Stress|stress
Finding|Functional Concept|SIMPLE_SEGMENT|4521,4530|false|false|false|C4281794;C4723760|Perfusion (biological);Perfusion route|perfusion
Finding|Organism Function|SIMPLE_SEGMENT|4521,4530|false|false|false|C4281794;C4723760|Perfusion (biological);Perfusion route|perfusion
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4521,4530|false|false|false|C0031001;C4721534|Chemotherapeutic Perfusion;Perfusion (procedure)|perfusion
Event|Event|SIMPLE_SEGMENT|4531,4537|false|false|false|||images
Event|Event|SIMPLE_SEGMENT|4547,4557|false|false|false|||reversible
Finding|Functional Concept|SIMPLE_SEGMENT|4547,4557|false|false|false|C0205343|Reversible|reversible
Event|Event|SIMPLE_SEGMENT|4559,4567|false|false|false|||moderate
Finding|Finding|SIMPLE_SEGMENT|4559,4567|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|SIMPLE_SEGMENT|4559,4567|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Event|Event|SIMPLE_SEGMENT|4569,4578|false|false|false|||reduction
Finding|Finding|SIMPLE_SEGMENT|4569,4578|false|false|false|C0392756|Reduced|reduction
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|4569,4578|false|false|false|C0301630|Reduction (chemical)|reduction
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4569,4578|false|false|false|C1293152;C4551656|Reduction procedure;Surgical reduction|reduction
Drug|Substance|SIMPLE_SEGMENT|4582,4588|false|false|false|C0086805|Photons|photon
Event|Event|SIMPLE_SEGMENT|4596,4605|false|false|false|||involving
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4653,4659|false|false|false|C4522154|Distal Resection Margin|distal
Event|Event|SIMPLE_SEGMENT|4680,4686|false|false|false|||images
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4702,4713|false|false|false|C1980023|Wall motion|wall motion
Event|Event|SIMPLE_SEGMENT|4707,4713|false|false|false|||motion
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|4707,4713|false|false|false|C0026597|Motion|motion
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4721,4766|false|false|false|C4525750|Calculated Left Ventricular Ejection Fraction|calculated left ventricular ejection fraction
Finding|Functional Concept|SIMPLE_SEGMENT|4732,4736|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Finding|Physiologic Function|SIMPLE_SEGMENT|4732,4757|false|false|false|C2733342|Left ventricular ejection|left ventricular ejection
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4732,4766|false|false|false|C0428772;C0488728|Left ventricular ejection fraction|left ventricular ejection fraction
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4737,4748|false|false|false|C0018827|Heart Ventricle|ventricular
Finding|Physiologic Function|SIMPLE_SEGMENT|4737,4757|false|false|false|C2733340|Ventricular ejection|ventricular ejection
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4737,4766|false|false|false|C0042508|Ventricular Ejection Fraction|ventricular ejection fraction
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4749,4757|false|false|false|C0812388|Ejection time|ejection
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|4749,4757|false|false|false|C0336969|Ejection as a Sports activity|ejection
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|4749,4757|false|false|false|C0302131|Ejection as a Circumstance of Injury|ejection
Finding|Finding|SIMPLE_SEGMENT|4749,4766|false|false|false|C2020641;C2700378|Ejection fraction;stress echo measurements ejection fraction|ejection fraction
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4749,4766|false|false|false|C0489482|Ejection fraction (procedure)|ejection fraction
Event|Event|SIMPLE_SEGMENT|4758,4766|false|false|false|||fraction
Finding|Intellectual Product|SIMPLE_SEGMENT|4758,4766|false|false|false|C1554103|MDFAttributeType - Fraction|fraction
Event|Event|SIMPLE_SEGMENT|4783,4786|false|false|false|||EDV
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4783,4786|false|false|false|C2986747|End Diastolic Volume Imaging|EDV
Event|Event|SIMPLE_SEGMENT|4798,4809|false|false|false|||reprocessed
Event|Event|SIMPLE_SEGMENT|4829,4839|false|false|false|||IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|4829,4839|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|4829,4839|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Event|Event|SIMPLE_SEGMENT|4845,4855|false|false|false|||Reversible
Finding|Functional Concept|SIMPLE_SEGMENT|4845,4855|false|false|false|C0205343|Reversible|Reversible
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|4857,4863|false|false|false|C0010454;C1705217|Culture Media;Medium (Substance)|medium
Drug|Substance|SIMPLE_SEGMENT|4857,4863|false|false|false|C0010454;C1705217|Culture Media;Medium (Substance)|medium
Event|Event|SIMPLE_SEGMENT|4857,4863|false|false|false|||medium
Finding|Finding|SIMPLE_SEGMENT|4857,4863|false|false|false|C0009458;C4522282;C4522283|A Medium Amount;A Medium Amount of Time;Communications Media|medium
Finding|Intellectual Product|SIMPLE_SEGMENT|4857,4863|false|false|false|C0009458;C4522282;C4522283|A Medium Amount;A Medium Amount of Time;Communications Media|medium
Finding|Finding|SIMPLE_SEGMENT|4871,4879|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|SIMPLE_SEGMENT|4871,4879|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Event|Event|SIMPLE_SEGMENT|4889,4898|false|false|false|||perfusion
Finding|Functional Concept|SIMPLE_SEGMENT|4889,4898|false|false|false|C4281794;C4723760|Perfusion (biological);Perfusion route|perfusion
Finding|Organism Function|SIMPLE_SEGMENT|4889,4898|false|false|false|C4281794;C4723760|Perfusion (biological);Perfusion route|perfusion
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4889,4898|false|false|false|C0031001;C4721534|Chemotherapeutic Perfusion;Perfusion (procedure)|perfusion
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4899,4905|false|false|false|C1861101|THYROID HORMONE PLASMA MEMBRANE TRANSPORT DEFECT|defect
Event|Event|SIMPLE_SEGMENT|4899,4905|false|false|false|||defect
Finding|Functional Concept|SIMPLE_SEGMENT|4899,4905|false|false|false|C1457869|Defect|defect
Event|Event|SIMPLE_SEGMENT|4907,4916|false|false|false|||involving
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4921,4924|false|false|false|C2987138|Methylcytosine Dioxygenase TET1|LCx
Drug|Enzyme|SIMPLE_SEGMENT|4921,4924|false|false|false|C2987138|Methylcytosine Dioxygenase TET1|LCx
Finding|Gene or Genome|SIMPLE_SEGMENT|4921,4924|false|false|false|C1428863;C2987137|TET1 gene;TET1 wt Allele|LCx
Event|Event|SIMPLE_SEGMENT|4925,4934|false|false|false|||territory
Event|Event|SIMPLE_SEGMENT|4940,4949|false|false|false|||Increased
Finding|Functional Concept|SIMPLE_SEGMENT|4950,4954|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4950,4973|false|false|false|C0503990|Cavity of left ventricle|left ventricular cavity
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4950,4978|false|false|false|C0455830|Left ventricular cavity size|left ventricular cavity size
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4955,4966|false|false|false|C0018827|Heart Ventricle|ventricular
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4955,4973|false|false|false|C0507083|Cavity of ventricle|ventricular cavity
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4967,4973|false|false|false|C0333343|Body cavities|cavity
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|4967,4973|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4967,4973|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Event|Event|SIMPLE_SEGMENT|4974,4978|false|false|false|||size
Event|Event|SIMPLE_SEGMENT|4991,4999|false|false|false|||systolic
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|4991,4999|false|false|false|C0039155|Systole|systolic
Event|Event|SIMPLE_SEGMENT|5001,5009|false|false|false|||function
Finding|Finding|SIMPLE_SEGMENT|5001,5009|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|SIMPLE_SEGMENT|5001,5009|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|SIMPLE_SEGMENT|5001,5009|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|SIMPLE_SEGMENT|5001,5009|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Event|Event|SIMPLE_SEGMENT|5034,5039|false|false|false|||study
Finding|Intellectual Product|SIMPLE_SEGMENT|5034,5039|false|false|false|C1705923|Study Object|study
Procedure|Research Activity|SIMPLE_SEGMENT|5034,5039|false|false|false|C0008972;C0947630;C2603343|Clinical Research;Scientific Study;Study|study
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5052,5058|false|false|false|C1861101|THYROID HORMONE PLASMA MEMBRANE TRANSPORT DEFECT|defect
Event|Event|SIMPLE_SEGMENT|5052,5058|false|false|false|||defect
Finding|Functional Concept|SIMPLE_SEGMENT|5052,5058|false|false|false|C1457869|Defect|defect
Event|Event|SIMPLE_SEGMENT|5062,5065|false|false|false|||new
Finding|Finding|SIMPLE_SEGMENT|5062,5065|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|5062,5065|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5070,5077|false|false|false|C0018787|Heart|Cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|5070,5077|false|false|false|C1314974|Cardiac attachment|Cardiac
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|5070,5093|false|false|false|C0261588|Cardiac catheterisation as the cause of abnormal reaction of the patient, or of later complication, without mention of misadventure at the time of the procedure|Cardiac catheterization
Finding|Intellectual Product|SIMPLE_SEGMENT|5070,5093|false|false|false|C1547981|Diagnostic Service Section ID - Cardiac Catheterization|Cardiac catheterization
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5070,5093|false|false|false|C0018795;C1548828|Cardiac Catheterization Procedures;Consent Type - Cardiac Catheterization|Cardiac catheterization
Procedure|Health Care Activity|SIMPLE_SEGMENT|5070,5093|false|false|false|C0018795;C1548828|Cardiac Catheterization Procedures;Consent Type - Cardiac Catheterization|Cardiac catheterization
Event|Event|SIMPLE_SEGMENT|5078,5093|false|false|false|||catheterization
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5078,5093|false|false|false|C0007430|Catheterization|catheterization
Event|Event|SIMPLE_SEGMENT|5095,5103|false|false|false|||COMMENTS
Finding|Intellectual Product|SIMPLE_SEGMENT|5095,5103|false|false|false|C0282411;C0947611|Comment;Published Comment|COMMENTS
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5124,5132|false|false|false|C0018787|Heart|coronary
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5124,5144|false|false|false|C0085532;C1548829|Consent Type - Coronary Angiography;Coronary angiography|coronary angiography
Procedure|Health Care Activity|SIMPLE_SEGMENT|5124,5144|false|false|false|C0085532;C1548829|Consent Type - Coronary Angiography;Coronary angiography|coronary angiography
Event|Event|SIMPLE_SEGMENT|5133,5144|false|false|false|||angiography
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5133,5144|false|false|false|C0002978|angiogram|angiography
Finding|Functional Concept|SIMPLE_SEGMENT|5153,5158|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Finding|Functional Concept|SIMPLE_SEGMENT|5159,5167|false|false|false|C1527180|Dominant|dominant
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5168,5174|false|false|false|C5671121|System (basic dose form)|system
Event|Event|SIMPLE_SEGMENT|5168,5174|false|false|false|||system
Finding|Functional Concept|SIMPLE_SEGMENT|5168,5174|false|false|false|C0449913;C5441654|System;System, LOINC Axis 4|system
Event|Event|SIMPLE_SEGMENT|5176,5188|false|false|false|||demonstrated
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5195,5201|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5195,5201|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5195,5210|false|false|false|C0010075|Coronary Vessels|vessel coronary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5202,5210|false|false|false|C0018787|Heart|coronary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5202,5217|false|false|false|C0205042|Coronary artery|coronary artery
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5202,5225|false|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|coronary artery disease
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5211,5217|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|SIMPLE_SEGMENT|5211,5217|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5211,5225|false|false|false|C0852949|Arteriopathic disease|artery disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5218,5225|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|5218,5225|false|false|false|||disease
Finding|Idea or Concept|SIMPLE_SEGMENT|5268,5276|false|false|false|C0750489|apparent|apparent
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|5277,5281|false|false|false|C0806140|Flow|flow
Event|Event|SIMPLE_SEGMENT|5291,5299|false|false|false|||stenoses
Finding|Pathologic Function|SIMPLE_SEGMENT|5291,5299|false|false|false|C1261287|Stenosis|stenoses
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5306,5309|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5306,5309|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|SIMPLE_SEGMENT|5306,5309|false|false|false|||LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|5306,5309|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Finding|Pathologic Function|SIMPLE_SEGMENT|5323,5339|false|false|false|C3272317|Stent restenosis|stent restenosis
Event|Event|SIMPLE_SEGMENT|5329,5339|false|false|false|||restenosis
Finding|Pathologic Function|SIMPLE_SEGMENT|5329,5339|false|false|false|C0333186|Restenosis|restenosis
Finding|Gene or Genome|SIMPLE_SEGMENT|5367,5373|false|false|false|C1423674;C5890874|LDB3 gene;LDB3 wt Allele|Cypher
Event|Event|SIMPLE_SEGMENT|5374,5379|false|false|false|||stent
Event|Event|SIMPLE_SEGMENT|5381,5387|false|false|false|||placed
Finding|Finding|SIMPLE_SEGMENT|5404,5407|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|5404,5407|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Event|Event|SIMPLE_SEGMENT|5415,5420|false|false|false|||stent
Event|Event|SIMPLE_SEGMENT|5421,5427|false|false|false|||placed
Drug|Chemical Viewed Structurally|SIMPLE_SEGMENT|5442,5448|false|false|false|C1881507|Macromolecular Branch|branch
Event|Event|SIMPLE_SEGMENT|5442,5448|false|false|false|||branch
Finding|Classification|SIMPLE_SEGMENT|5471,5477|false|false|false|C0079946;C1550512|National origin;Participation Type - origin|origin
Finding|Intellectual Product|SIMPLE_SEGMENT|5471,5477|false|false|false|C0079946;C1550512|National origin;Participation Type - origin|origin
Event|Event|SIMPLE_SEGMENT|5478,5486|false|false|false|||stenosis
Finding|Pathologic Function|SIMPLE_SEGMENT|5478,5486|false|false|false|C1261287|Stenosis|stenosis
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5493,5496|false|false|false|C2987138|Methylcytosine Dioxygenase TET1|LCx
Drug|Enzyme|SIMPLE_SEGMENT|5493,5496|false|false|false|C2987138|Methylcytosine Dioxygenase TET1|LCx
Finding|Gene or Genome|SIMPLE_SEGMENT|5493,5496|false|false|false|C1428863;C2987137|TET1 gene;TET1 wt Allele|LCx
Event|Event|SIMPLE_SEGMENT|5507,5515|false|false|false|||stenosis
Finding|Pathologic Function|SIMPLE_SEGMENT|5507,5515|false|false|false|C1261287|Stenosis|stenosis
Event|Event|SIMPLE_SEGMENT|5524,5530|false|false|false|||origin
Finding|Classification|SIMPLE_SEGMENT|5524,5530|false|false|false|C0079946;C1550512|National origin;Participation Type - origin|origin
Finding|Intellectual Product|SIMPLE_SEGMENT|5524,5530|false|false|false|C0079946;C1550512|National origin;Participation Type - origin|origin
Event|Event|SIMPLE_SEGMENT|5549,5557|false|false|false|||stenosis
Finding|Pathologic Function|SIMPLE_SEGMENT|5549,5557|false|false|false|C1261287|Stenosis|stenosis
Drug|Chemical Viewed Structurally|SIMPLE_SEGMENT|5569,5575|false|false|false|C1881507|Macromolecular Branch|branch
Event|Event|SIMPLE_SEGMENT|5569,5575|false|false|false|||branch
Event|Event|SIMPLE_SEGMENT|5602,5610|false|false|false|||stenosis
Finding|Pathologic Function|SIMPLE_SEGMENT|5602,5610|false|false|false|C1261287|Stenosis|stenosis
Finding|Functional Concept|SIMPLE_SEGMENT|5616,5623|false|false|false|C0439801;C3542948|Limited (extensiveness);Limited component (foundation metadata concept)|Limited
Finding|Intellectual Product|SIMPLE_SEGMENT|5616,5623|false|false|false|C0439801;C3542948|Limited (extensiveness);Limited component (foundation metadata concept)|Limited
Event|Event|SIMPLE_SEGMENT|5632,5644|false|false|false|||hemodynamics
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|5632,5644|false|false|false|C0019010|Hemodynamics|hemodynamics
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5632,5644|false|false|false|C4281788|hemodynamics (procedure)|hemodynamics
Event|Event|SIMPLE_SEGMENT|5645,5653|false|false|false|||revealed
Finding|Intellectual Product|SIMPLE_SEGMENT|5654,5658|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Functional Concept|SIMPLE_SEGMENT|5659,5667|false|false|false|C0205373;C5849094|Systemic;Systemic Route of Administration|systemic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5668,5676|false|false|false|C0003842|Arteries|arterial
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5678,5690|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|SIMPLE_SEGMENT|5678,5690|false|false|false|||hypertension
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5699,5706|false|false|false|C0719205|Central brand of multivitamin with minerals|central
Drug|Vitamin|SIMPLE_SEGMENT|5699,5706|false|false|false|C0719205|Central brand of multivitamin with minerals|central
Event|Event|SIMPLE_SEGMENT|5699,5706|false|false|false|||central
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5699,5706|false|false|false|C1879652|Central Minus|central
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5707,5713|false|false|false|C0003483|Aorta|aortic
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5707,5722|false|false|false|C0456180|Aortic Pressure|aortic pressure
Event|Event|SIMPLE_SEGMENT|5714,5722|false|false|false|||pressure
Finding|Finding|SIMPLE_SEGMENT|5714,5722|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|SIMPLE_SEGMENT|5714,5722|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|5714,5722|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|5714,5722|false|false|false|C0033095||pressure
Finding|Social Behavior|SIMPLE_SEGMENT|5743,5753|false|false|false|C0597535|Success|Successful
Event|Event|SIMPLE_SEGMENT|5754,5758|false|false|false|||PTCA
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5754,5758|false|false|false|C2936173|Percutaneous Transluminal Coronary Angioplasty|PTCA
Event|Event|SIMPLE_SEGMENT|5763,5771|false|false|false|||stenting
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5763,5771|false|false|false|C2348535|Stenting|stenting
Event|Event|SIMPLE_SEGMENT|5795,5801|false|false|false|||PROMUS
Event|Event|SIMPLE_SEGMENT|5820,5831|false|false|false|||postdilated
Finding|Idea or Concept|SIMPLE_SEGMENT|5842,5847|false|false|false|C1546485|Diagnosis Type - Final|Final
Event|Event|SIMPLE_SEGMENT|5848,5859|false|false|false|||angiography
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5848,5859|false|false|false|C0002978|angiogram|angiography
Event|Event|SIMPLE_SEGMENT|5860,5868|false|false|false|||revealed
Event|Event|SIMPLE_SEGMENT|5883,5891|false|false|false|||stenosis
Finding|Pathologic Function|SIMPLE_SEGMENT|5883,5891|false|false|false|C1261287|Stenosis|stenosis
Finding|Idea or Concept|SIMPLE_SEGMENT|5913,5921|false|false|false|C0750489|apparent|apparent
Event|Event|SIMPLE_SEGMENT|5922,5932|false|false|false|||dissection
Finding|Pathologic Function|SIMPLE_SEGMENT|5922,5932|false|false|false|C0333288|Dissecting hemorrhage|dissection
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5922,5932|false|false|false|C0012737|Tissue Dissection|dissection
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|5947,5951|false|false|false|C0806140|Flow|flow
Event|Activity|SIMPLE_SEGMENT|5953,5956|false|false|false|C1947903|See|see
Finding|Organism Function|SIMPLE_SEGMENT|5953,5956|false|false|false|C0042789|Vision|see
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5958,5962|false|false|false|C2936173|Percutaneous Transluminal Coronary Angioplasty|PTCA
Event|Event|SIMPLE_SEGMENT|5963,5971|false|false|false|||comments
Finding|Intellectual Product|SIMPLE_SEGMENT|5963,5971|false|false|false|C0282411;C0947611|Comment;Published Comment|comments
Finding|Idea or Concept|SIMPLE_SEGMENT|5975,5980|false|false|false|C1546485|Diagnosis Type - Final|FINAL
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5981,5990|false|false|false|C0945731||DIAGNOSIS
Event|Event|SIMPLE_SEGMENT|5981,5990|false|false|false|||DIAGNOSIS
Finding|Classification|SIMPLE_SEGMENT|5981,5990|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|DIAGNOSIS
Finding|Functional Concept|SIMPLE_SEGMENT|5981,5990|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|DIAGNOSIS
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5981,5990|false|false|false|C0011900|Diagnosis|DIAGNOSIS
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6006,6012|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6006,6012|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6006,6021|false|false|false|C0010075|Coronary Vessels|vessel coronary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6013,6021|false|false|false|C0018787|Heart|coronary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6013,6028|false|false|false|C0205042|Coronary artery|coronary artery
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6013,6036|false|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|coronary artery disease
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6022,6028|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|SIMPLE_SEGMENT|6022,6028|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6022,6036|false|false|false|C0852949|Arteriopathic disease|artery disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6029,6036|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|6029,6036|false|false|false|||disease
Finding|Social Behavior|SIMPLE_SEGMENT|6042,6052|false|false|false|C0597535|Success|Successful
Event|Event|SIMPLE_SEGMENT|6053,6057|false|false|false|||PTCA
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6053,6057|false|false|false|C2936173|Percutaneous Transluminal Coronary Angioplasty|PTCA
Event|Event|SIMPLE_SEGMENT|6062,6070|false|false|false|||stenting
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6062,6070|false|false|false|C2348535|Stenting|stenting
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6089,6092|false|false|false|C4551552|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|DES
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6089,6092|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6089,6092|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Hormone|SIMPLE_SEGMENT|6089,6092|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Organic Chemical|SIMPLE_SEGMENT|6089,6092|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6089,6092|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Event|Event|SIMPLE_SEGMENT|6089,6092|false|false|false|||DES
Finding|Gene or Genome|SIMPLE_SEGMENT|6089,6092|false|false|false|C1413980|DES gene|DES
Finding|Intellectual Product|SIMPLE_SEGMENT|6100,6105|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|Brief
Finding|Idea or Concept|SIMPLE_SEGMENT|6106,6114|false|false|false|C1547192|Organization unit type - Hospital|Hospital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6106,6121|false|false|false|C0488549||Hospital Course
Finding|Finding|SIMPLE_SEGMENT|6106,6121|false|false|false|C0489547|Hospital course|Hospital Course
Finding|Finding|SIMPLE_SEGMENT|6125,6133|false|false|false|C0443343|Unstable status|Unstable
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6125,6140|false|false|false|C0002965|Angina, Unstable|Unstable angina
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6134,6140|false|false|false|C2926611||angina
Event|Event|SIMPLE_SEGMENT|6134,6140|false|false|false|||angina
Finding|Finding|SIMPLE_SEGMENT|6134,6140|false|false|false|C0002962;C2024883|Angina Pectoris|angina
Finding|Sign or Symptom|SIMPLE_SEGMENT|6134,6140|false|false|false|C0002962;C2024883|Angina Pectoris|angina
Event|Event|SIMPLE_SEGMENT|6142,6153|false|false|false|||Description
Finding|Intellectual Product|SIMPLE_SEGMENT|6142,6153|false|false|false|C0678257|Description|Description
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6161,6165|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|6161,6165|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|6161,6165|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|6161,6165|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|SIMPLE_SEGMENT|6170,6178|false|false|false|C2984079|Somewhat|somewhat
Event|Event|SIMPLE_SEGMENT|6179,6187|false|false|false|||atypical
Finding|Finding|SIMPLE_SEGMENT|6179,6187|false|false|false|C0741302|atypia morphology|atypical
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6193,6199|false|false|false|C2926611||angina
Event|Event|SIMPLE_SEGMENT|6193,6199|false|false|false|||angina
Finding|Finding|SIMPLE_SEGMENT|6193,6199|false|false|false|C0002962;C2024883|Angina Pectoris|angina
Finding|Sign or Symptom|SIMPLE_SEGMENT|6193,6199|false|false|false|C0002962;C2024883|Angina Pectoris|angina
Event|Event|SIMPLE_SEGMENT|6212,6223|false|false|false|||experiences
Event|Event|SIMPLE_SEGMENT|6236,6240|false|false|false|||lays
Event|Event|SIMPLE_SEGMENT|6262,6274|false|false|false|||reproducible
Event|Event|SIMPLE_SEGMENT|6295,6302|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|6295,6302|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|6295,6302|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|6295,6302|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|6295,6305|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6306,6309|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6306,6309|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|6306,6309|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|6306,6309|false|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|6306,6309|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6306,6309|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|6306,6309|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6306,6309|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6310,6316|false|false|false|C5889824||status
Event|Event|SIMPLE_SEGMENT|6310,6316|false|false|false|||status
Finding|Idea or Concept|SIMPLE_SEGMENT|6310,6316|false|false|false|C1546481|What subject filter - Status|status
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|6332,6336|false|false|false|C0228147|Structure of cisterna pontis|PCIs
Finding|Idea or Concept|SIMPLE_SEGMENT|6346,6350|false|false|false|C0035647|Risk|risk
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6346,6358|false|false|false|C1830376||risk factors
Finding|Finding|SIMPLE_SEGMENT|6346,6358|false|false|false|C0035648;C0455624;C1553898|History of - risk factor;risk factors;risk factors - observation list|risk factors
Finding|Intellectual Product|SIMPLE_SEGMENT|6346,6358|false|false|false|C0035648;C0455624;C1553898|History of - risk factor;risk factors;risk factors - observation list|risk factors
Event|Event|SIMPLE_SEGMENT|6351,6358|false|false|false|||factors
Finding|Body Substance|SIMPLE_SEGMENT|6364,6371|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|6364,6371|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|6364,6371|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6383,6389|false|false|false|C1718621|W stress|stress
Drug|Organic Chemical|SIMPLE_SEGMENT|6383,6389|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6383,6389|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Event|Event|SIMPLE_SEGMENT|6383,6389|false|false|false|||stress
Finding|Finding|SIMPLE_SEGMENT|6383,6389|false|false|false|C0038435|Stress|stress
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6383,6394|false|false|false|C0015260;C3494508|Exercise stress test;Stress Test|stress test
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6390,6394|false|false|false|C4318744|Test - temporal region|test
Event|Event|SIMPLE_SEGMENT|6390,6394|false|false|false|||test
Finding|Functional Concept|SIMPLE_SEGMENT|6390,6394|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Finding|Intellectual Product|SIMPLE_SEGMENT|6390,6394|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6390,6394|false|false|false|C0456984|Test Result|test
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6390,6394|false|false|false|C0022885|Laboratory Procedures|test
Event|Event|SIMPLE_SEGMENT|6398,6402|false|false|false|||rule
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6407,6410|false|true|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6407,6410|false|true|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|6407,6410|false|true|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|6407,6410|false|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|6407,6410|false|true|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6407,6410|false|true|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|6407,6410|false|true|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6407,6410|false|true|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6412,6431|false|false|false|C2825165|Nuclear stress test|Nuclear stress test
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6420,6426|false|false|false|C1718621|W stress|stress
Drug|Organic Chemical|SIMPLE_SEGMENT|6420,6426|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6420,6426|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Finding|Finding|SIMPLE_SEGMENT|6420,6426|false|false|false|C0038435|Stress|stress
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6420,6431|false|false|false|C0015260;C3494508|Exercise stress test;Stress Test|stress test
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6427,6431|false|false|false|C4318744|Test - temporal region|test
Event|Event|SIMPLE_SEGMENT|6427,6431|false|false|false|||test
Finding|Functional Concept|SIMPLE_SEGMENT|6427,6431|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Finding|Intellectual Product|SIMPLE_SEGMENT|6427,6431|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6427,6431|false|false|false|C0456984|Test Result|test
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6427,6431|false|false|false|C0022885|Laboratory Procedures|test
Event|Event|SIMPLE_SEGMENT|6432,6438|false|false|false|||showed
Event|Event|SIMPLE_SEGMENT|6442,6452|false|false|false|||reversible
Finding|Functional Concept|SIMPLE_SEGMENT|6442,6452|false|false|false|C0205343|Reversible|reversible
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|6454,6460|false|false|false|C0010454;C1705217|Culture Media;Medium (Substance)|medium
Drug|Substance|SIMPLE_SEGMENT|6454,6460|false|false|false|C0010454;C1705217|Culture Media;Medium (Substance)|medium
Event|Event|SIMPLE_SEGMENT|6454,6460|false|false|false|||medium
Finding|Finding|SIMPLE_SEGMENT|6454,6460|false|false|false|C0009458;C4522282;C4522283|A Medium Amount;A Medium Amount of Time;Communications Media|medium
Finding|Intellectual Product|SIMPLE_SEGMENT|6454,6460|false|false|false|C0009458;C4522282;C4522283|A Medium Amount;A Medium Amount of Time;Communications Media|medium
Finding|Finding|SIMPLE_SEGMENT|6468,6476|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|SIMPLE_SEGMENT|6468,6476|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Event|Event|SIMPLE_SEGMENT|6486,6495|false|false|false|||perfusion
Finding|Functional Concept|SIMPLE_SEGMENT|6486,6495|false|false|false|C4281794;C4723760|Perfusion (biological);Perfusion route|perfusion
Finding|Organism Function|SIMPLE_SEGMENT|6486,6495|false|false|false|C4281794;C4723760|Perfusion (biological);Perfusion route|perfusion
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6486,6495|false|false|false|C0031001;C4721534|Chemotherapeutic Perfusion;Perfusion (procedure)|perfusion
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6496,6502|false|false|false|C1861101|THYROID HORMONE PLASMA MEMBRANE TRANSPORT DEFECT|defect
Event|Event|SIMPLE_SEGMENT|6496,6502|false|false|false|||defect
Finding|Functional Concept|SIMPLE_SEGMENT|6496,6502|false|false|false|C1457869|Defect|defect
Event|Event|SIMPLE_SEGMENT|6504,6513|false|false|false|||involving
Finding|Functional Concept|SIMPLE_SEGMENT|6518,6522|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Event|Event|SIMPLE_SEGMENT|6534,6543|false|false|false|||territory
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6548,6553|false|false|false|C1570446|TNFSF14 protein, human|light
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6548,6553|false|false|false|C1570446|TNFSF14 protein, human|light
Event|Event|SIMPLE_SEGMENT|6548,6553|false|false|false|||light
Finding|Finding|SIMPLE_SEGMENT|6548,6553|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Functional Concept|SIMPLE_SEGMENT|6548,6553|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Gene or Genome|SIMPLE_SEGMENT|6548,6553|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|6548,6553|false|false|false|C0023693|Light|light
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6548,6553|false|false|false|C0031765|Phototherapy|light
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6564,6570|false|false|false|C1718621|W stress|stress
Drug|Organic Chemical|SIMPLE_SEGMENT|6564,6570|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6564,6570|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Event|Event|SIMPLE_SEGMENT|6564,6570|false|false|false|||stress
Finding|Finding|SIMPLE_SEGMENT|6564,6570|false|false|false|C0038435|Stress|stress
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6564,6575|false|false|false|C0015260;C3494508|Exercise stress test;Stress Test|stress test
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6571,6575|false|false|false|C4318744|Test - temporal region|test
Finding|Functional Concept|SIMPLE_SEGMENT|6571,6575|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Finding|Intellectual Product|SIMPLE_SEGMENT|6571,6575|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6571,6575|false|false|false|C0456984|Test Result|test
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6571,6575|false|false|false|C0022885|Laboratory Procedures|test
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6576,6584|false|false|false|C2926606||findings
Event|Event|SIMPLE_SEGMENT|6576,6584|false|false|false|||findings
Finding|Functional Concept|SIMPLE_SEGMENT|6576,6584|false|false|false|C2607943|findings aspects|findings
Finding|Body Substance|SIMPLE_SEGMENT|6590,6597|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|6590,6597|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|6590,6597|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6608,6615|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|6608,6615|false|false|false|C1314974|Cardiac attachment|cardiac
Event|Event|SIMPLE_SEGMENT|6617,6632|false|false|false|||catheterization
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6617,6632|false|false|false|C0007430|Catheterization|catheterization
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6643,6650|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|6643,6650|false|false|false|C1314974|Cardiac attachment|cardiac
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|6643,6666|false|false|false|C0261588|Cardiac catheterisation as the cause of abnormal reaction of the patient, or of later complication, without mention of misadventure at the time of the procedure|cardiac catheterization
Finding|Intellectual Product|SIMPLE_SEGMENT|6643,6666|false|false|false|C1547981|Diagnostic Service Section ID - Cardiac Catheterization|cardiac catheterization
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6643,6666|false|false|false|C0018795;C1548828|Cardiac Catheterization Procedures;Consent Type - Cardiac Catheterization|cardiac catheterization
Procedure|Health Care Activity|SIMPLE_SEGMENT|6643,6666|false|false|false|C0018795;C1548828|Cardiac Catheterization Procedures;Consent Type - Cardiac Catheterization|cardiac catheterization
Event|Event|SIMPLE_SEGMENT|6651,6666|false|false|false|||catheterization
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6651,6666|false|false|false|C0007430|Catheterization|catheterization
Event|Event|SIMPLE_SEGMENT|6677,6688|false|false|false|||prehydrated
Finding|Intellectual Product|SIMPLE_SEGMENT|6699,6704|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6699,6718|false|false|false|C0022660;C2609414|Acute kidney injury;Kidney Failure, Acute|acute kidney injury
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|6699,6718|false|false|false|C0022660;C2609414|Acute kidney injury;Kidney Failure, Acute|acute kidney injury
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6705,6711|false|false|false|C0022646;C0227665|Both kidneys;Kidney|kidney
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6705,6711|false|false|false|C0496892;C0496927|Benign neoplasm of kidney;Neoplasm of uncertain or unknown behavior of kidney|kidney
Event|Event|SIMPLE_SEGMENT|6705,6711|false|false|false|||kidney
Finding|Sign or Symptom|SIMPLE_SEGMENT|6705,6711|false|false|false|C0812426|Kidney problem|kidney
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6705,6711|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6705,6711|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|6705,6718|false|false|false|C0160420|Injury of kidney|kidney injury
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|6712,6718|false|false|false|C3263722;C3263723|Traumatic AND/OR non-traumatic injury;Traumatic injury|injury
Event|Event|SIMPLE_SEGMENT|6712,6718|false|false|false|||injury
Finding|Body Substance|SIMPLE_SEGMENT|6724,6731|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|6724,6731|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|6724,6731|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6739,6743|false|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|drug
Event|Event|SIMPLE_SEGMENT|6739,6743|false|false|false|||drug
Finding|Finding|SIMPLE_SEGMENT|6739,6743|false|false|false|C0740721|Drug problem|drug
Event|Event|SIMPLE_SEGMENT|6752,6757|false|false|false|||stent
Event|Event|SIMPLE_SEGMENT|6758,6764|false|false|false|||placed
Finding|Finding|SIMPLE_SEGMENT|6779,6787|false|false|false|C1550517|Target Awareness - marginal|marginal
Drug|Chemical Viewed Structurally|SIMPLE_SEGMENT|6788,6794|false|false|false|C1881507|Macromolecular Branch|branch
Event|Event|SIMPLE_SEGMENT|6788,6794|false|false|false|||branch
Finding|Body Substance|SIMPLE_SEGMENT|6801,6808|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|6801,6808|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|6801,6808|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|6809,6815|false|false|false|||became
Event|Event|SIMPLE_SEGMENT|6824,6836|false|false|false|||hypertensive
Finding|Finding|SIMPLE_SEGMENT|6824,6836|false|false|false|C0857121|Hypertensive (finding)|hypertensive
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6844,6851|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|6844,6851|false|false|false|C1314974|Cardiac attachment|cardiac
Event|Event|SIMPLE_SEGMENT|6853,6868|false|false|false|||catheterization
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6853,6868|false|false|false|C0007430|Catheterization|catheterization
Event|Event|SIMPLE_SEGMENT|6877,6884|false|false|false|||started
Drug|Organic Chemical|SIMPLE_SEGMENT|6890,6903|false|false|false|C0017887|nitroglycerin|nitroglycerin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6890,6903|false|false|false|C0017887|nitroglycerin|nitroglycerin
Event|Event|SIMPLE_SEGMENT|6904,6908|false|false|false|||drip
Event|Event|SIMPLE_SEGMENT|6910,6913|false|false|false|||see
Event|Event|SIMPLE_SEGMENT|6915,6925|false|false|false|||discussion
Finding|Social Behavior|SIMPLE_SEGMENT|6915,6925|false|false|false|C2584313|Discussion (communication)|discussion
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6915,6925|false|false|false|C0557061|Discussion (procedure)|discussion
Finding|Body Substance|SIMPLE_SEGMENT|6938,6945|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|6938,6945|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|6938,6945|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|6950,6956|false|false|false|||weaned
Finding|Body Substance|SIMPLE_SEGMENT|6981,6988|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|6981,6988|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|6981,6988|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|6993,7002|false|false|false|||continued
Drug|Organic Chemical|SIMPLE_SEGMENT|7006,7013|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7006,7013|false|false|false|C0004057|aspirin|aspirin
Event|Event|SIMPLE_SEGMENT|7006,7013|false|false|false|||aspirin
Drug|Organic Chemical|SIMPLE_SEGMENT|7027,7033|false|false|false|C0633084|Plavix|plavix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7027,7033|false|false|false|C0633084|Plavix|plavix
Event|Event|SIMPLE_SEGMENT|7027,7033|false|false|false|||plavix
Drug|Organic Chemical|SIMPLE_SEGMENT|7036,7046|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7036,7046|false|false|false|C0025859|metoprolol|metoprolol
Event|Event|SIMPLE_SEGMENT|7036,7046|false|false|false|||metoprolol
Drug|Organic Chemical|SIMPLE_SEGMENT|7052,7057|false|false|false|C0590690|Imdur|imdur
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7052,7057|false|false|false|C0590690|Imdur|imdur
Event|Event|SIMPLE_SEGMENT|7052,7057|false|false|false|||imdur
Finding|Idea or Concept|SIMPLE_SEGMENT|7063,7067|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|7063,7067|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|7063,7067|false|false|false|C1553498|home health encounter|home
Event|Event|SIMPLE_SEGMENT|7068,7072|false|false|false|||dose
Drug|Organic Chemical|SIMPLE_SEGMENT|7076,7088|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7076,7088|false|false|false|C0286651|atorvastatin|atorvastatin
Event|Event|SIMPLE_SEGMENT|7076,7088|false|false|false|||atorvastatin
Event|Event|SIMPLE_SEGMENT|7094,7103|false|false|false|||increased
Event|Event|SIMPLE_SEGMENT|7110,7118|false|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|7110,7118|false|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|7110,7121|false|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7122,7130|false|false|false|C0018787|Heart|coronary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7122,7137|false|false|false|C0205042|Coronary artery|coronary artery
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7122,7145|false|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|coronary artery disease
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7131,7137|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|SIMPLE_SEGMENT|7131,7137|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7131,7145|false|false|false|C0852949|Arteriopathic disease|artery disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7138,7145|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|7138,7145|false|false|false|||disease
Finding|Intellectual Product|SIMPLE_SEGMENT|7147,7153|false|false|false|C0031082|Periodicals|Serial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7155,7162|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|7155,7162|false|false|false|C1314974|Cardiac attachment|cardiac
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7155,7170|false|false|false|C2926589||cardiac enzymes
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7155,7170|false|false|false|C0443763|Cardiac enzymes|cardiac enzymes
Drug|Enzyme|SIMPLE_SEGMENT|7155,7170|false|false|false|C0443763|Cardiac enzymes|cardiac enzymes
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7155,7170|false|false|false|C0201934|Cardiac enzymes/isoenzymes measurement|cardiac enzymes
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7163,7170|false|false|false|C0014442;C3540017;C3540048;C3540772;C3540790;C3541394;C3542456|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS;Enzymes;Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM;Enzymes for ALIMENTARY TRACT AND METABOLISM;Enzymes, antithrombotic;Enzymes, hematological;Enzymes, peripheral vasodilators|enzymes
Drug|Enzyme|SIMPLE_SEGMENT|7163,7170|false|false|false|C0014442;C3540017;C3540048;C3540772;C3540790;C3541394;C3542456|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS;Enzymes;Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM;Enzymes for ALIMENTARY TRACT AND METABOLISM;Enzymes, antithrombotic;Enzymes, hematological;Enzymes, peripheral vasodilators|enzymes
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7163,7170|false|false|false|C0014442;C3540017;C3540048;C3540772;C3540790;C3541394;C3542456|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS;Enzymes;Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM;Enzymes for ALIMENTARY TRACT AND METABOLISM;Enzymes, antithrombotic;Enzymes, hematological;Enzymes, peripheral vasodilators|enzymes
Event|Event|SIMPLE_SEGMENT|7163,7170|false|false|false|||enzymes
Finding|Functional Concept|SIMPLE_SEGMENT|7163,7170|false|false|false|C0014445|enzymology|enzymes
Event|Event|SIMPLE_SEGMENT|7176,7184|false|false|false|||negative
Finding|Classification|SIMPLE_SEGMENT|7176,7184|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|7176,7184|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|7176,7184|false|false|false|C5237010|Expression Negative|negative
Finding|Classification|SIMPLE_SEGMENT|7197,7207|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|OUTPATIENT
Finding|Idea or Concept|SIMPLE_SEGMENT|7197,7207|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|OUTPATIENT
Event|Event|SIMPLE_SEGMENT|7208,7214|false|false|false|||ISSUES
Finding|Body Substance|SIMPLE_SEGMENT|7216,7223|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|7216,7223|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|7216,7223|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|7230,7238|false|false|false|||continue
Drug|Organic Chemical|SIMPLE_SEGMENT|7246,7253|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7246,7253|false|false|false|C0004057|aspirin|aspirin
Event|Event|SIMPLE_SEGMENT|7246,7253|false|false|false|||aspirin
Drug|Organic Chemical|SIMPLE_SEGMENT|7265,7271|false|false|false|C0633084|Plavix|plavix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7265,7271|false|false|false|C0633084|Plavix|plavix
Finding|Idea or Concept|SIMPLE_SEGMENT|7291,7295|false|false|false|C1552851|next - HtmlLinkType|next
Finding|Idea or Concept|SIMPLE_SEGMENT|7296,7300|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|SIMPLE_SEGMENT|7296,7300|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Body Substance|SIMPLE_SEGMENT|7302,7309|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|7302,7309|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|7302,7309|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Anatomy|Body System|SIMPLE_SEGMENT|7321,7331|false|false|false|C0007226|Cardiovascular system|cardiology
Event|Event|SIMPLE_SEGMENT|7332,7338|false|false|false|||follow
Finding|Functional Concept|SIMPLE_SEGMENT|7332,7338|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|SIMPLE_SEGMENT|7332,7338|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|SIMPLE_SEGMENT|7332,7341|false|false|false|C0589120|Follow-up status|follow-up
Procedure|Health Care Activity|SIMPLE_SEGMENT|7332,7341|false|false|false|C1522577|follow-up|follow-up
Event|Event|SIMPLE_SEGMENT|7348,7358|false|false|false|||outpatient
Finding|Classification|SIMPLE_SEGMENT|7348,7358|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|7348,7358|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|SIMPLE_SEGMENT|7381,7386|false|false|false|||group
Finding|Body Substance|SIMPLE_SEGMENT|7381,7386|false|false|false|C0441833;C1519504;C1561557;C1705428|Group Object;Group Specimen;Groups;Stage Grouping|group
Finding|Conceptual Entity|SIMPLE_SEGMENT|7381,7386|false|false|false|C0441833;C1519504;C1561557;C1705428|Group Object;Group Specimen;Groups;Stage Grouping|group
Finding|Functional Concept|SIMPLE_SEGMENT|7381,7386|false|false|false|C0441833;C1519504;C1561557;C1705428|Group Object;Group Specimen;Groups;Stage Grouping|group
Finding|Idea or Concept|SIMPLE_SEGMENT|7381,7386|false|false|false|C0441833;C1519504;C1561557;C1705428|Group Object;Group Specimen;Groups;Stage Grouping|group
Finding|Intellectual Product|SIMPLE_SEGMENT|7402,7407|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|Acute
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7402,7421|false|false|false|C0022660;C2609414|Acute kidney injury;Kidney Failure, Acute|Acute kidney injury
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|7402,7421|false|false|false|C0022660;C2609414|Acute kidney injury;Kidney Failure, Acute|Acute kidney injury
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7408,7414|false|false|false|C0022646;C0227665|Both kidneys;Kidney|kidney
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7408,7414|false|false|false|C0496892;C0496927|Benign neoplasm of kidney;Neoplasm of uncertain or unknown behavior of kidney|kidney
Event|Event|SIMPLE_SEGMENT|7408,7414|false|false|false|||kidney
Finding|Sign or Symptom|SIMPLE_SEGMENT|7408,7414|false|false|false|C0812426|Kidney problem|kidney
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7408,7414|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7408,7414|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|7408,7421|false|false|false|C0160420|Injury of kidney|kidney injury
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|7415,7421|false|false|false|C3263722;C3263723|Traumatic AND/OR non-traumatic injury;Traumatic injury|injury
Event|Event|SIMPLE_SEGMENT|7415,7421|false|false|false|||injury
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7423,7433|false|false|false|C0010294|creatinine|Creatinine
Drug|Organic Chemical|SIMPLE_SEGMENT|7423,7433|false|false|false|C0010294|creatinine|Creatinine
Event|Event|SIMPLE_SEGMENT|7423,7433|false|false|false|||Creatinine
Finding|Physiologic Function|SIMPLE_SEGMENT|7423,7433|false|false|false|C4551889|Creatinine metabolic function|Creatinine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7423,7433|false|false|false|C0201975|Creatinine measurement|Creatinine
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7470,7475|false|false|false|C0022646|Kidney|Renal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7470,7475|false|false|false|C0042075|Urologic Diseases|Renal
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|7470,7484|false|false|false|C0232804|Renal function|Renal function
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7470,7484|false|false|false|C0022662|Kidney Function Tests|Renal function
Event|Event|SIMPLE_SEGMENT|7476,7484|false|false|false|||function
Finding|Finding|SIMPLE_SEGMENT|7476,7484|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|SIMPLE_SEGMENT|7476,7484|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|SIMPLE_SEGMENT|7476,7484|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|SIMPLE_SEGMENT|7476,7484|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Event|Event|SIMPLE_SEGMENT|7500,7506|false|false|false|||normal
Event|Event|SIMPLE_SEGMENT|7513,7522|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|7513,7522|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Body Substance|SIMPLE_SEGMENT|7529,7536|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|7529,7536|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|7529,7536|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7539,7549|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7539,7549|false|false|false|C0065374|lisinopril|lisinopril
Event|Event|SIMPLE_SEGMENT|7539,7549|false|false|false|||lisinopril
Drug|Organic Chemical|SIMPLE_SEGMENT|7554,7564|false|false|false|C0016860|furosemide|furosemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7554,7564|false|false|false|C0016860|furosemide|furosemide
Event|Event|SIMPLE_SEGMENT|7554,7564|false|false|false|||furosemide
Event|Event|SIMPLE_SEGMENT|7570,7582|false|false|false|||discontinued
Event|Event|SIMPLE_SEGMENT|7588,7592|false|false|false|||note
Finding|Gene or Genome|SIMPLE_SEGMENT|7594,7597|false|false|false|C1825832|ACOT8 gene|hte
Finding|Body Substance|SIMPLE_SEGMENT|7598,7605|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|7598,7605|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|7598,7605|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|7610,7617|false|false|false|||started
Drug|Organic Chemical|SIMPLE_SEGMENT|7621,7631|false|false|false|C0016860|furosemide|furosemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7621,7631|false|false|false|C0016860|furosemide|furosemide
Event|Event|SIMPLE_SEGMENT|7621,7631|false|false|false|||furosemide
Finding|Gene or Genome|SIMPLE_SEGMENT|7658,7661|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Event|Event|SIMPLE_SEGMENT|7669,7678|false|false|false|||coincides
Event|Event|SIMPLE_SEGMENT|7688,7699|false|false|false|||development
Finding|Functional Concept|SIMPLE_SEGMENT|7688,7699|false|false|false|C0018271;C0243107;C0678723;C1527148|Development;Growth and Development function;biological development;development aspects|development
Finding|Organism Function|SIMPLE_SEGMENT|7688,7699|false|false|false|C0018271;C0243107;C0678723;C1527148|Development;Growth and Development function;biological development;development aspects|development
Finding|Body Substance|SIMPLE_SEGMENT|7708,7715|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|7708,7715|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|7708,7715|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Finding|SIMPLE_SEGMENT|7718,7743|false|false|false|C0700225|Serum creatinine raised|elevated serum creatinine
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|7727,7732|false|false|false|C5575602|Cell Culture Serum|serum
Event|Event|SIMPLE_SEGMENT|7727,7732|false|false|false|||serum
Finding|Body Substance|SIMPLE_SEGMENT|7727,7732|false|false|false|C0229671;C1546774;C1550100|Serum;Serum specimen|serum
Finding|Intellectual Product|SIMPLE_SEGMENT|7727,7732|false|false|false|C0229671;C1546774;C1550100|Serum;Serum specimen|serum
Finding|Finding|SIMPLE_SEGMENT|7727,7743|false|false|false|C0600061|Serum creatinine level|serum creatinine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7727,7743|false|false|false|C0201976|Creatinine measurement, serum (procedure)|serum creatinine
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7733,7743|false|false|false|C0010294|creatinine|creatinine
Drug|Organic Chemical|SIMPLE_SEGMENT|7733,7743|false|false|false|C0010294|creatinine|creatinine
Event|Event|SIMPLE_SEGMENT|7733,7743|false|false|false|||creatinine
Finding|Physiologic Function|SIMPLE_SEGMENT|7733,7743|false|false|false|C4551889|Creatinine metabolic function|creatinine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7733,7743|false|false|false|C0201975|Creatinine measurement|creatinine
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|7745,7750|false|false|false|C5575602|Cell Culture Serum|Serum
Finding|Body Substance|SIMPLE_SEGMENT|7745,7750|false|false|false|C0229671;C1546774;C1550100|Serum;Serum specimen|Serum
Finding|Intellectual Product|SIMPLE_SEGMENT|7745,7750|false|false|false|C0229671;C1546774;C1550100|Serum;Serum specimen|Serum
Finding|Finding|SIMPLE_SEGMENT|7745,7761|false|false|false|C0600061|Serum creatinine level|Serum creatinine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7745,7761|false|false|false|C0201976|Creatinine measurement, serum (procedure)|Serum creatinine
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7751,7761|false|false|false|C0010294|creatinine|creatinine
Drug|Organic Chemical|SIMPLE_SEGMENT|7751,7761|false|false|false|C0010294|creatinine|creatinine
Event|Event|SIMPLE_SEGMENT|7751,7761|false|false|false|||creatinine
Finding|Physiologic Function|SIMPLE_SEGMENT|7751,7761|false|false|false|C4551889|Creatinine metabolic function|creatinine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7751,7761|false|false|false|C0201975|Creatinine measurement|creatinine
Event|Event|SIMPLE_SEGMENT|7767,7774|false|false|false|||trended
Event|Event|SIMPLE_SEGMENT|7787,7796|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|7787,7796|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|SIMPLE_SEGMENT|7801,7809|false|false|false|||improved
Finding|Body Substance|SIMPLE_SEGMENT|7815,7822|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|7815,7822|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|7815,7822|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|7828,7837|false|false|false|||restarted
Finding|Idea or Concept|SIMPLE_SEGMENT|7845,7849|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|7845,7849|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|7845,7849|false|false|false|C1553498|home health encounter|home
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7850,7860|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7850,7860|false|false|false|C0065374|lisinopril|lisinopril
Event|Event|SIMPLE_SEGMENT|7850,7860|false|false|false|||lisinopril
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|7873,7878|false|false|false|C5575602|Cell Culture Serum|serum
Finding|Body Substance|SIMPLE_SEGMENT|7873,7878|false|false|false|C0229671;C1546774;C1550100|Serum;Serum specimen|serum
Finding|Intellectual Product|SIMPLE_SEGMENT|7873,7878|false|false|false|C0229671;C1546774;C1550100|Serum;Serum specimen|serum
Finding|Finding|SIMPLE_SEGMENT|7873,7889|false|false|false|C0600061|Serum creatinine level|serum creatinine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7873,7889|false|false|false|C0201976|Creatinine measurement, serum (procedure)|serum creatinine
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7879,7889|false|false|false|C0010294|creatinine|creatinine
Drug|Organic Chemical|SIMPLE_SEGMENT|7879,7889|false|false|false|C0010294|creatinine|creatinine
Event|Event|SIMPLE_SEGMENT|7879,7889|false|false|false|||creatinine
Finding|Physiologic Function|SIMPLE_SEGMENT|7879,7889|false|false|false|C4551889|Creatinine metabolic function|creatinine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7879,7889|false|false|false|C0201975|Creatinine measurement|creatinine
Event|Event|SIMPLE_SEGMENT|7895,7902|false|false|false|||noticed
Event|Event|SIMPLE_SEGMENT|7909,7919|false|false|false|||increasing
Event|Event|SIMPLE_SEGMENT|7927,7939|false|false|false|||discontinued
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7946,7958|false|false|false|C3263700||instructions
Event|Event|SIMPLE_SEGMENT|7946,7958|false|false|false|||instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|7946,7958|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|instructions
Event|Event|SIMPLE_SEGMENT|7962,7969|false|false|false|||restart
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7975,7985|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|7975,7985|false|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|7975,7985|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|SIMPLE_SEGMENT|7992,7998|false|false|false|||follow
Finding|Functional Concept|SIMPLE_SEGMENT|7992,7998|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|SIMPLE_SEGMENT|7992,7998|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|SIMPLE_SEGMENT|7992,8001|false|false|false|C0589120|Follow-up status|follow-up
Procedure|Health Care Activity|SIMPLE_SEGMENT|7992,8001|false|false|false|C1522577|follow-up|follow-up
Event|Event|SIMPLE_SEGMENT|7999,8001|false|false|false|||up
Finding|Intellectual Product|SIMPLE_SEGMENT|8012,8024|false|false|false|C1547426|Location Service Code - Primary Care|primary care
Procedure|Health Care Activity|SIMPLE_SEGMENT|8012,8024|false|false|false|C0033137|Primary Health Care|primary care
Event|Activity|SIMPLE_SEGMENT|8020,8024|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|8020,8024|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|8020,8024|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|8020,8024|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8025,8034|false|false|false|C0804815||physician
Finding|Body Substance|SIMPLE_SEGMENT|8040,8047|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|8040,8047|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|8040,8047|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|8052,8062|false|false|false|||instructed
Drug|Chemical Viewed Functionally|SIMPLE_SEGMENT|8074,8079|false|false|false|C0178499|Base|basic
Event|Event|SIMPLE_SEGMENT|8074,8079|false|false|false|||basic
Finding|Functional Concept|SIMPLE_SEGMENT|8074,8079|false|false|false|C1527178|Basis - conceptual entity|basic
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8074,8095|false|false|false|C2237045|Basic metabolic panel|basic metabolic panel
Event|Event|SIMPLE_SEGMENT|8080,8089|false|false|false|||metabolic
Finding|Cell Function|SIMPLE_SEGMENT|8080,8089|false|false|false|C0311400;C1524026|Metabolic;Metabolic Process, Cellular|metabolic
Finding|Functional Concept|SIMPLE_SEGMENT|8080,8089|false|false|false|C0311400;C1524026|Metabolic;Metabolic Process, Cellular|metabolic
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8080,8089|false|false|false|C4263342|Multisection metabolic|metabolic
Event|Event|SIMPLE_SEGMENT|8090,8095|false|false|false|||panel
Finding|Idea or Concept|SIMPLE_SEGMENT|8090,8095|false|false|false|C0441833|Groups|panel
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8114,8123|false|false|false|C0012000|Diastole|Diastolic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8114,8137|false|false|false|C1135196|Heart Failure, Diastolic|Diastolic heart failure
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8124,8129|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|8124,8129|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|8124,8129|false|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8124,8137|false|false|false|C0018801;C0018802|Congestive heart failure;Heart failure|heart failure
Event|Event|SIMPLE_SEGMENT|8130,8137|false|false|false|||failure
Finding|Functional Concept|SIMPLE_SEGMENT|8130,8137|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|SIMPLE_SEGMENT|8130,8137|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|SIMPLE_SEGMENT|8130,8137|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Event|Event|SIMPLE_SEGMENT|8139,8146|false|false|false|||Patient
Finding|Body Substance|SIMPLE_SEGMENT|8139,8146|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|8139,8146|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|8139,8146|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|8151,8160|false|false|false|||euvolemic
Event|Event|SIMPLE_SEGMENT|8174,8183|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|8174,8183|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Idea or Concept|SIMPLE_SEGMENT|8189,8193|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|8189,8193|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|8189,8193|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|8194,8199|false|false|false|C0699992|Lasix|lasix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8194,8199|false|false|false|C0699992|Lasix|lasix
Event|Event|SIMPLE_SEGMENT|8194,8199|false|false|false|||lasix
Event|Event|SIMPLE_SEGMENT|8204,8216|false|false|false|||discontinued
Event|Event|SIMPLE_SEGMENT|8229,8238|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|8229,8238|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Intellectual Product|SIMPLE_SEGMENT|8250,8255|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8250,8269|false|false|false|C0022660;C2609414|Acute kidney injury;Kidney Failure, Acute|acute kidney injury
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|8250,8269|false|false|false|C0022660;C2609414|Acute kidney injury;Kidney Failure, Acute|acute kidney injury
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8256,8262|false|false|false|C0022646;C0227665|Both kidneys;Kidney|kidney
Disorder|Neoplastic Process|SIMPLE_SEGMENT|8256,8262|false|false|false|C0496892;C0496927|Benign neoplasm of kidney;Neoplasm of uncertain or unknown behavior of kidney|kidney
Event|Event|SIMPLE_SEGMENT|8256,8262|false|false|false|||kidney
Finding|Sign or Symptom|SIMPLE_SEGMENT|8256,8262|false|false|false|C0812426|Kidney problem|kidney
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8256,8262|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8256,8262|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|8256,8269|false|false|false|C0160420|Injury of kidney|kidney injury
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|8263,8269|false|false|false|C3263722;C3263723|Traumatic AND/OR non-traumatic injury;Traumatic injury|injury
Event|Event|SIMPLE_SEGMENT|8263,8269|false|false|false|||injury
Finding|Body Substance|SIMPLE_SEGMENT|8275,8282|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|8275,8282|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|8275,8282|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|8288,8294|false|false|false|||follow
Finding|Intellectual Product|SIMPLE_SEGMENT|8308,8320|false|false|false|C1547426|Location Service Code - Primary Care|primary care
Procedure|Health Care Activity|SIMPLE_SEGMENT|8308,8320|false|false|false|C0033137|Primary Health Care|primary care
Event|Activity|SIMPLE_SEGMENT|8316,8320|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|8316,8320|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|8316,8320|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|8316,8320|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8321,8330|false|false|false|C0804815||physician
Drug|Organic Chemical|SIMPLE_SEGMENT|8348,8353|false|false|false|C0699992|Lasix|lasix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8348,8353|false|false|false|C0699992|Lasix|lasix
Event|Event|SIMPLE_SEGMENT|8348,8353|false|false|false|||lasix
Finding|Classification|SIMPLE_SEGMENT|8359,8369|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|OUTPATIENT
Finding|Idea or Concept|SIMPLE_SEGMENT|8359,8369|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|OUTPATIENT
Event|Event|SIMPLE_SEGMENT|8370,8376|false|false|false|||ISSUES
Finding|Classification|SIMPLE_SEGMENT|8378,8388|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|Outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|8378,8388|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|Outpatient
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8389,8392|false|false|false|C0053932|Bone Morphogenetic Proteins|BMP
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8389,8392|false|false|false|C0053932|Bone Morphogenetic Proteins|BMP
Event|Event|SIMPLE_SEGMENT|8389,8392|false|false|false|||BMP
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8389,8392|false|false|false|C0279266|carmustine/methotrexate/procarbazine protocol|BMP
Event|Activity|SIMPLE_SEGMENT|8397,8407|false|false|false|C1283169||monitoring
Event|Event|SIMPLE_SEGMENT|8397,8407|false|false|false|||monitoring
Procedure|Health Care Activity|SIMPLE_SEGMENT|8397,8407|false|false|false|C0150369|Preventive monitoring|monitoring
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|8411,8416|false|false|false|C5575602|Cell Culture Serum|serum
Event|Event|SIMPLE_SEGMENT|8411,8416|false|false|false|||serum
Finding|Body Substance|SIMPLE_SEGMENT|8411,8416|false|false|false|C0229671;C1546774;C1550100|Serum;Serum specimen|serum
Finding|Intellectual Product|SIMPLE_SEGMENT|8411,8416|false|false|false|C0229671;C1546774;C1550100|Serum;Serum specimen|serum
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8418,8428|false|false|false|C0010294|creatinine|creatinine
Drug|Organic Chemical|SIMPLE_SEGMENT|8418,8428|false|false|false|C0010294|creatinine|creatinine
Event|Event|SIMPLE_SEGMENT|8418,8428|false|false|false|||creatinine
Finding|Physiologic Function|SIMPLE_SEGMENT|8418,8428|false|false|false|C4551889|Creatinine metabolic function|creatinine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8418,8428|false|false|false|C0201975|Creatinine measurement|creatinine
Event|Event|SIMPLE_SEGMENT|8433,8445|false|false|false|||reinitiation
Drug|Organic Chemical|SIMPLE_SEGMENT|8449,8454|false|false|false|C0699992|Lasix|lasix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8449,8454|false|false|false|C0699992|Lasix|lasix
Event|Event|SIMPLE_SEGMENT|8449,8454|false|false|false|||lasix
Finding|Intellectual Product|SIMPLE_SEGMENT|8462,8474|false|false|false|C1547426|Location Service Code - Primary Care|primary care
Procedure|Health Care Activity|SIMPLE_SEGMENT|8462,8474|false|false|false|C0033137|Primary Health Care|primary care
Event|Activity|SIMPLE_SEGMENT|8470,8474|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|8470,8474|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|8470,8474|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|8470,8474|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8476,8485|false|false|false|C0804815||physician
Finding|Gene or Genome|SIMPLE_SEGMENT|8494,8498|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|Type
Finding|Intellectual Product|SIMPLE_SEGMENT|8494,8498|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|Type
Finding|Classification|SIMPLE_SEGMENT|8494,8500|false|false|false|C0441730|Type 2|Type 2
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8494,8509|false|false|false|C0011860|Diabetes Mellitus, Non-Insulin-Dependent|Type 2 Diabetes
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8501,8509|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|Diabetes
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8520,8527|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|SIMPLE_SEGMENT|8520,8527|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8520,8527|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|SIMPLE_SEGMENT|8520,8527|false|false|false|||insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|8520,8527|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8520,8527|false|false|false|C0202098|Insulin measurement|insulin
Event|Event|SIMPLE_SEGMENT|8528,8537|false|false|false|||dependent
Finding|Functional Concept|SIMPLE_SEGMENT|8528,8537|false|false|false|C3244310|dependent|dependent
Finding|Finding|SIMPLE_SEGMENT|8539,8549|false|false|false|C4085643;C5201148;C5962468|Moderate;Moderate Effect;Moderate Response|Moderately
Event|Event|SIMPLE_SEGMENT|8551,8561|false|false|false|||controlled
Event|Event|SIMPLE_SEGMENT|8572,8575|false|false|false|||A1c
Finding|Classification|SIMPLE_SEGMENT|8572,8575|false|false|false|C4521595|United States Military enlisted E3 (qualifier value)|A1c
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8572,8575|false|false|false|C0474680|Hemoglobin A1c measurement|A1c
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8589,8595|false|false|false|C0876064|Lantus|Lantus
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8589,8595|false|false|false|C0876064|Lantus|Lantus
Event|Event|SIMPLE_SEGMENT|8589,8595|false|false|false|||Lantus
Event|Event|SIMPLE_SEGMENT|8600,8607|false|false|false|||sliding
Finding|Functional Concept|SIMPLE_SEGMENT|8600,8607|false|false|false|C0332246|Sliding|sliding
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8609,8614|false|false|false|C0222045|Integumentary scale|scale
Event|Activity|SIMPLE_SEGMENT|8609,8614|false|false|false|C1947916|Scaling|scale
Event|Event|SIMPLE_SEGMENT|8609,8614|false|false|false|||scale
Finding|Conceptual Entity|SIMPLE_SEGMENT|8609,8614|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|scale
Finding|Intellectual Product|SIMPLE_SEGMENT|8609,8614|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|scale
Event|Event|SIMPLE_SEGMENT|8619,8628|false|false|false|||continued
Event|Event|SIMPLE_SEGMENT|8641,8656|false|false|false|||hospitalization
Procedure|Health Care Activity|SIMPLE_SEGMENT|8641,8656|false|false|false|C0019993|Hospitalization|hospitalization
Event|Event|SIMPLE_SEGMENT|8667,8677|false|false|false|||discharged
Event|Event|SIMPLE_SEGMENT|8678,8682|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|8678,8682|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|8678,8682|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|8678,8682|false|false|false|C1553498|home health encounter|home
Finding|Idea or Concept|SIMPLE_SEGMENT|8690,8694|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|8690,8694|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|8690,8694|false|false|false|C1553498|home health encounter|home
Event|Event|SIMPLE_SEGMENT|8695,8700|false|false|false|||doses
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8704,8710|false|false|false|C0876064|Lantus|lantus
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8704,8710|false|false|false|C0876064|Lantus|lantus
Event|Event|SIMPLE_SEGMENT|8704,8710|false|false|false|||lantus
Finding|Idea or Concept|SIMPLE_SEGMENT|8719,8723|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|8719,8723|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|8719,8723|false|false|false|C1553498|home health encounter|home
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8724,8731|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|SIMPLE_SEGMENT|8724,8731|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8724,8731|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|SIMPLE_SEGMENT|8724,8731|false|false|false|||insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|8724,8731|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8724,8731|false|false|false|C0202098|Insulin measurement|insulin
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8741,8746|false|false|false|C0222045|Integumentary scale|scale
Event|Activity|SIMPLE_SEGMENT|8741,8746|false|false|false|C1947916|Scaling|scale
Event|Event|SIMPLE_SEGMENT|8741,8746|false|false|false|||scale
Finding|Conceptual Entity|SIMPLE_SEGMENT|8741,8746|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|scale
Finding|Intellectual Product|SIMPLE_SEGMENT|8741,8746|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|scale
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8755,8767|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|SIMPLE_SEGMENT|8755,8767|false|false|false|||Hypertension
Finding|Body Substance|SIMPLE_SEGMENT|8789,8796|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|8789,8796|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|8789,8796|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|8799,8808|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|8799,8808|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8815,8820|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|8815,8820|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|8815,8820|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Finding|SIMPLE_SEGMENT|8815,8829|false|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|blood pressure
Finding|Organism Function|SIMPLE_SEGMENT|8815,8829|false|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|blood pressure
Procedure|Health Care Activity|SIMPLE_SEGMENT|8815,8829|false|false|false|C0005824|Blood pressure determination|blood pressure
Event|Event|SIMPLE_SEGMENT|8821,8829|false|false|false|||pressure
Finding|Finding|SIMPLE_SEGMENT|8821,8829|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|SIMPLE_SEGMENT|8821,8829|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|8821,8829|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|8821,8829|false|false|false|C0033095||pressure
Finding|Finding|SIMPLE_SEGMENT|8835,8839|false|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|8840,8850|false|false|false|||controlled
Event|Event|SIMPLE_SEGMENT|8852,8856|false|false|false|||goal
Finding|Idea or Concept|SIMPLE_SEGMENT|8852,8856|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Finding|Intellectual Product|SIMPLE_SEGMENT|8852,8856|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Event|Event|SIMPLE_SEGMENT|8876,8885|false|false|false|||continued
Finding|Idea or Concept|SIMPLE_SEGMENT|8876,8885|false|false|false|C0549178|Continuous|continued
Drug|Organic Chemical|SIMPLE_SEGMENT|8889,8899|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8889,8899|false|false|false|C0025859|metoprolol|metoprolol
Event|Event|SIMPLE_SEGMENT|8889,8899|false|false|false|||metoprolol
Drug|Organic Chemical|SIMPLE_SEGMENT|8904,8909|false|false|false|C0590690|Imdur|imdur
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8904,8909|false|false|false|C0590690|Imdur|imdur
Event|Event|SIMPLE_SEGMENT|8904,8909|false|false|false|||imdur
Drug|Organic Chemical|SIMPLE_SEGMENT|8918,8928|false|false|false|C0016860|furosemide|furosemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8918,8928|false|false|false|C0016860|furosemide|furosemide
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8934,8944|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8934,8944|false|false|false|C0065374|lisinopril|lisinopril
Event|Event|SIMPLE_SEGMENT|8934,8944|false|false|false|||lisinopril
Event|Event|SIMPLE_SEGMENT|8950,8962|false|false|false|||discontinued
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8966,8971|false|false|false|C1570446|TNFSF14 protein, human|light
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8966,8971|false|false|false|C1570446|TNFSF14 protein, human|light
Event|Event|SIMPLE_SEGMENT|8966,8971|false|false|false|||light
Finding|Finding|SIMPLE_SEGMENT|8966,8971|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Functional Concept|SIMPLE_SEGMENT|8966,8971|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Gene or Genome|SIMPLE_SEGMENT|8966,8971|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|8966,8971|false|false|false|C0023693|Light|light
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8966,8971|false|false|false|C0031765|Phototherapy|light
Finding|Body Substance|SIMPLE_SEGMENT|8979,8986|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|8979,8986|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|8979,8986|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|8999,9004|false|false|false|C5575602|Cell Culture Serum|serum
Event|Event|SIMPLE_SEGMENT|8999,9004|false|false|false|||serum
Finding|Body Substance|SIMPLE_SEGMENT|8999,9004|false|false|false|C0229671;C1546774;C1550100|Serum;Serum specimen|serum
Finding|Intellectual Product|SIMPLE_SEGMENT|8999,9004|false|false|false|C0229671;C1546774;C1550100|Serum;Serum specimen|serum
Finding|Finding|SIMPLE_SEGMENT|8999,9015|false|false|false|C0600061|Serum creatinine level|serum creatinine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8999,9015|false|false|false|C0201976|Creatinine measurement, serum (procedure)|serum creatinine
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9005,9015|false|false|false|C0010294|creatinine|creatinine
Drug|Organic Chemical|SIMPLE_SEGMENT|9005,9015|false|false|false|C0010294|creatinine|creatinine
Event|Event|SIMPLE_SEGMENT|9005,9015|false|false|false|||creatinine
Finding|Physiologic Function|SIMPLE_SEGMENT|9005,9015|false|false|false|C4551889|Creatinine metabolic function|creatinine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9005,9015|false|false|false|C0201975|Creatinine measurement|creatinine
Finding|Body Substance|SIMPLE_SEGMENT|9037,9044|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|9037,9044|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|9037,9044|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9047,9054|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|9047,9054|false|false|false|C1314974|Cardiac attachment|cardiac
Event|Event|SIMPLE_SEGMENT|9056,9071|false|false|false|||catheterization
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9056,9071|false|false|false|C0007430|Catheterization|catheterization
Event|Event|SIMPLE_SEGMENT|9081,9086|false|false|false|||noted
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|9104,9112|false|false|false|C0039155|Systole|systolic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9113,9118|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|9113,9118|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|9113,9118|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Event|Event|SIMPLE_SEGMENT|9120,9129|false|false|false|||pressures
Finding|Finding|SIMPLE_SEGMENT|9120,9129|false|false|false|C0460139|Pressure (finding)|pressures
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|9120,9129|false|false|false|C0033095||pressures
Event|Event|SIMPLE_SEGMENT|9138,9145|false|false|false|||started
Drug|Organic Chemical|SIMPLE_SEGMENT|9151,9164|false|false|false|C0017887|nitroglycerin|nitroglycerin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9151,9164|false|false|false|C0017887|nitroglycerin|nitroglycerin
Event|Event|SIMPLE_SEGMENT|9151,9164|false|false|false|||nitroglycerin
Event|Event|SIMPLE_SEGMENT|9165,9169|false|false|false|||drip
Drug|Organic Chemical|SIMPLE_SEGMENT|9174,9181|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9174,9181|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Substance|SIMPLE_SEGMENT|9174,9181|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Event|Event|SIMPLE_SEGMENT|9174,9181|false|false|false|||control
Finding|Conceptual Entity|SIMPLE_SEGMENT|9174,9181|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Functional Concept|SIMPLE_SEGMENT|9174,9181|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Idea or Concept|SIMPLE_SEGMENT|9174,9181|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9186,9191|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|9186,9191|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|9186,9191|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Finding|SIMPLE_SEGMENT|9186,9201|false|false|false|C1272641|Systemic arterial pressure|blood pressures
Event|Event|SIMPLE_SEGMENT|9192,9201|false|false|false|||pressures
Finding|Finding|SIMPLE_SEGMENT|9192,9201|false|false|false|C0460139|Pressure (finding)|pressures
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|9192,9201|false|false|false|C0033095||pressures
Finding|Body Substance|SIMPLE_SEGMENT|9207,9214|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|9207,9214|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|9207,9214|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|9219,9225|false|false|false|||weaned
Drug|Organic Chemical|SIMPLE_SEGMENT|9235,9248|false|false|false|C0017887|nitroglycerin|nitroglycerin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9235,9248|false|false|false|C0017887|nitroglycerin|nitroglycerin
Event|Event|SIMPLE_SEGMENT|9235,9248|false|false|false|||nitroglycerin
Event|Event|SIMPLE_SEGMENT|9250,9254|false|false|false|||drip
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9277,9284|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|9277,9284|false|false|false|C1314974|Cardiac attachment|cardiac
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|9277,9300|false|false|false|C0261588|Cardiac catheterisation as the cause of abnormal reaction of the patient, or of later complication, without mention of misadventure at the time of the procedure|cardiac catheterization
Finding|Intellectual Product|SIMPLE_SEGMENT|9277,9300|false|false|false|C1547981|Diagnostic Service Section ID - Cardiac Catheterization|cardiac catheterization
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|9277,9300|false|false|false|C0018795;C1548828|Cardiac Catheterization Procedures;Consent Type - Cardiac Catheterization|cardiac catheterization
Procedure|Health Care Activity|SIMPLE_SEGMENT|9277,9300|false|false|false|C0018795;C1548828|Cardiac Catheterization Procedures;Consent Type - Cardiac Catheterization|cardiac catheterization
Event|Event|SIMPLE_SEGMENT|9285,9300|false|false|false|||catheterization
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9285,9300|false|false|false|C0007430|Catheterization|catheterization
Finding|Body Substance|SIMPLE_SEGMENT|9306,9313|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|9306,9313|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|9306,9313|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|9326,9330|false|false|false|||dose
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9334,9344|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9334,9344|false|false|false|C0065374|lisinopril|lisinopril
Event|Event|SIMPLE_SEGMENT|9334,9344|false|false|false|||lisinopril
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|9368,9373|false|false|false|C5575602|Cell Culture Serum|serum
Event|Event|SIMPLE_SEGMENT|9368,9373|false|false|false|||serum
Finding|Body Substance|SIMPLE_SEGMENT|9368,9373|false|false|false|C0229671;C1546774;C1550100|Serum;Serum specimen|serum
Finding|Intellectual Product|SIMPLE_SEGMENT|9368,9373|false|false|false|C0229671;C1546774;C1550100|Serum;Serum specimen|serum
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9375,9385|false|false|false|C0010294|creatinine|creatinine
Drug|Organic Chemical|SIMPLE_SEGMENT|9375,9385|false|false|false|C0010294|creatinine|creatinine
Event|Event|SIMPLE_SEGMENT|9375,9385|false|false|false|||creatinine
Finding|Physiologic Function|SIMPLE_SEGMENT|9375,9385|false|false|false|C4551889|Creatinine metabolic function|creatinine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9375,9385|false|false|false|C0201975|Creatinine measurement|creatinine
Finding|Body Substance|SIMPLE_SEGMENT|9391,9398|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|9391,9398|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|9391,9398|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|9401,9405|false|false|false|C1552851|next - HtmlLinkType|next
Event|Event|SIMPLE_SEGMENT|9406,9410|false|false|false|||dose
Event|Event|SIMPLE_SEGMENT|9415,9419|false|false|false|||held
Finding|Classification|SIMPLE_SEGMENT|9425,9435|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|OUTPATIENT
Finding|Idea or Concept|SIMPLE_SEGMENT|9425,9435|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|OUTPATIENT
Event|Event|SIMPLE_SEGMENT|9436,9442|false|false|false|||ISSUES
Event|Event|SIMPLE_SEGMENT|9444,9450|false|false|false|||Follow
Finding|Intellectual Product|SIMPLE_SEGMENT|9459,9471|false|false|false|C1547426|Location Service Code - Primary Care|primary care
Procedure|Health Care Activity|SIMPLE_SEGMENT|9459,9471|false|false|false|C0033137|Primary Health Care|primary care
Event|Activity|SIMPLE_SEGMENT|9467,9471|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|9467,9471|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|9467,9471|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|9467,9471|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9472,9481|false|false|false|C0804815||physician
Finding|Finding|SIMPLE_SEGMENT|9493,9515|false|false|false|C0745043|History of recent hospitalization|recent hospitalization
Event|Event|SIMPLE_SEGMENT|9500,9515|false|false|false|||hospitalization
Procedure|Health Care Activity|SIMPLE_SEGMENT|9500,9515|false|false|false|C0019993|Hospitalization|hospitalization
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9520,9537|false|false|false|C0003364|Antihypertensive Agents|anti-hypertensive
Event|Event|SIMPLE_SEGMENT|9538,9545|false|false|false|||regimen
Finding|Intellectual Product|SIMPLE_SEGMENT|9538,9545|false|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9538,9545|false|false|false|C0040808|Treatment Protocols|regimen
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9550,9555|false|false|false|C1570446|TNFSF14 protein, human|light
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9550,9555|false|false|false|C1570446|TNFSF14 protein, human|light
Event|Event|SIMPLE_SEGMENT|9550,9555|false|false|false|||light
Finding|Finding|SIMPLE_SEGMENT|9550,9555|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Functional Concept|SIMPLE_SEGMENT|9550,9555|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Gene or Genome|SIMPLE_SEGMENT|9550,9555|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|9550,9555|false|false|false|C0023693|Light|light
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9550,9555|false|false|false|C0031765|Phototherapy|light
Finding|Finding|SIMPLE_SEGMENT|9559,9584|false|false|false|C0700225|Serum creatinine raised|elevated serum creatinine
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|9568,9573|false|false|false|C5575602|Cell Culture Serum|serum
Event|Event|SIMPLE_SEGMENT|9568,9573|false|false|false|||serum
Finding|Body Substance|SIMPLE_SEGMENT|9568,9573|false|false|false|C0229671;C1546774;C1550100|Serum;Serum specimen|serum
Finding|Intellectual Product|SIMPLE_SEGMENT|9568,9573|false|false|false|C0229671;C1546774;C1550100|Serum;Serum specimen|serum
Finding|Finding|SIMPLE_SEGMENT|9568,9584|false|false|false|C0600061|Serum creatinine level|serum creatinine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9568,9584|false|false|false|C0201976|Creatinine measurement, serum (procedure)|serum creatinine
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9574,9584|false|false|false|C0010294|creatinine|creatinine
Drug|Organic Chemical|SIMPLE_SEGMENT|9574,9584|false|false|false|C0010294|creatinine|creatinine
Event|Event|SIMPLE_SEGMENT|9574,9584|false|false|false|||creatinine
Finding|Physiologic Function|SIMPLE_SEGMENT|9574,9584|false|false|false|C4551889|Creatinine metabolic function|creatinine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9574,9584|false|false|false|C0201975|Creatinine measurement|creatinine
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9592,9606|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|Hyperlipidemia
Event|Event|SIMPLE_SEGMENT|9592,9606|false|false|false|||Hyperlipidemia
Finding|Finding|SIMPLE_SEGMENT|9592,9606|false|false|false|C0428465|Serum lipids high (finding)|Hyperlipidemia
Finding|Finding|SIMPLE_SEGMENT|9608,9612|false|false|false|C5575035|Well (answer to question)|Well
Event|Event|SIMPLE_SEGMENT|9613,9623|false|false|false|||controlled
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9634,9637|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Drug|Organic Chemical|SIMPLE_SEGMENT|9634,9637|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Event|Event|SIMPLE_SEGMENT|9634,9637|false|false|false|||LDL
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9634,9637|false|false|false|C0202117|Low density lipoprotein cholesterol measurement|LDL
Finding|Idea or Concept|SIMPLE_SEGMENT|9650,9654|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Finding|Intellectual Product|SIMPLE_SEGMENT|9650,9654|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9655,9658|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Drug|Organic Chemical|SIMPLE_SEGMENT|9655,9658|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Event|Event|SIMPLE_SEGMENT|9655,9658|false|false|false|||LDL
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9655,9658|false|false|false|C0202117|Low density lipoprotein cholesterol measurement|LDL
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9671,9684|false|false|false|C0041004|Triglycerides|triglycerides
Drug|Organic Chemical|SIMPLE_SEGMENT|9671,9684|false|false|false|C0041004|Triglycerides|triglycerides
Event|Event|SIMPLE_SEGMENT|9671,9684|false|false|false|||triglycerides
Finding|Physiologic Function|SIMPLE_SEGMENT|9671,9684|false|false|false|C4554056|Triglycerides metabolic function|triglycerides
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9671,9684|false|false|false|C0202236|Triglycerides measurement|triglycerides
Event|Event|SIMPLE_SEGMENT|9692,9700|false|false|false|||elevated
Drug|Organic Chemical|SIMPLE_SEGMENT|9704,9716|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9704,9716|false|false|false|C0286651|atorvastatin|Atorvastatin
Event|Event|SIMPLE_SEGMENT|9704,9716|false|false|false|||Atorvastatin
Event|Event|SIMPLE_SEGMENT|9721,9730|false|false|false|||increased
Finding|Finding|SIMPLE_SEGMENT|9755,9758|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|9755,9758|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9759,9762|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9759,9762|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|9759,9762|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|9759,9762|false|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|9759,9762|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|9759,9762|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|9759,9762|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9759,9762|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Event|Event|SIMPLE_SEGMENT|9764,9771|false|false|false|||lesions
Finding|Finding|SIMPLE_SEGMENT|9764,9771|false|false|false|C0221198|Lesion|lesions
Finding|Body Substance|SIMPLE_SEGMENT|9773,9780|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|9773,9780|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|9773,9780|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Finding|SIMPLE_SEGMENT|9792,9799|false|false|false|C0015663|Fasting|fasting
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9792,9799|false|false|false|C5203658|Fasting (regime/therapy)|fasting
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9792,9811|false|false|false|C0430044|Fasting lipid profile|fasting lipid panel
Drug|Organic Chemical|SIMPLE_SEGMENT|9800,9805|false|false|false|C0023779|Lipids|lipid
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9800,9811|false|false|false|C5671281||lipid panel
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9800,9811|false|false|false|C0200382;C5574763|Lipid panel|lipid panel
Event|Event|SIMPLE_SEGMENT|9806,9811|false|false|false|||panel
Finding|Idea or Concept|SIMPLE_SEGMENT|9806,9811|false|false|false|C0441833|Groups|panel
Event|Event|SIMPLE_SEGMENT|9839,9846|false|false|false|||pending
Finding|Idea or Concept|SIMPLE_SEGMENT|9839,9846|false|false|false|C1691786;C1704475|Pending - Allergy Clinical Status;Pending - referral status|pending
Finding|Finding|SIMPLE_SEGMENT|9850,9854|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|9850,9854|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|9850,9854|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|SIMPLE_SEGMENT|9858,9867|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|9858,9867|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|9858,9867|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|9858,9867|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|9858,9867|false|false|false|C0030685|Patient Discharge|discharge
Finding|Classification|SIMPLE_SEGMENT|9872,9882|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|OUTPATIENT
Finding|Idea or Concept|SIMPLE_SEGMENT|9872,9882|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|OUTPATIENT
Event|Event|SIMPLE_SEGMENT|9883,9889|false|false|false|||ISSUES
Event|Event|SIMPLE_SEGMENT|9891,9897|false|false|false|||Follow
Finding|Idea or Concept|SIMPLE_SEGMENT|9904,9911|false|false|false|C1691786;C1704475|Pending - Allergy Clinical Status;Pending - referral status|pending
Finding|Finding|SIMPLE_SEGMENT|9912,9919|false|false|false|C0015663|Fasting|fasting
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9912,9919|false|false|false|C5203658|Fasting (regime/therapy)|fasting
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9912,9931|false|false|false|C0430044|Fasting lipid profile|fasting lipid panel
Drug|Organic Chemical|SIMPLE_SEGMENT|9920,9925|false|false|false|C0023779|Lipids|lipid
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9920,9931|false|false|false|C5671281||lipid panel
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9920,9931|false|false|false|C0200382;C5574763|Lipid panel|lipid panel
Event|Event|SIMPLE_SEGMENT|9926,9931|false|false|false|||panel
Finding|Idea or Concept|SIMPLE_SEGMENT|9926,9931|false|false|false|C0441833|Groups|panel
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9941,9945|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9941,9945|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|SIMPLE_SEGMENT|9941,9945|false|false|false|||COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|9941,9945|false|false|false|C1412502|ARCN1 gene|COPD
Event|Event|SIMPLE_SEGMENT|9957,9969|false|false|false|||asymptomatic
Finding|Finding|SIMPLE_SEGMENT|9957,9969|false|false|false|C0231221;C0332151|Asymptomatic (finding);Asymptomatic diagnosis of|asymptomatic
Finding|Body Substance|SIMPLE_SEGMENT|9971,9978|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|9971,9978|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|9971,9978|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|9983,9991|false|false|false|||continue
Drug|Organic Chemical|SIMPLE_SEGMENT|9992,10003|false|false|false|C0082607|fluticasone|fluticasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9992,10003|false|false|false|C0082607|fluticasone|fluticasone
Event|Event|SIMPLE_SEGMENT|9992,10003|false|false|false|||fluticasone
Drug|Organic Chemical|SIMPLE_SEGMENT|10009,10018|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10009,10018|false|false|false|C0001927|albuterol|albuterol
Event|Event|SIMPLE_SEGMENT|10009,10018|false|false|false|||albuterol
Event|Event|SIMPLE_SEGMENT|10022,10028|false|false|false|||needed
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10036,10047|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10036,10047|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|10036,10047|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|10036,10047|false|false|false|C4284232|Medications|Medications
Finding|Finding|SIMPLE_SEGMENT|10036,10060|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|SIMPLE_SEGMENT|10051,10060|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|10051,10060|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Organic Chemical|SIMPLE_SEGMENT|10064,10075|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10064,10075|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Organic Chemical|SIMPLE_SEGMENT|10116,10128|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10116,10128|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10145,10155|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10145,10155|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Organic Chemical|SIMPLE_SEGMENT|10172,10182|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10172,10182|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Organic Chemical|SIMPLE_SEGMENT|10172,10192|false|false|false|C0724633|metoprolol succinate|Metoprolol succinate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10172,10192|false|false|false|C0724633|metoprolol succinate|Metoprolol succinate
Drug|Organic Chemical|SIMPLE_SEGMENT|10183,10192|false|false|false|C0038617;C0220918|Succinates;succinate|succinate
Event|Event|SIMPLE_SEGMENT|10183,10192|false|false|false|||succinate
Drug|Organic Chemical|SIMPLE_SEGMENT|10210,10220|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10210,10220|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Organic Chemical|SIMPLE_SEGMENT|10210,10232|false|false|false|C0064079|isosorbide mononitrate|Isosorbide mononitrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10210,10232|false|false|false|C0064079|isosorbide mononitrate|Isosorbide mononitrate
Event|Event|SIMPLE_SEGMENT|10221,10232|false|false|false|||mononitrate
Drug|Organic Chemical|SIMPLE_SEGMENT|10249,10259|false|false|false|C0016860|furosemide|Furosemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10249,10259|false|false|false|C0016860|furosemide|Furosemide
Drug|Organic Chemical|SIMPLE_SEGMENT|10276,10289|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10276,10289|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Finding|Gene or Genome|SIMPLE_SEGMENT|10300,10303|false|false|false|C1422467|CIAO3 gene|prn
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10308,10316|false|false|false|C0907402|insulin glargine|Glargine
Drug|Hormone|SIMPLE_SEGMENT|10308,10316|false|false|false|C0907402|insulin glargine|Glargine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10308,10316|false|false|false|C0907402|insulin glargine|Glargine
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10308,10324|false|false|false|C0907402|insulin glargine|Glargine insulin
Drug|Hormone|SIMPLE_SEGMENT|10308,10324|false|false|false|C0907402|insulin glargine|Glargine insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10308,10324|false|false|false|C0907402|insulin glargine|Glargine insulin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10317,10324|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|SIMPLE_SEGMENT|10317,10324|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10317,10324|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|SIMPLE_SEGMENT|10317,10324|false|false|false|||insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|10317,10324|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10317,10324|false|false|false|C0202098|Insulin measurement|insulin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10342,10348|false|false|false|C0293359|insulin lispro|Lispro
Drug|Hormone|SIMPLE_SEGMENT|10342,10348|false|false|false|C0293359|insulin lispro|Lispro
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10342,10348|false|false|false|C0293359|insulin lispro|Lispro
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10342,10356|false|false|false|C0293359|insulin lispro|Lispro insulin
Drug|Hormone|SIMPLE_SEGMENT|10342,10356|false|false|false|C0293359|insulin lispro|Lispro insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10342,10356|false|false|false|C0293359|insulin lispro|Lispro insulin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10349,10356|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|SIMPLE_SEGMENT|10349,10356|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10349,10356|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|SIMPLE_SEGMENT|10349,10356|false|false|false|||insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|10349,10356|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10349,10356|false|false|false|C0202098|Insulin measurement|insulin
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10365,10370|false|false|false|C0222045|Integumentary scale|scale
Event|Activity|SIMPLE_SEGMENT|10365,10370|false|false|false|C1947916|Scaling|scale
Finding|Conceptual Entity|SIMPLE_SEGMENT|10365,10370|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|scale
Finding|Intellectual Product|SIMPLE_SEGMENT|10365,10370|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|scale
Drug|Organic Chemical|SIMPLE_SEGMENT|10375,10384|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10375,10384|false|false|false|C0001927|albuterol|Albuterol
Event|Event|SIMPLE_SEGMENT|10395,10400|false|false|false|||puffs
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10406,10409|false|false|false|C0751781|Dentatorubral-Pallidoluysian Atrophy|hrs
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10406,10409|false|false|false|C1568891|HGS protein, human|hrs
Drug|Biologically Active Substance|SIMPLE_SEGMENT|10406,10409|false|false|false|C1568891|HGS protein, human|hrs
Event|Event|SIMPLE_SEGMENT|10406,10409|false|false|false|||hrs
Finding|Gene or Genome|SIMPLE_SEGMENT|10406,10409|false|false|false|C1366514;C1415473;C1419996;C1708271;C5575450;C5780798|ATN1 wt Allele;HARS1 gene;HARS1 wt Allele;HGS gene;HGS wt Allele;SRSF5 gene|hrs
Finding|Gene or Genome|SIMPLE_SEGMENT|10410,10413|false|false|false|C1422467|CIAO3 gene|prn
Drug|Organic Chemical|SIMPLE_SEGMENT|10418,10429|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10418,10429|false|false|false|C0082607|fluticasone|Fluticasone
Event|Event|SIMPLE_SEGMENT|10418,10429|false|false|false|||Fluticasone
Event|Event|SIMPLE_SEGMENT|10434,10437|false|false|false|||mcg
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|10447,10450|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10447,10450|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|10447,10450|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|10447,10450|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|10447,10450|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|10455,10467|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10455,10467|false|false|false|C0081876|pantoprazole|Pantoprazole
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|10474,10477|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10474,10477|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|10474,10477|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|10474,10477|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|10474,10477|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|10490,10503|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10490,10503|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|SIMPLE_SEGMENT|10490,10503|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10490,10503|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|SIMPLE_SEGMENT|10520,10523|false|false|false|C1422467|CIAO3 gene|prn
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10524,10528|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|10524,10528|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|10524,10528|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|10524,10528|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Biologically Active Substance|SIMPLE_SEGMENT|10533,10542|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|10533,10542|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Food|SIMPLE_SEGMENT|10533,10542|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|10533,10542|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10533,10542|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Event|Event|SIMPLE_SEGMENT|10533,10542|false|false|false|||Potassium
Finding|Physiologic Function|SIMPLE_SEGMENT|10533,10542|false|false|false|C4553027|Potassium metabolic function|Potassium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10533,10542|false|false|false|C0202194|Potassium measurement|Potassium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|10533,10551|false|false|false|C0032825|potassium chloride|Potassium chloride
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10533,10551|false|false|false|C0032825|potassium chloride|Potassium chloride
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|10543,10551|false|false|false|C0008203;C0596019|Chlorides;chloride ion|chloride
Event|Event|SIMPLE_SEGMENT|10543,10551|false|false|false|||chloride
Finding|Physiologic Function|SIMPLE_SEGMENT|10543,10551|false|false|false|C4553021|Chloride metabolic function|chloride
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10543,10551|false|false|false|C0201952|Chloride measurement|chloride
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|10559,10562|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10559,10562|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|10559,10562|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|10559,10562|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|10559,10562|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|10567,10582|false|false|false|C0008318|cholecalciferol|Cholecalciferol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10567,10582|false|false|false|C0008318|cholecalciferol|Cholecalciferol
Drug|Vitamin|SIMPLE_SEGMENT|10567,10582|false|false|false|C0008318|cholecalciferol|Cholecalciferol
Drug|Organic Chemical|SIMPLE_SEGMENT|10604,10617|false|false|false|C0025872|metronidazole|Metronidazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10604,10617|false|false|false|C0025872|metronidazole|Metronidazole
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10624,10630|false|false|false|C0544341|Lotion|lotion
Event|Event|SIMPLE_SEGMENT|10624,10630|false|false|false|||lotion
Event|Event|SIMPLE_SEGMENT|10644,10653|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|10644,10653|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|10644,10653|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|10644,10653|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|10644,10653|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|10644,10665|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10654,10665|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10654,10665|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|10654,10665|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|10654,10665|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|SIMPLE_SEGMENT|10670,10681|false|false|false|C0070166|clopidogrel|clopidogrel
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10670,10681|false|false|false|C0070166|clopidogrel|clopidogrel
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10688,10694|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10708,10714|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|10708,10714|false|false|false|||Tablet
Drug|Organic Chemical|SIMPLE_SEGMENT|10739,10746|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10739,10746|false|false|false|C0004057|aspirin|aspirin
Event|Event|SIMPLE_SEGMENT|10739,10746|false|false|false|||aspirin
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10754,10760|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10774,10780|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|10774,10780|false|false|false|||Tablet
Drug|Organic Chemical|SIMPLE_SEGMENT|10804,10816|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10804,10816|false|false|false|C0286651|atorvastatin|atorvastatin
Event|Event|SIMPLE_SEGMENT|10804,10816|false|false|false|||atorvastatin
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10823,10829|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10843,10849|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|10843,10849|false|false|false|||Tablet
Drug|Organic Chemical|SIMPLE_SEGMENT|10874,10884|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10874,10884|false|false|false|C0025859|metoprolol|metoprolol
Event|Event|SIMPLE_SEGMENT|10874,10884|false|false|false|||metoprolol
Drug|Organic Chemical|SIMPLE_SEGMENT|10874,10894|false|false|false|C0724633|metoprolol succinate|metoprolol succinate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10874,10894|false|false|false|C0724633|metoprolol succinate|metoprolol succinate
Drug|Organic Chemical|SIMPLE_SEGMENT|10885,10894|false|false|false|C0038617;C0220918|Succinates;succinate|succinate
Event|Event|SIMPLE_SEGMENT|10885,10894|false|false|false|||succinate
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10902,10908|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Finding|SIMPLE_SEGMENT|10909,10917|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|SIMPLE_SEGMENT|10909,10917|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|SIMPLE_SEGMENT|10918,10925|false|false|false|||Release
Finding|Functional Concept|SIMPLE_SEGMENT|10918,10925|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|10918,10925|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10918,10925|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Event|Event|SIMPLE_SEGMENT|10933,10936|false|false|false|||Sig
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10946,10952|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Finding|SIMPLE_SEGMENT|10953,10961|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|SIMPLE_SEGMENT|10953,10961|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|SIMPLE_SEGMENT|10962,10969|false|false|false|||Release
Finding|Functional Concept|SIMPLE_SEGMENT|10962,10969|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|10962,10969|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10962,10969|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Finding|Intellectual Product|SIMPLE_SEGMENT|10979,10983|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10979,10989|false|false|false|C3537736|Once A Day|once a day
Finding|Idea or Concept|SIMPLE_SEGMENT|10986,10989|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|10986,10989|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|SIMPLE_SEGMENT|10996,11006|false|false|false|C0022251|isosorbide|isosorbide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10996,11006|false|false|false|C0022251|isosorbide|isosorbide
Event|Event|SIMPLE_SEGMENT|10996,11006|false|false|false|||isosorbide
Drug|Organic Chemical|SIMPLE_SEGMENT|10996,11018|false|false|false|C0064079|isosorbide mononitrate|isosorbide mononitrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10996,11018|false|false|false|C0064079|isosorbide mononitrate|isosorbide mononitrate
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|11025,11031|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Finding|SIMPLE_SEGMENT|11032,11040|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|SIMPLE_SEGMENT|11032,11040|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|SIMPLE_SEGMENT|11041,11048|false|false|false|||Release
Finding|Functional Concept|SIMPLE_SEGMENT|11041,11048|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|11041,11048|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11041,11048|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Event|Event|SIMPLE_SEGMENT|11056,11059|false|false|false|||Sig
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|11069,11075|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Finding|SIMPLE_SEGMENT|11076,11084|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|SIMPLE_SEGMENT|11076,11084|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|SIMPLE_SEGMENT|11085,11092|false|false|false|||Release
Finding|Functional Concept|SIMPLE_SEGMENT|11085,11092|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|11085,11092|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11085,11092|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|SIMPLE_SEGMENT|11122,11135|false|false|false|C0017887|nitroglycerin|nitroglycerin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11122,11135|false|false|false|C0017887|nitroglycerin|nitroglycerin
Event|Event|SIMPLE_SEGMENT|11122,11135|false|false|false|||nitroglycerin
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|11143,11149|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|11143,11161|false|false|false|C0991582|Sublingual Tablet|Tablet, Sublingual
Finding|Finding|SIMPLE_SEGMENT|11151,11161|false|false|false|C0001565;C4521982|Sublingual (intended site);Sublingual Route of Administration|Sublingual
Finding|Functional Concept|SIMPLE_SEGMENT|11151,11161|false|false|false|C0001565;C4521982|Sublingual (intended site);Sublingual Route of Administration|Sublingual
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11162,11165|false|false|false|C0262329|Short insular gyrus|Sig
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|11162,11165|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Drug|Immunologic Factor|SIMPLE_SEGMENT|11162,11165|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Finding|Receptor|SIMPLE_SEGMENT|11162,11165|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|11175,11181|false|false|false|C0039225|Tablet Dosage Form|tablet
Event|Event|SIMPLE_SEGMENT|11175,11181|false|false|false|||tablet
Finding|Finding|SIMPLE_SEGMENT|11184,11194|false|false|false|C0001565;C4521982|Sublingual (intended site);Sublingual Route of Administration|Sublingual
Finding|Functional Concept|SIMPLE_SEGMENT|11184,11194|false|false|false|C0001565;C4521982|Sublingual (intended site);Sublingual Route of Administration|Sublingual
Finding|Gene or Genome|SIMPLE_SEGMENT|11195,11198|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|SIMPLE_SEGMENT|11203,11209|false|false|false|||needed
Anatomy|Body Location or Region|SIMPLE_SEGMENT|11214,11219|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|11214,11219|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11214,11224|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|11214,11224|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11220,11224|false|true|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|11220,11224|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|11220,11224|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|11220,11224|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|11231,11238|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|SIMPLE_SEGMENT|11231,11238|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11231,11238|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|SIMPLE_SEGMENT|11231,11238|false|false|false|||insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|11231,11238|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|11231,11238|false|false|false|C0202098|Insulin measurement|insulin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|11231,11247|false|false|false|C0907402|insulin glargine|insulin glargine
Drug|Hormone|SIMPLE_SEGMENT|11231,11247|false|false|false|C0907402|insulin glargine|insulin glargine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11231,11247|false|false|false|C0907402|insulin glargine|insulin glargine
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|11239,11247|false|false|false|C0907402|insulin glargine|glargine
Drug|Hormone|SIMPLE_SEGMENT|11239,11247|false|false|false|C0907402|insulin glargine|glargine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11239,11247|false|false|false|C0907402|insulin glargine|glargine
Event|Event|SIMPLE_SEGMENT|11239,11247|false|false|false|||glargine
Event|Event|SIMPLE_SEGMENT|11252,11256|false|false|false|||unit
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|11260,11268|false|false|false|C0037633;C0525069;C1382100|Pharmaceutical Solutions;Solution Dosage Form;Solutions|Solution
Drug|Substance|SIMPLE_SEGMENT|11260,11268|false|false|false|C0037633;C0525069;C1382100|Pharmaceutical Solutions;Solution Dosage Form;Solutions|Solution
Event|Event|SIMPLE_SEGMENT|11260,11268|false|false|false|||Solution
Finding|Conceptual Entity|SIMPLE_SEGMENT|11260,11268|false|false|false|C2699488|Resolution|Solution
Event|Event|SIMPLE_SEGMENT|11269,11272|false|false|false|||Sig
Event|Event|SIMPLE_SEGMENT|11293,11305|false|false|false|||Subcutaneous
Finding|Functional Concept|SIMPLE_SEGMENT|11293,11305|false|false|false|C1522438|Subcutaneous Route of Administration|Subcutaneous
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|11323,11330|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|SIMPLE_SEGMENT|11323,11330|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11323,11330|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|SIMPLE_SEGMENT|11323,11330|false|false|false|||insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|11323,11330|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|11323,11330|false|false|false|C0202098|Insulin measurement|insulin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|11323,11337|false|false|false|C0293359|insulin lispro|insulin lispro
Drug|Hormone|SIMPLE_SEGMENT|11323,11337|false|false|false|C0293359|insulin lispro|insulin lispro
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11323,11337|false|false|false|C0293359|insulin lispro|insulin lispro
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|11331,11337|false|false|false|C0293359|insulin lispro|lispro
Drug|Hormone|SIMPLE_SEGMENT|11331,11337|false|false|false|C0293359|insulin lispro|lispro
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11331,11337|false|false|false|C0293359|insulin lispro|lispro
Event|Event|SIMPLE_SEGMENT|11331,11337|false|false|false|||lispro
Event|Event|SIMPLE_SEGMENT|11342,11346|false|false|false|||unit
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|11350,11358|false|false|false|C0037633;C0525069;C1382100|Pharmaceutical Solutions;Solution Dosage Form;Solutions|Solution
Drug|Substance|SIMPLE_SEGMENT|11350,11358|false|false|false|C0037633;C0525069;C1382100|Pharmaceutical Solutions;Solution Dosage Form;Solutions|Solution
Event|Event|SIMPLE_SEGMENT|11350,11358|false|false|false|||Solution
Finding|Conceptual Entity|SIMPLE_SEGMENT|11350,11358|false|false|false|C2699488|Resolution|Solution
Finding|Functional Concept|SIMPLE_SEGMENT|11364,11371|false|false|false|C0332246|Sliding|Sliding
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11364,11377|false|false|false|C2937251|sliding scale|Sliding scale
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11372,11377|false|false|false|C0222045|Integumentary scale|scale
Event|Activity|SIMPLE_SEGMENT|11372,11377|false|false|false|C1947916|Scaling|scale
Finding|Conceptual Entity|SIMPLE_SEGMENT|11372,11377|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|scale
Finding|Intellectual Product|SIMPLE_SEGMENT|11372,11377|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|scale
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|11388,11395|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|SIMPLE_SEGMENT|11388,11395|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11388,11395|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|SIMPLE_SEGMENT|11388,11395|false|false|false|||insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|11388,11395|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|11388,11395|false|false|false|C0202098|Insulin measurement|insulin
Finding|Functional Concept|SIMPLE_SEGMENT|11396,11408|false|false|false|C1522438|Subcutaneous Route of Administration|Subcutaneous
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11415,11420|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|SIMPLE_SEGMENT|11423,11426|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|11423,11426|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|11431,11439|false|false|false|||directed
Finding|Classification|SIMPLE_SEGMENT|11444,11454|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|11444,11454|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|SIMPLE_SEGMENT|11455,11463|false|false|false|||provider
Finding|Functional Concept|SIMPLE_SEGMENT|11455,11463|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|provider
Finding|Intellectual Product|SIMPLE_SEGMENT|11455,11463|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|provider
Drug|Organic Chemical|SIMPLE_SEGMENT|11471,11480|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11471,11480|false|false|false|C0001927|albuterol|albuterol
Event|Event|SIMPLE_SEGMENT|11471,11480|false|false|false|||albuterol
Drug|Organic Chemical|SIMPLE_SEGMENT|11471,11488|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11471,11488|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|11481,11488|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Inorganic Chemical|SIMPLE_SEGMENT|11481,11488|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11481,11488|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Event|Event|SIMPLE_SEGMENT|11481,11488|false|false|false|||sulfate
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11506,11509|false|false|false|C0015458|Facial Hemiatrophy|HFA
Event|Event|SIMPLE_SEGMENT|11506,11509|false|false|false|||HFA
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|11506,11509|false|false|false|C0430649|High frequency audiometry|HFA
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|11510,11517|false|false|false|C1112870|Aerosol Dose Form|Aerosol
Event|Event|SIMPLE_SEGMENT|11518,11525|false|false|false|||Inhaler
Finding|Functional Concept|SIMPLE_SEGMENT|11518,11525|false|false|false|C4319647|Inhaler (unit of presentation)|Inhaler
Event|Event|SIMPLE_SEGMENT|11545,11555|false|false|false|||Inhalation
Finding|Functional Concept|SIMPLE_SEGMENT|11545,11555|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Finding|Organism Function|SIMPLE_SEGMENT|11545,11555|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Event|Event|SIMPLE_SEGMENT|11575,11581|false|false|false|||needed
Event|Event|SIMPLE_SEGMENT|11586,11589|false|false|false|||SOB
Finding|Sign or Symptom|SIMPLE_SEGMENT|11586,11589|false|false|false|C0013404|Dyspnea|SOB
Event|Event|SIMPLE_SEGMENT|11592,11600|false|false|false|||wheezing
Finding|Sign or Symptom|SIMPLE_SEGMENT|11592,11600|false|false|false|C0043144|Wheezing|wheezing
Drug|Organic Chemical|SIMPLE_SEGMENT|11608,11619|false|false|false|C0082607|fluticasone|fluticasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11608,11619|false|false|false|C0082607|fluticasone|fluticasone
Event|Event|SIMPLE_SEGMENT|11608,11619|false|false|false|||fluticasone
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|11638,11645|false|false|false|C1112870|Aerosol Dose Form|Aerosol
Event|Event|SIMPLE_SEGMENT|11646,11649|false|false|false|||Sig
Event|Event|SIMPLE_SEGMENT|11665,11675|false|false|false|||Inhalation
Finding|Functional Concept|SIMPLE_SEGMENT|11665,11675|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Finding|Organism Function|SIMPLE_SEGMENT|11665,11675|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|11676,11679|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|11676,11679|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|11676,11679|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|11676,11679|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|11676,11679|false|false|false|C1332410|BID gene|BID
Finding|Finding|SIMPLE_SEGMENT|11681,11688|false|false|false|C4035627|2 times|2 times
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11683,11688|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|SIMPLE_SEGMENT|11691,11694|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|11691,11694|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|SIMPLE_SEGMENT|11703,11715|false|false|false|C0081876|pantoprazole|pantoprazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11703,11715|false|false|false|C0081876|pantoprazole|pantoprazole
Event|Event|SIMPLE_SEGMENT|11703,11715|false|false|false|||pantoprazole
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|11722,11728|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|11722,11728|false|false|false|||Tablet
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11730,11737|false|false|false|C1545665|Views delayed|Delayed
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|11730,11745|false|false|false|C1707664|Delayed Release Dosage Form|Delayed Release
Event|Event|SIMPLE_SEGMENT|11738,11745|false|false|false|||Release
Finding|Functional Concept|SIMPLE_SEGMENT|11738,11745|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|11738,11745|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11738,11745|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Event|Event|SIMPLE_SEGMENT|11753,11756|false|false|false|||Sig
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|11767,11773|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|11767,11773|false|false|false|||Tablet
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11775,11782|false|false|false|C1545665|Views delayed|Delayed
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|11775,11790|false|false|false|C1707664|Delayed Release Dosage Form|Delayed Release
Event|Event|SIMPLE_SEGMENT|11783,11790|false|false|false|||Release
Finding|Functional Concept|SIMPLE_SEGMENT|11783,11790|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|11783,11790|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11783,11790|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|SIMPLE_SEGMENT|11830,11839|false|false|false|C0030049|oxycodone|oxycodone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11830,11839|false|false|false|C0030049|oxycodone|oxycodone
Event|Event|SIMPLE_SEGMENT|11830,11839|false|false|false|||oxycodone
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|11830,11839|false|false|false|C0524222|Oxycodone measurement|oxycodone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11830,11853|false|false|false|C0717368|acetaminophen / oxycodone|oxycodone-acetaminophen
Drug|Organic Chemical|SIMPLE_SEGMENT|11840,11853|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11840,11853|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Event|Event|SIMPLE_SEGMENT|11840,11853|false|false|false|||acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|11840,11853|false|false|false|C0373527|Acetaminophen measurement|acetaminophen
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|11861,11867|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|11881,11887|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|11915,11921|false|false|false|||needed
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11926,11930|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|11926,11930|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|11926,11930|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|11926,11930|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|SIMPLE_SEGMENT|11938,11953|false|false|false|C0008318|cholecalciferol|cholecalciferol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11938,11953|false|false|false|C0008318|cholecalciferol|cholecalciferol
Drug|Vitamin|SIMPLE_SEGMENT|11938,11953|false|false|false|C0008318|cholecalciferol|cholecalciferol
Event|Event|SIMPLE_SEGMENT|11938,11953|false|false|false|||cholecalciferol
Drug|Organic Chemical|SIMPLE_SEGMENT|11938,11966|false|false|false|C0008318|cholecalciferol|cholecalciferol (vitamin D3)
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11938,11966|false|false|false|C0008318|cholecalciferol|cholecalciferol (vitamin D3)
Drug|Vitamin|SIMPLE_SEGMENT|11938,11966|false|false|false|C0008318|cholecalciferol|cholecalciferol (vitamin D3)
Drug|Organic Chemical|SIMPLE_SEGMENT|11955,11962|false|false|false|C0042890|Vitamins|vitamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11955,11962|false|false|false|C0042890|Vitamins|vitamin
Drug|Vitamin|SIMPLE_SEGMENT|11955,11962|false|false|false|C0042890|Vitamins|vitamin
Event|Event|SIMPLE_SEGMENT|11955,11962|false|false|false|||vitamin
Drug|Organic Chemical|SIMPLE_SEGMENT|11955,11965|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11955,11965|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Drug|Vitamin|SIMPLE_SEGMENT|11955,11965|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11978,11985|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|SIMPLE_SEGMENT|11978,11985|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|11978,11985|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|12000,12007|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|SIMPLE_SEGMENT|12000,12007|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|12000,12007|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Event|Event|SIMPLE_SEGMENT|12008,12010|false|false|false|||PO
Finding|Intellectual Product|SIMPLE_SEGMENT|12011,12015|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12011,12021|false|false|false|C3537736|Once A Day|once a day
Finding|Idea or Concept|SIMPLE_SEGMENT|12018,12021|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|12018,12021|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|SIMPLE_SEGMENT|12029,12042|false|false|false|C0025872|metronidazole|metronidazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12029,12042|false|false|false|C0025872|metronidazole|metronidazole
Event|Event|SIMPLE_SEGMENT|12029,12042|false|false|false|||metronidazole
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|12050,12056|false|false|false|C0544341|Lotion|Lotion
Event|Event|SIMPLE_SEGMENT|12070,12081|false|false|false|||application
Finding|Functional Concept|SIMPLE_SEGMENT|12070,12081|false|false|false|C0870325;C1547755;C1947919;C2347934;C4048755|Application Document;Apply;Computer Application;HL7 Version 2.5 - Application;Regulatory Application|application
Finding|Idea or Concept|SIMPLE_SEGMENT|12070,12081|false|false|false|C0870325;C1547755;C1947919;C2347934;C4048755|Application Document;Apply;Computer Application;HL7 Version 2.5 - Application;Regulatory Application|application
Finding|Intellectual Product|SIMPLE_SEGMENT|12070,12081|false|false|false|C0870325;C1547755;C1947919;C2347934;C4048755|Application Document;Apply;Computer Application;HL7 Version 2.5 - Application;Regulatory Application|application
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|12070,12081|false|false|false|C0185125|Application procedure|application
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|12084,12091|false|false|false|C1710439|Topical Dosage Form|Topical
Event|Event|SIMPLE_SEGMENT|12084,12091|false|false|false|||Topical
Finding|Functional Concept|SIMPLE_SEGMENT|12084,12091|false|false|false|C1522168|Topical Route of Administration|Topical
Event|Event|SIMPLE_SEGMENT|12095,12103|false|false|false|||directed
Event|Event|SIMPLE_SEGMENT|12111,12120|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|12111,12120|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|12111,12120|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|12111,12120|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|12111,12120|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12111,12132|false|false|false|C4019243||Discharge Disposition
Finding|Finding|SIMPLE_SEGMENT|12111,12132|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12121,12132|false|false|false|C2926604||Disposition
Event|Event|SIMPLE_SEGMENT|12121,12132|false|false|false|||Disposition
Procedure|Health Care Activity|SIMPLE_SEGMENT|12121,12132|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|SIMPLE_SEGMENT|12134,12138|false|false|false|||Home
Finding|Idea or Concept|SIMPLE_SEGMENT|12134,12138|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|SIMPLE_SEGMENT|12134,12138|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|SIMPLE_SEGMENT|12134,12138|false|false|false|C1553498|home health encounter|Home
Event|Event|SIMPLE_SEGMENT|12141,12150|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|12141,12150|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|12141,12150|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|12141,12150|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|12141,12150|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|12141,12160|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12151,12160|false|false|false|C0945731||Diagnosis
Event|Event|SIMPLE_SEGMENT|12151,12160|false|false|false|||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|12151,12160|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|12151,12160|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|12151,12160|false|false|false|C0011900|Diagnosis|Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12162,12179|false|false|false|C0801658||Primary diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12170,12179|false|false|false|C0945731||diagnosis
Event|Event|SIMPLE_SEGMENT|12170,12179|false|false|false|||diagnosis
Finding|Classification|SIMPLE_SEGMENT|12170,12179|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|12170,12179|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|12170,12179|false|false|false|C0011900|Diagnosis|diagnosis
Finding|Finding|SIMPLE_SEGMENT|12181,12189|false|false|false|C0741302|atypia morphology|Atypical
Finding|Sign or Symptom|SIMPLE_SEGMENT|12181,12200|false|false|false|C0262384|Atypical chest pain|Atypical chest pain
Anatomy|Body Location or Region|SIMPLE_SEGMENT|12190,12195|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|12190,12195|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12190,12200|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|12190,12200|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12196,12200|false|true|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|12196,12200|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|12196,12200|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|12196,12200|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Disorder|Neoplastic Process|SIMPLE_SEGMENT|12202,12211|false|false|false|C0027627|Neoplasm Metastasis|Secondary
Event|Event|SIMPLE_SEGMENT|12202,12211|false|false|false|||Secondary
Finding|Functional Concept|SIMPLE_SEGMENT|12202,12211|false|false|false|C1522484|metastatic qualifier|Secondary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12202,12221|false|false|false|C4255018||Secondary diagnosis
Finding|Finding|SIMPLE_SEGMENT|12202,12221|false|false|false|C0332138|Secondary diagnosis|Secondary diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12212,12221|false|false|false|C0945731||diagnosis
Event|Event|SIMPLE_SEGMENT|12212,12221|false|false|false|||diagnosis
Finding|Classification|SIMPLE_SEGMENT|12212,12221|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|12212,12221|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|12212,12221|false|false|false|C0011900|Diagnosis|diagnosis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|12223,12231|false|false|false|C0018787|Heart|Coronary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|12223,12238|false|false|false|C0205042|Coronary artery|Coronary artery
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12223,12246|false|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|Coronary artery disease
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|12232,12238|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|SIMPLE_SEGMENT|12232,12238|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12232,12246|false|false|false|C0852949|Arteriopathic disease|artery disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12239,12246|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|12239,12246|false|false|false|||disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12248,12260|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|SIMPLE_SEGMENT|12248,12260|false|false|false|||Hypertension
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12261,12275|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|Hyperlipidemia
Event|Event|SIMPLE_SEGMENT|12261,12275|false|false|false|||Hyperlipidemia
Finding|Finding|SIMPLE_SEGMENT|12261,12275|false|false|false|C0428465|Serum lipids high (finding)|Hyperlipidemia
Finding|Gene or Genome|SIMPLE_SEGMENT|12276,12280|false|true|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|Type
Finding|Intellectual Product|SIMPLE_SEGMENT|12276,12280|false|true|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|Type
Finding|Classification|SIMPLE_SEGMENT|12276,12282|false|false|false|C0441730|Type 2|Type 2
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12276,12291|false|false|false|C0011860|Diabetes Mellitus, Non-Insulin-Dependent|Type 2 Diabetes
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12276,12300|false|false|false|C0011860|Diabetes Mellitus, Non-Insulin-Dependent|Type 2 Diabetes Mellitus
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12283,12291|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|Diabetes
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12283,12300|false|false|false|C0011849|Diabetes Mellitus|Diabetes Mellitus
Event|Event|SIMPLE_SEGMENT|12292,12300|false|false|false|||Mellitus
Event|Event|SIMPLE_SEGMENT|12304,12313|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|12304,12313|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|12304,12313|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|12304,12313|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|12304,12313|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12314,12323|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12314,12323|false|false|false|C0012634|Disease|Condition
Event|Event|SIMPLE_SEGMENT|12314,12323|false|false|false|||Condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|12314,12323|false|false|false|C1705253|Logical Condition|Condition
Finding|Mental Process|SIMPLE_SEGMENT|12325,12331|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12325,12338|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|SIMPLE_SEGMENT|12325,12338|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12332,12338|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|12332,12338|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|12340,12345|false|false|false|||Clear
Finding|Idea or Concept|SIMPLE_SEGMENT|12340,12345|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|SIMPLE_SEGMENT|12350,12358|false|false|false|||coherent
Finding|Finding|SIMPLE_SEGMENT|12350,12358|false|false|false|C4068804|Coherent|coherent
Event|Event|SIMPLE_SEGMENT|12360,12365|false|false|false|||Level
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12360,12382|false|false|false|C4050479||Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|12360,12382|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|SIMPLE_SEGMENT|12369,12382|false|false|false|||Consciousness
Finding|Finding|SIMPLE_SEGMENT|12369,12382|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|SIMPLE_SEGMENT|12369,12382|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12384,12389|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|12384,12389|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12384,12389|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|SIMPLE_SEGMENT|12384,12389|false|false|false|||Alert
Finding|Finding|SIMPLE_SEGMENT|12384,12389|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|12384,12389|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|12384,12389|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|SIMPLE_SEGMENT|12394,12405|false|false|false|||interactive
Finding|Functional Concept|SIMPLE_SEGMENT|12394,12405|false|false|false|C1704675|Interaction|interactive
Event|Activity|SIMPLE_SEGMENT|12407,12415|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|12407,12415|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|SIMPLE_SEGMENT|12407,12415|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12416,12422|false|false|false|C5889824||Status
Event|Event|SIMPLE_SEGMENT|12416,12422|false|false|false|||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|12416,12422|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|12424,12434|false|false|false|||Ambulatory
Finding|Functional Concept|SIMPLE_SEGMENT|12424,12434|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|SIMPLE_SEGMENT|12424,12434|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|SIMPLE_SEGMENT|12424,12434|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|SIMPLE_SEGMENT|12424,12434|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|SIMPLE_SEGMENT|12437,12448|false|false|false|||Independent
Finding|Finding|SIMPLE_SEGMENT|12437,12448|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|SIMPLE_SEGMENT|12437,12448|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Event|Event|SIMPLE_SEGMENT|12453,12462|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|12453,12462|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|12453,12462|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|12453,12462|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|12453,12462|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12453,12475|false|false|false|C3669312||Discharge Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|12453,12475|false|false|false|C4282220|Discharge instructions|Discharge Instructions
Procedure|Health Care Activity|SIMPLE_SEGMENT|12453,12475|false|false|false|C2266673|hospital discharge instructions (treatment)|Discharge Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12463,12475|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|12463,12475|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|12463,12475|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Event|Event|SIMPLE_SEGMENT|12486,12494|false|false|false|||pleasure
Finding|Intellectual Product|SIMPLE_SEGMENT|12486,12494|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|SIMPLE_SEGMENT|12486,12494|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|SIMPLE_SEGMENT|12502,12506|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|12502,12506|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|12502,12506|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|12502,12506|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|12502,12509|false|false|false|C1555558|care of - AddressPartType|care of
Event|Event|SIMPLE_SEGMENT|12526,12541|false|false|false|||hospitalization
Procedure|Health Care Activity|SIMPLE_SEGMENT|12526,12541|false|false|false|C0019993|Hospitalization|hospitalization
Event|Event|SIMPLE_SEGMENT|12562,12574|false|false|false|||hospitalized
Anatomy|Body Location or Region|SIMPLE_SEGMENT|12580,12585|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|12580,12585|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12580,12590|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|12580,12590|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12586,12590|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|12586,12590|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|12586,12590|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|12586,12590|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12609,12615|false|false|false|C1718621|W stress|stress
Drug|Organic Chemical|SIMPLE_SEGMENT|12609,12615|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12609,12615|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Event|Event|SIMPLE_SEGMENT|12609,12615|false|false|false|||stress
Finding|Finding|SIMPLE_SEGMENT|12609,12615|false|false|false|C0038435|Stress|stress
Anatomy|Body Location or Region|SIMPLE_SEGMENT|12617,12621|false|false|false|C4318744|Test - temporal region|test
Event|Event|SIMPLE_SEGMENT|12617,12621|false|false|false|||test
Finding|Functional Concept|SIMPLE_SEGMENT|12617,12621|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Finding|Intellectual Product|SIMPLE_SEGMENT|12617,12621|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|12617,12621|false|false|false|C0456984|Test Result|test
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|12617,12621|false|false|false|C0022885|Laboratory Procedures|test
Event|Event|SIMPLE_SEGMENT|12631,12639|false|false|false|||abnormal
Finding|Finding|SIMPLE_SEGMENT|12631,12639|false|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Finding|Idea or Concept|SIMPLE_SEGMENT|12631,12639|false|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|12664,12671|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|12664,12671|false|false|false|C1314974|Cardiac attachment|cardiac
Event|Event|SIMPLE_SEGMENT|12673,12688|false|false|false|||catheterization
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|12673,12688|false|false|false|C0007430|Catheterization|catheterization
Event|Event|SIMPLE_SEGMENT|12702,12707|false|false|false|||found
Event|Event|SIMPLE_SEGMENT|12718,12726|false|false|false|||blockage
Finding|Finding|SIMPLE_SEGMENT|12718,12726|false|false|false|C1706968;C1879887;C2237319|Blockage (obstruction - finding);Partial Blockage within Medical Device|blockage
Finding|Functional Concept|SIMPLE_SEGMENT|12735,12739|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|12735,12766|false|false|false|C0226037|Structure of circumflex branch of left coronary artery|left circumflex coronary artery
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|12740,12766|false|false|false|C0226037|Structure of circumflex branch of left coronary artery|circumflex coronary artery
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|12751,12759|false|false|false|C0018787|Heart|coronary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|12751,12766|false|false|false|C0205042|Coronary artery|coronary artery
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|12760,12766|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|SIMPLE_SEGMENT|12760,12766|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|12779,12784|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|12779,12784|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|12779,12784|false|false|false|C0795691|HEART PROBLEM|heart
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|12785,12792|false|false|false|C0005847|Blood Vessel|vessels
Event|Event|SIMPLE_SEGMENT|12797,12801|false|false|false|||Take
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12806,12816|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|12806,12816|false|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|12806,12816|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|SIMPLE_SEGMENT|12820,12830|false|false|false|||instructed
Event|Event|SIMPLE_SEGMENT|12839,12843|false|false|false|||note
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12859,12869|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|12859,12869|false|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|12859,12869|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|SIMPLE_SEGMENT|12870,12877|false|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|12870,12877|false|false|false|C0392747|Changing|changes
Event|Event|SIMPLE_SEGMENT|12882,12886|false|false|false|||Stop
Drug|Biologically Active Substance|SIMPLE_SEGMENT|12899,12908|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|12899,12908|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Food|SIMPLE_SEGMENT|12899,12908|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|12899,12908|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12899,12908|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Event|Event|SIMPLE_SEGMENT|12899,12908|false|false|false|||potassium
Finding|Physiologic Function|SIMPLE_SEGMENT|12899,12908|false|false|false|C4553027|Potassium metabolic function|potassium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|12899,12908|false|false|false|C0202194|Potassium measurement|potassium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|12899,12919|false|false|false|C0304475|Potassium supplement|potassium supplement
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12899,12919|false|false|false|C0304475|Potassium supplement|potassium supplement
Drug|Food|SIMPLE_SEGMENT|12909,12919|false|false|false|C0242295|Dietary Supplements|supplement
Event|Event|SIMPLE_SEGMENT|12909,12919|false|false|false|||supplement
Finding|Functional Concept|SIMPLE_SEGMENT|12909,12919|false|false|false|C1549514;C1947943;C2348609|Supplement;Supplement (document);Supplement - Diet Code Specification Type|supplement
Finding|Idea or Concept|SIMPLE_SEGMENT|12909,12919|false|false|false|C1549514;C1947943;C2348609|Supplement;Supplement (document);Supplement - Diet Code Specification Type|supplement
Finding|Intellectual Product|SIMPLE_SEGMENT|12909,12919|false|false|false|C1549514;C1947943;C2348609|Supplement;Supplement (document);Supplement - Diet Code Specification Type|supplement
Drug|Biologically Active Substance|SIMPLE_SEGMENT|12938,12947|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|12938,12947|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Food|SIMPLE_SEGMENT|12938,12947|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|12938,12947|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12938,12947|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Event|Event|SIMPLE_SEGMENT|12938,12947|false|false|false|||potassium
Finding|Physiologic Function|SIMPLE_SEGMENT|12938,12947|false|false|false|C4553027|Potassium metabolic function|potassium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|12938,12947|false|false|false|C0202194|Potassium measurement|potassium
Event|Event|SIMPLE_SEGMENT|12948,12954|false|false|false|||levels
Event|Event|SIMPLE_SEGMENT|12960,12966|false|false|false|||normal
Finding|Idea or Concept|SIMPLE_SEGMENT|12974,12982|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|SIMPLE_SEGMENT|12987,12995|false|false|false|||Increase
Drug|Organic Chemical|SIMPLE_SEGMENT|13001,13013|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13001,13013|false|false|false|C0286651|atorvastatin|atorvastatin
Event|Event|SIMPLE_SEGMENT|13001,13013|false|false|false|||atorvastatin
Drug|Organic Chemical|SIMPLE_SEGMENT|13015,13022|false|false|false|C0593906|Lipitor|lipitor
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13015,13022|false|false|false|C0593906|Lipitor|lipitor
Event|Event|SIMPLE_SEGMENT|13015,13022|false|false|false|||lipitor
Event|Event|SIMPLE_SEGMENT|13024,13028|false|false|false|||dose
Event|Event|SIMPLE_SEGMENT|13058,13062|false|false|false|||Stop
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|13068,13078|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13068,13078|false|false|false|C0065374|lisinopril|lisinopril
Event|Event|SIMPLE_SEGMENT|13068,13078|false|false|false|||lisinopril
Drug|Organic Chemical|SIMPLE_SEGMENT|13083,13088|false|false|false|C0699992|Lasix|lasix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13083,13088|false|false|false|C0699992|Lasix|lasix
Event|Event|SIMPLE_SEGMENT|13083,13088|false|false|false|||lasix
Drug|Organic Chemical|SIMPLE_SEGMENT|13090,13100|false|false|false|C0016860|furosemide|furosemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13090,13100|false|false|false|C0016860|furosemide|furosemide
Event|Event|SIMPLE_SEGMENT|13090,13100|false|false|false|||furosemide
Event|Event|SIMPLE_SEGMENT|13119,13129|false|false|false|||instructed
Finding|Intellectual Product|SIMPLE_SEGMENT|13138,13150|false|false|false|C1547426|Location Service Code - Primary Care|primary care
Procedure|Health Care Activity|SIMPLE_SEGMENT|13138,13150|false|false|false|C0033137|Primary Health Care|primary care
Event|Activity|SIMPLE_SEGMENT|13146,13150|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|13146,13150|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|13146,13150|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|13146,13150|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13151,13160|false|false|false|C0804815||physician
Event|Event|SIMPLE_SEGMENT|13171,13175|false|false|false|||need
Event|Event|SIMPLE_SEGMENT|13176,13182|false|false|false|||repeat
Finding|Functional Concept|SIMPLE_SEGMENT|13176,13182|false|false|false|C0205341;C1705914|Repeat;Repeat Object|repeat
Event|Event|SIMPLE_SEGMENT|13184,13193|false|false|false|||bloodwork
Event|Event|SIMPLE_SEGMENT|13218,13222|false|false|false|||sent
Finding|Intellectual Product|SIMPLE_SEGMENT|13232,13244|false|false|false|C1547426|Location Service Code - Primary Care|primary care
Procedure|Health Care Activity|SIMPLE_SEGMENT|13232,13244|false|false|false|C0033137|Primary Health Care|primary care
Event|Activity|SIMPLE_SEGMENT|13240,13244|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|13240,13244|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|13240,13244|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|13240,13244|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13245,13254|false|false|false|C0804815||physician
Event|Event|SIMPLE_SEGMENT|13262,13266|false|false|false|||Keep
Finding|Idea or Concept|SIMPLE_SEGMENT|13271,13279|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|SIMPLE_SEGMENT|13280,13286|false|false|false|||follow
Event|Activity|SIMPLE_SEGMENT|13290,13302|false|false|false|C0003629|Appointments|appointments
Event|Event|SIMPLE_SEGMENT|13290,13302|false|false|false|||appointments
Event|Event|SIMPLE_SEGMENT|13312,13318|false|false|false|||coming
Event|Activity|SIMPLE_SEGMENT|13320,13332|false|false|false|C0003629|Appointments|appointments
Event|Event|SIMPLE_SEGMENT|13320,13332|false|false|false|||appointments
Event|Event|SIMPLE_SEGMENT|13337,13343|false|false|false|||listed
Procedure|Health Care Activity|SIMPLE_SEGMENT|13354,13362|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13363,13375|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|13363,13375|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|13363,13375|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

