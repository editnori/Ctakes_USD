 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Procedure|Health Care Activity|SIMPLE_SEGMENT|47,56|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|47,61|false|false|false|C2598112||Admission Date
Finding|Body Substance|SIMPLE_SEGMENT|81,90|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|81,90|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|81,90|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|81,90|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|81,95|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|113,118|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|113,118|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|113,118|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|137,140|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|137,140|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|137,140|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|137,140|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|137,140|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|148,155|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|148,155|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|157,165|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|Allergies|189,198|false|false|false|C1717415||Allergies
Finding|Pathologic Function|Allergies|189,198|false|false|false|C0020517|Hypersensitivity|Allergies
Finding|Pathologic Function|Allergies|201,223|true|false|false|C0041755|Adverse reaction to drug|Adverse Drug Reactions
Drug|Pharmacologic Substance|Allergies|209,213|false|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|Drug
Finding|Finding|Allergies|209,213|false|false|false|C0740721|Drug problem|Drug
Finding|Pathologic Function|Allergies|209,223|true|false|false|C0041755|Adverse reaction to drug|Drug Reactions
Finding|Functional Concept|Allergies|226,235|false|false|false|C1999232|Attending (action)|Attending
Disorder|Disease or Syndrome|Chief Complaint|278,284|false|false|false|C4255010||NSTEMI
Finding|Finding|Chief Complaint|278,284|false|false|false|C3537184||NSTEMI
Finding|Classification|Chief Complaint|287,292|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|293,301|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|293,301|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|305,323|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|314,323|false|false|false|C0945766||Procedure
Event|Occupational Activity|Chief Complaint|314,323|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|314,323|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|314,323|false|false|false|C0184661|Interventional procedure|Procedure
Anatomy|Body Part, Organ, or Organ Component|Chief Complaint|327,334|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|Chief Complaint|327,334|false|false|false|C1314974|Cardiac attachment|cardiac
Disorder|Injury or Poisoning|Chief Complaint|327,350|false|false|false|C0261588|Cardiac catheterisation as the cause of abnormal reaction of the patient, or of later complication, without mention of misadventure at the time of the procedure|cardiac catheterization
Finding|Intellectual Product|Chief Complaint|327,350|false|false|false|C1547981|Diagnostic Service Section ID - Cardiac Catheterization|cardiac catheterization
Procedure|Diagnostic Procedure|Chief Complaint|327,350|false|false|false|C0018795;C1548828|Cardiac Catheterization Procedures;Consent Type - Cardiac Catheterization|cardiac catheterization
Procedure|Health Care Activity|Chief Complaint|327,350|false|false|false|C0018795;C1548828|Cardiac Catheterization Procedures;Consent Type - Cardiac Catheterization|cardiac catheterization
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|335,350|false|false|false|C0007430|Catheterization|catheterization
Disorder|Disease or Syndrome|Chief Complaint|356,359|false|false|false|C4551552|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|DES
Drug|Amino Acid, Peptide, or Protein|Chief Complaint|356,359|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Biologically Active Substance|Chief Complaint|356,359|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Hormone|Chief Complaint|356,359|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Organic Chemical|Chief Complaint|356,359|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Pharmacologic Substance|Chief Complaint|356,359|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Finding|Gene or Genome|Chief Complaint|356,359|false|false|false|C1413980|DES gene|DES
Disorder|Acquired Abnormality|Chief Complaint|371,380|false|false|false|C0001168|Complete obstruction|occlusion
Finding|Finding|Chief Complaint|371,380|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Functional Concept|Chief Complaint|371,380|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Organ or Tissue Function|Chief Complaint|371,380|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Pathologic Function|Chief Complaint|371,380|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Conceptual Entity|Chief Complaint|388,394|false|false|false|C0442038;C0920847|Circumpennate;Radial|radial
Finding|Functional Concept|Chief Complaint|395,401|false|false|false|C1554204|Role Class - access|access
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|404,408|false|false|false|C0021860|Intra-Aortic Balloon Pumping|IABP
Procedure|Health Care Activity|Chief Complaint|409,418|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|409,418|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Event|Activity|Chief Complaint|423,430|false|false|false|C1883720|Removing (action)|removal
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|423,430|false|false|false|C0015252;C0185115;C0728940|Excision;Extraction;removal technique|removal
Disorder|Disease or Syndrome|History of Present Illness|485,488|false|false|false|C0020538|Hypertensive disease|HTN
Finding|Functional Concept|History of Present Illness|520,527|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Idea or Concept|History of Present Illness|520,527|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Intellectual Product|History of Present Illness|520,527|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Procedure|Health Care Activity|History of Present Illness|520,527|false|false|false|C0199168|Medical service|medical
Event|Occupational Activity|History of Present Illness|528,538|false|false|false|C0001554;C1273870|Administration occupational activities;Management procedure|management
Procedure|Health Care Activity|History of Present Illness|528,538|false|false|false|C0376636|Disease Management|management
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|543,547|false|false|false|C0007430|Catheterization|cath
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|598,613|false|false|false|C0007430|Catheterization|catheterization
Finding|Idea or Concept|History of Present Illness|618,625|false|false|false|C2699424|Concern|concern
Disorder|Disease or Syndrome|History of Present Illness|630,635|false|false|false|C1536220|ST segment elevation myocardial infarction|STEMI
Finding|Finding|History of Present Illness|630,635|false|false|false|C3538872|ST Elevation Myocardial Infarction by ECG Finding|STEMI
Finding|Body Substance|History of Present Illness|639,646|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|639,646|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|639,646|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Functional Concept|History of Present Illness|639,650|false|false|false|C0332310|Has patient|Patient has
Attribute|Clinical Attribute|History of Present Illness|665,671|false|false|false|C2926611||angina
Finding|Finding|History of Present Illness|665,671|false|false|false|C0002962;C2024883|Angina Pectoris|angina
Finding|Sign or Symptom|History of Present Illness|665,671|false|false|false|C0002962;C2024883|Angina Pectoris|angina
Finding|Sign or Symptom|History of Present Illness|665,676|false|false|false|C0002962|Angina Pectoris|angina pain
Attribute|Clinical Attribute|History of Present Illness|672,676|false|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|672,676|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|672,676|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Organism Function|History of Present Illness|680,688|false|false|false|C0015264|Exertion|exertion
Finding|Intellectual Product|History of Present Illness|708,713|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Intellectual Product|History of Present Illness|708,719|false|false|false|C1272517|Sudden onset (contextual qualifier) (qualifier value)|acute onset
Finding|Finding|History of Present Illness|767,770|false|false|false|C1417953;C1847730;C5575300|GLAUCOMA, NORMAL TENSION, SUSCEPTIBILITY TO;OPA1 gene;OPA1 wt Allele|NTG
Finding|Gene or Genome|History of Present Illness|767,770|false|false|false|C1417953;C1847730;C5575300|GLAUCOMA, NORMAL TENSION, SUSCEPTIBILITY TO;OPA1 gene;OPA1 wt Allele|NTG
Finding|Functional Concept|History of Present Illness|805,813|false|false|false|C0332287;C1883712|Add - instruction imperative;In addition to|addition
Finding|Finding|History of Present Illness|833,841|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|History of Present Illness|833,841|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|History of Present Illness|846,854|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Finding|Sign or Symptom|History of Present Illness|855,862|false|false|false|C0231218|Malaise|malaise
Finding|Finding|History of Present Illness|886,895|false|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Finding|Sign or Symptom|History of Present Illness|886,895|false|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Disorder|Disease or Syndrome|History of Present Illness|897,900|false|false|false|C1956415|Paroxysmal nocturnal dyspnea|PND
Finding|Gene or Genome|History of Present Illness|897,900|false|false|false|C1417807;C4552608|NPPA gene;NPPA wt Allele|PND
Attribute|Clinical Attribute|History of Present Illness|906,911|false|false|false|C1717255||edema
Finding|Pathologic Function|History of Present Illness|906,911|false|false|false|C0013604|Edema|edema
Finding|Finding|History of Present Illness|913,925|false|false|false|C0030252|Palpitations|palpitations
Finding|Sign or Symptom|History of Present Illness|930,933|false|false|false|C0013404|Dyspnea|SOB
Finding|Idea or Concept|History of Present Illness|948,955|false|false|false|C1555582|Initial (abbreviation)|initial
Finding|Functional Concept|History of Present Illness|971,975|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|History of Present Illness|971,975|false|false|false|C0582103|Medical Examination|Exam
Anatomy|Body Location or Region|History of Present Illness|977,982|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|History of Present Illness|977,982|false|false|false|C0741025|Chest problem|Chest
Attribute|Clinical Attribute|History of Present Illness|977,987|false|false|false|C2926613||Chest pain
Finding|Sign or Symptom|History of Present Illness|977,987|false|false|false|C0008031|Chest Pain|Chest pain
Attribute|Clinical Attribute|History of Present Illness|983,987|false|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|983,987|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|983,987|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Lab|Laboratory or Test Result|History of Present Illness|1005,1009|false|false|false|C0587081|Laboratory test finding|Labs
Anatomy|Cell|History of Present Illness|1024,1027|false|false|false|C0023516|Leukocytes|WBC
Procedure|Laboratory Procedure|History of Present Illness|1034,1037|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1034,1037|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Laboratory Procedure|History of Present Illness|1044,1047|false|false|false|C0201617|Primed lymphocyte test|Plt
Attribute|Clinical Attribute|History of Present Illness|1053,1056|false|false|false|C0368980|Coagulation tissue factor induced.INR|INR
Procedure|Laboratory Procedure|History of Present Illness|1053,1056|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1053,1056|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Drug|Biologically Active Substance|History of Present Illness|1080,1083|false|false|false|C0600137|Blood Urea Nitrogen|BUN
Drug|Inorganic Chemical|History of Present Illness|1080,1083|false|false|false|C0600137|Blood Urea Nitrogen|BUN
Procedure|Laboratory Procedure|History of Present Illness|1080,1083|false|false|false|C0005845|Blood urea nitrogen measurement|BUN
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1087,1090|false|false|false|C0056182;C1721462|CR1 protein, human;Complement 3b Receptor|Cr1
Drug|Immunologic Factor|History of Present Illness|1087,1090|false|false|false|C0056182;C1721462|CR1 protein, human;Complement 3b Receptor|Cr1
Finding|Gene or Genome|History of Present Illness|1087,1090|false|false|false|C0056182;C1413694;C1721462|CR1 gene;CR1 protein, human;Complement 3b Receptor|Cr1
Finding|Receptor|History of Present Illness|1087,1090|false|false|false|C0056182;C1413694;C1721462|CR1 gene;CR1 protein, human;Complement 3b Receptor|Cr1
Finding|Finding|History of Present Illness|1094,1101|false|false|false|C0740845|Imaging problem|Imaging
Procedure|Diagnostic Procedure|History of Present Illness|1094,1101|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|Imaging
Finding|Intellectual Product|History of Present Illness|1103,1106|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|History of Present Illness|1103,1106|false|false|false|C1623258|Electrocardiography|EKG
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1154,1163|false|false|false|C0439775|Elevation procedure|elevation
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|1196,1207|false|false|false|C0011570|Mental Depression|depressions
Procedure|Health Care Activity|History of Present Illness|1218,1222|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1218,1222|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Attribute|Clinical Attribute|History of Present Illness|1233,1244|false|false|false|C1980023|Wall motion|wall motion
Phenomenon|Natural Phenomenon or Process|History of Present Illness|1238,1244|false|false|false|C0026597|Motion|motion
Disorder|Congenital Abnormality|History of Present Illness|1245,1258|false|false|false|C0000768|Congenital Abnormality|abnormalities
Finding|Functional Concept|History of Present Illness|1245,1258|false|false|false|C0000769|teratologic|abnormalities
Procedure|Diagnostic Procedure|History of Present Illness|1260,1263|false|false|false|C0039985|Plain chest X-ray|CXR
Finding|Intellectual Product|History of Present Illness|1272,1277|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Disorder|Congenital Abnormality|History of Present Illness|1279,1292|false|false|false|C0000768|Congenital Abnormality|abnormalities
Finding|Functional Concept|History of Present Illness|1279,1292|false|false|false|C0000769|teratologic|abnormalities
Finding|Body Substance|History of Present Illness|1295,1302|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|1295,1302|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|1295,1302|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Biologically Active Substance|History of Present Illness|1314,1321|false|false|false|C0019134;C0770546|heparin;heparin, porcine|Heparin
Drug|Organic Chemical|History of Present Illness|1314,1321|false|false|false|C0019134;C0770546|heparin;heparin, porcine|Heparin
Drug|Pharmacologic Substance|History of Present Illness|1314,1321|false|false|false|C0019134;C0770546|heparin;heparin, porcine|Heparin
Disorder|Neoplastic Process|History of Present Illness|1322,1325|false|false|false|C1135868|Gestational Trophoblastic Neoplasms|gtt
Drug|Biomedical or Dental Material|History of Present Illness|1322,1325|false|false|false|C0991568|Drops - Drug Form|gtt
Procedure|Laboratory Procedure|History of Present Illness|1322,1325|false|false|false|C0017741|Glucose tolerance test|gtt
Disorder|Neoplastic Process|History of Present Illness|1333,1336|false|false|false|C1135868|Gestational Trophoblastic Neoplasms|gtt
Drug|Biomedical or Dental Material|History of Present Illness|1333,1336|false|false|false|C0991568|Drops - Drug Form|gtt
Procedure|Laboratory Procedure|History of Present Illness|1333,1336|false|false|false|C0017741|Glucose tolerance test|gtt
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1338,1341|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Enzyme|History of Present Illness|1338,1341|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Organic Chemical|History of Present Illness|1338,1341|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Pharmacologic Substance|History of Present Illness|1338,1341|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Finding|Gene or Genome|History of Present Illness|1338,1341|false|false|false|C1412553|ARSA gene|ASA
Drug|Nucleic Acid, Nucleoside, or Nucleotide|History of Present Illness|1349,1359|false|false|false|C1999375|ticagrelor|Ticagrelor
Drug|Pharmacologic Substance|History of Present Illness|1349,1359|false|false|false|C1999375|ticagrelor|Ticagrelor
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1375,1380|false|false|false|C0042313|vancomycin|Vanco
Drug|Antibiotic|History of Present Illness|1375,1380|false|false|false|C0042313|vancomycin|Vanco
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1419,1426|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|History of Present Illness|1419,1426|false|false|false|C1314974|Cardiac attachment|cardiac
Procedure|Diagnostic Procedure|History of Present Illness|1419,1431|false|false|false|C0018795|Cardiac Catheterization Procedures|cardiac cath
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1427,1431|false|false|false|C0007430|Catheterization|cath
Finding|Functional Concept|History of Present Illness|1443,1451|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|History of Present Illness|1443,1451|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|History of Present Illness|1443,1451|false|false|false|C4706767|Transfer (immobility management)|transfer
Finding|Finding|History of Present Illness|1483,1491|false|false|false|C0277797|Apyrexial|afebrile
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1492,1496|false|false|false|C0007430|Catheterization|Cath
Finding|Gene or Genome|History of Present Illness|1497,1500|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|lab
Finding|Intellectual Product|History of Present Illness|1497,1500|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|lab
Disorder|Disease or Syndrome|History of Present Illness|1510,1515|false|false|false|C1410088|Still|still
Attribute|Clinical Attribute|History of Present Illness|1524,1528|false|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|1524,1528|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1524,1528|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Biologically Active Substance|History of Present Illness|1532,1539|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Organic Chemical|History of Present Illness|1532,1539|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Pharmacologic Substance|History of Present Illness|1532,1539|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Disorder|Neoplastic Process|History of Present Illness|1550,1553|false|false|false|C1135868|Gestational Trophoblastic Neoplasms|gtt
Drug|Biomedical or Dental Material|History of Present Illness|1550,1553|false|false|false|C0991568|Drops - Drug Form|gtt
Procedure|Laboratory Procedure|History of Present Illness|1550,1553|false|false|false|C0017741|Glucose tolerance test|gtt
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1556,1571|false|false|false|C0007430|Catheterization|Catheterization
Disorder|Acquired Abnormality|History of Present Illness|1594,1603|false|false|false|C0001168|Complete obstruction|occlusion
Finding|Finding|History of Present Illness|1594,1603|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Functional Concept|History of Present Illness|1594,1603|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Organ or Tissue Function|History of Present Illness|1594,1603|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Pathologic Function|History of Present Illness|1594,1603|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Disorder|Disease or Syndrome|History of Present Illness|1613,1620|false|false|false|C0012634|Disease|disease
Drug|Organic Chemical|History of Present Illness|1638,1646|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|History of Present Illness|1638,1646|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|History of Present Illness|1638,1646|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Finding|Functional Concept|History of Present Illness|1638,1646|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|History of Present Illness|1638,1646|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Disorder|Acquired Abnormality|History of Present Illness|1647,1656|false|false|false|C0001168|Complete obstruction|occlusion
Finding|Finding|History of Present Illness|1647,1656|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Functional Concept|History of Present Illness|1647,1656|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Organ or Tissue Function|History of Present Illness|1647,1656|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Pathologic Function|History of Present Illness|1647,1656|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Pathologic Function|History of Present Illness|1696,1704|false|false|false|C1261287|Stenosis|stenosis
Disorder|Disease or Syndrome|History of Present Illness|1716,1719|false|false|false|C4551552|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|DES
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1716,1719|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Biologically Active Substance|History of Present Illness|1716,1719|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Hormone|History of Present Illness|1716,1719|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Organic Chemical|History of Present Illness|1716,1719|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Pharmacologic Substance|History of Present Illness|1716,1719|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Finding|Gene or Genome|History of Present Illness|1716,1719|false|false|false|C1413980|DES gene|DES
Disorder|Acquired Abnormality|History of Present Illness|1731,1740|false|false|false|C0001168|Complete obstruction|occlusion
Finding|Finding|History of Present Illness|1731,1740|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Functional Concept|History of Present Illness|1731,1740|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Organ or Tissue Function|History of Present Illness|1731,1740|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Pathologic Function|History of Present Illness|1731,1740|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Conceptual Entity|History of Present Illness|1748,1754|false|false|false|C0442038;C0920847|Circumpennate;Radial|radial
Finding|Functional Concept|History of Present Illness|1755,1761|false|false|false|C1554204|Role Class - access|access
Finding|Pathologic Function|History of Present Illness|1763,1774|false|false|false|C0857353|Hypotensive|Hypotensive
Anatomy|Body Space or Junction|History of Present Illness|1801,1804|false|false|false|C0016520|Structure of interventricular foramen|IVF
Disorder|Disease or Syndrome|History of Present Illness|1801,1804|false|false|false|C2751898|Ventricular Fibrillation, Paroxysmal Familial, 1|IVF
Finding|Gene or Genome|History of Present Illness|1801,1804|false|false|false|C1419864;C4321334|SCN5A gene;SCN5A wt Allele|IVF
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1801,1804|false|false|false|C0015915;C0872104|Assisted Reproductive Technologies;Fertilization in Vitro|IVF
Finding|Sign or Symptom|History of Present Illness|1807,1815|false|false|false|C0010200|Coughing|Coughing
Finding|Finding|History of Present Illness|1836,1841|false|false|false|C0456190|Left ventricular end-diastolic pressure|LVEDP
Drug|Organic Chemical|History of Present Illness|1854,1859|false|false|false|C0699992|Lasix|Lasix
Drug|Pharmacologic Substance|History of Present Illness|1854,1859|false|false|false|C0699992|Lasix|Lasix
Finding|Intellectual Product|History of Present Illness|1874,1878|false|false|false|C1720594|Then - dosing instruction fragment|then
Finding|Finding|History of Present Illness|1879,1891|false|false|false|C0857121|Hypertensive (finding)|hypertensive
Drug|Organic Chemical|History of Present Illness|1916,1921|false|false|false|C0699992|Lasix|Lasix
Drug|Pharmacologic Substance|History of Present Illness|1916,1921|false|false|false|C0699992|Lasix|Lasix
Finding|Finding|History of Present Illness|1952,1963|false|false|false|C0020649|Hypotension|hypotension
Attribute|Clinical Attribute|History of Present Illness|1975,1984|false|false|false|C0945766||procedure
Event|Occupational Activity|History of Present Illness|1975,1984|false|false|false|C1546467|Act Class - procedure|procedure
Finding|Functional Concept|History of Present Illness|1975,1984|false|false|false|C2700391|Procedure (set of actions)|procedure
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1975,1984|false|false|false|C0184661|Interventional procedure|procedure
Anatomy|Cell|History of Present Illness|1986,1989|false|false|false|C0023516|Leukocytes|WBC
Finding|Body Substance|History of Present Illness|2029,2036|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|2029,2036|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|2029,2036|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Anatomy|Body Location or Region|History of Present Illness|2048,2053|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|2048,2053|true|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|History of Present Illness|2048,2058|true|false|false|C2926613||chest pain
Finding|Sign or Symptom|History of Present Illness|2048,2058|true|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|History of Present Illness|2054,2058|true|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|2054,2058|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|2054,2058|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|History of Present Illness|2082,2098|false|false|false|C0239134|Productive Cough|productive cough
Drug|Organic Chemical|History of Present Illness|2093,2098|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|History of Present Illness|2093,2098|false|false|false|C3815497|Cough (guaifenesin)|cough
Finding|Sign or Symptom|History of Present Illness|2093,2098|false|false|false|C0010200|Coughing|cough
Finding|Finding|History of Present Illness|2103,2111|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|History of Present Illness|2103,2111|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Gene or Genome|History of Present Illness|2133,2136|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Procedure|Diagnostic Procedure|History of Present Illness|2141,2150|false|false|false|C0014245;C0079278|Endoscopy (procedure);Endoscopy, Gastrointestinal|endoscopy
Drug|Antibiotic|History of Present Illness|2194,2208|false|false|false|C0055856|clarithromycin|clarithromycin
Drug|Organic Chemical|History of Present Illness|2194,2208|false|false|false|C0055856|clarithromycin|clarithromycin
Drug|Antibiotic|History of Present Illness|2213,2224|false|false|false|C0002645|amoxicillin|amoxicillin
Drug|Organic Chemical|History of Present Illness|2213,2224|false|false|false|C0002645|amoxicillin|amoxicillin
Finding|Finding|History of Present Illness|2250,2258|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|History of Present Illness|2250,2258|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Attribute|Clinical Attribute|History of Present Illness|2274,2280|false|false|false|C0944911||weight
Finding|Finding|History of Present Illness|2274,2280|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|History of Present Illness|2274,2280|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|History of Present Illness|2274,2280|false|false|false|C1305866|Weighing patient|weight
Finding|Finding|History of Present Illness|2274,2285|false|false|false|C1262477;C3540682|Losing Weight (question);Weight Loss|weight loss
Finding|Intellectual Product|History of Present Illness|2274,2285|false|false|false|C1262477;C3540682|Losing Weight (question);Weight Loss|weight loss
Finding|Finding|History of Present Illness|2281,2285|false|false|false|C5890125|Loss (adaptation)|loss
Disorder|Disease or Syndrome|Past Medical History|2333,2336|false|false|false|C0020538|Hypertensive disease|HTN
Disorder|Disease or Syndrome|Past Medical History|2355,2358|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Past Medical History|2355,2358|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Past Medical History|2355,2358|false|false|false|C1504769|DFFB protein, human|CAD
Finding|Gene or Genome|Past Medical History|2355,2358|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Past Medical History|2355,2358|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Past Medical History|2355,2358|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2355,2358|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Event|Occupational Activity|Past Medical History|2378,2385|false|false|false|C1273870|Management procedure|managed
Disorder|Acquired Abnormality|Past Medical History|2402,2417|false|false|false|C0037944;C1861329|Spinal Stenosis;Spinal canal stenosis|Spinal stenosis
Disorder|Anatomical Abnormality|Past Medical History|2402,2417|false|false|false|C0037944;C1861329|Spinal Stenosis;Spinal canal stenosis|Spinal stenosis
Finding|Pathologic Function|Past Medical History|2409,2417|false|false|false|C1261287|Stenosis|stenosis
Finding|Conceptual Entity|Family Medical History|2456,2462|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Idea or Concept|Family Medical History|2456,2462|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Finding|Family Medical History|2464,2472|false|false|false|C0332149|Possible|possible
Disorder|Disease or Syndrome|Family Medical History|2481,2495|false|true|false|C0878544|Cardiomyopathies|cardiomyopathy
Finding|Classification|Family Medical History|2499,2505|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|Family Medical History|2499,2505|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|Family Medical History|2499,2505|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|Family Medical History|2499,2505|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Finding|Family Medical History|2499,2513|true|false|false|C0241889|Family Medical History|family history
Finding|Finding|Family Medical History|2499,2516|true|false|false|C0241889|Family Medical History|family history of
Finding|Conceptual Entity|Family Medical History|2506,2513|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|2506,2513|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Family Medical History|2506,2513|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|2506,2516|true|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|Family Medical History|2527,2537|true|false|false|C0003811|Cardiac Arrhythmia|arrhythmia
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2549,2556|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|Family Medical History|2549,2556|false|false|false|C1314974|Cardiac attachment|cardiac
Finding|Finding|Family Medical History|2558,2563|false|false|false|C0011065;C1306577;C1546949|Cessation of life;Death (finding);Event Consequence - Death|death
Finding|Idea or Concept|Family Medical History|2558,2563|false|false|false|C0011065;C1306577;C1546949|Cessation of life;Death (finding);Event Consequence - Death|death
Finding|Organism Function|Family Medical History|2558,2563|false|false|false|C0011065;C1306577;C1546949|Cessation of life;Death (finding);Event Consequence - Death|death
Procedure|Health Care Activity|General Exam|2615,2624|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Finding|General Exam|2646,2654|false|false|false|C0277797|Apyrexial|afebrile
Attribute|Clinical Attribute|General Exam|2695,2701|false|false|false|C0944911||Weight
Finding|Finding|General Exam|2695,2701|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|Weight
Finding|Sign or Symptom|General Exam|2695,2701|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|Weight
Procedure|Health Care Activity|General Exam|2695,2701|false|false|false|C1305866|Weighing patient|Weight
Finding|Gene or Genome|General Exam|2708,2712|false|false|false|C1420621;C1515258|TCAP gene;Telephone Number|Tele
Finding|Intellectual Product|General Exam|2708,2712|false|false|false|C1420621;C1515258|TCAP gene;Telephone Number|Tele
Finding|Molecular Function|General Exam|2714,2717|false|false|false|C1704493;C2700623|Neutral Sidebent Rotated|NSR
Finding|Pathologic Function|General Exam|2714,2717|false|false|false|C1704493;C2700623|Neutral Sidebent Rotated|NSR
Finding|Classification|General Exam|2718,2721|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Finding|Gene or Genome|General Exam|2718,2721|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Finding|Finding|General Exam|2732,2742|false|false|false|C0231835|Tachypnea|tachypneic
Finding|Sign or Symptom|General Exam|2761,2769|false|false|false|C0043144|Wheezing|wheezing
Finding|Intellectual Product|General Exam|2797,2806|false|false|false|C0876929|Sentence|sentences
Anatomy|Body Location or Region|General Exam|2808,2813|false|false|false|C1512338|HEENT|HEENT
Finding|Finding|General Exam|2821,2827|false|false|false|C2143306|PERRLA|PERRLA
Anatomy|Body Location or Region|General Exam|2829,2833|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|General Exam|2829,2833|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|General Exam|2829,2833|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Finding|Finding|General Exam|2838,2841|true|false|false|C0425687|Jugular venous engorgement|JVD
Finding|Finding|General Exam|2859,2868|false|false|false|C0332218|Difficult (qualifier value)|difficult
Anatomy|Body Part, Organ, or Organ Component|General Exam|2883,2888|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|General Exam|2883,2888|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|General Exam|2883,2888|false|false|false|C0795691|HEART PROBLEM|heart
Attribute|Clinical Attribute|General Exam|2883,2895|false|false|false|C4050434||heart sounds
Finding|Organ or Tissue Function|General Exam|2883,2895|false|false|false|C0018820|Heart Sounds|heart sounds
Procedure|Diagnostic Procedure|General Exam|2883,2895|false|false|false|C2230284|auscultation of heart sounds|heart sounds
Phenomenon|Natural Phenomenon or Process|General Exam|2889,2895|false|false|false|C0037709||sounds
Finding|Idea or Concept|General Exam|2904,2915|false|false|false|C0750502|Significant|significant
Finding|Finding|General Exam|2916,2923|false|false|false|C0035508|Rhonchi|rhonchi
Anatomy|Body Part, Organ, or Organ Component|General Exam|2925,2930|false|false|false|C0024109|Lung|LUNGS
Finding|Finding|General Exam|2936,2943|false|false|false|C0035508|Rhonchi|rhonchi
Finding|Intellectual Product|General Exam|2958,2962|false|false|false|C1547225|Mild Severity of Illness Code|mild
Drug|Amino Acid, Peptide, or Protein|General Exam|2963,2966|false|false|false|C0082420|Endoglin, human|end
Drug|Immunologic Factor|General Exam|2963,2966|false|false|false|C0082420|Endoglin, human|end
Finding|Functional Concept|General Exam|2963,2966|false|false|false|C1366583;C1561490;C1704837|ENG gene;ENG wt Allele;end - ActRelationshipCheckpoint|end
Finding|Gene or Genome|General Exam|2963,2966|false|false|false|C1366583;C1561490;C1704837|ENG gene;ENG wt Allele;end - ActRelationshipCheckpoint|end
Finding|Organism Function|General Exam|2967,2977|false|false|false|C0231800|Expiration, Respiratory|expiratory
Finding|Sign or Symptom|General Exam|2967,2986|false|false|false|C0231875|Expiratory wheezing|expiratory wheezing
Finding|Sign or Symptom|General Exam|2978,2986|false|false|false|C0043144|Wheezing|wheezing
Anatomy|Body Location or Region|General Exam|2994,2998|false|false|false|C2987514|Anatomical base|base
Drug|Biomedical or Dental Material|General Exam|2994,2998|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Chemical Viewed Functionally|General Exam|2994,2998|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|2994,2998|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Finding|Gene or Genome|General Exam|2994,2998|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Finding|Idea or Concept|General Exam|2994,2998|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Finding|Finding|General Exam|2999,3007|false|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Anatomy|Body Location or Region|General Exam|3008,3011|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|ABD
Disorder|Cell or Molecular Dysfunction|General Exam|3008,3011|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|ABD
Disorder|Disease or Syndrome|General Exam|3013,3017|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Disorder|Congenital Abnormality|General Exam|3045,3048|false|false|false|C0015306|Hereditary Multiple Exostoses|EXT
Finding|Gene or Genome|General Exam|3045,3048|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|EXT
Finding|Conceptual Entity|General Exam|3055,3061|false|false|false|C0442038;C0920847|Circumpennate;Radial|radial
Drug|Food|General Exam|3062,3068|false|false|false|C5890763||pulses
Finding|Physiologic Function|General Exam|3062,3068|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|General Exam|3062,3068|false|false|false|C0034107|Pulse taking|pulses
Anatomy|Body Part, Organ, or Organ Component|General Exam|3070,3075|false|false|false|C4048756|Right arm|R arm
Anatomy|Body Part, Organ, or Organ Component|General Exam|3072,3075|false|false|false|C0446516;C1140618;C1269078|Upper Extremity;Upper arm|arm
Disorder|Anatomical Abnormality|General Exam|3072,3075|false|false|false|C3495676|Anorectal Malformations|arm
Finding|Gene or Genome|General Exam|3072,3075|false|false|false|C1824218;C3715044|AKR1A1 wt Allele;ARMC9 gene|arm
Procedure|Diagnostic Procedure|General Exam|3072,3075|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Research Activity|General Exam|3072,3075|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Therapeutic or Preventive Procedure|General Exam|3072,3075|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Event|Activity|General Exam|3087,3092|false|false|false|C1882509|put - instruction imperative|place
Finding|Functional Concept|General Exam|3087,3092|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|General Exam|3087,3092|false|false|false|C1533810||place
Finding|Functional Concept|General Exam|3105,3110|false|false|false|C1513492|motor movement|motor
Finding|Organ or Tissue Function|General Exam|3111,3127|false|false|false|C0036658|Sensory perception|sensory function
Finding|Finding|General Exam|3119,3127|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|General Exam|3119,3127|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|General Exam|3119,3127|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|General Exam|3119,3127|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Finding|General Exam|3128,3134|false|false|false|C1554187|Gender Status - Intact|intact
Disorder|Disease or Syndrome|General Exam|3211,3215|false|false|false|C0009443;C0024117|Chronic Obstructive Airway Disease;Common Cold|cold
Drug|Organic Chemical|General Exam|3211,3215|false|false|false|C0719425|Cold brand of chlorpheniramine-phenylpropanolamine|cold
Drug|Pharmacologic Substance|General Exam|3211,3215|false|false|false|C0719425|Cold brand of chlorpheniramine-phenylpropanolamine|cold
Finding|Organism Function|General Exam|3211,3215|false|false|false|C0234192|Cold Sensation|cold
Phenomenon|Natural Phenomenon or Process|General Exam|3211,3215|false|false|false|C0009264|Cold Temperature|cold
Procedure|Therapeutic or Preventive Procedure|General Exam|3211,3215|false|false|false|C0010412|Cold Therapy|cold
Finding|Finding|General Exam|3228,3237|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|General Exam|3228,3237|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|General Exam|3228,3237|false|false|false|C2229507|sensory exam|sensation
Finding|Functional Concept|General Exam|3246,3251|false|false|false|C1513492|motor movement|motor
Finding|Idea or Concept|General Exam|3252,3260|false|false|false|C0808080|Strength (attribute)|strength
Finding|Finding|General Exam|3265,3268|false|false|false|C0948106;C1419600|ROM1 gene;Rupture of Membranes|ROM
Finding|Gene or Genome|General Exam|3265,3268|false|false|false|C0948106;C1419600|ROM1 gene;Rupture of Membranes|ROM
Procedure|Laboratory Procedure|General Exam|3265,3268|false|false|false|C1562926|Range of motion technique (procedure)|ROM
Anatomy|Body System|General Exam|3269,3273|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|General Exam|3269,3273|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|General Exam|3269,3273|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Finding|Body Substance|General Exam|3269,3273|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|General Exam|3269,3273|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Sign or Symptom|General Exam|3278,3284|true|false|false|C0015230;C5779628|Exanthema;Skin rash|rashes
Finding|Intellectual Product|General Exam|3288,3295|true|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|General Exam|3288,3295|true|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Finding|Pathologic Function|General Exam|3296,3305|false|false|false|C0013604|Edema|edematous
Finding|Functional Concept|General Exam|3306,3313|true|false|false|C0392747|Changing|changes
Attribute|Clinical Attribute|General Exam|3321,3326|false|false|false|C5890168||Alert
Drug|Organic Chemical|General Exam|3321,3326|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|General Exam|3321,3326|false|false|false|C0718338|Alert brand of caffeine|Alert
Finding|Finding|General Exam|3321,3326|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|General Exam|3321,3326|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|General Exam|3321,3326|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Anatomy|Body Part, Organ, or Organ Component|General Exam|3355,3370|false|false|false|C0278454|All extremities|all extremities
Anatomy|Body Part, Organ, or Organ Component|General Exam|3359,3370|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Finding|Body Substance|General Exam|3375,3384|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|General Exam|3375,3384|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|General Exam|3375,3384|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|General Exam|3375,3384|false|false|false|C0030685|Patient Discharge|discharge
Attribute|Clinical Attribute|General Exam|3401,3407|false|false|false|C0944911||Weight
Finding|Finding|General Exam|3401,3407|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|Weight
Finding|Sign or Symptom|General Exam|3401,3407|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|Weight
Procedure|Health Care Activity|General Exam|3401,3407|false|false|false|C1305866|Weighing patient|Weight
Finding|Classification|General Exam|3506,3509|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Finding|Gene or Genome|General Exam|3506,3509|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Finding|Finding|General Exam|3511,3516|false|false|false|C0234422|Awake (finding)|awake
Attribute|Clinical Attribute|General Exam|3518,3523|false|false|false|C5890168||alert
Drug|Organic Chemical|General Exam|3518,3523|false|false|false|C0718338|Alert brand of caffeine|alert
Drug|Pharmacologic Substance|General Exam|3518,3523|false|false|false|C0718338|Alert brand of caffeine|alert
Finding|Finding|General Exam|3518,3523|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Functional Concept|General Exam|3518,3523|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Intellectual Product|General Exam|3518,3523|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Finding|General Exam|3525,3533|false|false|false|C1961028|Oriented to place|oriented
Finding|Idea or Concept|General Exam|3537,3541|false|false|false|C0036588;C1551994|Self;subscriber - self|self
Finding|Intellectual Product|General Exam|3537,3541|false|false|false|C0036588;C1551994|Self;subscriber - self|self
Finding|Idea or Concept|General Exam|3549,3557|false|false|false|C1547192|Organization unit type - Hospital|hospital
Anatomy|Body Location or Region|General Exam|3558,3563|false|false|false|C1512338|HEENT|HEENT
Finding|Finding|General Exam|3571,3577|false|false|false|C2143306|PERRLA|PERRLA
Anatomy|Body Location or Region|General Exam|3579,3583|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|General Exam|3579,3583|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|General Exam|3579,3583|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Finding|Finding|General Exam|3588,3591|true|false|false|C0425687|Jugular venous engorgement|JVD
Finding|Finding|General Exam|3609,3618|false|false|false|C0332218|Difficult (qualifier value)|difficult
Anatomy|Body Part, Organ, or Organ Component|General Exam|3633,3638|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|General Exam|3633,3638|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|General Exam|3633,3638|false|false|false|C0795691|HEART PROBLEM|heart
Attribute|Clinical Attribute|General Exam|3633,3645|false|false|false|C4050434||heart sounds
Finding|Organ or Tissue Function|General Exam|3633,3645|false|false|false|C0018820|Heart Sounds|heart sounds
Procedure|Diagnostic Procedure|General Exam|3633,3645|false|false|false|C2230284|auscultation of heart sounds|heart sounds
Phenomenon|Natural Phenomenon or Process|General Exam|3639,3645|false|false|false|C0037709||sounds
Anatomy|Body Part, Organ, or Organ Component|General Exam|3647,3652|false|false|false|C0024109|Lung|LUNGS
Finding|Finding|General Exam|3665,3673|false|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Anatomy|Body Location or Region|General Exam|3674,3677|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|ABD
Disorder|Cell or Molecular Dysfunction|General Exam|3674,3677|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|ABD
Disorder|Disease or Syndrome|General Exam|3679,3683|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Disorder|Congenital Abnormality|General Exam|3711,3714|false|false|false|C0015306|Hereditary Multiple Exostoses|EXT
Finding|Gene or Genome|General Exam|3711,3714|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|EXT
Finding|Conceptual Entity|General Exam|3723,3729|false|false|false|C0442038;C0920847|Circumpennate;Radial|radial
Drug|Food|General Exam|3730,3736|false|false|false|C5890763||pulses
Finding|Physiologic Function|General Exam|3730,3736|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|General Exam|3730,3736|false|false|false|C0034107|Pulse taking|pulses
Anatomy|Body Part, Organ, or Organ Component|General Exam|3738,3743|false|false|false|C4048756|Right arm|R arm
Anatomy|Body Part, Organ, or Organ Component|General Exam|3740,3743|false|false|false|C0446516;C1140618;C1269078|Upper Extremity;Upper arm|arm
Disorder|Anatomical Abnormality|General Exam|3740,3743|false|false|false|C3495676|Anorectal Malformations|arm
Finding|Gene or Genome|General Exam|3740,3743|false|false|false|C1824218;C3715044|AKR1A1 wt Allele;ARMC9 gene|arm
Procedure|Diagnostic Procedure|General Exam|3740,3743|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Research Activity|General Exam|3740,3743|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Therapeutic or Preventive Procedure|General Exam|3740,3743|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Finding|Functional Concept|General Exam|3752,3757|false|false|false|C1513492|motor movement|motor
Finding|Organ or Tissue Function|General Exam|3758,3774|false|true|false|C0036658|Sensory perception|sensory function
Finding|Finding|General Exam|3766,3774|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|General Exam|3766,3774|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|General Exam|3766,3774|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|General Exam|3766,3774|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Finding|General Exam|3776,3782|false|false|false|C1554187|Gender Status - Intact|intact
Finding|Functional Concept|General Exam|3830,3835|false|false|false|C1883002|Sequence Chromatogram|trace
Attribute|Clinical Attribute|General Exam|3837,3842|false|false|false|C1717255||edema
Finding|Pathologic Function|General Exam|3837,3842|false|false|false|C0013604|Edema|edema
Disorder|Disease or Syndrome|General Exam|3865,3869|false|false|false|C0009443;C0024117|Chronic Obstructive Airway Disease;Common Cold|cold
Drug|Organic Chemical|General Exam|3865,3869|false|false|false|C0719425|Cold brand of chlorpheniramine-phenylpropanolamine|cold
Drug|Pharmacologic Substance|General Exam|3865,3869|false|false|false|C0719425|Cold brand of chlorpheniramine-phenylpropanolamine|cold
Finding|Organism Function|General Exam|3865,3869|false|false|false|C0234192|Cold Sensation|cold
Phenomenon|Natural Phenomenon or Process|General Exam|3865,3869|false|false|false|C0009264|Cold Temperature|cold
Procedure|Therapeutic or Preventive Procedure|General Exam|3865,3869|false|false|false|C0010412|Cold Therapy|cold
Finding|Finding|General Exam|3881,3890|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|General Exam|3881,3890|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|General Exam|3881,3890|false|false|false|C2229507|sensory exam|sensation
Finding|Functional Concept|General Exam|3900,3905|false|false|false|C1513492|motor movement|motor
Finding|Idea or Concept|General Exam|3906,3914|false|false|false|C0808080|Strength (attribute)|strength
Finding|Finding|General Exam|3919,3922|false|false|false|C0948106;C1419600|ROM1 gene;Rupture of Membranes|ROM
Finding|Gene or Genome|General Exam|3919,3922|false|false|false|C0948106;C1419600|ROM1 gene;Rupture of Membranes|ROM
Procedure|Laboratory Procedure|General Exam|3919,3922|false|false|false|C1562926|Range of motion technique (procedure)|ROM
Anatomy|Body System|General Exam|3923,3927|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|General Exam|3923,3927|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|General Exam|3923,3927|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Finding|Body Substance|General Exam|3923,3927|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|General Exam|3923,3927|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Sign or Symptom|General Exam|3932,3938|true|false|false|C0015230;C5779628|Exanthema;Skin rash|rashes
Finding|Intellectual Product|General Exam|3942,3949|true|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|General Exam|3942,3949|true|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Finding|Pathologic Function|General Exam|3950,3959|false|false|false|C0013604|Edema|edematous
Finding|Functional Concept|General Exam|3960,3967|true|false|false|C0392747|Changing|changes
Attribute|Clinical Attribute|General Exam|3975,3980|false|false|false|C5890168||Alert
Drug|Organic Chemical|General Exam|3975,3980|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|General Exam|3975,3980|false|false|false|C0718338|Alert brand of caffeine|Alert
Finding|Finding|General Exam|3975,3980|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|General Exam|3975,3980|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|General Exam|3975,3980|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Anatomy|Body Part, Organ, or Organ Component|General Exam|4009,4024|false|false|false|C0278454|All extremities|all extremities
Anatomy|Body Part, Organ, or Organ Component|General Exam|4013,4024|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Lab|Laboratory or Test Result|General Exam|4047,4051|false|false|false|C0587081|Laboratory test finding|Labs
Procedure|Health Care Activity|General Exam|4055,4064|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Anatomy|Cell|General Exam|4100,4103|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|4110,4113|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|4110,4113|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|4110,4113|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|4120,4123|false|false|false|C0019046|Hemoglobin|HGB
Drug|Biologically Active Substance|General Exam|4120,4123|false|false|false|C0019046|Hemoglobin|HGB
Finding|Gene or Genome|General Exam|4120,4123|false|false|false|C1424337|CYGB gene|HGB
Lab|Laboratory or Test Result|General Exam|4120,4123|false|false|false|C0019029|Hemoglobin concentration|HGB
Procedure|Laboratory Procedure|General Exam|4129,4132|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Procedure|Therapeutic or Preventive Procedure|General Exam|4129,4132|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Disorder|Virus|General Exam|4138,4141|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|General Exam|4138,4141|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|4138,4141|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|4138,4141|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|4146,4149|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|4146,4149|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|General Exam|4146,4149|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|4146,4149|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|4146,4149|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|General Exam|4155,4159|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|4199,4202|false|false|false|C0201617|Primed lymphocyte test|PLT
Drug|Amino Acid, Peptide, or Protein|General Exam|4203,4206|false|false|false|C5441956|Megakaryocyte-Potentiating Factor, human|SMR
Drug|Immunologic Factor|General Exam|4203,4206|false|false|false|C5441956|Megakaryocyte-Potentiating Factor, human|SMR
Finding|Gene or Genome|General Exam|4203,4206|false|false|false|C1334533;C1704868|MSLN gene;MSLN wt Allele|SMR
Procedure|Laboratory Procedure|General Exam|4214,4217|false|false|false|C0201617|Primed lymphocyte test|PLT
Finding|Body Substance|General Exam|4262,4268|false|false|false|C0024202|Lymph|LYMPHS
Drug|Antibiotic|General Exam|4272,4277|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Biomedical or Dental Material|General Exam|4272,4277|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Organic Chemical|General Exam|4272,4277|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Disorder|Disease or Syndrome|General Exam|4280,4283|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|EOS
Finding|Gene or Genome|General Exam|4280,4283|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|EOS
Disorder|Neoplastic Process|General Exam|4397,4400|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Procedure|Laboratory Procedure|General Exam|4397,4400|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Drug|Biologically Active Substance|General Exam|4425,4432|false|false|false|C0017725|glucose|GLUCOSE
Drug|Organic Chemical|General Exam|4425,4432|false|false|false|C0017725|glucose|GLUCOSE
Drug|Pharmacologic Substance|General Exam|4425,4432|false|false|false|C0017725|glucose|GLUCOSE
Lab|Laboratory or Test Result|General Exam|4425,4432|false|false|false|C5781949|Glucose^1.5H post dose glucagon|GLUCOSE
Procedure|Laboratory Procedure|General Exam|4425,4432|false|false|false|C0337438|Glucose measurement|GLUCOSE
Drug|Biologically Active Substance|General Exam|4438,4442|false|false|false|C0041942|urea|UREA
Drug|Organic Chemical|General Exam|4438,4442|false|false|false|C0041942|urea|UREA
Drug|Pharmacologic Substance|General Exam|4438,4442|false|false|false|C0041942|urea|UREA
Procedure|Laboratory Procedure|General Exam|4438,4442|false|false|false|C0523961|Urea measurement|UREA
Drug|Biologically Active Substance|General Exam|4461,4467|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Element, Ion, or Isotope|General Exam|4461,4467|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Pharmacologic Substance|General Exam|4461,4467|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Finding|Physiologic Function|General Exam|4461,4467|false|false|false|C4553025|Sodium metabolic function|SODIUM
Procedure|Laboratory Procedure|General Exam|4461,4467|false|false|false|C0337443|Sodium measurement|SODIUM
Drug|Biologically Active Substance|General Exam|4473,4482|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Element, Ion, or Isotope|General Exam|4473,4482|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Food|General Exam|4473,4482|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Inorganic Chemical|General Exam|4473,4482|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Pharmacologic Substance|General Exam|4473,4482|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Finding|Physiologic Function|General Exam|4473,4482|false|false|false|C4553027|Potassium metabolic function|POTASSIUM
Procedure|Laboratory Procedure|General Exam|4473,4482|false|false|false|C0202194|Potassium measurement|POTASSIUM
Drug|Element, Ion, or Isotope|General Exam|4487,4495|false|false|false|C0008203;C0596019|Chlorides;chloride ion|CHLORIDE
Finding|Physiologic Function|General Exam|4487,4495|false|false|false|C4553021|Chloride metabolic function|CHLORIDE
Procedure|Laboratory Procedure|General Exam|4487,4495|false|false|false|C0201952|Chloride measurement|CHLORIDE
Drug|Biologically Active Substance|General Exam|4505,4508|false|false|false|C0007012|carbon dioxide|CO2
Drug|Inorganic Chemical|General Exam|4505,4508|false|false|false|C0007012|carbon dioxide|CO2
Finding|Finding|General Exam|4505,4508|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Finding|Gene or Genome|General Exam|4505,4508|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Drug|Element, Ion, or Isotope|General Exam|4513,4518|false|false|false|C0003075|Anions|ANION
Drug|Amino Acid, Peptide, or Protein|General Exam|4520,4523|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Drug|Biologically Active Substance|General Exam|4520,4523|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Finding|Gene or Genome|General Exam|4520,4523|false|false|false|C1419277;C2984552|RASA1 gene;RASA1 wt Allele|GAP
Drug|Biologically Active Substance|General Exam|4542,4549|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Element, Ion, or Isotope|General Exam|4542,4549|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Inorganic Chemical|General Exam|4542,4549|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Pharmacologic Substance|General Exam|4542,4549|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Vitamin|General Exam|4542,4549|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Finding|Physiologic Function|General Exam|4542,4549|false|false|false|C4553026|Calcium metabolic function|CALCIUM
Procedure|Laboratory Procedure|General Exam|4542,4549|false|false|false|C0201925|Calcium measurement|CALCIUM
Drug|Element, Ion, or Isotope|General Exam|4555,4564|false|false|false|C0031603;C1601799|Phosphates;phosphate ion|PHOSPHATE
Drug|Inorganic Chemical|General Exam|4555,4564|false|false|false|C0031603;C1601799|Phosphates;phosphate ion|PHOSPHATE
Drug|Pharmacologic Substance|General Exam|4555,4564|false|false|false|C0031603;C1601799|Phosphates;phosphate ion|PHOSPHATE
Procedure|Laboratory Procedure|General Exam|4555,4564|false|false|false|C0523826|Phosphate measurement|PHOSPHATE
Drug|Biologically Active Substance|General Exam|4569,4578|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Drug|Element, Ion, or Isotope|General Exam|4569,4578|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Drug|Inorganic Chemical|General Exam|4569,4578|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Drug|Pharmacologic Substance|General Exam|4569,4578|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Procedure|Laboratory Procedure|General Exam|4569,4578|false|false|false|C0373675|Magnesium measurement|MAGNESIUM
Drug|Amino Acid, Peptide, or Protein|General Exam|4611,4616|false|false|false|C0019018|Glycosylated hemoglobin A|HbA1c
Drug|Biologically Active Substance|General Exam|4611,4616|false|false|false|C0019018|Glycosylated hemoglobin A|HbA1c
Procedure|Laboratory Procedure|General Exam|4611,4616|false|false|false|C0202054|Glucohemoglobin measurement|HbA1c
Finding|Gene or Genome|General Exam|4621,4624|false|false|false|C1416571|KCNH1 gene|eAG
Drug|Amino Acid, Peptide, or Protein|General Exam|4643,4648|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|General Exam|4643,4648|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|General Exam|4643,4648|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|General Exam|4643,4648|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Drug|Amino Acid, Peptide, or Protein|General Exam|4694,4697|false|false|false|C0023821|High Density Lipoproteins|HDL
Drug|Biologically Active Substance|General Exam|4694,4697|false|false|false|C0023821|High Density Lipoproteins|HDL
Finding|Gene or Genome|General Exam|4694,4697|false|false|false|C3715113|HSD11B1 wt Allele|HDL
Procedure|Laboratory Procedure|General Exam|4694,4697|false|false|false|C0392885|High density lipoprotein measurement|HDL
Drug|Amino Acid, Peptide, or Protein|General Exam|4711,4714|false|false|false|C0023821|High Density Lipoproteins|HDL
Drug|Biologically Active Substance|General Exam|4711,4714|false|false|false|C0023821|High Density Lipoproteins|HDL
Finding|Gene or Genome|General Exam|4711,4714|false|false|false|C3715113|HSD11B1 wt Allele|HDL
Procedure|Laboratory Procedure|General Exam|4711,4714|false|false|false|C0392885|High density lipoprotein measurement|HDL
Drug|Biologically Active Substance|General Exam|4720,4723|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Drug|Organic Chemical|General Exam|4720,4723|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Procedure|Laboratory Procedure|General Exam|4720,4723|false|false|false|C0202117|Low density lipoprotein cholesterol measurement|LDL
Anatomy|Body Part, Organ, or Organ Component|General Exam|4724,4728|false|false|false|C4084820|Intracalcarine cortex|CALC
Finding|Gene or Genome|General Exam|4724,4728|false|false|false|C1413147|MICU1 gene|CALC
Lab|Laboratory or Test Result|General Exam|4852,4856|false|false|false|C0587081|Laboratory test finding|Labs
Finding|Body Substance|General Exam|4860,4869|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|General Exam|4860,4869|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|General Exam|4860,4869|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|General Exam|4860,4869|false|false|false|C0030685|Patient Discharge|Discharge
Disorder|Disease or Syndrome|General Exam|4903,4908|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4903,4908|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|4909,4912|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|4919,4922|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|4919,4922|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|4919,4922|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|4929,4932|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|4929,4932|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|4929,4932|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|4929,4932|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|4939,4942|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|4939,4942|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|4950,4953|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|General Exam|4950,4953|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|4950,4953|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|4950,4953|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|4957,4960|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|4957,4960|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|General Exam|4957,4960|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|4957,4960|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|4957,4960|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|General Exam|4966,4970|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|4997,5000|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|5017,5022|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|5017,5022|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Finding|Body Substance|General Exam|5041,5047|false|false|false|C0024202|Lymph|Lymphs
Drug|Antibiotic|General Exam|5052,5057|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|General Exam|5052,5057|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|General Exam|5052,5057|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|General Exam|5061,5064|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|Eos
Finding|Gene or Genome|General Exam|5061,5064|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|Eos
Disorder|Disease or Syndrome|General Exam|5175,5180|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|5175,5180|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|5185,5188|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Procedure|Laboratory Procedure|General Exam|5185,5188|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|General Exam|5210,5215|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|5210,5215|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|5210,5223|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|5210,5223|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|5210,5223|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|5216,5223|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|5216,5223|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|5216,5223|false|false|false|C0017725|glucose|Glucose
Lab|Laboratory or Test Result|General Exam|5216,5223|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|5216,5223|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|General Exam|5270,5274|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|5270,5274|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|General Exam|5270,5274|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|General Exam|5299,5304|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|5299,5304|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|5305,5308|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|General Exam|5305,5308|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|General Exam|5305,5308|false|false|false|C0001899|Alanine Transaminase|ALT
Finding|Gene or Genome|General Exam|5305,5308|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|General Exam|5305,5308|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|General Exam|5305,5308|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|General Exam|5305,5308|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|General Exam|5312,5315|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|General Exam|5312,5315|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|5312,5315|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|General Exam|5312,5315|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|General Exam|5312,5315|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Finding|Gene or Genome|General Exam|5312,5315|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|5322,5325|false|false|false|C0022917|Lactate Dehydrogenase|LDH
Drug|Enzyme|General Exam|5322,5325|false|false|false|C0022917|Lactate Dehydrogenase|LDH
Finding|Finding|General Exam|5322,5325|false|false|false|C0851148|Lifetime Drinking History|LDH
Procedure|Laboratory Procedure|General Exam|5322,5325|false|false|false|C0202113|Lactate dehydrogenase measurement|LDH
Drug|Amino Acid, Peptide, or Protein|General Exam|5332,5339|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|General Exam|5332,5339|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Disorder|Disease or Syndrome|General Exam|5368,5373|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|5368,5373|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|5368,5381|false|false|false|C0853248|Blood albumin|BLOOD Albumin
Drug|Amino Acid, Peptide, or Protein|General Exam|5374,5381|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Biologically Active Substance|General Exam|5374,5381|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Pharmacologic Substance|General Exam|5374,5381|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Finding|Gene or Genome|General Exam|5374,5381|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Finding|Physiologic Function|General Exam|5374,5381|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Procedure|Laboratory Procedure|General Exam|5374,5381|false|false|false|C0201838|Albumin measurement|Albumin
Drug|Biologically Active Substance|General Exam|5387,5394|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|General Exam|5387,5394|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|General Exam|5387,5394|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|General Exam|5387,5394|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|General Exam|5387,5394|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Finding|Physiologic Function|General Exam|5387,5394|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|General Exam|5387,5394|false|false|false|C0201925|Calcium measurement|Calcium
Finding|Finding|General Exam|5425,5432|false|false|false|C0740845|Imaging problem|Imaging
Procedure|Diagnostic Procedure|General Exam|5425,5432|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|Imaging
Procedure|Diagnostic Procedure|General Exam|5452,5455|false|false|false|C0430462|Transthoracic echocardiography|TTE
Finding|Functional Concept|General Exam|5465,5469|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|General Exam|5465,5476|false|false|false|C0225860|Left atrial structure|left atrium
Anatomy|Body Part, Organ, or Organ Component|General Exam|5470,5476|false|false|false|C0018792|Heart Atrium|atrium
Finding|Functional Concept|General Exam|5510,5515|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|General Exam|5516,5522|false|false|false|C0018792|Heart Atrium|atrial
Finding|Finding|General Exam|5524,5532|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|General Exam|5524,5532|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|General Exam|5524,5532|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|General Exam|5524,5532|false|false|false|C0033095||pressure
Finding|Functional Concept|General Exam|5546,5550|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|General Exam|5546,5567|false|false|false|C0504053|Wall of left ventricle|Left ventricular wall
Anatomy|Body Part, Organ, or Organ Component|General Exam|5551,5562|false|false|false|C0018827|Heart Ventricle|ventricular
Anatomy|Body Part, Organ, or Organ Component|General Exam|5551,5567|false|false|false|C0507618|Wall of ventricle|ventricular wall
Anatomy|Body Space or Junction|General Exam|5585,5591|false|false|false|C0333343|Body cavities|cavity
Disorder|Anatomical Abnormality|General Exam|5585,5591|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Disorder|Disease or Syndrome|General Exam|5585,5591|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Finding|Intellectual Product|General Exam|5609,5616|false|false|false|C0282416|Overall Publication Type|Overall
Finding|Functional Concept|General Exam|5617,5621|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|General Exam|5622,5633|false|false|false|C0018827|Heart Ventricle|ventricular
Finding|Organ or Tissue Function|General Exam|5634,5642|false|false|false|C0039155|Systole|systolic
Finding|Finding|General Exam|5644,5652|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|General Exam|5644,5652|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|General Exam|5644,5652|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|General Exam|5644,5652|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Finding|General Exam|5656,5666|false|false|false|C4085643;C5201148;C5962468|Moderate;Moderate Effect;Moderate Response|moderately
Disorder|Mental or Behavioral Dysfunction|General Exam|5667,5676|false|false|false|C0344315|Depressed mood|depressed
Attribute|Clinical Attribute|General Exam|5678,5682|false|false|false|C0428772|Left ventricular ejection fraction|LVEF
Procedure|Diagnostic Procedure|General Exam|5678,5682|false|false|false|C3837267|LVEF (procedure)|LVEF
Event|Activity|General Exam|5695,5705|false|false|false|C1516048|Assessed|assessment
Finding|Intellectual Product|General Exam|5695,5705|false|false|false|C0679207|Knowledge acquisition using a method of assessment|assessment
Procedure|Diagnostic Procedure|General Exam|5695,5705|false|false|false|C0028708;C0031809;C0220825;C0542573;C0549068;C0549070;C0549071;C0549072;C0549073;C0549074;C0549075;C0549076;C0549078;C0549079;C0549080;C1161151;C1261322;C2237115|Evaluation;Evaluation procedure;Nutrition Assessment;Personal care assessment;Physical Examination;assessment of cognitive functions|assessment
Procedure|Health Care Activity|General Exam|5695,5705|false|false|false|C0028708;C0031809;C0220825;C0542573;C0549068;C0549070;C0549071;C0549072;C0549073;C0549074;C0549075;C0549076;C0549078;C0549079;C0549080;C1161151;C1261322;C2237115|Evaluation;Evaluation procedure;Nutrition Assessment;Personal care assessment;Physical Examination;assessment of cognitive functions|assessment
Finding|Finding|General Exam|5718,5734|false|false|false|C2828075|Suboptimal Image Reason|suboptimal image
Disorder|Disease or Syndrome|General Exam|5729,5734|false|false|false|C1846009|Intrauterine growth restriction, metaphyseal dysplasia, adrenal hypoplasia congenita, and genital anomaly syndrome|image
Finding|Intellectual Product|General Exam|5729,5734|false|false|false|C1696103;C1704254;C1704922;C3542466|Image;Image (foundation metadata concept);Medical Image;image - dosage form|image
Finding|Idea or Concept|General Exam|5747,5758|false|false|false|C0750502|Significant|significant
Finding|Conceptual Entity|General Exam|5773,5784|false|false|false|C2827666|Variability|variability
Finding|Finding|General Exam|5796,5807|false|false|false|C0086439|Hypokinesia|hypokinesis
Anatomy|Cell Component|General Exam|5843,5847|false|false|false|C3890171|dinoflagellate apex|apex
Drug|Amino Acid, Peptide, or Protein|General Exam|5843,5847|false|false|false|C0140145|APEX1 protein, human|apex
Drug|Enzyme|General Exam|5843,5847|false|false|false|C0140145|APEX1 protein, human|apex
Finding|Gene or Genome|General Exam|5843,5847|false|false|false|C1332102|APEX1 gene|apex
Anatomy|Body Part, Organ, or Organ Component|General Exam|5861,5872|false|false|false|C0018827|Heart Ventricle|ventricular
Disorder|Congenital Abnormality|General Exam|5861,5886|true|false|false|C0018818|Ventricular Septal Defects|ventricular septal defect
Disorder|Anatomical Abnormality|General Exam|5873,5886|true|false|false|C0018816;C5779791|Congenital septal defect of heart;Heart Septal Defects|septal defect
Disorder|Congenital Abnormality|General Exam|5873,5886|true|false|false|C0018816;C5779791|Congenital septal defect of heart;Heart Septal Defects|septal defect
Disorder|Disease or Syndrome|General Exam|5880,5886|true|false|false|C1861101|THYROID HORMONE PLASMA MEMBRANE TRANSPORT DEFECT|defect
Finding|Functional Concept|General Exam|5880,5886|true|false|false|C1457869|Defect|defect
Finding|Functional Concept|General Exam|5888,5893|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Anatomy|Body Part, Organ, or Organ Component|General Exam|5895,5906|false|false|false|C0018827|Heart Ventricle|ventricular
Anatomy|Body Part, Organ, or Organ Component|General Exam|5907,5914|false|false|false|C0935616|chamber [body part]|chamber
Finding|Functional Concept|General Exam|5924,5928|false|false|false|C0332296|Free of (attribute)|free
Attribute|Clinical Attribute|General Exam|5929,5940|false|false|false|C1980023|Wall motion|wall motion
Phenomenon|Natural Phenomenon or Process|General Exam|5934,5940|false|false|false|C0026597|Motion|motion
Finding|Functional Concept|General Exam|5958,5967|false|false|false|C1547175;C1962987|Ascend (action);Sequencing - Ascending|ascending
Anatomy|Body Part, Organ, or Organ Component|General Exam|5958,5973|false|false|false|C0003956|Ascending aorta structure|ascending aorta
Anatomy|Body Part, Organ, or Organ Component|General Exam|5968,5973|false|false|false|C0003483;C4037978|Aorta;Chest+Abdomen>Aorta|aorta
Procedure|Health Care Activity|General Exam|5968,5973|false|false|false|C0869784|Procedure on aorta|aorta
Finding|Idea or Concept|General Exam|5997,6003|false|false|false|C1554106|MDF AttributeType - Number|number
Anatomy|Body Part, Organ, or Organ Component|General Exam|6007,6013|false|false|false|C0003483|Aorta|aortic
Anatomy|Body Part, Organ, or Organ Component|General Exam|6007,6019|false|false|false|C0003501;C4533215|Aortic valve structure;Chest>Aortic valve|aortic valve
Anatomy|Body Part, Organ, or Organ Component|General Exam|6014,6019|false|false|false|C1186983|Anatomical valve|valve
Finding|Intellectual Product|General Exam|6061,6065|false|false|false|C1547225|Mild Severity of Illness Code|mild
Anatomy|Body Part, Organ, or Organ Component|General Exam|6066,6072|false|false|false|C0003483|Aorta|aortic
Anatomy|Body Part, Organ, or Organ Component|General Exam|6066,6078|false|false|false|C0003501;C4533215|Aortic valve structure;Chest>Aortic valve|aortic valve
Anatomy|Body Part, Organ, or Organ Component|General Exam|6073,6078|false|false|false|C1186983|Anatomical valve|valve
Finding|Pathologic Function|General Exam|6080,6088|false|false|false|C1261287|Stenosis|stenosis
Anatomy|Body Part, Organ, or Organ Component|General Exam|6090,6095|false|false|false|C1186983|Anatomical valve|valve
Finding|Finding|General Exam|6090,6100|false|false|false|C4687749|Valve Area|valve area
Event|Governmental or Regulatory Activity|General Exam|6096,6100|false|false|false|C1510751|Academic Research Enhancement Awards|area
Disorder|Congenital Abnormality|General Exam|6108,6111|false|false|false|C0555206|Chiari malformation type II|cm2
Anatomy|Body Part, Organ, or Organ Component|General Exam|6117,6123|false|false|false|C0003483|Aorta|aortic
Disorder|Disease or Syndrome|General Exam|6117,6137|true|false|false|C0003504|Aortic Valve Insufficiency|aortic regurgitation
Finding|Finding|General Exam|6124,6137|true|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|General Exam|6124,6137|true|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|General Exam|6124,6137|true|false|false|C0460152|Regurgitation - mechanism|regurgitation
Anatomy|Body Part, Organ, or Organ Component|General Exam|6152,6164|false|false|false|C0026264|Mitral Valve|mitral valve
Anatomy|Body Part, Organ, or Organ Component|General Exam|6159,6164|false|false|false|C1186983|Anatomical valve|valve
Disorder|Disease or Syndrome|General Exam|6207,6227|false|false|false|C0026266|Mitral Valve Insufficiency|mitral regurgitation
Finding|Finding|General Exam|6214,6227|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|General Exam|6214,6227|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|General Exam|6214,6227|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Anatomy|Body Part, Organ, or Organ Component|General Exam|6233,6242|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|General Exam|6233,6242|false|false|false|C2707265||pulmonary
Finding|Finding|General Exam|6233,6242|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Anatomy|Body Part, Organ, or Organ Component|General Exam|6233,6249|false|false|false|C0034052|Pulmonary artery structure|pulmonary artery
Finding|Finding|General Exam|6233,6267|false|false|false|C0428643|Pulmonary artery systolic pressure|pulmonary artery systolic pressure
Anatomy|Body Part, Organ, or Organ Component|General Exam|6243,6249|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|General Exam|6243,6249|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Finding|Organ or Tissue Function|General Exam|6250,6258|false|false|false|C0039155|Systole|systolic
Attribute|Clinical Attribute|General Exam|6250,6267|false|false|false|C0871470|Systolic Pressure|systolic pressure
Finding|Finding|General Exam|6259,6267|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|General Exam|6259,6267|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|General Exam|6259,6267|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|General Exam|6259,6267|false|false|false|C0033095||pressure
Finding|Functional Concept|General Exam|6313,6324|false|false|false|C0205463|Physiological|physiologic
Anatomy|Body Location or Region|General Exam|6326,6337|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Anatomy|Body Part, Organ, or Organ Component|General Exam|6326,6337|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Disorder|Disease or Syndrome|General Exam|6326,6346|false|false|false|C0031039|Pericardial effusion|pericardial effusion
Finding|Body Substance|General Exam|6326,6346|false|false|false|C1253937|Pericardial effusion body substance|pericardial effusion
Finding|Body Substance|General Exam|6338,6346|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|General Exam|6338,6346|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|General Exam|6338,6346|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|General Exam|6382,6387|false|false|false|C1705923|Study Object|study
Procedure|Research Activity|General Exam|6382,6387|false|false|false|C0008972;C0947630;C2603343|Clinical Research;Scientific Study;Study|study
Finding|Functional Concept|General Exam|6415,6419|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|General Exam|6420,6431|false|false|false|C0018827|Heart Ventricle|ventricular
Finding|Organ or Tissue Function|General Exam|6432,6440|false|false|false|C0039155|Systole|systolic
Finding|Finding|General Exam|6441,6449|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|General Exam|6441,6449|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|General Exam|6441,6449|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|General Exam|6441,6449|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Finding|General Exam|6453,6461|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|probably
Finding|Idea or Concept|General Exam|6453,6461|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|probably
Finding|Finding|General Exam|6481,6497|false|false|false|C2828075|Suboptimal Image Reason|suboptimal image
Disorder|Disease or Syndrome|General Exam|6492,6497|false|false|false|C1846009|Intrauterine growth restriction, metaphyseal dysplasia, adrenal hypoplasia congenita, and genital anomaly syndrome|image
Finding|Intellectual Product|General Exam|6492,6497|false|false|false|C1696103;C1704254;C1704922;C3542466|Image;Image (foundation metadata concept);Medical Image;image - dosage form|image
Procedure|Research Activity|General Exam|6514,6521|false|false|false|C0947630|Scientific Study|studies
Event|Activity|General Exam|6542,6552|false|false|false|C1707455|Comparison|comparison
Procedure|Diagnostic Procedure|General Exam|6561,6564|false|false|false|C0039985|Plain chest X-ray|CXR
Finding|Conceptual Entity|Impression|6596,6607|false|false|false|C2986411|Improvement|improvement
Anatomy|Body Part, Organ, or Organ Component|Impression|6611,6621|false|false|false|C0225754|Bilateral lungs|both lungs
Anatomy|Body Part, Organ, or Organ Component|Impression|6616,6621|false|false|false|C0024109|Lung|lungs
Finding|Finding|Impression|6625,6633|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|probably
Finding|Idea or Concept|Impression|6625,6633|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|probably
Finding|Finding|Impression|6642,6650|false|false|false|C0392756|Reduced|decrease
Anatomy|Body Part, Organ, or Organ Component|Impression|6654,6663|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Impression|6654,6663|false|false|false|C2707265||pulmonary
Finding|Finding|Impression|6654,6663|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Attribute|Clinical Attribute|Impression|6665,6670|false|false|false|C1717255||edema
Finding|Pathologic Function|Impression|6665,6670|false|false|false|C0013604|Edema|edema
Finding|Intellectual Product|Impression|6676,6680|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Finding|Impression|6686,6694|false|false|false|C0392756|Reduced|decrease
Finding|Finding|Impression|6707,6715|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|Impression|6707,6715|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Functional Concept|Impression|6716,6721|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Tissue|Impression|6722,6729|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|Impression|6722,6729|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Body Substance|Impression|6731,6739|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|Impression|6731,6739|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|Impression|6731,6739|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Disorder|Disease or Syndrome|Impression|6752,6757|false|false|false|C1410088|Still|still
Disorder|Disease or Syndrome|Impression|6770,6783|false|false|false|C0521530|Lung consolidation|consolidation
Finding|Functional Concept|Impression|6791,6796|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|Impression|6791,6807|false|false|false|C1261074|Structure of right upper lobe of lung|right upper lobe
Anatomy|Body Part, Organ, or Organ Component|Impression|6797,6807|false|false|false|C0225756|Structure of upper lobe of lung|upper lobe
Anatomy|Body Part, Organ, or Organ Component|Impression|6803,6807|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|Impression|6803,6807|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Finding|Finding|Impression|6809,6817|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|probably
Finding|Idea or Concept|Impression|6809,6817|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|probably
Disorder|Disease or Syndrome|Impression|6819,6828|false|false|false|C0032285|Pneumonia|pneumonia
Anatomy|Body Location or Region|Impression|6847,6852|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|Impression|6847,6852|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|Impression|6847,6857|false|false|false|C0225758|Structure of lower lobe of lung|lower lobe
Anatomy|Body Part, Organ, or Organ Component|Impression|6853,6857|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|Impression|6853,6857|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Anatomy|Body Part, Organ, or Organ Component|Impression|6886,6891|false|false|false|C0018787;C4037974|Chest>Heart;Heart|Heart
Disorder|Neoplastic Process|Impression|6886,6891|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|Heart
Finding|Sign or Symptom|Impression|6886,6891|false|false|false|C0795691|HEART PROBLEM|Heart
Finding|Finding|Impression|6886,6896|false|false|false|C0744689|heart size|Heart size
Disorder|Disease or Syndrome|Impression|6914,6926|true|false|false|C0032326|Pneumothorax|pneumothorax
Finding|Conceptual Entity|Impression|6930,6935|false|false|false|C3811161;C4049106|Micro (prefix);Microbiology - Laboratory Class|MICRO
Finding|Intellectual Product|Impression|6930,6935|false|false|false|C3811161;C4049106|Micro (prefix);Microbiology - Laboratory Class|MICRO
Procedure|Laboratory Procedure|Impression|6930,6935|false|false|false|C0085672|Microbiology procedure|MICRO
Finding|Idea or Concept|Impression|6945,6950|false|false|false|C1546485|Diagnosis Type - Final|FINAL
Finding|Intellectual Product|Impression|6945,6957|false|false|false|C0460114|Final report|FINAL REPORT
Attribute|Clinical Attribute|Impression|6951,6957|false|false|false|C4255046||REPORT
Finding|Intellectual Product|Impression|6951,6957|false|false|false|C0684224|Report (document)|REPORT
Procedure|Health Care Activity|Impression|6951,6957|false|false|false|C0700287|Reporting|REPORT
Drug|Biologically Active Substance|Impression|6979,6982|false|false|false|C0012854|DNA|DNA
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Impression|6979,6982|false|false|false|C0012854|DNA|DNA
Finding|Genetic Function|Impression|6979,6996|false|false|false|C0683230|dna amplification|DNA amplification
Disorder|Cell or Molecular Dysfunction|Impression|6983,6996|false|false|false|C1705759|Gene Amplification Abnormality|amplification
Phenomenon|Phenomenon or Process|Impression|6983,6996|false|false|false|C1521871|Amplification|amplification
Procedure|Molecular Biology Research Technique|Impression|6983,6996|false|false|false|C1517480|Gene Amplification Technique|amplification
Procedure|Laboratory Procedure|Impression|6997,7002|false|false|false|C0005507;C1510438|Assay;Biological Assay|assay
Finding|Idea or Concept|Impression|7004,7009|false|false|false|C1546485|Diagnosis Type - Final|Final
Disorder|Cell or Molecular Dysfunction|Impression|7055,7063|false|false|false|C4727483|BRAF Gene Rearrangement|Positive
Finding|Classification|Impression|7055,7063|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|Positive
Finding|Finding|Impression|7055,7063|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|Positive
Finding|Finding|Impression|7055,7067|false|false|false|C1446409|Positive|Positive for
Finding|Intellectual Product|Impression|7068,7077|false|false|false|C0445332|Toxigenic|toxigenic
Drug|Biologically Active Substance|Impression|7110,7113|false|false|false|C0012854|DNA|DNA
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Impression|7110,7113|false|false|false|C0012854|DNA|DNA
Disorder|Cell or Molecular Dysfunction|Impression|7123,7136|false|false|false|C1705759|Gene Amplification Abnormality|amplification
Phenomenon|Phenomenon or Process|Impression|7123,7136|false|false|false|C1521871|Amplification|amplification
Procedure|Molecular Biology Research Technique|Impression|7123,7136|false|false|false|C1517480|Gene Amplification Technique|amplification
Finding|Conceptual Entity|Impression|7150,7159|false|false|false|C1514811;C1561577;C1706462;C3244318;C4266518|Bibliographic Reference;Reference - HL7UpdateMode;Reference - MdfHmdMetSourceType;Reference Object;Reference source|Reference
Finding|Idea or Concept|Impression|7150,7159|false|false|false|C1514811;C1561577;C1706462;C3244318;C4266518|Bibliographic Reference;Reference - HL7UpdateMode;Reference - MdfHmdMetSourceType;Reference Object;Reference source|Reference
Finding|Intellectual Product|Impression|7150,7159|false|false|false|C1514811;C1561577;C1706462;C3244318;C4266518|Bibliographic Reference;Reference - HL7UpdateMode;Reference - MdfHmdMetSourceType;Reference Object;Reference source|Reference
Finding|Intellectual Product|Impression|7160,7165|false|false|false|C3542016|Concept model range (foundation metadata concept)|Range
Finding|Classification|Impression|7166,7174|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|Negative
Finding|Finding|Impression|7166,7174|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|Negative
Lab|Laboratory or Test Result|Impression|7166,7174|false|false|false|C5237010|Expression Negative|Negative
Finding|Body Substance|Impression|7192,7198|false|false|false|C0038056;C1546789;C1576419|Specimen Type - Sputum;Sputum|SPUTUM
Finding|Intellectual Product|Impression|7192,7198|false|false|false|C0038056;C1546789;C1576419|Specimen Type - Sputum;Sputum|SPUTUM
Finding|Finding|Impression|7204,7210|false|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|Source
Finding|Functional Concept|Impression|7204,7210|false|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|Source
Finding|Intellectual Product|Impression|7204,7210|false|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|Source
Finding|Finding|Impression|7212,7224|false|false|false|C0566528|Does expectorate|Expectorated
Drug|Indicator, Reagent, or Diagnostic Aid|Impression|7231,7241|false|false|false|C0061856|Gram's stain|GRAM STAIN
Drug|Organic Chemical|Impression|7231,7241|false|false|false|C0061856|Gram's stain|GRAM STAIN
Procedure|Laboratory Procedure|Impression|7231,7241|false|false|false|C0200966|Bacterial stain, routine|GRAM STAIN
Drug|Indicator, Reagent, or Diagnostic Aid|Impression|7236,7241|false|false|false|C0038128|Stains|STAIN
Procedure|Laboratory Procedure|Impression|7236,7241|false|false|false|C0487602|Staining method|STAIN
Finding|Idea or Concept|Impression|7243,7248|false|false|false|C1546485|Diagnosis Type - Final|Final
Anatomy|Cell|Impression|7278,7294|false|false|false|C0014597|Epithelial Cells|epithelial cells
Anatomy|Cell|Impression|7289,7294|false|false|false|C0007634|Cells|cells
Finding|Conceptual Entity|Impression|7300,7305|false|false|false|C1521738;C2346620;C2349184|Field;Force Field;Knowledge Field|field
Procedure|Health Care Activity|Impression|7300,7305|false|false|false|C1553496|field - patient encounter|field
Finding|Conceptual Entity|Impression|7333,7338|true|false|false|C1521738;C2346620;C2349184|Field;Force Field;Knowledge Field|FIELD
Procedure|Health Care Activity|Impression|7333,7338|true|false|false|C1553496|field - patient encounter|FIELD
Finding|Classification|Impression|7348,7356|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|NEGATIVE
Finding|Finding|Impression|7348,7356|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|NEGATIVE
Lab|Laboratory or Test Result|Impression|7348,7356|false|false|false|C5237010|Expression Negative|NEGATIVE
Anatomy|Cell|Impression|7357,7360|false|false|false|C0206427|Rod Photoreceptors|ROD
Disorder|Disease or Syndrome|Impression|7357,7360|true|false|false|C0035086|Renal Osteodystrophy|ROD
Finding|Gene or Genome|Impression|7357,7360|true|false|false|C1424852|KNTC1 gene|ROD
Finding|Conceptual Entity|Impression|7391,7396|false|false|false|C1521738;C2346620;C2349184|Field;Force Field;Knowledge Field|FIELD
Procedure|Health Care Activity|Impression|7391,7396|false|false|false|C1553496|field - patient encounter|FIELD
Finding|Cell Function|Impression|7401,7408|false|false|false|C1155616|Cell budding|BUDDING
Drug|Food|Impression|7409,7414|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Drug|Immunologic Factor|Impression|7409,7414|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Drug|Indicator, Reagent, or Diagnostic Aid|Impression|7409,7414|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Drug|Pharmacologic Substance|Impression|7409,7414|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Drug|Substance|Impression|7434,7442|false|false|false|C0370003|Specimen|SPECIMEN
Finding|Body Substance|Impression|7434,7442|false|false|false|C1561495;C2347026|Biospecimen;Role Class - specimen|SPECIMEN
Finding|Functional Concept|Impression|7434,7442|false|false|false|C1561495;C2347026|Biospecimen;Role Class - specimen|SPECIMEN
Attribute|Clinical Attribute|Impression|7468,7479|false|false|false|C0231832|Respiratory rate|RESPIRATORY
Finding|Body Substance|Impression|7468,7479|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|RESPIRATORY
Finding|Functional Concept|Impression|7468,7479|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|RESPIRATORY
Finding|Intellectual Product|Impression|7468,7479|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|RESPIRATORY
Procedure|Laboratory Procedure|Impression|7468,7487|false|false|false|C4282127|Respiratory culture|RESPIRATORY CULTURE
Drug|Biomedical or Dental Material|Impression|7480,7487|false|false|false|C1706355|Culture Dose Form|CULTURE
Finding|Functional Concept|Impression|7480,7487|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|Impression|7480,7487|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|Impression|7480,7487|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Procedure|Laboratory Procedure|Impression|7518,7528|false|false|false|C5453732|Incubation|incubation
Procedure|Therapeutic or Preventive Procedure|Impression|7555,7563|false|false|false|C0392148|Providing presence (regime/therapy)|presence
Disorder|Anatomical Abnormality|Impression|7568,7575|false|false|false|C1689985|Absence (morphologic abnormality)|absence
Finding|Functional Concept|Impression|7568,7575|false|false|false|C0332197|Absent|absence
Finding|Functional Concept|Impression|7568,7578|false|false|false|C0332197|Absent|absence of
Finding|Functional Concept|Impression|7585,7594|false|false|false|C0231202|Symbiotic|commensal
Attribute|Clinical Attribute|Impression|7595,7606|false|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|Impression|7595,7606|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|Impression|7595,7606|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|Impression|7595,7606|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Disorder|Disease or Syndrome|Impression|7621,7631|false|false|false|C0519030|Pneumonia due to Klebsiella pneumoniae|KLEBSIELLA
Disorder|Disease or Syndrome|Impression|7621,7642|false|false|false|C2712605|Infection by Klebsiella pneumoniae in conditions classified elsewhere and of unspecified site|KLEBSIELLA PNEUMONIAE
Finding|Finding|Impression|7654,7660|false|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organ or Tissue Function|Impression|7654,7660|false|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organism Function|Impression|7654,7660|false|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Physiologic Function|Impression|7654,7660|false|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Phenomenon|Phenomenon or Process|Impression|7654,7660|false|false|false|C2911660|Growth action|GROWTH
Drug|Antibiotic|Impression|7672,7681|false|false|false|C0007546|cefazolin|Cefazolin
Drug|Organic Chemical|Impression|7672,7681|false|false|false|C0007546|cefazolin|Cefazolin
Finding|Idea or Concept|Impression|7697,7705|false|false|false|C0243161|criteria|criteria
Finding|Intellectual Product|Impression|7729,7736|false|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|Impression|7729,7736|false|false|false|C0040808|Treatment Protocols|regimen
Finding|Classification|Impression|7774,7782|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|NEGATIVE
Finding|Finding|Impression|7774,7782|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|NEGATIVE
Lab|Laboratory or Test Result|Impression|7774,7782|false|false|false|C5237010|Expression Negative|NEGATIVE
Anatomy|Cell|Impression|7783,7786|false|false|false|C0206427|Rod Photoreceptors|ROD
Disorder|Disease or Syndrome|Impression|7783,7786|false|false|false|C0035086|Renal Osteodystrophy|ROD
Finding|Gene or Genome|Impression|7783,7786|false|false|false|C1424852|KNTC1 gene|ROD
Finding|Finding|Impression|7801,7807|false|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organ or Tissue Function|Impression|7801,7807|false|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organism Function|Impression|7801,7807|false|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Physiologic Function|Impression|7801,7807|false|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Phenomenon|Phenomenon or Process|Impression|7801,7807|false|false|false|C2911660|Growth action|GROWTH
Finding|Finding|Impression|7841,7854|false|false|false|C0427965|Antimicrobial susceptibility|SENSITIVITIES
Disorder|Neoplastic Process|Impression|7856,7859|false|false|false|C2732473|Ductal Carcinoma In Situ with Microinvasion|MIC
Drug|Hazardous or Poisonous Substance|Impression|7856,7859|false|false|false|C0066256|methyl isocyanate|MIC
Drug|Organic Chemical|Impression|7856,7859|false|false|false|C0066256|methyl isocyanate|MIC
Procedure|Laboratory Procedure|Impression|7856,7859|false|false|false|C0281162;C0427978|Minimum Inhibitory Concentration Test;cisplatin/ifosfamide/mitomycin protocol|MIC
Procedure|Therapeutic or Preventive Procedure|Impression|7856,7859|false|false|false|C0281162;C0427978|Minimum Inhibitory Concentration Test;cisplatin/ifosfamide/mitomycin protocol|MIC
Disorder|Disease or Syndrome|Impression|7991,8001|false|false|false|C0519030|Pneumonia due to Klebsiella pneumoniae|KLEBSIELLA
Disorder|Disease or Syndrome|Impression|7991,8012|false|false|false|C2712605|Infection by Klebsiella pneumoniae in conditions classified elsewhere and of unspecified site|KLEBSIELLA PNEUMONIAE
Drug|Antibiotic|Impression|8047,8057|false|false|false|C0002680;C2095775|ampicillin;ampicillins|AMPICILLIN
Drug|Organic Chemical|Impression|8047,8057|false|false|false|C0002680;C2095775|ampicillin;ampicillins|AMPICILLIN
Drug|Pharmacologic Substance|Impression|8047,8067|false|false|false|C2930041|Ampicillin / Sulbactam|AMPICILLIN/SULBACTAM
Drug|Antibiotic|Impression|8058,8067|false|false|false|C0038665|sulbactam|SULBACTAM
Drug|Organic Chemical|Impression|8058,8067|false|false|false|C0038665|sulbactam|SULBACTAM
Drug|Antibiotic|Impression|8078,8087|false|false|false|C0007546|cefazolin|CEFAZOLIN
Drug|Organic Chemical|Impression|8078,8087|false|false|false|C0007546|cefazolin|CEFAZOLIN
Drug|Antibiotic|Impression|8109,8117|false|false|false|C0055003|cefepime|CEFEPIME
Drug|Organic Chemical|Impression|8109,8117|false|false|false|C0055003|cefepime|CEFEPIME
Drug|Antibiotic|Impression|8140,8151|false|false|false|C0007559|ceftazidime|CEFTAZIDIME
Drug|Organic Chemical|Impression|8140,8151|false|false|false|C0007559|ceftazidime|CEFTAZIDIME
Drug|Antibiotic|Impression|8171,8182|false|false|false|C0007561|ceftriaxone|CEFTRIAXONE
Drug|Organic Chemical|Impression|8171,8182|false|false|false|C0007561|ceftriaxone|CEFTRIAXONE
Drug|Organic Chemical|Impression|8202,8215|false|false|false|C0008809|ciprofloxacin|CIPROFLOXACIN
Drug|Pharmacologic Substance|Impression|8202,8215|false|false|false|C0008809|ciprofloxacin|CIPROFLOXACIN
Drug|Antibiotic|Impression|8233,8243|false|false|false|C3854019|gentamicin|GENTAMICIN
Drug|Organic Chemical|Impression|8233,8243|false|false|false|C3854019|gentamicin|GENTAMICIN
Procedure|Laboratory Procedure|Impression|8233,8243|false|false|false|C0202391|Gentamicin measurement|GENTAMICIN
Drug|Antibiotic|Impression|8264,8273|false|false|false|C0066005;C1314417|INJECTION, MEROPENEM, 100 MG ADMINISTERED;meropenem|MEROPENEM
Drug|Clinical Drug|Impression|8264,8273|false|false|false|C0066005;C1314417|INJECTION, MEROPENEM, 100 MG ADMINISTERED;meropenem|MEROPENEM
Drug|Organic Chemical|Impression|8264,8273|false|false|false|C0066005;C1314417|INJECTION, MEROPENEM, 100 MG ADMINISTERED;meropenem|MEROPENEM
Drug|Antibiotic|Impression|8295,8307|false|false|false|C0031955|piperacillin|PIPERACILLIN
Drug|Organic Chemical|Impression|8295,8307|false|false|false|C0031955|piperacillin|PIPERACILLIN
Drug|Antibiotic|Impression|8308,8312|false|false|false|C0075870|tazobactam|TAZO
Drug|Organic Chemical|Impression|8308,8312|false|false|false|C0075870|tazobactam|TAZO
Drug|Antibiotic|Impression|8326,8336|false|false|false|C0040341|tobramycin|TOBRAMYCIN
Drug|Organic Chemical|Impression|8326,8336|false|false|false|C0040341|tobramycin|TOBRAMYCIN
Procedure|Laboratory Procedure|Impression|8326,8336|false|false|false|C0202490|Tobramycin measurement|TOBRAMYCIN
Drug|Antibiotic|Impression|8357,8369|false|false|false|C0041041|trimethoprim|TRIMETHOPRIM
Drug|Organic Chemical|Impression|8357,8369|false|false|false|C0041041|trimethoprim|TRIMETHOPRIM
Drug|Pharmacologic Substance|Impression|8370,8375|false|false|false|C0749139|sulfa|SULFA
Disorder|Disease or Syndrome|Hospital Course|8436,8439|false|false|false|C0020538|Hypertensive disease|HTN
Disorder|Disease or Syndrome|Hospital Course|8488,8494|false|false|false|C4255010||NSTEMI
Finding|Finding|Hospital Course|8488,8494|false|false|false|C3537184||NSTEMI
Anatomy|Body Location or Region|Hospital Course|8508,8514|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8508,8514|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Disorder|Disease or Syndrome|Hospital Course|8515,8522|false|false|false|C0012634|Disease|disease
Disorder|Disease or Syndrome|Hospital Course|8527,8530|false|false|false|C4551552|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|DES
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8527,8530|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Biologically Active Substance|Hospital Course|8527,8530|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Hormone|Hospital Course|8527,8530|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Organic Chemical|Hospital Course|8527,8530|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Pharmacologic Substance|Hospital Course|8527,8530|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Finding|Gene or Genome|Hospital Course|8527,8530|false|false|false|C1413980|DES gene|DES
Disorder|Acquired Abnormality|Hospital Course|8543,8552|false|false|false|C0001168|Complete obstruction|occlusion
Finding|Finding|Hospital Course|8543,8552|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Functional Concept|Hospital Course|8543,8552|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Organ or Tissue Function|Hospital Course|8543,8552|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Pathologic Function|Hospital Course|8543,8552|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Finding|Hospital Course|8567,8573|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|Hospital Course|8567,8573|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Disorder|Disease or Syndrome|Hospital Course|8613,8619|false|false|false|C4255010||NSTEMI
Finding|Finding|Hospital Course|8613,8619|false|false|false|C3537184||NSTEMI
Disorder|Disease or Syndrome|Hospital Course|8621,8627|false|false|false|C4255010||NSTEMI
Finding|Finding|Hospital Course|8621,8627|false|false|false|C3537184||NSTEMI
Finding|Gene or Genome|Hospital Course|8637,8640|false|false|false|C1420459;C3811127|SULT1E1 gene;SULT1E1 wt Allele|STE
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8663,8674|false|false|false|C0011570|Mental Depression|depressions
Finding|Idea or Concept|Hospital Course|8679,8690|false|false|false|C0750502|Significant|significant
Anatomy|Body Location or Region|Hospital Course|8697,8703|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8697,8703|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Disorder|Disease or Syndrome|Hospital Course|8704,8711|false|false|false|C0012634|Disease|disease
Finding|Idea or Concept|Hospital Course|8716,8727|false|true|false|C0750502|Significant|significant
Finding|Pathologic Function|Hospital Course|8728,8736|false|true|false|C1261287|Stenosis|stenosis
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8740,8743|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|Hospital Course|8740,8743|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Finding|Gene or Genome|Hospital Course|8740,8743|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Disorder|Disease or Syndrome|Hospital Course|8749,8752|false|false|false|C4551552|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|DES
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8749,8752|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Biologically Active Substance|Hospital Course|8749,8752|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Hormone|Hospital Course|8749,8752|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Organic Chemical|Hospital Course|8749,8752|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Pharmacologic Substance|Hospital Course|8749,8752|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Finding|Gene or Genome|Hospital Course|8749,8752|false|false|false|C1413980|DES gene|DES
Finding|Finding|Hospital Course|8758,8766|false|false|false|C0028778;C1947917|Obstruction;Occluded|occluded
Finding|Functional Concept|Hospital Course|8758,8766|false|false|false|C0028778;C1947917|Obstruction;Occluded|occluded
Finding|Functional Concept|Hospital Course|8778,8784|false|false|false|C0205341;C1705914|Repeat;Repeat Object|Repeat
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8785,8789|false|false|false|C0007430|Catheterization|cath
Finding|Finding|Hospital Course|8790,8799|false|false|false|C0442739||unchanged
Drug|Organic Chemical|Hospital Course|8820,8826|false|false|false|C0633084|Plavix|plavix
Drug|Pharmacologic Substance|Hospital Course|8820,8826|false|false|false|C0633084|Plavix|plavix
Drug|Organic Chemical|Hospital Course|8828,8840|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|Hospital Course|8828,8840|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8842,8845|false|false|false|C1452534|ACE protein, human|ACE
Drug|Biologically Active Substance|Hospital Course|8842,8845|false|false|false|C1452534|ACE protein, human|ACE
Finding|Gene or Genome|Hospital Course|8842,8845|false|false|false|C1413931;C4284014|ACE gene;Adverse Childhood Experience questionnaire|ACE
Finding|Intellectual Product|Hospital Course|8842,8845|false|false|false|C1413931;C4284014|ACE gene;Adverse Childhood Experience questionnaire|ACE
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8842,8845|false|false|false|C0050385;C0108844;C0279078;C1879921|CDE Regimen;CDE protocol;cisplatin, cytarabine, and etoposide chemotherapy protocol;cyclophosphamide/doxorubicin protocol|ACE
Drug|Organic Chemical|Hospital Course|8853,8863|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|Hospital Course|8853,8863|false|false|false|C0025859|metoprolol|metoprolol
Procedure|Health Care Activity|Hospital Course|8865,8869|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|Echo
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8865,8869|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|Echo
Attribute|Clinical Attribute|Hospital Course|8878,8882|false|false|false|C0428772|Left ventricular ejection fraction|LVEF
Procedure|Diagnostic Procedure|Hospital Course|8878,8882|false|false|false|C3837267|LVEF (procedure)|LVEF
Finding|Finding|Hospital Course|8895,8906|false|false|false|C0086439|Hypokinesia|hypokinesis
Anatomy|Cell Component|Hospital Course|8938,8942|false|false|false|C3890171|dinoflagellate apex|apex
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8938,8942|false|false|false|C0140145|APEX1 protein, human|apex
Drug|Enzyme|Hospital Course|8938,8942|false|false|false|C0140145|APEX1 protein, human|apex
Finding|Gene or Genome|Hospital Course|8938,8942|false|false|false|C1332102|APEX1 gene|apex
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8959,8970|false|false|false|C0851145|on warfarin|on warfarin
Drug|Hazardous or Poisonous Substance|Hospital Course|8962,8970|false|false|false|C0043031|warfarin|warfarin
Drug|Organic Chemical|Hospital Course|8962,8970|false|false|false|C0043031|warfarin|warfarin
Drug|Pharmacologic Substance|Hospital Course|8962,8970|false|false|false|C0043031|warfarin|warfarin
Finding|Finding|Hospital Course|8979,8990|false|false|false|C0086439|Hypokinesia|hypokinetic
Finding|Finding|Hospital Course|8998,9002|false|false|false|C5575035|Well (answer to question)|well
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9010,9016|false|false|false|C0018792|Heart Atrium|atrial
Attribute|Clinical Attribute|Hospital Course|9010,9029|false|false|false|C2926591||atrial fibrillation
Disorder|Disease or Syndrome|Hospital Course|9010,9029|false|false|false|C0004238|Atrial Fibrillation|atrial fibrillation
Lab|Laboratory or Test Result|Hospital Course|9010,9029|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|atrial fibrillation
Disorder|Disease or Syndrome|Hospital Course|9017,9029|false|false|false|C0232197|Fibrillation|fibrillation
Finding|Finding|Hospital Course|9057,9065|false|false|false|C0332149|Possible|Possibly
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9109,9115|false|false|false|C0042449|Veins|venous
Attribute|Clinical Attribute|Hospital Course|9133,9137|false|false|false|C0034094|Pulmonary Wedge Pressure|PCWP
Drug|Pharmacologic Substance|Hospital Course|9164,9172|false|false|false|C0237795|Pressors|pressors
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9177,9184|false|false|false|C0004704|Balloon Dilatation|balloon
Finding|Molecular Function|Hospital Course|9186,9190|false|false|false|C1150186|matrix metalloproteinase 7 activity|pump
Finding|Intellectual Product|Hospital Course|9199,9203|false|false|false|C1720594|Then - dosing instruction fragment|then
Finding|Finding|Hospital Course|9247,9269|false|false|false|C0578150|Hemodynamically stable|hemodynamically stable
Finding|Intellectual Product|Hospital Course|9263,9269|false|false|false|C1547311|Patient Condition Code - Stable|stable
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9277,9281|false|false|false|C1742913|REST protein, human|rest
Drug|Biologically Active Substance|Hospital Course|9277,9281|false|false|false|C1742913|REST protein, human|rest
Finding|Daily or Recreational Activity|Hospital Course|9277,9281|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Gene or Genome|Hospital Course|9277,9281|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Molecular Function|Hospital Course|9277,9281|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Idea or Concept|Hospital Course|9285,9293|false|false|false|C1547192|Organization unit type - Hospital|hospital
Attribute|Clinical Attribute|Hospital Course|9285,9300|false|false|false|C0488549||hospital course
Finding|Finding|Hospital Course|9285,9300|false|false|false|C0489547|Hospital course|hospital course
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9306,9312|false|false|false|C0018792|Heart Atrium|Atrial
Attribute|Clinical Attribute|Hospital Course|9306,9325|false|false|false|C2926591||Atrial Fibrillation
Disorder|Disease or Syndrome|Hospital Course|9306,9325|false|false|false|C0004238|Atrial Fibrillation|Atrial Fibrillation
Lab|Laboratory or Test Result|Hospital Course|9306,9325|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Atrial Fibrillation
Disorder|Disease or Syndrome|Hospital Course|9313,9325|false|false|false|C0232197|Fibrillation|Fibrillation
Finding|Body Substance|Hospital Course|9326,9333|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|9326,9333|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|9326,9333|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Conceptual Entity|Hospital Course|9350,9357|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|9350,9357|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Hospital Course|9350,9357|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|9350,9360|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|Hospital Course|9372,9376|false|false|false|C0004238|Atrial Fibrillation|afib
Lab|Laboratory or Test Result|Hospital Course|9372,9376|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|afib
Disorder|Disease or Syndrome|Hospital Course|9385,9388|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9385,9388|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|Hospital Course|9385,9388|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9385,9388|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|Hospital Course|9385,9388|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|Hospital Course|9385,9388|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|Hospital Course|9385,9388|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|Hospital Course|9385,9388|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Finding|Gene or Genome|Hospital Course|9385,9388|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|Hospital Course|9385,9388|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Drug|Organic Chemical|Hospital Course|9421,9428|false|false|false|C0012265|digoxin|digoxin
Drug|Pharmacologic Substance|Hospital Course|9421,9428|false|false|false|C0012265|digoxin|digoxin
Procedure|Laboratory Procedure|Hospital Course|9421,9428|false|false|false|C0337449|Digoxin measurement|digoxin
Finding|Finding|Hospital Course|9432,9436|false|false|false|C5575035|Well (answer to question)|well
Drug|Organic Chemical|Hospital Course|9440,9447|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|Hospital Course|9440,9447|false|false|false|C0004057|aspirin|aspirin
Procedure|Health Care Activity|Hospital Course|9473,9482|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9507,9513|false|false|false|C0018792|Heart Atrium|atrial
Disorder|Disease or Syndrome|Hospital Course|9515,9527|false|false|false|C0232197|Fibrillation|fibrillation
Procedure|Health Care Activity|Hospital Course|9535,9544|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Mental Process|Hospital Course|9553,9561|false|false|false|C0679006|Decision|decision
Drug|Organic Chemical|Hospital Course|9594,9602|false|false|false|C0699129|Coumadin|Coumadin
Drug|Pharmacologic Substance|Hospital Course|9594,9602|false|false|false|C0699129|Coumadin|Coumadin
Finding|Idea or Concept|Hospital Course|9625,9629|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|9625,9629|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|9625,9629|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Hospital Course|9636,9643|false|false|false|C0012265|digoxin|digoxin
Drug|Pharmacologic Substance|Hospital Course|9636,9643|false|false|false|C0012265|digoxin|digoxin
Procedure|Laboratory Procedure|Hospital Course|9636,9643|false|false|false|C0337449|Digoxin measurement|digoxin
Finding|Idea or Concept|Hospital Course|9650,9654|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|9650,9654|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|9650,9654|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Hospital Course|9660,9667|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|Hospital Course|9660,9667|false|false|false|C0004057|aspirin|aspirin
Finding|Idea or Concept|Hospital Course|9695,9700|false|false|false|C1552828|Table Frame - above|above
Finding|Functional Concept|Hospital Course|9707,9717|false|false|false|C0589507;C1158830;C1704686|Initiation;Transcription Initiation|initiation
Finding|Genetic Function|Hospital Course|9707,9717|false|false|false|C0589507;C1158830;C1704686|Initiation;Transcription Initiation|initiation
Finding|Mental Process|Hospital Course|9707,9717|false|false|false|C0589507;C1158830;C1704686|Initiation;Transcription Initiation|initiation
Drug|Organic Chemical|Hospital Course|9721,9729|false|false|false|C0699129|Coumadin|Coumadin
Drug|Pharmacologic Substance|Hospital Course|9721,9729|false|false|false|C0699129|Coumadin|Coumadin
Disorder|Disease or Syndrome|Hospital Course|9734,9743|false|false|false|C0018965|Hematuria|Hematuria
Finding|Finding|Hospital Course|9746,9752|false|true|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Finding|Idea or Concept|Hospital Course|9746,9752|false|true|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Finding|Functional Concept|Hospital Course|9753,9762|false|true|false|C0332663|Traumatic|traumatic
Finding|Functional Concept|Hospital Course|9777,9785|false|false|false|C0205373;C5849094|Systemic;Systemic Route of Administration|systemic
Finding|Finding|Hospital Course|9786,9801|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Finding|Physiologic Function|Hospital Course|9786,9801|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9786,9801|false|false|false|C0003281|Anticoagulation Therapy|anticoagulation
Finding|Body Substance|Hospital Course|9807,9814|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|9807,9814|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|9807,9814|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Procedure|Laboratory Procedure|Hospital Course|9830,9838|false|false|false|C0010818;C1305671|Cytological Techniques;Cytology--Technique|Cytology
Finding|Classification|Hospital Course|9843,9851|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|9843,9851|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|9843,9851|false|false|false|C5237010|Expression Negative|negative
Finding|Classification|Hospital Course|9871,9881|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|9871,9881|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Finding|Hospital Course|9899,9906|false|false|false|C0013404;C2024878|Dyspnea|Dyspnea
Finding|Sign or Symptom|Hospital Course|9899,9906|false|false|false|C0013404;C2024878|Dyspnea|Dyspnea
Finding|Body Substance|Hospital Course|9909,9916|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|9909,9916|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|9909,9916|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|9921,9926|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Finding|Hospital Course|9939,9946|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|Hospital Course|9939,9946|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9980,9989|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Hospital Course|9980,9989|false|false|false|C2707265||pulmonary
Finding|Finding|Hospital Course|9980,9989|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|Hospital Course|9980,9995|false|false|false|C0034063|Pulmonary Edema|pulmonary edema
Attribute|Clinical Attribute|Hospital Course|9990,9995|false|false|false|C1717255||edema
Finding|Pathologic Function|Hospital Course|9990,9995|false|false|false|C0013604|Edema|edema
Finding|Finding|Hospital Course|10000,10008|false|false|false|C0184511;C1561611;C4084203|Admission Level of Care Code - Improved;Improved;Improved - answer to question|improved
Finding|Intellectual Product|Hospital Course|10000,10008|false|false|false|C0184511;C1561611;C4084203|Admission Level of Care Code - Improved;Improved;Improved - answer to question|improved
Procedure|Diagnostic Procedure|Hospital Course|10040,10043|false|false|false|C0039985|Plain chest X-ray|CXR
Finding|Finding|Hospital Course|10051,10059|false|false|false|C0332149|Possible|possible
Disorder|Disease or Syndrome|Hospital Course|10060,10073|false|true|false|C0521530|Lung consolidation|consolidation
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10077,10080|false|false|false|C1261074|Structure of right upper lobe of lung|RUL
Disorder|Injury or Poisoning|Hospital Course|10098,10108|false|false|false|C1720922|Respiratory Aspiration|aspiration
Finding|Finding|Hospital Course|10098,10108|false|false|false|C0220787;C0700198;C2712334|Aspiration into respiratory tract;Endotracheal aspiration;Pulmonary aspiration|aspiration
Finding|Organ or Tissue Function|Hospital Course|10098,10108|false|false|false|C0220787;C0700198;C2712334|Aspiration into respiratory tract;Endotracheal aspiration;Pulmonary aspiration|aspiration
Finding|Pathologic Function|Hospital Course|10098,10108|false|false|false|C0220787;C0700198;C2712334|Aspiration into respiratory tract;Endotracheal aspiration;Pulmonary aspiration|aspiration
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10098,10108|false|false|false|C0349707||aspiration
Disorder|Disease or Syndrome|Hospital Course|10098,10118|false|false|false|C0032290;C1761609|Aspiration Pneumonia;Aspiration pneumonitis|aspiration pneumonia
Disorder|Disease or Syndrome|Hospital Course|10109,10118|false|false|false|C0032285|Pneumonia|pneumonia
Finding|Conceptual Entity|Hospital Course|10129,10138|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|Hospital Course|10129,10138|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|Hospital Course|10129,10138|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10129,10138|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Finding|Finding|Hospital Course|10178,10183|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|Hospital Course|10178,10183|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Disorder|Disease or Syndrome|Hospital Course|10187,10197|false|false|false|C0009450|Communicable Diseases|infectious
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Hospital Course|10198,10201|false|false|false|C0600500|Peptide Nucleic Acids|pna
Finding|Body Substance|Hospital Course|10217,10223|false|false|false|C0038056;C1546789;C1576419|Specimen Type - Sputum;Sputum|sputum
Finding|Intellectual Product|Hospital Course|10217,10223|false|false|false|C0038056;C1546789;C1576419|Specimen Type - Sputum;Sputum|sputum
Finding|Idea or Concept|Hospital Course|10224,10232|false|true|false|C0010453|Culture (Anthropological)|cultures
Disorder|Disease or Syndrome|Hospital Course|10244,10254|false|false|false|C0519030|Pneumonia due to Klebsiella pneumoniae|Klebsiella
Disorder|Disease or Syndrome|Hospital Course|10244,10264|false|false|false|C0519030|Pneumonia due to Klebsiella pneumoniae|Klebsiella pneumonia
Disorder|Disease or Syndrome|Hospital Course|10255,10264|false|false|false|C0032285|Pneumonia|pneumonia
Finding|Social Behavior|Hospital Course|10273,10283|false|false|false|C2584313|Discussion (communication)|discussion
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10273,10283|false|false|false|C0557061|Discussion (procedure)|discussion
Finding|Conceptual Entity|Hospital Course|10323,10332|true|false|true|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|Hospital Course|10323,10332|true|false|true|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|Hospital Course|10323,10332|true|false|true|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10323,10332|true|false|true|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Finding|Finding|Hospital Course|10344,10356|false|false|false|C0231221;C0332151|Asymptomatic (finding);Asymptomatic diagnosis of|asymptomatic
Drug|Organic Chemical|Hospital Course|10383,10388|false|false|false|C0699992|Lasix|lasix
Drug|Pharmacologic Substance|Hospital Course|10383,10388|false|false|false|C0699992|Lasix|lasix
Finding|Idea or Concept|Hospital Course|10407,10411|false|false|false|C1552851|next - HtmlLinkType|next
Drug|Inorganic Chemical|Hospital Course|10412,10424|false|false|false|C0013832;C3536863|Electrolyte [EPC];Electrolytes|electrolytes
Drug|Pharmacologic Substance|Hospital Course|10412,10424|false|false|false|C0013832;C3536863|Electrolyte [EPC];Electrolytes|electrolytes
Finding|Finding|Hospital Course|10457,10463|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|Hospital Course|10457,10463|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Sign or Symptom|Hospital Course|10470,10481|false|false|false|C2129214|Loose stool|loose stool
Finding|Body Substance|Hospital Course|10476,10481|false|true|false|C0015733|Feces|stool
Finding|Mental Process|Hospital Course|10485,10492|false|false|false|C0542559|contextual factors|setting
Drug|Antibiotic|Hospital Course|10496,10506|false|false|false|C0003232|Antibiotics|antibiotic
Finding|Classification|Hospital Course|10534,10544|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|10534,10544|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Anatomy|Cell|Hospital Course|10553,10556|false|false|false|C0023516|Leukocytes|WBC
Attribute|Clinical Attribute|Hospital Course|10567,10570|false|false|false|C1114365||age
Drug|Biologically Active Substance|Hospital Course|10567,10570|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|Hospital Course|10567,10570|false|false|false|C0162574|Glycation End Products, Advanced|age
Finding|Finding|Hospital Course|10588,10594|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|Hospital Course|10588,10594|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Body Substance|Hospital Course|10596,10603|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|10596,10603|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|10596,10603|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10619,10629|false|false|false|C0042313|vancomycin|vancomycin
Drug|Antibiotic|Hospital Course|10619,10629|false|false|false|C0042313|vancomycin|vancomycin
Procedure|Laboratory Procedure|Hospital Course|10619,10629|false|false|false|C0489941|Vancomycin measurement|vancomycin
Finding|Idea or Concept|Hospital Course|10651,10654|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|10651,10654|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Idea or Concept|Hospital Course|10663,10666|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|10663,10666|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Idea or Concept|Hospital Course|10677,10680|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|10677,10680|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Anatomy|Body Location or Region|Hospital Course|10691,10707|false|false|false|C0744316|gastroesophageal|GASTROESOPHAGEAL
Disorder|Disease or Syndrome|Hospital Course|10691,10714|false|false|false|C0017168|Gastroesophageal reflux disease|GASTROESOPHAGEAL REFLUX
Finding|Finding|Hospital Course|10691,10714|false|false|false|C3813607;C4317146|Acid reflux;Infantile Gastroesophageal Reflux|GASTROESOPHAGEAL REFLUX
Disorder|Disease or Syndrome|Hospital Course|10691,10722|false|false|false|C0017168|Gastroesophageal reflux disease|GASTROESOPHAGEAL REFLUX DISEASE
Disorder|Disease or Syndrome|Hospital Course|10691,10729|false|false|false|C0017168|Gastroesophageal reflux disease|GASTROESOPHAGEAL REFLUX DISEASE (GERD)
Finding|Pathologic Function|Hospital Course|10708,10714|false|false|false|C0232483|Reflux|REFLUX
Disorder|Disease or Syndrome|Hospital Course|10715,10722|false|false|false|C0012634|Disease|DISEASE
Disorder|Disease or Syndrome|Hospital Course|10724,10728|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Procedure|Diagnostic Procedure|Hospital Course|10732,10741|false|false|false|C0014245;C0079278|Endoscopy (procedure);Endoscopy, Gastrointestinal|Endoscopy
Drug|Pharmacologic Substance|Hospital Course|10774,10777|false|false|false|C0358591|Proton Pump Inhibitors|PPI
Finding|Physiologic Function|Hospital Course|10774,10777|false|false|false|C0871125|Prepulse Inhibition|PPI
Drug|Antibiotic|Hospital Course|10781,10795|false|false|false|C0055856|clarithromycin|clarithromycin
Drug|Organic Chemical|Hospital Course|10781,10795|false|false|false|C0055856|clarithromycin|clarithromycin
Drug|Antibiotic|Hospital Course|10796,10807|false|false|false|C0002645|amoxicillin|amoxicillin
Drug|Organic Chemical|Hospital Course|10796,10807|false|false|false|C0002645|amoxicillin|amoxicillin
Drug|Organic Chemical|Hospital Course|10831,10841|false|false|false|C0028978|omeprazole|Omeprazole
Drug|Pharmacologic Substance|Hospital Course|10831,10841|false|false|false|C0028978|omeprazole|Omeprazole
Drug|Antibiotic|Hospital Course|10858,10869|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|Antibiotics
Finding|Mental Process|Hospital Course|10878,10885|false|false|false|C0542559|contextual factors|setting
Disorder|Disease or Syndrome|Hospital Course|10889,10905|false|false|false|C0343386|Clostridium difficile infection|c.diff infection
Disorder|Disease or Syndrome|Hospital Course|10896,10905|false|false|false|C0009450|Communicable Diseases|infection
Finding|Pathologic Function|Hospital Course|10896,10905|false|false|false|C3714514|Infection|infection
Disorder|Mental or Behavioral Dysfunction|Hospital Course|10911,10919|false|false|false|C0011206|Delirium|Delirium
Finding|Body Substance|Hospital Course|10922,10929|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|10922,10929|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|10922,10929|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Disorder|Mental or Behavioral Dysfunction|Hospital Course|10944,10954|false|false|false|C1142436|Sundowning|sundowning
Procedure|Health Care Activity|Hospital Course|10962,10977|false|false|false|C0019993|Hospitalization|hospitalization
Drug|Organic Chemical|Hospital Course|10989,10997|false|false|false|C0287163|Seroquel|Seroquel
Drug|Pharmacologic Substance|Hospital Course|10989,10997|false|false|false|C0287163|Seroquel|Seroquel
Finding|Intellectual Product|Hospital Course|11003,11010|false|false|false|C1547296|Chronic - Admission Level of Care Code|CHRONIC
Procedure|Health Care Activity|Hospital Course|11003,11010|false|false|false|C1555457|Provision of recurring care for chronic illness|CHRONIC
Disorder|Acquired Abnormality|Hospital Course|11036,11051|false|false|false|C0037944;C1861329|Spinal Stenosis;Spinal canal stenosis|Spinal Stenosis
Disorder|Anatomical Abnormality|Hospital Course|11036,11051|false|false|false|C0037944;C1861329|Spinal Stenosis;Spinal canal stenosis|Spinal Stenosis
Finding|Pathologic Function|Hospital Course|11043,11051|false|false|false|C1261287|Stenosis|Stenosis
Drug|Organic Chemical|Hospital Course|11063,11073|false|false|false|C0060926|gabapentin|gabapentin
Drug|Pharmacologic Substance|Hospital Course|11063,11073|false|false|false|C0060926|gabapentin|gabapentin
Disorder|Disease or Syndrome|Hospital Course|11077,11080|false|false|false|C0011989;C4551571|Camurati-Engelmann Syndrome;Cranioectodermal dysplasia|ced
Drug|Antibiotic|Hospital Course|11077,11080|false|false|false|C0007738|cephradine|ced
Drug|Organic Chemical|Hospital Course|11077,11080|false|false|false|C0007738|cephradine|ced
Finding|Functional Concept|Hospital Course|11077,11080|false|false|false|C1366557;C1704974;C3890738|Convection-Enhanced Delivery;TGFB1 gene;TGFB1 wt Allele|ced
Finding|Gene or Genome|Hospital Course|11077,11080|false|false|false|C1366557;C1704974;C3890738|Convection-Enhanced Delivery;TGFB1 gene;TGFB1 wt Allele|ced
Procedure|Therapeutic or Preventive Procedure|Hospital Course|11077,11080|false|false|false|C0108844;C0280001|CDE protocol;cisplatin/dexamethasone/etoposide protocol|ced
Drug|Organic Chemical|Hospital Course|11081,11089|false|false|false|C0027396|naproxen|naproxen
Drug|Pharmacologic Substance|Hospital Course|11081,11089|false|false|false|C0027396|naproxen|naproxen
Attribute|Clinical Attribute|Hospital Course|11113,11117|false|true|false|C2598155||pain
Finding|Functional Concept|Hospital Course|11113,11117|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|11113,11117|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Idea or Concept|Hospital Course|11129,11137|false|false|false|C1547192|Organization unit type - Hospital|hospital
Attribute|Clinical Attribute|Hospital Course|11129,11144|true|false|false|C0488549||hospital course
Finding|Finding|Hospital Course|11129,11144|true|false|false|C0489547|Hospital course|hospital course
Drug|Pharmacologic Substance|Hospital Course|11186,11192|false|true|false|C0003211;C0358845|Analgesics and non-steroidal anti-inflammatory drugs;Anti-Inflammatory Agents, Non-Steroidal|NSAIDS
Finding|Mental Process|Hospital Course|11196,11203|false|false|false|C0542559|contextual factors|setting
Anatomy|Body Space or Junction|Hospital Course|11214,11217|false|false|false|C0262187|anterior calcarine sulcus (human only)|ACS
Disorder|Disease or Syndrome|Hospital Course|11214,11217|false|false|false|C0742343;C0796147|Acrocallosal Syndrome;Acute Chest Syndrome|ACS
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11214,11217|false|false|false|C4042561|ACSS2 protein, human|ACS
Drug|Enzyme|Hospital Course|11214,11217|false|false|false|C4042561|ACSS2 protein, human|ACS
Finding|Gene or Genome|Hospital Course|11214,11217|false|false|false|C1150760;C1424787;C1825842;C1842089;C2266615;C4318612;C5400867;C5551036|ACCS gene;ACS - Activity Card Sort;ACSS2 gene;ACSS2 wt Allele;American Community Survey;CO-methylating acetyl-CoA synthase activity;PLA2G15 gene;acetate-CoA ligase activity|ACS
Finding|Intellectual Product|Hospital Course|11214,11217|false|false|false|C1150760;C1424787;C1825842;C1842089;C2266615;C4318612;C5400867;C5551036|ACCS gene;ACS - Activity Card Sort;ACSS2 gene;ACSS2 wt Allele;American Community Survey;CO-methylating acetyl-CoA synthase activity;PLA2G15 gene;acetate-CoA ligase activity|ACS
Finding|Molecular Function|Hospital Course|11214,11217|false|false|false|C1150760;C1424787;C1825842;C1842089;C2266615;C4318612;C5400867;C5551036|ACCS gene;ACS - Activity Card Sort;ACSS2 gene;ACSS2 wt Allele;American Community Survey;CO-methylating acetyl-CoA synthase activity;PLA2G15 gene;acetate-CoA ligase activity|ACS
Drug|Organic Chemical|Hospital Course|11230,11238|false|false|false|C0699129|Coumadin|Coumadin
Drug|Pharmacologic Substance|Hospital Course|11230,11238|false|false|false|C0699129|Coumadin|Coumadin
Drug|Organic Chemical|Hospital Course|11240,11246|false|false|false|C0633084|Plavix|Plavix
Drug|Pharmacologic Substance|Hospital Course|11240,11246|false|false|false|C0633084|Plavix|Plavix
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11251,11254|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|asa
Drug|Enzyme|Hospital Course|11251,11254|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|asa
Drug|Organic Chemical|Hospital Course|11251,11254|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|asa
Drug|Pharmacologic Substance|Hospital Course|11251,11254|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|asa
Finding|Gene or Genome|Hospital Course|11251,11254|false|false|false|C1412553|ARSA gene|asa
Disorder|Congenital Abnormality|Hospital Course|11277,11280|false|false|false|C1845118|SHORT STATURE, IDIOPATHIC, X-LINKED|ISS
Procedure|Health Care Activity|Hospital Course|11288,11297|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Idea or Concept|Hospital Course|11316,11320|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|11316,11320|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|11316,11320|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Hospital Course|11322,11331|false|false|false|C0017642|glipizide|glipizide
Drug|Pharmacologic Substance|Hospital Course|11322,11331|false|false|false|C0017642|glipizide|glipizide
Drug|Organic Chemical|Hospital Course|11336,11345|false|false|false|C0025598|metformin|metformin
Drug|Pharmacologic Substance|Hospital Course|11336,11345|false|false|false|C0025598|metformin|metformin
Disorder|Disease or Syndrome|Hospital Course|11348,11351|false|false|false|C0020538|Hypertensive disease|HTN
Finding|Idea or Concept|Hospital Course|11353,11357|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|11353,11357|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|11353,11357|false|false|false|C1553498|home health encounter|Home
Drug|Organic Chemical|Hospital Course|11363,11373|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|Hospital Course|11363,11373|false|false|false|C0025859|metoprolol|metoprolol
Finding|Idea or Concept|Hospital Course|11387,11391|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|11387,11391|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|11387,11391|false|false|false|C1553498|home health encounter|Home
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11397,11407|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|Hospital Course|11397,11407|false|false|false|C0065374|lisinopril|lisinopril
Finding|Idea or Concept|Hospital Course|11421,11425|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|11421,11425|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|11421,11425|false|false|false|C1553498|home health encounter|Home
Drug|Organic Chemical|Hospital Course|11431,11436|false|false|false|C0590690|Imdur|imdur
Drug|Pharmacologic Substance|Hospital Course|11431,11436|false|false|false|C0590690|Imdur|imdur
Finding|Idea or Concept|Hospital Course|11471,11475|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|11471,11475|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|11471,11475|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Hospital Course|11481,11492|false|false|false|C0074554|simvastatin|simvastatin
Drug|Pharmacologic Substance|Hospital Course|11481,11492|false|false|false|C0074554|simvastatin|simvastatin
Drug|Organic Chemical|Hospital Course|11496,11508|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|Hospital Course|11496,11508|false|false|false|C0286651|atorvastatin|atorvastatin
Finding|Idea or Concept|Hospital Course|11510,11522|false|false|false|C1548597|Marketing basis - Transitional|TRANSITIONAL
Finding|Body Substance|Hospital Course|11554,11563|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|11554,11563|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|11554,11563|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|11554,11563|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|11564,11570|false|false|false|C0944911||weight
Finding|Finding|Hospital Course|11564,11570|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|Hospital Course|11564,11570|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|Hospital Course|11564,11570|false|false|false|C1305866|Weighing patient|weight
Finding|Body Substance|Hospital Course|11582,11589|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|11582,11589|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|11582,11589|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Procedure|Health Care Activity|Hospital Course|11611,11619|false|false|false|C1522577|follow-up|followup
Disorder|Disease or Syndrome|Hospital Course|11626,11635|false|false|false|C0018965|Hematuria|hematuria
Procedure|Health Care Activity|Hospital Course|11644,11653|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Body Substance|Hospital Course|11656,11661|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Finding|Functional Concept|Hospital Course|11656,11661|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Finding|Intellectual Product|Hospital Course|11656,11661|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Finding|Finding|Hospital Course|11656,11670|false|false|false|C0587953|Urine cytology (finding)|Urine cytology
Procedure|Laboratory Procedure|Hospital Course|11656,11670|false|false|false|C2979983|Urine cytology|Urine cytology
Procedure|Laboratory Procedure|Hospital Course|11662,11670|false|false|false|C0010818;C1305671|Cytological Techniques;Cytology--Technique|cytology
Finding|Classification|Hospital Course|11671,11679|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|11671,11679|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|11671,11679|false|false|false|C5237010|Expression Negative|negative
Finding|Body Substance|Hospital Course|11683,11690|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|11683,11690|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|11683,11690|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11761,11771|false|false|false|C0042313|vancomycin|Vancomycin
Drug|Antibiotic|Hospital Course|11761,11771|false|false|false|C0042313|vancomycin|Vancomycin
Procedure|Laboratory Procedure|Hospital Course|11761,11771|false|false|false|C0489941|Vancomycin measurement|Vancomycin
Finding|Finding|Hospital Course|11776,11782|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|Severe
Finding|Intellectual Product|Hospital Course|11776,11782|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|Severe
Drug|Inorganic Chemical|Hospital Course|11804,11816|false|false|false|C0013832;C3536863|Electrolyte [EPC];Electrolytes|electrolytes
Drug|Pharmacologic Substance|Hospital Course|11804,11816|false|false|false|C0013832;C3536863|Electrolyte [EPC];Electrolytes|electrolytes
Drug|Organic Chemical|Hospital Course|11835,11843|false|false|false|C0699129|Coumadin|Coumadin
Drug|Pharmacologic Substance|Hospital Course|11835,11843|false|false|false|C0699129|Coumadin|Coumadin
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11860,11866|false|false|false|C0018792|Heart Atrium|atrial
Attribute|Clinical Attribute|Hospital Course|11860,11879|false|false|false|C2926591||atrial fibrillation
Disorder|Disease or Syndrome|Hospital Course|11860,11879|false|false|false|C0004238|Atrial Fibrillation|atrial fibrillation
Lab|Laboratory or Test Result|Hospital Course|11860,11879|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|atrial fibrillation
Disorder|Disease or Syndrome|Hospital Course|11867,11879|false|false|false|C0232197|Fibrillation|fibrillation
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11881,11884|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Enzyme|Hospital Course|11881,11884|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Organic Chemical|Hospital Course|11881,11884|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Pharmacologic Substance|Hospital Course|11881,11884|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Finding|Gene or Genome|Hospital Course|11881,11884|false|false|false|C1412553|ARSA gene|ASA
Drug|Organic Chemical|Hospital Course|11936,11942|false|false|false|C0633084|Plavix|Plavix
Drug|Pharmacologic Substance|Hospital Course|11936,11942|false|false|false|C0633084|Plavix|Plavix
Procedure|Therapeutic or Preventive Procedure|Hospital Course|11956,11971|false|false|false|C2348535|Stenting|stent placement
Procedure|Health Care Activity|Hospital Course|11962,11971|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|Hospital Course|11962,11971|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Drug|Organic Chemical|Hospital Course|11973,11985|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|Hospital Course|11973,11985|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Organic Chemical|Hospital Course|12002,12013|false|false|false|C0074554|simvastatin|simvastatin
Drug|Pharmacologic Substance|Hospital Course|12002,12013|false|false|false|C0074554|simvastatin|simvastatin
Drug|Organic Chemical|Hospital Course|12020,12025|false|false|false|C0699992|Lasix|Lasix
Drug|Pharmacologic Substance|Hospital Course|12020,12025|false|false|false|C0699992|Lasix|Lasix
Finding|Idea or Concept|Hospital Course|12043,12047|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|12043,12047|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|12043,12047|false|false|false|C1553498|home health encounter|Home
Drug|Organic Chemical|Hospital Course|12048,12058|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|Hospital Course|12048,12058|false|false|false|C0025859|metoprolol|metoprolol
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12107,12117|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|Hospital Course|12107,12117|false|false|false|C0065374|lisinopril|lisinopril
Finding|Idea or Concept|Hospital Course|12151,12155|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|12151,12155|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|12151,12155|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Hospital Course|12156,12161|false|false|false|C0590690|Imdur|imdur
Drug|Pharmacologic Substance|Hospital Course|12156,12161|false|false|false|C0590690|Imdur|imdur
Finding|Body Substance|Hospital Course|12182,12189|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|12182,12189|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|12182,12189|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|12217,12220|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|12217,12220|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Idea or Concept|Hospital Course|12240,12243|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|12240,12243|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Idea or Concept|Hospital Course|12259,12262|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|12259,12262|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Disorder|Disease or Syndrome|Hospital Course|12277,12286|false|false|false|C0009450|Communicable Diseases|infection
Finding|Pathologic Function|Hospital Course|12277,12286|false|false|false|C3714514|Infection|infection
Finding|Body Substance|Hospital Course|12289,12296|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|12289,12296|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|12289,12296|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Pharmacologic Substance|Hospital Course|12324,12330|true|false|false|C0003211;C0358845|Analgesics and non-steroidal anti-inflammatory drugs;Anti-Inflammatory Agents, Non-Steroidal|NSAIDS
Finding|Gene or Genome|Hospital Course|12333,12336|false|false|false|C1412999;C4283853|C4A gene;C4A wt Allele|SLP
Finding|Conceptual Entity|Hospital Course|12337,12346|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|Hospital Course|12337,12346|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|Hospital Course|12337,12346|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|Hospital Course|12337,12346|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|Hospital Course|12350,12355|false|false|false|C0034991|Rehabilitation therapy|rehab
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|12360,12370|false|false|false|C0031354|Pharyngeal structure|pharyngeal
Procedure|Therapeutic or Preventive Procedure|Hospital Course|12371,12394|false|false|false|C0452260|Muscular strength development exercise|strengthening exercises
Finding|Daily or Recreational Activity|Hospital Course|12385,12394|false|false|false|C0015259|Exercise|exercises
Procedure|Therapeutic or Preventive Procedure|Hospital Course|12385,12394|false|false|false|C0452240|Physical therapy exercises|exercises
Attribute|Clinical Attribute|Hospital Course|12397,12408|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|12397,12408|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|Hospital Course|12397,12408|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|12397,12421|false|false|false|C1627937|Medications on admission|Medications on Admission
Procedure|Health Care Activity|Hospital Course|12412,12421|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|Hospital Course|12440,12450|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|Hospital Course|12440,12450|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|Hospital Course|12440,12455|false|false|false|C0746470|MEDICATION LIST|Medication list
Finding|Intellectual Product|Hospital Course|12451,12455|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Drug|Organic Chemical|Hospital Course|12472,12480|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|Hospital Course|12472,12480|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|Hospital Course|12472,12480|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Finding|Functional Concept|Hospital Course|12472,12480|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|Hospital Course|12472,12480|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Organic Chemical|Hospital Course|12485,12495|false|false|false|C0060926|gabapentin|Gabapentin
Drug|Pharmacologic Substance|Hospital Course|12485,12495|false|false|false|C0060926|gabapentin|Gabapentin
Drug|Organic Chemical|Hospital Course|12514,12522|false|false|false|C0027396|naproxen|Naproxen
Drug|Pharmacologic Substance|Hospital Course|12514,12522|false|false|false|C0027396|naproxen|Naproxen
Drug|Organic Chemical|Hospital Course|12543,12552|false|false|false|C0025598|metformin|MetFORMIN
Drug|Pharmacologic Substance|Hospital Course|12543,12552|false|false|false|C0025598|metformin|MetFORMIN
Drug|Organic Chemical|Hospital Course|12554,12564|false|false|false|C0591573|Glucophage|Glucophage
Drug|Pharmacologic Substance|Hospital Course|12554,12564|false|false|false|C0591573|Glucophage|Glucophage
Disorder|Mental or Behavioral Dysfunction|Hospital Course|12576,12579|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12576,12579|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|12576,12579|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|12576,12579|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|12584,12594|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|Hospital Course|12584,12594|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Organic Chemical|Hospital Course|12584,12604|false|false|false|C0724633|metoprolol succinate|Metoprolol Succinate
Drug|Pharmacologic Substance|Hospital Course|12584,12604|false|false|false|C0724633|metoprolol succinate|Metoprolol Succinate
Drug|Organic Chemical|Hospital Course|12595,12604|false|false|false|C0038617;C0220918|Succinates;succinate|Succinate
Drug|Organic Chemical|Hospital Course|12627,12636|false|false|false|C0017642|glipizide|GlipiZIDE
Drug|Pharmacologic Substance|Hospital Course|12627,12636|false|false|false|C0017642|glipizide|GlipiZIDE
Disorder|Mental or Behavioral Dysfunction|Hospital Course|12647,12650|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12647,12650|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|12647,12650|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|12647,12650|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|12655,12666|false|false|false|C0074554|simvastatin|Simvastatin
Drug|Pharmacologic Substance|Hospital Course|12655,12666|false|false|false|C0074554|simvastatin|Simvastatin
Drug|Organic Chemical|Hospital Course|12684,12694|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Pharmacologic Substance|Hospital Course|12684,12694|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Organic Chemical|Hospital Course|12684,12706|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Drug|Pharmacologic Substance|Hospital Course|12684,12706|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Finding|Finding|Hospital Course|12708,12716|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|12708,12716|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|12717,12724|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|12717,12724|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|12717,12724|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12745,12755|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Pharmacologic Substance|Hospital Course|12745,12755|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Organic Chemical|Hospital Course|12775,12782|false|false|false|C0012265|digoxin|Digoxin
Drug|Pharmacologic Substance|Hospital Course|12775,12782|false|false|false|C0012265|digoxin|Digoxin
Procedure|Laboratory Procedure|Hospital Course|12775,12782|false|false|false|C0337449|Digoxin measurement|Digoxin
Drug|Organic Chemical|Hospital Course|12806,12813|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|Hospital Course|12806,12813|false|false|false|C0004057|aspirin|Aspirin
Finding|Body Substance|Hospital Course|12834,12843|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|12834,12843|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|12834,12843|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|12834,12843|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|12834,12855|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|12844,12855|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|12844,12855|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|Hospital Course|12844,12855|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Hospital Course|12860,12867|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|Hospital Course|12860,12867|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|Hospital Course|12860,12870|false|false|false|C5874014|Aspirin EC|Aspirin EC
Drug|Pharmacologic Substance|Hospital Course|12860,12870|false|false|false|C5874014|Aspirin EC|Aspirin EC
Drug|Organic Chemical|Hospital Course|12890,12897|false|false|false|C0012265|digoxin|Digoxin
Drug|Pharmacologic Substance|Hospital Course|12890,12897|false|false|false|C0012265|digoxin|Digoxin
Procedure|Laboratory Procedure|Hospital Course|12890,12897|false|false|false|C0337449|Digoxin measurement|Digoxin
Drug|Organic Chemical|Hospital Course|12920,12930|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|Hospital Course|12920,12930|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Organic Chemical|Hospital Course|12920,12940|false|false|false|C0724633|metoprolol succinate|Metoprolol Succinate
Drug|Pharmacologic Substance|Hospital Course|12920,12940|false|false|false|C0724633|metoprolol succinate|Metoprolol Succinate
Drug|Organic Chemical|Hospital Course|12931,12940|false|false|false|C0038617;C0220918|Succinates;succinate|Succinate
Drug|Organic Chemical|Hospital Course|12963,12975|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|Hospital Course|12963,12975|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Hazardous or Poisonous Substance|Hospital Course|12993,13001|false|false|false|C0043031|warfarin|Warfarin
Drug|Organic Chemical|Hospital Course|12993,13001|false|false|false|C0043031|warfarin|Warfarin
Drug|Pharmacologic Substance|Hospital Course|12993,13001|false|false|false|C0043031|warfarin|Warfarin
Drug|Organic Chemical|Hospital Course|13022,13031|false|false|false|C0017642|glipizide|GlipiZIDE
Drug|Pharmacologic Substance|Hospital Course|13022,13031|false|false|false|C0017642|glipizide|GlipiZIDE
Disorder|Mental or Behavioral Dysfunction|Hospital Course|13042,13045|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|13042,13045|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|13042,13045|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|13042,13045|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|13050,13061|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Pharmacologic Substance|Hospital Course|13050,13061|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Organic Chemical|Hospital Course|13081,13091|false|false|false|C0028978|omeprazole|Omeprazole
Drug|Pharmacologic Substance|Hospital Course|13081,13091|false|false|false|C0028978|omeprazole|Omeprazole
Disorder|Mental or Behavioral Dysfunction|Hospital Course|13101,13104|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|13101,13104|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|13101,13104|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|13101,13104|false|false|false|C1332410|BID gene|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|13109,13119|false|false|false|C0042313|vancomycin|Vancomycin
Drug|Antibiotic|Hospital Course|13109,13119|false|false|false|C0042313|vancomycin|Vancomycin
Procedure|Laboratory Procedure|Hospital Course|13109,13119|false|false|false|C0489941|Vancomycin measurement|Vancomycin
Drug|Clinical Drug|Hospital Course|13109,13124|false|false|false|C0360373||Vancomycin Oral
Anatomy|Body Space or Junction|Hospital Course|13120,13124|false|false|false|C0226896|Oral cavity|Oral
Drug|Biomedical or Dental Material|Hospital Course|13120,13124|false|false|false|C1272919|Oral Dosage Form|Oral
Finding|Finding|Hospital Course|13120,13124|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Finding|Functional Concept|Hospital Course|13120,13124|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Drug|Biomedical or Dental Material|Hospital Course|13120,13131|false|false|false|C1273619|Oral Liquid Product|Oral Liquid
Drug|Biomedical or Dental Material|Hospital Course|13125,13131|false|false|false|C0302908;C1697794|Liquid Dosage Form;Liquid substance|Liquid
Drug|Substance|Hospital Course|13125,13131|false|false|false|C0302908;C1697794|Liquid Dosage Form;Liquid substance|Liquid
Finding|Finding|Hospital Course|13125,13131|false|false|false|C1304698|Liquid (finding)|Liquid
Procedure|Therapeutic or Preventive Procedure|Hospital Course|13125,13131|false|false|false|C0301571|Liquid diet|Liquid
Drug|Organic Chemical|Hospital Course|13151,13160|false|false|false|C0025598|metformin|MetFORMIN
Drug|Pharmacologic Substance|Hospital Course|13151,13160|false|false|false|C0025598|metformin|MetFORMIN
Drug|Organic Chemical|Hospital Course|13162,13172|false|false|false|C0591573|Glucophage|Glucophage
Drug|Pharmacologic Substance|Hospital Course|13162,13172|false|false|false|C0591573|Glucophage|Glucophage
Disorder|Mental or Behavioral Dysfunction|Hospital Course|13184,13187|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|13184,13187|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|13184,13187|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|13184,13187|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|13193,13203|false|false|false|C0060926|gabapentin|Gabapentin
Drug|Pharmacologic Substance|Hospital Course|13193,13203|false|false|false|C0060926|gabapentin|Gabapentin
Drug|Amino Acid, Peptide, or Protein|Hospital Course|13223,13233|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Pharmacologic Substance|Hospital Course|13223,13233|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Organic Chemical|Hospital Course|13255,13265|false|false|false|C0016860|furosemide|Furosemide
Drug|Pharmacologic Substance|Hospital Course|13255,13265|false|false|false|C0016860|furosemide|Furosemide
Finding|Body Substance|Hospital Course|13285,13294|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|13285,13294|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|13285,13294|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|13285,13294|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|13285,13306|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|13285,13306|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|13295,13306|false|false|false|C2926604||Disposition
Procedure|Health Care Activity|Hospital Course|13295,13306|false|false|false|C0184758|Patient disposition|Disposition
Finding|Finding|Hospital Course|13308,13316|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|13308,13316|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Procedure|Health Care Activity|Hospital Course|13308,13321|false|false|false|C0023977|long-term care|Extended Care
Event|Activity|Hospital Course|13317,13321|false|false|false|C1947933|care activity|Care
Finding|Finding|Hospital Course|13317,13321|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|Hospital Course|13317,13321|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|Hospital Course|13324,13332|false|false|false|C4695111|ADMIN.FACILITY|Facility
Finding|Body Substance|Hospital Course|13340,13349|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|13340,13349|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|13340,13349|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|13340,13349|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|13340,13359|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|13350,13359|false|false|false|C0945731||Diagnosis
Finding|Classification|Hospital Course|13350,13359|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|13350,13359|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|13350,13359|false|false|false|C0011900|Diagnosis|Diagnosis
Disorder|Disease or Syndrome|Hospital Course|13361,13367|false|false|false|C4255010||NSTEMI
Finding|Finding|Hospital Course|13361,13367|false|false|false|C3537184||NSTEMI
Finding|Finding|Hospital Course|13377,13383|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Hospital Course|13377,13383|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Finding|Hospital Course|13384,13389|false|true|false|C0205430;C3160715|Mixed (Normal and Tumor);Mixed (qualifier value)|mixed
Finding|Functional Concept|Hospital Course|13384,13389|false|true|false|C0205430;C3160715|Mixed (Normal and Tumor);Mixed (qualifier value)|mixed
Disorder|Disease or Syndrome|Hospital Course|13416,13425|false|false|false|C0018965|Hematuria|Hematuria
Finding|Finding|Hospital Course|13426,13433|false|false|false|C0013404;C2024878|Dyspnea|Dyspnea
Finding|Sign or Symptom|Hospital Course|13426,13433|false|false|false|C0013404;C2024878|Dyspnea|Dyspnea
Finding|Gene or Genome|Hospital Course|13437,13440|false|false|false|C0812246;C1710304|TNF gene;TNF wt Allele|dif
Finding|Finding|Hospital Course|13442,13448|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|Hospital Course|13442,13448|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Disorder|Disease or Syndrome|Hospital Course|13449,13453|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Disorder|Mental or Behavioral Dysfunction|Hospital Course|13454,13462|false|false|false|C0011206|Delirium|Delirium
Finding|Mental Process|Discharge Condition|13487,13493|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|13487,13500|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|13487,13500|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|13494,13500|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|13494,13500|false|false|false|C1546481|What subject filter - Status|Status
Finding|Idea or Concept|Discharge Condition|13502,13507|false|false|false|C1550016|Remote control command - Clear|Clear
Finding|Finding|Discharge Condition|13512,13520|false|false|false|C4068804|Coherent|coherent
Attribute|Clinical Attribute|Discharge Condition|13522,13544|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|13522,13544|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Finding|Finding|Discharge Condition|13531,13544|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|13531,13544|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|13546,13551|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|13546,13551|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|13546,13551|false|false|false|C0718338|Alert brand of caffeine|Alert
Finding|Finding|Discharge Condition|13546,13551|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|13546,13551|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|13546,13551|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|13556,13567|false|false|false|C1704675|Interaction|interactive
Finding|Gene or Genome|Discharge Instructions|13595,13599|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Anatomy|Body Location or Region|Discharge Instructions|13665,13670|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Discharge Instructions|13665,13670|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Discharge Instructions|13672,13676|false|false|false|C2598155||pain
Finding|Functional Concept|Discharge Instructions|13672,13676|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|13672,13676|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|13686,13691|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Discharge Instructions|13686,13691|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Discharge Instructions|13686,13691|false|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|Discharge Instructions|13686,13698|false|false|false|C0027051|Myocardial Infarction|heart attack
Finding|Finding|Discharge Instructions|13692,13698|false|false|false|C1261512;C1304680|Attack (finding);Attack behavior|attack
Finding|Social Behavior|Discharge Instructions|13692,13698|false|false|false|C1261512;C1304680|Attack (finding);Attack behavior|attack
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|13707,13711|false|false|false|C0007430|Catheterization|cath
Finding|Gene or Genome|Discharge Instructions|13712,13715|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|lab
Finding|Intellectual Product|Discharge Instructions|13712,13715|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|lab
Finding|Finding|Discharge Instructions|13740,13748|false|false|false|C1706968;C1879887;C2237319|Blockage (obstruction - finding);Partial Blockage within Medical Device|blockage
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|13757,13765|false|false|false|C0003842;C0226004|Arterial system;Arteries|arteries
Anatomy|Body System|Discharge Instructions|13757,13765|false|false|false|C0003842;C0226004|Arterial system;Arteries|arteries
Procedure|Health Care Activity|Discharge Instructions|13757,13765|false|false|false|C0397581|Procedure on artery|arteries
Finding|Finding|Discharge Instructions|13813,13816|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|Discharge Instructions|13813,13816|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Finding|Discharge Instructions|13813,13831|false|false|false|C0020649|Hypotension|low blood pressure
Disorder|Disease or Syndrome|Discharge Instructions|13817,13822|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|Discharge Instructions|13817,13822|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Finding|Discharge Instructions|13817,13831|false|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|blood pressure
Finding|Organism Function|Discharge Instructions|13817,13831|false|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|blood pressure
Procedure|Health Care Activity|Discharge Instructions|13817,13831|false|false|false|C0005824|Blood pressure determination|blood pressure
Finding|Finding|Discharge Instructions|13823,13831|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|Discharge Instructions|13823,13831|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|Discharge Instructions|13823,13831|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|Discharge Instructions|13823,13831|false|false|false|C0033095||pressure
Disorder|Disease or Syndrome|Discharge Instructions|13833,13843|false|false|false|C0009450|Communicable Diseases|infectious
Disorder|Disease or Syndrome|Discharge Instructions|13833,13852|false|false|false|C0013369|Dysentery|infectious diarrhea
Finding|Finding|Discharge Instructions|13844,13852|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|Discharge Instructions|13844,13852|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Disorder|Injury or Poisoning|Discharge Instructions|13858,13864|false|false|false|C1368081;C3263723;C3714660|Physical trauma;Trauma;Traumatic injury|trauma
Procedure|Health Care Activity|Discharge Instructions|13858,13864|false|false|false|C0548346|Trauma assessment and care|trauma
Procedure|Health Care Activity|Discharge Instructions|13877,13886|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|13877,13886|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Finding|Finding|Discharge Instructions|13902,13906|false|false|false|C5575035|Well (answer to question)|well
Attribute|Clinical Attribute|Discharge Instructions|13938,13949|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|13938,13949|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|Discharge Instructions|13938,13949|false|false|false|C4284232|Medications|medications
Drug|Organic Chemical|Discharge Instructions|13992,14000|false|false|false|C0699129|Coumadin|coumadin
Drug|Pharmacologic Substance|Discharge Instructions|13992,14000|false|false|false|C0699129|Coumadin|coumadin
Drug|Pharmacologic Substance|Discharge Instructions|14041,14057|false|false|false|C0003209|Anti-Inflammatory Agents|antiinflammatory
Drug|Pharmacologic Substance|Discharge Instructions|14058,14063|false|false|false|C0013227|Pharmaceutical Preparations|drugs
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|14058,14063|false|false|false|C3687832|Drugs - dental services|drugs
Drug|Pharmacologic Substance|Discharge Instructions|14065,14071|false|false|false|C0003211;C0358845|Analgesics and non-steroidal anti-inflammatory drugs;Anti-Inflammatory Agents, Non-Steroidal|NSAIDS
Drug|Organic Chemical|Discharge Instructions|14081,14090|false|false|false|C0020740|ibuprofen|ibuprofen
Drug|Pharmacologic Substance|Discharge Instructions|14081,14090|false|false|false|C0020740|ibuprofen|ibuprofen
Drug|Organic Chemical|Discharge Instructions|14092,14097|false|false|false|C0593507|Advil|advil
Drug|Pharmacologic Substance|Discharge Instructions|14092,14097|false|false|false|C0593507|Advil|advil
Finding|Gene or Genome|Discharge Instructions|14092,14097|false|false|false|C1422473|AVIL gene|advil
Drug|Organic Chemical|Discharge Instructions|14100,14106|false|false|false|C0699203|Motrin|motrin
Drug|Pharmacologic Substance|Discharge Instructions|14100,14106|false|false|false|C0699203|Motrin|motrin
Drug|Organic Chemical|Discharge Instructions|14108,14113|false|false|false|C0718343|Aleve|aleve
Drug|Pharmacologic Substance|Discharge Instructions|14108,14113|false|false|false|C0718343|Aleve|aleve
Drug|Organic Chemical|Discharge Instructions|14115,14123|false|false|false|C0027396|naproxen|naproxen
Drug|Pharmacologic Substance|Discharge Instructions|14115,14123|false|false|false|C0027396|naproxen|naproxen
Anatomy|Body System|Discharge Instructions|14159,14169|false|false|false|C0007226|Cardiovascular system|cardiology
Disorder|Disease or Syndrome|Discharge Instructions|14174,14177|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|Discharge Instructions|14174,14177|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|Discharge Instructions|14174,14177|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|Discharge Instructions|14174,14177|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|Discharge Instructions|14174,14177|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|Discharge Instructions|14174,14177|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|Discharge Instructions|14174,14177|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|Discharge Instructions|14174,14177|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Finding|Gene or Genome|Discharge Instructions|14174,14177|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|Discharge Instructions|14174,14177|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Activity|Discharge Instructions|14178,14190|false|false|false|C0003629|Appointments|appointments
Finding|Intellectual Product|Discharge Instructions|14214,14222|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|Discharge Instructions|14214,14222|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|Discharge Instructions|14230,14234|false|false|false|C1947933|care activity|care
Finding|Finding|Discharge Instructions|14230,14234|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|14230,14234|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|14230,14237|false|false|false|C1555558|care of - AddressPartType|care of
Event|Activity|Discharge Instructions|14252,14256|false|false|false|C1947933|care activity|Care
Finding|Finding|Discharge Instructions|14252,14256|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|Discharge Instructions|14252,14256|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Attribute|Clinical Attribute|Discharge Instructions|14252,14261|false|false|false|C4321316||Care Team
Finding|Finding|Discharge Instructions|14252,14261|false|false|false|C4321315|Care team|Care Team
Procedure|Health Care Activity|Discharge Instructions|14264,14272|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|14273,14285|false|false|false|C3263700||Instructions
Finding|Intellectual Product|Discharge Instructions|14273,14285|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

