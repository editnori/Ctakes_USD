 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Procedure|Health Care Activity|SIMPLE_SEGMENT|49,58|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|49,63|false|false|false|C2598112||Admission Date
Finding|Body Substance|SIMPLE_SEGMENT|83,92|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|83,92|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|83,92|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|83,92|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|83,97|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|115,120|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|115,120|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|115,120|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|139,142|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|139,142|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|139,142|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|139,142|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|139,142|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|150,157|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|150,157|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|159,167|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Disorder|Injury or Poisoning|Allergies|182,193|false|false|false|C0161486;C2876539|Poisoning by penicillin;Poisoning by, adverse effect of and underdosing of penicillins|Penicillins
Drug|Antibiotic|Allergies|182,193|false|false|false|C0030842|penicillins|Penicillins
Drug|Organic Chemical|Allergies|182,193|false|false|false|C0030842|penicillins|Penicillins
Finding|Pathologic Function|Allergies|182,193|false|false|false|C0413443|Adverse reaction to penicillins|Penicillins
Drug|Organic Chemical|Allergies|196,204|false|false|false|C0699512|Dilantin|Dilantin
Drug|Pharmacologic Substance|Allergies|196,204|false|false|false|C0699512|Dilantin|Dilantin
Drug|Organic Chemical|Allergies|215,221|false|false|false|C0206046|Zofran|Zofran
Drug|Pharmacologic Substance|Allergies|215,221|false|false|false|C0206046|Zofran|Zofran
Drug|Inorganic Chemical|Allergies|226,239|false|false|false|C1512523|hydrochloride|hydrochloride
Drug|Pharmacologic Substance|Allergies|226,239|false|false|false|C1512523|hydrochloride|hydrochloride
Finding|Functional Concept|Allergies|243,252|false|false|false|C1999232|Attending (action)|Attending
Finding|Functional Concept|Chief Complaint|278,283|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Anatomy|Body Location or Region|Chief Complaint|278,287|false|false|false|C0524470|Right hip region structure|Right hip
Finding|Sign or Symptom|Chief Complaint|278,292|false|false|false|C2202100|Pain of right hip joint|Right hip pain
Anatomy|Body Part, Organ, or Organ Component|Chief Complaint|284,287|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|hip
Drug|Amino Acid, Peptide, or Protein|Chief Complaint|284,287|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Biologically Active Substance|Chief Complaint|284,287|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Pharmacologic Substance|Chief Complaint|284,287|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Finding|Gene or Genome|Chief Complaint|284,287|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|hip
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|284,287|false|false|false|C1292890|Procedure on hip|hip
Attribute|Clinical Attribute|Chief Complaint|284,292|false|false|false|C1716793||hip pain
Finding|Sign or Symptom|Chief Complaint|284,292|false|false|false|C0019559;C4551516|Hip joint pain;Hip pain|hip pain
Attribute|Clinical Attribute|Chief Complaint|288,292|false|false|false|C2598155||pain
Finding|Functional Concept|Chief Complaint|288,292|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Chief Complaint|288,292|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Classification|Chief Complaint|296,301|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|302,310|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|302,310|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|314,332|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|323,332|false|false|false|C0945766||Procedure
Event|Occupational Activity|Chief Complaint|323,332|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|323,332|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|323,332|false|false|false|C0184661|Interventional procedure|Procedure
Anatomy|Body Space or Junction|History of Present Illness|399,402|false|false|false|C0262212|Choroidal fissure|CHF
Disorder|Disease or Syndrome|History of Present Illness|399,402|false|false|false|C0018802|Congestive heart failure|CHF
Disorder|Disease or Syndrome|History of Present Illness|404,408|false|false|false|C0004238|Atrial Fibrillation|Afib
Lab|Laboratory or Test Result|History of Present Illness|404,408|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Afib
Finding|Finding|History of Present Illness|417,432|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Finding|Physiologic Function|History of Present Illness|417,432|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|417,432|false|false|false|C0003281|Anticoagulation Therapy|anticoagulation
Finding|Finding|History of Present Illness|434,440|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|History of Present Illness|434,440|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Disorder|Disease or Syndrome|History of Present Illness|450,459|false|false|false|C0002395|Alzheimer's Disease|Alzheimer
Disorder|Disease or Syndrome|History of Present Illness|450,470|false|false|false|C0002395|Alzheimer's Disease|Alzheimer's dementia
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|462,470|false|false|false|C0011265;C0497327|Dementia;Presenile dementia|dementia
Disorder|Disease or Syndrome|History of Present Illness|473,485|false|false|false|C0029456|Osteoporosis|osteoporosis
Finding|Finding|History of Present Illness|473,485|false|false|false|C2911643|Encounter due to family history of osteoporosis|osteoporosis
Disorder|Disease or Syndrome|History of Present Illness|487,490|false|false|false|C0020538|Hypertensive disease|HTN
Procedure|Health Care Activity|History of Present Illness|510,525|false|false|false|C1456630|Assisted Living|assisted living
Finding|Conceptual Entity|History of Present Illness|519,525|false|false|false|C0595998;C4520849;C4551704|Alive;Household composition;Living|living
Finding|Finding|History of Present Illness|519,525|false|false|false|C0595998;C4520849;C4551704|Alive;Household composition;Living|living
Finding|Intellectual Product|History of Present Illness|526,534|false|false|false|C4695111|ADMIN.FACILITY|facility
Anatomy|Body Location or Region|History of Present Illness|541,546|false|false|false|C0524470|Right hip region structure|R hip
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|543,546|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|hip
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|543,546|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Biologically Active Substance|History of Present Illness|543,546|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Pharmacologic Substance|History of Present Illness|543,546|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Finding|Gene or Genome|History of Present Illness|543,546|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|hip
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|543,546|false|false|false|C1292890|Procedure on hip|hip
Attribute|Clinical Attribute|History of Present Illness|543,551|false|false|false|C1716793||hip pain
Finding|Sign or Symptom|History of Present Illness|543,551|false|false|false|C0019559;C4551516|Hip joint pain;Hip pain|hip pain
Attribute|Clinical Attribute|History of Present Illness|547,551|false|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|547,551|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|547,551|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Body Substance|History of Present Illness|558,565|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|558,565|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|558,565|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|History of Present Illness|558,569|false|false|false|C0332310|Has patient|patient has
Finding|Finding|History of Present Illness|570,576|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|History of Present Illness|570,576|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|570,585|false|false|false|C3494652|Severe dementia|severe dementia
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|577,585|false|false|false|C0011265;C0497327|Dementia;Presenile dementia|dementia
Finding|Mental Process|History of Present Illness|592,609|false|false|false|C0025265|Memory, Short-Term|short term memory
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|592,614|false|false|false|C0701811|Poor short-term memory|short term memory loss
Finding|Idea or Concept|History of Present Illness|598,602|false|false|false|C0233324;C1705313|Term (lexical);Term Birth|term
Finding|Organism Function|History of Present Illness|598,602|false|false|false|C0233324;C1705313|Term (lexical);Term Birth|term
Finding|Finding|History of Present Illness|603,609|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Finding|Intellectual Product|History of Present Illness|603,609|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Finding|Mental Process|History of Present Illness|603,609|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|603,614|false|false|false|C0002622|Amnesia|memory loss
Finding|Sign or Symptom|History of Present Illness|603,614|false|false|false|C0751295|Memory Loss|memory loss
Finding|Finding|History of Present Illness|610,614|false|false|false|C5890125|Loss (adaptation)|loss
Finding|Finding|History of Present Illness|622,628|false|false|false|C1299582|Unable|unable
Finding|Conceptual Entity|History of Present Illness|640,647|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|640,647|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|History of Present Illness|640,647|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|649,653|false|false|false|C4281574|Much|Much
Finding|Conceptual Entity|History of Present Illness|661,668|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|661,668|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|History of Present Illness|661,668|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Classification|History of Present Illness|696,702|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|History of Present Illness|696,702|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|History of Present Illness|696,702|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|History of Present Illness|696,702|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Classification|History of Present Illness|742,748|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|History of Present Illness|742,748|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|History of Present Illness|742,748|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|History of Present Illness|742,748|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Finding|History of Present Illness|766,771|false|false|false|C0587267;C3810854|Close;Closed|close
Finding|Functional Concept|History of Present Illness|766,771|false|false|false|C0587267;C3810854|Close;Closed|close
Event|Activity|History of Present Illness|811,815|false|false|false|C1947933|care activity|care
Finding|Finding|History of Present Illness|811,815|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|History of Present Illness|811,815|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Procedure|Health Care Activity|History of Present Illness|843,858|false|false|false|C1456630|Assisted Living|assisted living
Finding|Conceptual Entity|History of Present Illness|852,858|false|false|false|C0595998;C4520849;C4551704|Alive;Household composition;Living|living
Finding|Finding|History of Present Illness|852,858|false|false|false|C0595998;C4520849;C4551704|Alive;Household composition;Living|living
Finding|Intellectual Product|History of Present Illness|859,867|false|false|false|C4695111|ADMIN.FACILITY|facility
Finding|Body Substance|History of Present Illness|891,898|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|891,898|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|891,898|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|History of Present Illness|910,915|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|History of Present Illness|910,919|false|false|false|C0524470|Right hip region structure|right hip
Finding|Sign or Symptom|History of Present Illness|910,924|false|false|false|C2202100|Pain of right hip joint|right hip pain
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|916,919|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|hip
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|916,919|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Biologically Active Substance|History of Present Illness|916,919|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Pharmacologic Substance|History of Present Illness|916,919|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Finding|Gene or Genome|History of Present Illness|916,919|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|hip
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|916,919|false|false|false|C1292890|Procedure on hip|hip
Attribute|Clinical Attribute|History of Present Illness|916,924|false|false|false|C1716793||hip pain
Finding|Sign or Symptom|History of Present Illness|916,924|false|false|false|C0019559;C4551516|Hip joint pain;Hip pain|hip pain
Attribute|Clinical Attribute|History of Present Illness|920,924|false|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|920,924|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|920,924|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Disorder|Injury or Poisoning|History of Present Illness|954,960|true|false|false|C1368081;C3263723;C3714660|Physical trauma;Trauma;Traumatic injury|trauma
Procedure|Health Care Activity|History of Present Illness|954,960|true|false|false|C0548346|Trauma assessment and care|trauma
Disorder|Injury or Poisoning|History of Present Illness|974,979|true|false|false|C0000921|Accidental Falls|falls
Finding|Finding|History of Present Illness|974,979|true|false|false|C0085639|Falls|falls
Finding|Functional Concept|History of Present Illness|1015,1023|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|History of Present Illness|1015,1023|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Body Substance|History of Present Illness|1074,1081|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|1074,1081|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|1074,1081|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Procedure|Health Care Activity|History of Present Illness|1102,1117|false|false|false|C1456630|Assisted Living|Assisted living
Finding|Conceptual Entity|History of Present Illness|1111,1117|false|false|false|C0595998;C4520849;C4551704|Alive;Household composition;Living|living
Finding|Finding|History of Present Illness|1111,1117|false|false|false|C0595998;C4520849;C4551704|Alive;Household composition;Living|living
Finding|Intellectual Product|History of Present Illness|1119,1127|false|false|false|C4695111|ADMIN.FACILITY|facility
Finding|Idea or Concept|History of Present Illness|1148,1157|false|false|false|C1546960|Patient Outcome - Worsening|worsening
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|1166,1174|false|false|false|C0011265;C0497327|Dementia;Presenile dementia|dementia
Finding|Functional Concept|History of Present Illness|1221,1227|false|false|false|C0728831|Social|social
Finding|Intellectual Product|History of Present Illness|1259,1264|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Sign or Symptom|History of Present Illness|1265,1268|false|false|false|C0013404|Dyspnea|SOB
Finding|Daily or Recreational Activity|History of Present Illness|1274,1284|false|false|false|C0080331;C0945826|Ambulation;Walking (function)|ambulation
Finding|Functional Concept|History of Present Illness|1274,1284|false|false|false|C0080331;C0945826|Ambulation;Walking (function)|ambulation
Procedure|Health Care Activity|History of Present Illness|1296,1305|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Disorder|Disease or Syndrome|History of Present Illness|1343,1347|false|false|false|C0004238|Atrial Fibrillation|Afib
Lab|Laboratory or Test Result|History of Present Illness|1343,1347|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Afib
Finding|Intellectual Product|History of Present Illness|1359,1363|false|false|false|C1561540|Transaction counts and value totals - week|week
Finding|Idea or Concept|History of Present Illness|1369,1377|false|false|false|C1547192|Organization unit type - Hospital|hospital
Anatomy|Body Space or Junction|History of Present Illness|1402,1405|false|false|false|C0228479|Structure of intraculminate fissure|ICU
Finding|Intellectual Product|History of Present Illness|1402,1405|false|false|false|C4554035|Inventory of Callous-Unemotional Traits|ICU
Finding|Functional Concept|History of Present Illness|1420,1428|false|false|false|C0700624|Allergic|allergic
Finding|Pathologic Function|History of Present Illness|1420,1437|false|false|false|C0020517;C1527304|Allergic Reaction;Hypersensitivity|allergic reaction
Finding|Functional Concept|History of Present Illness|1429,1437|false|false|false|C0443286|Reaction|reaction
Drug|Pharmacologic Substance|History of Present Illness|1443,1453|false|false|false|C0013227|Pharmaceutical Preparations|medication
Finding|Intellectual Product|History of Present Illness|1443,1453|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Finding|Classification|History of Present Illness|1455,1461|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|History of Present Illness|1455,1461|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|History of Present Illness|1455,1461|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|History of Present Illness|1455,1461|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Drug|Organic Chemical|History of Present Illness|1470,1476|false|false|false|C0206046|Zofran|Zofran
Drug|Pharmacologic Substance|History of Present Illness|1470,1476|false|false|false|C0206046|Zofran|Zofran
Procedure|Health Care Activity|History of Present Illness|1505,1520|false|false|false|C0019993|Hospitalization|hospitalization
Drug|Biomedical or Dental Material|History of Present Illness|1548,1556|false|false|false|C0168634|BaseLine dental cement|baseline
Finding|Idea or Concept|History of Present Illness|1548,1556|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Finding|Finding|History of Present Illness|1594,1598|false|false|false|C4281574|Much|much
Finding|Finding|History of Present Illness|1606,1610|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|History of Present Illness|1606,1610|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|History of Present Illness|1606,1610|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Finding|History of Present Illness|1611,1621|false|false|false|C2135586;C4321408|Wheelchair Usually Used;has wheelchair at home (history)|wheelchair
Finding|Finding|History of Present Illness|1611,1627|false|false|false|C0558195|Wheelchair bound|wheelchair bound
Event|Activity|History of Present Illness|1622,1627|false|false|false|C1145667|Binding action|bound
Finding|Conceptual Entity|History of Present Illness|1622,1627|false|false|false|C2349209;C2825311|Bound (value);XML Bound|bound
Finding|Finding|History of Present Illness|1669,1675|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Finding|Intellectual Product|History of Present Illness|1669,1675|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Finding|Mental Process|History of Present Illness|1669,1675|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Finding|Mental Process|History of Present Illness|1669,1684|false|false|false|C0025260|Memory|memory function
Finding|Finding|History of Present Illness|1676,1684|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|History of Present Illness|1676,1684|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|History of Present Illness|1676,1684|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|History of Present Illness|1676,1684|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Finding|History of Present Illness|1695,1701|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|History of Present Illness|1695,1701|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Idea or Concept|History of Present Illness|1708,1712|false|false|false|C0233324;C1705313|Term (lexical);Term Birth|term
Finding|Organism Function|History of Present Illness|1708,1712|false|false|false|C0233324;C1705313|Term (lexical);Term Birth|term
Finding|Finding|History of Present Illness|1714,1720|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Finding|Intellectual Product|History of Present Illness|1714,1720|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Finding|Mental Process|History of Present Illness|1714,1720|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|1714,1725|false|false|false|C0002622|Amnesia|memory loss
Finding|Sign or Symptom|History of Present Illness|1714,1725|false|false|false|C0751295|Memory Loss|memory loss
Finding|Finding|History of Present Illness|1721,1725|false|false|false|C5890125|Loss (adaptation)|loss
Finding|Sign or Symptom|History of Present Illness|1727,1745|false|false|false|C0232462|Decrease in appetite|Decreased appetite
Finding|Organism Function|History of Present Illness|1737,1745|false|false|false|C0003618|Desire for food|appetite
Finding|Functional Concept|History of Present Illness|1753,1759|false|false|false|C1512806|Intake|intake
Procedure|Health Care Activity|History of Present Illness|1753,1759|false|false|false|C3251814;C4521161|Intake (treatment);Measurement of fluid intake|intake
Finding|Finding|History of Present Illness|1809,1812|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|History of Present Illness|1809,1812|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Finding|History of Present Illness|1809,1822|false|false|false|C2585997|New diagnosis (finding)|new diagnosis
Procedure|Diagnostic Procedure|History of Present Illness|1809,1822|false|false|false|C1882082|New Diagnosis Procedure|new diagnosis
Attribute|Clinical Attribute|History of Present Illness|1813,1822|false|false|false|C0945731||diagnosis
Finding|Classification|History of Present Illness|1813,1822|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Finding|Functional Concept|History of Present Illness|1813,1822|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Procedure|Diagnostic Procedure|History of Present Illness|1813,1822|false|false|false|C0011900|Diagnosis|diagnosis
Anatomy|Body Space or Junction|History of Present Illness|1826,1829|false|false|false|C0262212|Choroidal fissure|CHF
Disorder|Disease or Syndrome|History of Present Illness|1826,1829|false|false|false|C0018802|Congestive heart failure|CHF
Procedure|Diagnostic Procedure|History of Present Illness|1849,1852|false|false|false|C0430462|Transthoracic echocardiography|TTE
Finding|Organ or Tissue Function|History of Present Illness|1891,1899|false|false|false|C0039155|Systole|systolic
Finding|Finding|History of Present Illness|1900,1908|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|History of Present Illness|1900,1908|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|History of Present Illness|1900,1908|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|History of Present Illness|1900,1908|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Idea or Concept|History of Present Illness|1924,1931|false|false|false|C1555582|Initial (abbreviation)|initial
Finding|Functional Concept|History of Present Illness|1978,1982|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|History of Present Illness|1978,1982|false|false|false|C0582103|Medical Examination|Exam
Finding|Idea or Concept|History of Present Illness|1987,1998|false|false|false|C0750502|Significant|significant
Anatomy|Body Location or Region|History of Present Illness|2005,2010|false|false|false|C0524470|Right hip region structure|R hip
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2007,2010|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|hip
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|2007,2010|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Biologically Active Substance|History of Present Illness|2007,2010|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Pharmacologic Substance|History of Present Illness|2007,2010|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Finding|Gene or Genome|History of Present Illness|2007,2010|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|hip
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|2007,2010|false|false|false|C1292890|Procedure on hip|hip
Disorder|Disease or Syndrome|History of Present Illness|2011,2014|false|false|false|C0034155;C1268935|Congenital Thrombotic Thrombocytopenic Purpura;Purpura, Thrombotic Thrombocytopenic|TTP
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|2011,2014|false|false|false|C1506603;C4723973|ZFP36 protein, human;thiamine triphosphorate|TTP
Drug|Biologically Active Substance|History of Present Illness|2011,2014|false|false|false|C1506603;C4723973|ZFP36 protein, human;thiamine triphosphorate|TTP
Drug|Organic Chemical|History of Present Illness|2011,2014|false|false|false|C1506603;C4723973|ZFP36 protein, human;thiamine triphosphorate|TTP
Drug|Vitamin|History of Present Illness|2011,2014|false|false|false|C1506603;C4723973|ZFP36 protein, human;thiamine triphosphorate|TTP
Finding|Gene or Genome|History of Present Illness|2011,2014|false|false|false|C1413036;C1421571;C3539814|ADAMTS13 gene;ZFP36 gene;ZFP36 wt Allele|TTP
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2015,2033|false|false|false|C0223865|Structure of greater trochanter of femur|greater trochanter
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2023,2033|false|false|false|C0162370|Trochanter|trochanter
Finding|Finding|History of Present Illness|2035,2038|false|false|false|C5848551|Neg - answer|neg
Finding|Social Behavior|History of Present Illness|2039,2047|false|false|false|C0019421|Heterosexuality|straight
Finding|Finding|History of Present Illness|2039,2057|false|true|false|C0422926|Straight leg raise test response|straight leg raise
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2048,2051|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Drug|Food|History of Present Illness|2064,2070|false|false|false|C5890763||pulses
Finding|Physiologic Function|History of Present Illness|2064,2070|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|History of Present Illness|2064,2070|false|false|false|C0034107|Pulse taking|pulses
Attribute|Clinical Attribute|History of Present Illness|2081,2086|false|true|false|C1717255||edema
Finding|Pathologic Function|History of Present Illness|2081,2086|false|true|false|C0013604|Edema|edema
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|2088,2095|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Immunologic Factor|History of Present Illness|2088,2095|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Pharmacologic Substance|History of Present Illness|2088,2095|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Finding|Finding|History of Present Illness|2088,2095|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Functional Concept|History of Present Illness|2088,2095|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Idea or Concept|History of Present Illness|2088,2095|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Intellectual Product|History of Present Illness|2088,2095|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Drug|Pharmacologic Substance|History of Present Illness|2096,2104|false|false|false|C0720099|Duration brand of oxymetazoline|duration
Lab|Laboratory or Test Result|History of Present Illness|2105,2109|false|false|false|C0587081|Laboratory test finding|Labs
Finding|Idea or Concept|History of Present Illness|2115,2126|false|false|false|C0750502|Significant|significant
Anatomy|Cell Component|History of Present Illness|2148,2151|false|false|false|C2263086|Nuclear cap binding complex location|CBC
Procedure|Laboratory Procedure|History of Present Illness|2148,2151|false|false|false|C0009555|Complete Blood Count|CBC
Anatomy|Cell|History of Present Illness|2176,2179|false|false|false|C0023516|Leukocytes|WBC
Finding|Finding|History of Present Illness|2184,2192|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|History of Present Illness|2184,2192|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Classification|History of Present Illness|2200,2208|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|History of Present Illness|2200,2208|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|History of Present Illness|2200,2208|false|false|false|C5237010|Expression Negative|negative
Drug|Biologically Active Substance|History of Present Illness|2209,2217|false|false|false|C0028137|Nitrites|nitrites
Drug|Inorganic Chemical|History of Present Illness|2209,2217|false|false|false|C0028137|Nitrites|nitrites
Drug|Pharmacologic Substance|History of Present Illness|2209,2217|false|false|false|C0028137|Nitrites|nitrites
Procedure|Research Activity|History of Present Illness|2220,2227|false|false|false|C0947630|Scientific Study|Studies
Anatomy|Body Location or Region|History of Present Illness|2230,2235|false|false|false|C1548802|Body Site Modifier - Lower|Lower
Event|Activity|History of Present Illness|2230,2235|false|false|false|C2003888|Lower (action)|Lower
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2230,2245|false|false|false|C0023216|Lower Extremity|Lower extremity
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2236,2245|false|false|false|C0015385|Limb structure|extremity
Finding|Functional Concept|History of Present Illness|2246,2256|false|false|false|C0220934|Ultrasonic|ultrasound
Phenomenon|Natural Phenomenon or Process|History of Present Illness|2246,2256|false|false|false|C0041621;C1456803|Ultrasonic Shockwave;Ultrasonics (sound)|ultrasound
Procedure|Diagnostic Procedure|History of Present Illness|2246,2256|false|false|false|C0041618;C1315081|Ultrasonography;Urological ultrasound|ultrasound
Attribute|Clinical Attribute|History of Present Illness|2261,2265|false|false|false|C4318566|Deep Resection Margin|Deep
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2261,2270|false|false|false|C0226514|Structure of deep vein|Deep vein
Disorder|Disease or Syndrome|History of Present Illness|2261,2281|false|false|false|C0149871;C0340708|Deep Vein Thrombosis;Deep vein thrombosis of lower limb|Deep vein thrombosis
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2266,2270|false|false|false|C0042449|Veins|vein
Finding|Pathologic Function|History of Present Illness|2266,2281|false|false|false|C0042487|Venous Thrombosis|vein thrombosis
Finding|Pathologic Function|History of Present Illness|2271,2281|false|false|false|C0040053|Thrombosis|thrombosis
Finding|Functional Concept|History of Present Illness|2289,2293|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Finding|Functional Concept|History of Present Illness|2295,2301|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Finding|Intellectual Product|History of Present Illness|2295,2301|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2295,2314|false|false|false|C1275667|Common femoral vein|common femoral vein
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2302,2309|false|false|false|C0015811|Femur|femoral
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2302,2314|false|false|false|C0015809|Femoral vein|femoral vein
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2310,2314|false|false|false|C0042449|Veins|vein
Anatomy|Body Location or Region|History of Present Illness|2343,2352|false|false|false|C0442037|popliteal|popliteal
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2343,2357|false|false|false|C0032652|Structure of popliteal vein|popliteal vein
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2353,2357|false|false|false|C0042449|Veins|vein
Finding|Functional Concept|History of Present Illness|2360,2364|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Location or Region|History of Present Illness|2360,2369|false|false|false|C0489800|Posterior part of left leg|Left calf
Anatomy|Body Location or Region|History of Present Illness|2365,2369|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2365,2369|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2370,2375|false|false|false|C0042449|Veins|veins
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|2370,2375|false|false|false|C0398102|Procedure on vein|veins
Finding|Finding|History of Present Illness|2408,2416|false|false|false|C0332149|Possible|possibly
Finding|Finding|History of Present Illness|2423,2431|false|false|false|C0028778;C1947917|Obstruction;Occluded|occluded
Finding|Functional Concept|History of Present Illness|2423,2431|false|false|false|C0028778;C1947917|Obstruction;Occluded|occluded
Anatomy|Body Location or Region|History of Present Illness|2439,2442|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|History of Present Illness|2439,2442|true|false|false|C2926618||DVT
Disorder|Disease or Syndrome|History of Present Illness|2439,2442|true|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Finding|Functional Concept|History of Present Illness|2450,2455|true|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2450,2471|false|false|false|C0230415|Right lower extremity|right lower extremity
Anatomy|Body Location or Region|History of Present Illness|2456,2461|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|History of Present Illness|2456,2461|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2456,2471|false|false|false|C0023216|Lower Extremity|lower extremity
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2462,2471|false|false|false|C0015385|Limb structure|extremity
Procedure|Diagnostic Procedure|History of Present Illness|2474,2477|false|false|false|C0039985|Plain chest X-ray|CXR
Anatomy|Tissue|History of Present Illness|2488,2495|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|History of Present Illness|2488,2495|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Pathologic Function|History of Present Illness|2488,2505|false|false|false|C0032227|Pleural effusion (disorder)|pleural effusions
Finding|Pathologic Function|History of Present Illness|2496,2505|false|false|false|C0013687|effusion|effusions
Finding|Gene or Genome|History of Present Illness|2507,2512|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Finding|Functional Concept|History of Present Illness|2520,2525|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Finding|Functional Concept|History of Present Illness|2544,2548|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Disorder|Disease or Syndrome|History of Present Illness|2568,2581|true|false|false|C0521530|Lung consolidation|consolidation
Finding|Idea or Concept|History of Present Illness|2604,2614|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|History of Present Illness|2604,2614|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Disorder|Neoplastic Process|History of Present Illness|2626,2635|false|false|false|C0027627|Neoplasm Metastasis|secondary
Finding|Functional Concept|History of Present Illness|2626,2635|false|false|false|C1522484|metastatic qualifier|secondary
Finding|Pathologic Function|History of Present Illness|2645,2654|false|false|false|C0013687|effusion|effusions
Drug|Organic Chemical|History of Present Illness|2693,2703|false|false|false|C0206460|enoxaparin|Enoxaparin
Drug|Pharmacologic Substance|History of Present Illness|2693,2703|false|false|false|C0206460|enoxaparin|Enoxaparin
Drug|Organic Chemical|History of Present Illness|2693,2710|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Pharmacologic Substance|History of Present Illness|2693,2710|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Biologically Active Substance|History of Present Illness|2704,2710|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|History of Present Illness|2704,2710|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|History of Present Illness|2704,2710|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Finding|Physiologic Function|History of Present Illness|2704,2710|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|History of Present Illness|2704,2710|false|false|false|C0337443|Sodium measurement|Sodium
Finding|Functional Concept|History of Present Illness|2726,2734|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|History of Present Illness|2726,2734|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|History of Present Illness|2726,2734|false|false|false|C4706767|Transfer (immobility management)|transfer
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2768,2773|false|false|false|C0028429||Nasal
Drug|Biomedical or Dental Material|History of Present Illness|2768,2773|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Organic Chemical|History of Present Illness|2768,2773|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Pharmacologic Substance|History of Present Illness|2768,2773|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Finding|Finding|History of Present Illness|2768,2773|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Finding|Functional Concept|History of Present Illness|2768,2773|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2775,2782|false|false|false|C1550232|Body Parts - Cannula|Cannula
Finding|Body Substance|History of Present Illness|2775,2782|false|false|false|C1546577;C1550622|Specimen Type - Cannula|Cannula
Finding|Intellectual Product|History of Present Illness|2775,2782|false|false|false|C1546577;C1550622|Specimen Type - Cannula|Cannula
Anatomy|Anatomical Structure|History of Present Illness|2794,2799|false|false|false|C3714591|Floor (anatomic)|floor
Disorder|Disease or Syndrome|History of Present Illness|2831,2834|false|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Finding|Intellectual Product|History of Present Illness|2831,2834|false|false|false|C2346952|Bachelor of Education|bed
Finding|Conceptual Entity|History of Present Illness|2836,2843|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|History of Present Illness|2836,2843|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|History of Present Illness|2836,2843|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Idea or Concept|History of Present Illness|2860,2865|false|false|false|C1552828|Table Frame - above|above
Finding|Classification|History of Present Illness|2871,2877|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|History of Present Illness|2871,2877|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|History of Present Illness|2871,2877|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|History of Present Illness|2871,2877|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Finding|History of Present Illness|2914,2921|false|false|false|C4534363|At home|at home
Finding|Idea or Concept|History of Present Illness|2917,2921|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|History of Present Illness|2917,2921|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|History of Present Illness|2917,2921|false|false|false|C1553498|home health encounter|home
Finding|Sign or Symptom|History of Present Illness|2930,2933|false|false|false|C0231807|Dyspnea on exertion|DOE
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2953,2958|false|false|false|C0021853|Intestines|bowel
Finding|Organism Function|History of Present Illness|2953,2967|true|false|false|C0011135|Defecation|bowel movement
Finding|Organism Function|History of Present Illness|2959,2967|false|false|false|C0026649|Movement|movement
Finding|Idea or Concept|History of Present Illness|2982,2988|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|Review
Finding|Intellectual Product|History of Present Illness|2982,2988|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|Review
Finding|Functional Concept|History of Present Illness|2982,2991|false|false|false|C0699752|Review of|Review of
Attribute|Clinical Attribute|History of Present Illness|2982,2999|false|false|false|C0488564;C0488565||Review of systems
Procedure|Health Care Activity|History of Present Illness|2982,2999|false|false|false|C0489633|Review of systems (procedure)|Review of systems
Finding|Functional Concept|History of Present Illness|2992,2999|false|false|false|C0449913|System|systems
Disorder|Disease or Syndrome|History of Present Illness|3011,3014|false|false|false|C0268529|Proline dehydrogenase deficiency|HPI
Finding|Finding|History of Present Illness|3011,3014|false|false|false|C0262512;C1323983|History of present illness (finding);allene oxide synthase activity|HPI
Finding|Molecular Function|History of Present Illness|3011,3014|false|false|false|C0262512;C1323983|History of present illness (finding);allene oxide synthase activity|HPI
Finding|Finding|History of Present Illness|3028,3033|true|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|History of Present Illness|3028,3033|true|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|History of Present Illness|3035,3041|true|false|false|C0085593|Chills|chills
Finding|Sign or Symptom|History of Present Illness|3043,3055|true|false|false|C0028081|Night sweats|night sweats
Finding|Body Substance|History of Present Illness|3049,3055|true|false|false|C0038984;C0038990|Sweat;Sweating|sweats
Finding|Finding|History of Present Illness|3049,3055|true|false|false|C0038984;C0038990|Sweat;Sweating|sweats
Finding|Sign or Symptom|History of Present Illness|3064,3072|true|false|false|C0018681|Headache|headache
Anatomy|Body Space or Junction|History of Present Illness|3074,3079|false|false|false|C0030471;C1305231|Nasal sinus;Sinus - general anatomical term|sinus
Disorder|Anatomical Abnormality|History of Present Illness|3074,3079|true|false|false|C0016169|pathologic fistula|sinus
Drug|Organic Chemical|History of Present Illness|3074,3079|true|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Drug|Pharmacologic Substance|History of Present Illness|3074,3079|true|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Finding|Mental Process|History of Present Illness|3081,3091|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|History of Present Illness|3081,3091|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|History of Present Illness|3093,3103|false|false|false|C1260880|Rhinorrhea|rhinorrhea
Finding|Pathologic Function|History of Present Illness|3107,3117|false|false|false|C0700148|Congestion|congestion
Drug|Organic Chemical|History of Present Illness|3126,3131|true|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|History of Present Illness|3126,3131|true|false|false|C3815497|Cough (guaifenesin)|cough
Finding|Sign or Symptom|History of Present Illness|3126,3131|true|false|false|C0010200|Coughing|cough
Attribute|Clinical Attribute|History of Present Illness|3141,3147|false|false|false|C4255480||nausea
Finding|Sign or Symptom|History of Present Illness|3141,3147|false|false|false|C0027497|Nausea|nausea
Finding|Sign or Symptom|History of Present Illness|3149,3157|false|false|false|C0042963|Vomiting|vomiting
Finding|Finding|History of Present Illness|3159,3167|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|History of Present Illness|3159,3167|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|History of Present Illness|3169,3181|false|false|false|C0009806|Constipation|constipation
Anatomy|Body Location or Region|History of Present Illness|3185,3194|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|History of Present Illness|3185,3199|false|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|History of Present Illness|3195,3199|false|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|3195,3199|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|3195,3199|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|3205,3212|false|false|false|C0013428|Dysuria|dysuria
Finding|Sign or Symptom|History of Present Illness|3221,3232|true|false|false|C0003862|Arthralgia|arthralgias
Finding|Sign or Symptom|History of Present Illness|3236,3244|true|false|false|C0231528|Myalgia|myalgias
Disorder|Disease or Syndrome|Past Medical History|3273,3285|false|false|false|C0020538|Hypertensive disease|Hypertension
Disorder|Mental or Behavioral Dysfunction|Past Medical History|3286,3294|false|false|false|C0011265;C0497327|Dementia;Presenile dementia|Dementia
Disorder|Disease or Syndrome|Past Medical History|3295,3307|false|false|false|C0029456|Osteoporosis|Osteoporosis
Finding|Finding|Past Medical History|3295,3307|false|false|false|C2911643|Encounter due to family history of osteoporosis|Osteoporosis
Finding|Finding|Past Medical History|3308,3317|false|false|false|C0022107;C2700617|Irritability - emotion;Irritable Mood|Irritable
Finding|Mental Process|Past Medical History|3308,3317|false|false|false|C0022107;C2700617|Irritability - emotion;Irritable Mood|Irritable
Disorder|Disease or Syndrome|Past Medical History|3308,3323|false|false|false|C0022104|Irritable Bowel Syndrome|Irritable bowel
Disorder|Disease or Syndrome|Past Medical History|3308,3332|false|false|false|C0022104|Irritable Bowel Syndrome|Irritable bowel syndrome
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|3318,3323|false|false|false|C0021853|Intestines|bowel
Disorder|Disease or Syndrome|Past Medical History|3324,3332|false|false|false|C0039082|Syndrome|syndrome
Disorder|Cell or Molecular Dysfunction|Past Medical History|3333,3345|false|false|false|C0085662;C2004480|Macrocytosis;Macrocytosis (morphologic abnormality)|Macrocytosis
Disorder|Disease or Syndrome|Past Medical History|3333,3345|false|false|false|C0085662;C2004480|Macrocytosis;Macrocytosis (morphologic abnormality)|Macrocytosis
Lab|Laboratory or Test Result|Past Medical History|3333,3345|false|false|false|C0684332|Macrocytosis (finding)|Macrocytosis
Finding|Conceptual Entity|Past Medical History|3357,3365|false|false|false|C0015127;C1314792;C1524003|Etiology;Etiology aspects;Science of Etiology|etiology
Finding|Functional Concept|Past Medical History|3357,3365|false|false|false|C0015127;C1314792;C1524003|Etiology;Etiology aspects;Science of Etiology|etiology
Finding|Functional Concept|Past Medical History|3366,3370|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|3366,3374|false|false|false|C0229299|Left ear structure|Left ear
Finding|Sign or Symptom|Past Medical History|3366,3374|false|false|false|C2127178|left ear symptoms (symptom)|Left ear
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|3371,3374|false|false|false|C0013443;C0521421|Ear structure|ear
Disorder|Disease or Syndrome|Past Medical History|3371,3374|false|false|false|C0851354|Ear and labyrinth disorders|ear
Finding|Body Substance|Past Medical History|3371,3374|false|false|false|C1546608;C1550629|SpecimenType - Ear|ear
Finding|Intellectual Product|Past Medical History|3371,3374|false|false|false|C1546608;C1550629|SpecimenType - Ear|ear
Finding|Finding|Past Medical History|3375,3382|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|hearing
Finding|Physiologic Function|Past Medical History|3375,3382|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|hearing
Disorder|Disease or Syndrome|Past Medical History|3375,3387|false|false|false|C1384666|hearing impairment|hearing loss
Finding|Finding|Past Medical History|3375,3387|false|false|false|C0011053;C0018772;C2029884;C3887873|Deafness;Hearing Loss;Partial Hearing Loss;hearing loss by exam|hearing loss
Finding|Finding|Past Medical History|3383,3387|false|false|false|C5890125|Loss (adaptation)|loss
Attribute|Clinical Attribute|Past Medical History|3388,3394|false|false|false|C5889824||Status
Finding|Idea or Concept|Past Medical History|3388,3394|false|false|false|C1546481|What subject filter - Status|Status
Finding|Finding|Past Medical History|3400,3412|false|false|false|C1548863|Consent Type - Hysterectomy|hysterectomy
Procedure|Therapeutic or Preventive Procedure|Past Medical History|3400,3412|false|false|false|C0020699|Hysterectomy|hysterectomy
Attribute|Clinical Attribute|Past Medical History|3413,3419|false|false|false|C5889824||Status
Finding|Idea or Concept|Past Medical History|3413,3419|false|false|false|C1546481|What subject filter - Status|Status
Procedure|Therapeutic or Preventive Procedure|Past Medical History|3425,3437|false|false|false|C0003611;C0003612|Appendectomy;Appendectomy; for ruptured appendix with abscess or generalized peritonitis|appendectomy
Attribute|Clinical Attribute|Past Medical History|3438,3444|false|false|false|C5889824||Status
Finding|Idea or Concept|Past Medical History|3438,3444|false|false|false|C1546481|What subject filter - Status|Status
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|3450,3457|false|false|false|C0205065|Ovarian|ovarian
Disorder|Disease or Syndrome|Past Medical History|3450,3462|false|false|false|C0029927|Ovarian Cysts|ovarian cyst
Procedure|Therapeutic or Preventive Procedure|Past Medical History|3450,3470|false|false|false|C0195488|Removal of ovarian cyst|ovarian cyst removal
Disorder|Anatomical Abnormality|Past Medical History|3458,3462|false|false|false|C0010709|Cyst|cyst
Finding|Body Substance|Past Medical History|3458,3462|false|false|false|C1546594;C1550626|SpecimenType - Cyst|cyst
Finding|Intellectual Product|Past Medical History|3458,3462|false|false|false|C1546594;C1550626|SpecimenType - Cyst|cyst
Procedure|Therapeutic or Preventive Procedure|Past Medical History|3458,3470|false|false|false|C0742962|Cyst removal|cyst removal
Event|Activity|Past Medical History|3463,3470|false|false|false|C1883720|Removing (action)|removal
Procedure|Therapeutic or Preventive Procedure|Past Medical History|3463,3470|false|false|false|C0015252;C0185115;C0728940|Excision;Extraction;removal technique|removal
Disorder|Disease or Syndrome|Past Medical History|3471,3479|false|false|false|C0086543|Cataract|Cataract
Finding|Finding|Past Medical History|3471,3479|false|false|false|C1690964|cataract on exam (physical finding)|Cataract
Finding|Finding|Past Medical History|3471,3487|false|false|false|C1548833;C2186377|Consent Type - Cataract Surgery;reported history of cataract surgery|Cataract surgery
Finding|Intellectual Product|Past Medical History|3471,3487|false|false|false|C1548833;C2186377|Consent Type - Cataract Surgery;reported history of cataract surgery|Cataract surgery
Procedure|Therapeutic or Preventive Procedure|Past Medical History|3471,3487|false|false|false|C0007389;C2939459|Cataract Extraction;Cataract surgery|Cataract surgery
Finding|Finding|Past Medical History|3480,3487|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|Past Medical History|3480,3487|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|Past Medical History|3480,3487|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|Past Medical History|3480,3487|false|false|false|C0543467|Operative Surgical Procedures|surgery
Disorder|Disease or Syndrome|Past Medical History|3488,3496|false|false|false|C0017601|Glaucoma|Glaucoma
Phenomenon|Natural Phenomenon or Process|Family Medical History|3555,3562|false|false|false|C1705970|Electrical Current|current
Procedure|Health Care Activity|Family Medical History|3563,3572|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Procedure|Health Care Activity|General Exam|3591,3600|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Finding|Functional Concept|General Exam|3601,3605|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|General Exam|3601,3605|false|false|false|C0582103|Medical Examination|EXAM
Drug|Food|General Exam|3622,3627|false|false|false|C1875856|Vital High Nitrogen Enteral Nutrition|Vital
Attribute|Clinical Attribute|General Exam|3622,3633|false|false|false|C0488614;C0518766|Vital signs|Vital Signs
Procedure|Health Care Activity|General Exam|3622,3633|false|false|false|C0150404|Taking vital signs|Vital Signs
Finding|Finding|General Exam|3628,3633|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|Signs
Finding|Functional Concept|General Exam|3628,3633|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|Signs
Finding|Classification|General Exam|3668,3675|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|General Exam|3668,3675|false|false|false|C3812897|General medical service|General
Finding|Gene or Genome|General Exam|3677,3681|false|false|false|C1412433|AOX1 gene|AOx1
Finding|Mental Process|General Exam|3683,3691|false|false|false|C2987187|Pleasant|pleasant
Finding|Social Behavior|General Exam|3693,3700|false|false|false|C0037363|Smiling|smiling
Drug|Biomedical or Dental Material|General Exam|3705,3713|false|false|false|C0168634|BaseLine dental cement|baseline
Finding|Idea or Concept|General Exam|3705,3713|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Finding|Classification|General Exam|3718,3724|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|General Exam|3718,3724|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|General Exam|3718,3724|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|General Exam|3718,3724|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Anatomy|Body Part, Organ, or Organ Component|General Exam|3751,3757|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|General Exam|3751,3757|false|false|false|C0036412|Scleral Diseases|Sclera
Procedure|Health Care Activity|General Exam|3751,3757|false|false|false|C2228481|examination of sclera|Sclera
Finding|Finding|General Exam|3758,3767|false|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Part, Organ, or Organ Component|General Exam|3769,3772|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|General Exam|3769,3772|false|false|false|C0026987|Myelofibrosis|MMM
Anatomy|Body Location or Region|General Exam|3774,3784|false|false|false|C0521367|Oropharyngeal|oropharynx
Finding|Idea or Concept|General Exam|3785,3790|false|false|false|C1550016|Remote control command - Clear|clear
Finding|Finding|General Exam|3798,3803|false|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Anatomy|Body Location or Region|General Exam|3806,3810|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|General Exam|3806,3810|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|General Exam|3806,3810|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Finding|Finding|General Exam|3806,3817|false|false|false|C2230237|Supple neck|neck supple
Finding|Functional Concept|General Exam|3811,3817|false|false|false|C0332254|Supple|supple
Finding|Finding|General Exam|3819,3822|false|false|false|C0428897|Jugular venous pressure|JVP
Anatomy|Body Part, Organ, or Organ Component|General Exam|3840,3843|true|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|General Exam|3840,3843|true|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Finding|Gene or Genome|General Exam|3840,3843|true|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Event|Activity|General Exam|3858,3862|false|false|false|C0871208|Rating (action)|rate
Finding|Idea or Concept|General Exam|3858,3862|false|false|false|C1549480|Amount type - Rate|rate
Finding|Finding|General Exam|3867,3873|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|General Exam|3867,3873|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Disorder|Disease or Syndrome|General Exam|3891,3895|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Finding|Organ or Tissue Function|General Exam|3900,3908|false|false|false|C0039155|Systole|systolic
Finding|Finding|General Exam|3910,3916|false|false|false|C0018808|Heart murmur|murmur
Anatomy|Body Part, Organ, or Organ Component|General Exam|3921,3926|false|false|false|C0024109|Lung|Lungs
Finding|Finding|General Exam|3928,3936|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Intellectual Product|General Exam|3928,3936|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Organism Function|General Exam|3937,3948|false|false|false|C0004048|Inspiration (function)|inspiratory
Finding|Organism Function|General Exam|3949,3955|false|false|false|C0015264|Exertion|effort
Finding|Finding|General Exam|3957,3980|false|false|false|C0238844|Decreased breath sounds|decreased breath sounds
Finding|Body Substance|General Exam|3967,3973|false|false|false|C0225386|Breath|breath
Attribute|Clinical Attribute|General Exam|3967,3980|false|false|false|C0035234;C3484186|Respiratory Sounds|breath sounds
Phenomenon|Natural Phenomenon or Process|General Exam|3974,3980|false|false|false|C0037709||sounds
Drug|Chemical Viewed Functionally|General Exam|3997,4002|false|false|false|C0178499|Base|bases
Finding|Sign or Symptom|General Exam|4011,4018|true|false|false|C0043144|Wheezing|wheezes
Finding|Finding|General Exam|4020,4025|true|false|false|C0034642;C0240859|Basilar Rales;Rales|rales
Finding|Finding|General Exam|4027,4034|true|false|false|C0035508|Rhonchi|rhonchi
Anatomy|Body Location or Region|General Exam|4037,4044|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|General Exam|4037,4044|false|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Finding|Finding|General Exam|4037,4044|false|false|false|C0941288|Abdomen problem|Abdomen
Disorder|Disease or Syndrome|General Exam|4046,4050|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Anatomy|Body Part, Organ, or Organ Component|General Exam|4079,4084|false|false|false|C0021853|Intestines|bowel
Finding|Finding|General Exam|4079,4091|false|false|false|C0232693|Bowel sounds|bowel sounds
Phenomenon|Natural Phenomenon or Process|General Exam|4085,4091|false|false|false|C0037709||sounds
Finding|Finding|General Exam|4092,4099|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|General Exam|4092,4099|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Finding|General Exam|4105,4117|true|false|false|C4054315|Organomegaly|organomegaly
Finding|Finding|General Exam|4133,4141|true|false|false|C0427198|Protective muscle spasm|guarding
Disorder|Congenital Abnormality|General Exam|4159,4162|false|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Finding|Gene or Genome|General Exam|4159,4162|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Finding|Finding|General Exam|4164,4168|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|General Exam|4164,4168|false|false|false|C0687712|warming process|Warm
Finding|Finding|General Exam|4170,4174|false|false|false|C5575035|Well (answer to question)|well
Drug|Food|General Exam|4188,4194|false|false|false|C5890763||pulses
Finding|Physiologic Function|General Exam|4188,4194|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|General Exam|4188,4194|false|false|false|C0034107|Pulse taking|pulses
Anatomy|Body Location or Region|General Exam|4200,4205|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|General Exam|4200,4205|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|General Exam|4200,4215|false|false|false|C0023216|Lower Extremity|lower extremity
Anatomy|Body Part, Organ, or Organ Component|General Exam|4206,4215|false|false|false|C0015385|Limb structure|extremity
Finding|Finding|General Exam|4217,4225|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|General Exam|4217,4225|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Functional Concept|General Exam|4231,4235|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|General Exam|4231,4239|false|false|false|C0230416;C0230443|Left lower extremity;Structure of left lower leg|left leg
Anatomy|Body Part, Organ, or Organ Component|General Exam|4236,4239|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Finding|Functional Concept|General Exam|4240,4252|false|false|false|C0332476|erythematous|erythematous
Procedure|Diagnostic Procedure|General Exam|4267,4276|false|false|false|C0030247|Palpation|palpation
Finding|Functional Concept|General Exam|4282,4289|false|false|false|C0205323|Pitting|pitting
Finding|Finding|General Exam|4282,4295|false|false|false|C0333243|Pitting edema|pitting edema
Attribute|Clinical Attribute|General Exam|4290,4295|false|false|false|C1717255||edema
Finding|Pathologic Function|General Exam|4290,4295|false|false|false|C0013604|Edema|edema
Finding|Functional Concept|General Exam|4304,4309|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|General Exam|4304,4325|false|false|false|C0230415|Right lower extremity|right lower extremity
Anatomy|Body Location or Region|General Exam|4310,4315|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|General Exam|4310,4315|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|General Exam|4310,4325|false|false|false|C0023216|Lower Extremity|lower extremity
Anatomy|Body Part, Organ, or Organ Component|General Exam|4316,4325|false|false|false|C0015385|Limb structure|extremity
Finding|Intellectual Product|General Exam|4335,4342|false|true|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|General Exam|4335,4342|false|true|false|C1555457|Provision of recurring care for chronic illness|chronic
Anatomy|Body Part, Organ, or Organ Component|General Exam|4344,4350|false|false|false|C0042449|Veins|venous
Disorder|Disease or Syndrome|General Exam|4344,4357|false|false|false|C0042344|Varicose Ulcer|venous stasis
Finding|Pathologic Function|General Exam|4344,4357|false|false|false|C4551518|Venous stasis|venous stasis
Finding|Pathologic Function|General Exam|4351,4357|false|false|false|C0333138|Stasis|stasis
Finding|Functional Concept|General Exam|4358,4365|false|false|false|C0392747|Changing|changes
Finding|Finding|General Exam|4367,4383|false|false|false|C1720243|1+ pitting edema|1+ pitting edema
Finding|Functional Concept|General Exam|4370,4377|false|false|false|C0205323|Pitting|pitting
Finding|Finding|General Exam|4370,4383|false|false|false|C0333243|Pitting edema|pitting edema
Attribute|Clinical Attribute|General Exam|4378,4383|false|false|false|C1717255||edema
Finding|Pathologic Function|General Exam|4378,4383|false|false|false|C0013604|Edema|edema
Finding|Gene or Genome|General Exam|4405,4409|false|false|false|C1412433|AOX1 gene|AOx1
Finding|Idea or Concept|General Exam|4411,4419|false|false|false|C0808080|Strength (attribute)|strength
Anatomy|Body Location or Region|General Exam|4434,4439|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|General Exam|4434,4439|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Location or Region|General Exam|4459,4465|false|false|false|C0015450|Face|facial
Finding|Organism Function|General Exam|4466,4475|false|false|false|C0026649|Movement|movements
Drug|Amino Acid, Peptide, or Protein|General Exam|4479,4483|false|false|false|C0618927;C5239612|Tact;bis(tetraheptylammonium)tetraiodocyclopentane tellurate(IV)|tact
Drug|Element, Ion, or Isotope|General Exam|4479,4483|false|false|false|C0618927;C5239612|Tact;bis(tetraheptylammonium)tetraiodocyclopentane tellurate(IV)|tact
Drug|Immunologic Factor|General Exam|4479,4483|false|false|false|C0618927;C5239612|Tact;bis(tetraheptylammonium)tetraiodocyclopentane tellurate(IV)|tact
Drug|Pharmacologic Substance|General Exam|4479,4483|false|false|false|C0618927;C5239612|Tact;bis(tetraheptylammonium)tetraiodocyclopentane tellurate(IV)|tact
Finding|Finding|General Exam|4485,4494|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|General Exam|4485,4494|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|General Exam|4485,4494|false|false|false|C2229507|sensory exam|sensation
Drug|Amino Acid, Peptide, or Protein|General Exam|4506,4510|false|false|false|C0618927;C5239612|Tact;bis(tetraheptylammonium)tetraiodocyclopentane tellurate(IV)|tact
Drug|Element, Ion, or Isotope|General Exam|4506,4510|false|false|false|C0618927;C5239612|Tact;bis(tetraheptylammonium)tetraiodocyclopentane tellurate(IV)|tact
Drug|Immunologic Factor|General Exam|4506,4510|false|false|false|C0618927;C5239612|Tact;bis(tetraheptylammonium)tetraiodocyclopentane tellurate(IV)|tact
Drug|Pharmacologic Substance|General Exam|4506,4510|false|false|false|C0618927;C5239612|Tact;bis(tetraheptylammonium)tetraiodocyclopentane tellurate(IV)|tact
Finding|Finding|General Exam|4512,4516|false|false|false|C0016928|Gait|gait
Finding|Body Substance|General Exam|4532,4541|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|General Exam|4532,4541|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|General Exam|4532,4541|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|General Exam|4532,4541|false|false|false|C0030685|Patient Discharge|DISCHARGE
Finding|Functional Concept|General Exam|4542,4546|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|General Exam|4542,4546|false|false|false|C0582103|Medical Examination|EXAM
Finding|Classification|General Exam|4603,4610|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|General Exam|4603,4610|false|false|false|C3812897|General medical service|General
Finding|Gene or Genome|General Exam|4612,4616|false|false|false|C1412433|AOX1 gene|AOx1
Finding|Mental Process|General Exam|4618,4626|false|false|false|C2987187|Pleasant|pleasant
Finding|Social Behavior|General Exam|4628,4635|false|false|false|C0037363|Smiling|smiling
Drug|Biomedical or Dental Material|General Exam|4640,4648|false|false|false|C0168634|BaseLine dental cement|baseline
Finding|Idea or Concept|General Exam|4640,4648|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Finding|Classification|General Exam|4653,4659|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|General Exam|4653,4659|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|General Exam|4653,4659|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|General Exam|4653,4659|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Anatomy|Body Part, Organ, or Organ Component|General Exam|4686,4692|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|General Exam|4686,4692|false|false|false|C0036412|Scleral Diseases|Sclera
Procedure|Health Care Activity|General Exam|4686,4692|false|false|false|C2228481|examination of sclera|Sclera
Finding|Finding|General Exam|4693,4702|false|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Part, Organ, or Organ Component|General Exam|4704,4707|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|General Exam|4704,4707|false|false|false|C0026987|Myelofibrosis|MMM
Disorder|Disease or Syndrome|General Exam|4753,4757|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Finding|Organ or Tissue Function|General Exam|4762,4770|false|false|false|C0039155|Systole|systolic
Finding|Finding|General Exam|4772,4778|false|false|false|C0018808|Heart murmur|murmur
Anatomy|Body Part, Organ, or Organ Component|General Exam|4783,4788|false|false|false|C0024109|Lung|Lungs
Finding|Finding|General Exam|4790,4798|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Intellectual Product|General Exam|4790,4798|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Organism Function|General Exam|4799,4810|false|false|false|C0004048|Inspiration (function)|inspiratory
Finding|Organism Function|General Exam|4811,4817|false|false|false|C0015264|Exertion|effort
Finding|Finding|General Exam|4819,4842|false|false|false|C0238844|Decreased breath sounds|decreased breath sounds
Finding|Body Substance|General Exam|4829,4835|false|false|false|C0225386|Breath|breath
Attribute|Clinical Attribute|General Exam|4829,4842|false|false|false|C0035234;C3484186|Respiratory Sounds|breath sounds
Phenomenon|Natural Phenomenon or Process|General Exam|4836,4842|false|false|false|C0037709||sounds
Drug|Chemical Viewed Functionally|General Exam|4854,4859|false|false|false|C0178499|Base|bases
Disorder|Congenital Abnormality|General Exam|4861,4864|false|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Finding|Gene or Genome|General Exam|4861,4864|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Finding|Finding|General Exam|4866,4870|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|General Exam|4866,4870|false|false|false|C0687712|warming process|Warm
Finding|Finding|General Exam|4872,4876|false|false|false|C5575035|Well (answer to question)|well
Drug|Food|General Exam|4890,4896|false|false|false|C5890763||pulses
Finding|Physiologic Function|General Exam|4890,4896|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|General Exam|4890,4896|false|false|false|C0034107|Pulse taking|pulses
Anatomy|Body Location or Region|General Exam|4902,4907|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|General Exam|4902,4907|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|General Exam|4902,4917|false|false|false|C0023216|Lower Extremity|lower extremity
Anatomy|Body Part, Organ, or Organ Component|General Exam|4908,4917|false|false|false|C0015385|Limb structure|extremity
Finding|Finding|General Exam|4919,4927|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|General Exam|4919,4927|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Functional Concept|General Exam|4933,4937|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|General Exam|4933,4941|false|false|false|C0230416;C0230443|Left lower extremity;Structure of left lower leg|left leg
Anatomy|Body Part, Organ, or Organ Component|General Exam|4938,4941|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Finding|Functional Concept|General Exam|4942,4954|false|false|false|C0332476|erythematous|erythematous
Procedure|Diagnostic Procedure|General Exam|4978,4987|false|false|false|C0030247|Palpation|palpation
Finding|Finding|General Exam|4989,5005|false|false|false|C1720371|2+ pitting edema|2+ pitting edema
Finding|Functional Concept|General Exam|4992,4999|false|false|false|C0205323|Pitting|pitting
Finding|Finding|General Exam|4992,5005|false|false|false|C0333243|Pitting edema|pitting edema
Attribute|Clinical Attribute|General Exam|5000,5005|false|false|false|C1717255||edema
Finding|Pathologic Function|General Exam|5000,5005|false|false|false|C0013604|Edema|edema
Finding|Functional Concept|General Exam|5014,5019|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|General Exam|5014,5035|false|false|false|C0230415|Right lower extremity|right lower extremity
Anatomy|Body Location or Region|General Exam|5020,5025|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|General Exam|5020,5025|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|General Exam|5020,5035|false|false|false|C0023216|Lower Extremity|lower extremity
Anatomy|Body Part, Organ, or Organ Component|General Exam|5026,5035|false|false|false|C0015385|Limb structure|extremity
Finding|Intellectual Product|General Exam|5046,5053|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|General Exam|5046,5053|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Anatomy|Body Part, Organ, or Organ Component|General Exam|5054,5060|false|false|false|C0042449|Veins|venous
Disorder|Disease or Syndrome|General Exam|5054,5067|false|false|false|C0042344|Varicose Ulcer|venous stasis
Finding|Pathologic Function|General Exam|5054,5067|false|false|false|C4551518|Venous stasis|venous stasis
Finding|Pathologic Function|General Exam|5061,5067|false|false|false|C0333138|Stasis|stasis
Finding|Functional Concept|General Exam|5068,5075|false|false|false|C0392747|Changing|changes
Finding|Finding|General Exam|5077,5093|false|false|false|C1720243|1+ pitting edema|1+ pitting edema
Finding|Functional Concept|General Exam|5080,5087|false|false|false|C0205323|Pitting|pitting
Finding|Finding|General Exam|5080,5093|false|false|false|C0333243|Pitting edema|pitting edema
Attribute|Clinical Attribute|General Exam|5088,5093|false|false|false|C1717255||edema
Finding|Pathologic Function|General Exam|5088,5093|false|false|false|C0013604|Edema|edema
Finding|Gene or Genome|General Exam|5116,5120|false|false|false|C1412433|AOX1 gene|AOx1
Procedure|Health Care Activity|General Exam|5145,5154|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Lab|Laboratory or Test Result|General Exam|5155,5159|false|false|false|C0587081|Laboratory test finding|LABS
Finding|Body Substance|General Exam|5187,5192|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|5187,5192|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|5187,5192|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Lab|Laboratory or Test Result|General Exam|5187,5197|false|false|false|C0221752;C2188659|Red blood cells urine positive|URINE  RBC
Anatomy|Cell|General Exam|5194,5197|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|5194,5197|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|5194,5197|false|false|false|C0014792|Erythrocytes|RBC
Anatomy|Cell|General Exam|5200,5203|false|false|false|C0023516|Leukocytes|WBC
Finding|Functional Concept|General Exam|5208,5216|false|false|false|C1510439|bacteria aspects|BACTERIA
Drug|Food|General Exam|5222,5227|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Drug|Immunologic Factor|General Exam|5222,5227|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|5222,5227|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Drug|Pharmacologic Substance|General Exam|5222,5227|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Disorder|Disease or Syndrome|General Exam|5234,5237|false|false|false|C0267963|Exocrine pancreatic insufficiency|EPI
Drug|Amino Acid, Peptide, or Protein|General Exam|5234,5237|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Drug|Biologically Active Substance|General Exam|5234,5237|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Drug|Hormone|General Exam|5234,5237|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Drug|Organic Chemical|General Exam|5234,5237|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Drug|Pharmacologic Substance|General Exam|5234,5237|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Finding|Gene or Genome|General Exam|5234,5237|false|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|EPI
Finding|Intellectual Product|General Exam|5234,5237|false|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|EPI
Procedure|Diagnostic Procedure|General Exam|5234,5237|false|false|false|C0162734;C3641909|Echo-Planar Imaging;Electronic Portal Imaging|EPI
Finding|Finding|General Exam|5241,5246|false|false|false|C0558141|Transsexual (finding)|TRANS
Disorder|Disease or Syndrome|General Exam|5247,5250|false|false|false|C0267963|Exocrine pancreatic insufficiency|EPI
Drug|Amino Acid, Peptide, or Protein|General Exam|5247,5250|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Drug|Biologically Active Substance|General Exam|5247,5250|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Drug|Hormone|General Exam|5247,5250|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Drug|Organic Chemical|General Exam|5247,5250|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Drug|Pharmacologic Substance|General Exam|5247,5250|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Finding|Gene or Genome|General Exam|5247,5250|false|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|EPI
Finding|Intellectual Product|General Exam|5247,5250|false|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|EPI
Procedure|Diagnostic Procedure|General Exam|5247,5250|false|false|false|C0162734;C3641909|Echo-Planar Imaging;Electronic Portal Imaging|EPI
Finding|Body Substance|General Exam|5266,5271|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|5266,5271|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|5266,5271|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Disorder|Disease or Syndrome|General Exam|5266,5278|false|false|false|C0018965|Hematuria|URINE  BLOOD
Disorder|Disease or Syndrome|General Exam|5273,5278|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|5273,5278|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Finding|Finding|General Exam|5279,5282|false|false|false|C5848551|Neg - answer|NEG
Drug|Biologically Active Substance|General Exam|5283,5290|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|NITRITE
Drug|Inorganic Chemical|General Exam|5283,5290|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|NITRITE
Drug|Pharmacologic Substance|General Exam|5283,5290|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|NITRITE
Finding|Finding|General Exam|5291,5294|false|false|false|C5848551|Neg - answer|NEG
Drug|Amino Acid, Peptide, or Protein|General Exam|5295,5302|false|false|false|C0033684|Proteins|PROTEIN
Drug|Biologically Active Substance|General Exam|5295,5302|false|false|false|C0033684|Proteins|PROTEIN
Finding|Conceptual Entity|General Exam|5295,5302|false|false|false|C1521746|Protein Info|PROTEIN
Procedure|Laboratory Procedure|General Exam|5295,5302|false|false|false|C0202202|Protein measurement|PROTEIN
Finding|Finding|General Exam|5303,5306|false|false|false|C5848551|Neg - answer|NEG
Drug|Biologically Active Substance|General Exam|5308,5315|false|false|false|C0017725|glucose|GLUCOSE
Drug|Organic Chemical|General Exam|5308,5315|false|false|false|C0017725|glucose|GLUCOSE
Drug|Pharmacologic Substance|General Exam|5308,5315|false|false|false|C0017725|glucose|GLUCOSE
Lab|Laboratory or Test Result|General Exam|5308,5315|false|false|false|C5781949|Glucose^1.5H post dose glucagon|GLUCOSE
Procedure|Laboratory Procedure|General Exam|5308,5315|false|false|false|C0337438|Glucose measurement|GLUCOSE
Finding|Finding|General Exam|5316,5319|false|false|false|C5848551|Neg - answer|NEG
Drug|Organic Chemical|General Exam|5320,5326|false|false|false|C0022634|Ketones|KETONE
Finding|Finding|General Exam|5327,5330|false|false|false|C5848551|Neg - answer|NEG
Drug|Biologically Active Substance|General Exam|5331,5340|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|BILIRUBIN
Drug|Organic Chemical|General Exam|5331,5340|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|BILIRUBIN
Drug|Pharmacologic Substance|General Exam|5331,5340|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|BILIRUBIN
Procedure|Laboratory Procedure|General Exam|5331,5340|false|false|false|C0201913;C0863174|Bilirubin, total measurement;blood bilirubin level test|BILIRUBIN
Finding|Finding|General Exam|5341,5344|false|false|false|C5848551|Neg - answer|NEG
Finding|Finding|General Exam|5355,5358|false|false|false|C5848551|Neg - answer|NEG
Disorder|Disease or Syndrome|General Exam|5372,5375|false|false|false|C0011860|Diabetes Mellitus, Non-Insulin-Dependent|MOD
Procedure|Laboratory Procedure|General Exam|5390,5393|false|false|false|C0201617|Primed lymphocyte test|PLT
Finding|Body Substance|General Exam|5430,5436|false|false|false|C0024202|Lymph|LYMPHS
Drug|Antibiotic|General Exam|5443,5448|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Biomedical or Dental Material|General Exam|5443,5448|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Organic Chemical|General Exam|5443,5448|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Disorder|Disease or Syndrome|General Exam|5453,5456|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|EOS
Finding|Gene or Genome|General Exam|5453,5456|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|EOS
Anatomy|Cell|General Exam|5563,5566|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|5573,5576|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|5573,5576|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|5573,5576|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|5583,5586|false|false|false|C0019046|Hemoglobin|HGB
Drug|Biologically Active Substance|General Exam|5583,5586|false|false|false|C0019046|Hemoglobin|HGB
Finding|Gene or Genome|General Exam|5583,5586|false|false|false|C1424337|CYGB gene|HGB
Lab|Laboratory or Test Result|General Exam|5583,5586|false|false|false|C0019029|Hemoglobin concentration|HGB
Procedure|Laboratory Procedure|General Exam|5592,5595|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Procedure|Therapeutic or Preventive Procedure|General Exam|5592,5595|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Disorder|Virus|General Exam|5602,5605|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|General Exam|5602,5605|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|5602,5605|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|5602,5605|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|5611,5614|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|5611,5614|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|General Exam|5611,5614|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|5611,5614|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|5611,5614|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|General Exam|5621,5625|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Drug|Biologically Active Substance|General Exam|5667,5674|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Element, Ion, or Isotope|General Exam|5667,5674|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Inorganic Chemical|General Exam|5667,5674|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Pharmacologic Substance|General Exam|5667,5674|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Vitamin|General Exam|5667,5674|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Finding|Physiologic Function|General Exam|5667,5674|false|false|false|C4553026|Calcium metabolic function|CALCIUM
Procedure|Laboratory Procedure|General Exam|5667,5674|false|false|false|C0201925|Calcium measurement|CALCIUM
Drug|Element, Ion, or Isotope|General Exam|5680,5689|false|false|false|C0031603;C1601799|Phosphates;phosphate ion|PHOSPHATE
Drug|Inorganic Chemical|General Exam|5680,5689|false|false|false|C0031603;C1601799|Phosphates;phosphate ion|PHOSPHATE
Drug|Pharmacologic Substance|General Exam|5680,5689|false|false|false|C0031603;C1601799|Phosphates;phosphate ion|PHOSPHATE
Procedure|Laboratory Procedure|General Exam|5680,5689|false|false|false|C0523826|Phosphate measurement|PHOSPHATE
Drug|Biologically Active Substance|General Exam|5694,5703|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Drug|Element, Ion, or Isotope|General Exam|5694,5703|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Drug|Inorganic Chemical|General Exam|5694,5703|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Drug|Pharmacologic Substance|General Exam|5694,5703|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Procedure|Laboratory Procedure|General Exam|5694,5703|false|false|false|C0373675|Magnesium measurement|MAGNESIUM
Drug|Amino Acid, Peptide, or Protein|General Exam|5736,5742|false|false|false|C5574646|Natriuretic Peptides B, human|proBNP
Drug|Hormone|General Exam|5736,5742|false|false|false|C5574646|Natriuretic Peptides B, human|proBNP
Drug|Biologically Active Substance|General Exam|5763,5770|false|false|false|C0017725|glucose|GLUCOSE
Drug|Organic Chemical|General Exam|5763,5770|false|false|false|C0017725|glucose|GLUCOSE
Drug|Pharmacologic Substance|General Exam|5763,5770|false|false|false|C0017725|glucose|GLUCOSE
Lab|Laboratory or Test Result|General Exam|5763,5770|false|false|false|C5781949|Glucose^1.5H post dose glucagon|GLUCOSE
Procedure|Laboratory Procedure|General Exam|5763,5770|false|false|false|C0337438|Glucose measurement|GLUCOSE
Drug|Biologically Active Substance|General Exam|5776,5780|false|false|false|C0041942|urea|UREA
Drug|Organic Chemical|General Exam|5776,5780|false|false|false|C0041942|urea|UREA
Drug|Pharmacologic Substance|General Exam|5776,5780|false|false|false|C0041942|urea|UREA
Procedure|Laboratory Procedure|General Exam|5776,5780|false|false|false|C0523961|Urea measurement|UREA
Drug|Biologically Active Substance|General Exam|5797,5803|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Element, Ion, or Isotope|General Exam|5797,5803|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Pharmacologic Substance|General Exam|5797,5803|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Finding|Physiologic Function|General Exam|5797,5803|false|false|false|C4553025|Sodium metabolic function|SODIUM
Procedure|Laboratory Procedure|General Exam|5797,5803|false|false|false|C0337443|Sodium measurement|SODIUM
Drug|Biologically Active Substance|General Exam|5809,5818|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Element, Ion, or Isotope|General Exam|5809,5818|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Food|General Exam|5809,5818|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Inorganic Chemical|General Exam|5809,5818|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Pharmacologic Substance|General Exam|5809,5818|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Finding|Physiologic Function|General Exam|5809,5818|false|false|false|C4553027|Potassium metabolic function|POTASSIUM
Procedure|Laboratory Procedure|General Exam|5809,5818|false|false|false|C0202194|Potassium measurement|POTASSIUM
Drug|Element, Ion, or Isotope|General Exam|5824,5832|false|false|false|C0008203;C0596019|Chlorides;chloride ion|CHLORIDE
Finding|Physiologic Function|General Exam|5824,5832|false|false|false|C4553021|Chloride metabolic function|CHLORIDE
Procedure|Laboratory Procedure|General Exam|5824,5832|false|false|false|C0201952|Chloride measurement|CHLORIDE
Drug|Biologically Active Substance|General Exam|5843,5846|false|false|false|C0007012|carbon dioxide|CO2
Drug|Inorganic Chemical|General Exam|5843,5846|false|false|false|C0007012|carbon dioxide|CO2
Finding|Finding|General Exam|5843,5846|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Finding|Gene or Genome|General Exam|5843,5846|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Drug|Element, Ion, or Isotope|General Exam|5851,5856|false|false|false|C0003075|Anions|ANION
Attribute|Clinical Attribute|General Exam|5851,5860|false|false|false|C0003074|Anion Gap|ANION GAP
Lab|Laboratory or Test Result|General Exam|5851,5860|false|false|false|C1509129|Anion gap result|ANION GAP
Procedure|Laboratory Procedure|General Exam|5851,5860|false|false|false|C0201889;C2189246|Anion gap measurement;blood anion gap (lab test)|ANION GAP
Drug|Amino Acid, Peptide, or Protein|General Exam|5857,5860|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Drug|Biologically Active Substance|General Exam|5857,5860|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Finding|Gene or Genome|General Exam|5857,5860|false|false|false|C1419277;C2984552|RASA1 gene;RASA1 wt Allele|GAP
Procedure|Research Activity|General Exam|5865,5872|false|false|false|C0947630|Scientific Study|STUDIES
Procedure|Diagnostic Procedure|General Exam|5882,5885|false|false|false|C0039985|Plain chest X-ray|CXR
Anatomy|Tissue|General Exam|5897,5904|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|General Exam|5897,5904|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Pathologic Function|General Exam|5897,5914|false|false|false|C0032227|Pleural effusion (disorder)|pleural effusions
Finding|Pathologic Function|General Exam|5905,5914|false|false|false|C0013687|effusion|effusions
Finding|Gene or Genome|General Exam|5916,5921|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Finding|Functional Concept|General Exam|5929,5934|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Finding|Functional Concept|General Exam|5953,5957|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Disorder|Disease or Syndrome|General Exam|5979,5992|false|false|false|C0521530|Lung consolidation|consolidation
Finding|Idea or Concept|General Exam|6014,6024|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|General Exam|6014,6024|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Finding|Functional Concept|General Exam|6029,6036|false|false|false|C0439801;C3542948|Limited (extensiveness);Limited component (foundation metadata concept)|limited
Finding|Intellectual Product|General Exam|6029,6036|false|false|false|C0439801;C3542948|Limited (extensiveness);Limited component (foundation metadata concept)|limited
Disorder|Neoplastic Process|General Exam|6038,6047|false|false|false|C0027627|Neoplasm Metastasis|secondary
Finding|Functional Concept|General Exam|6038,6047|false|false|false|C1522484|metastatic qualifier|secondary
Finding|Pathologic Function|General Exam|6057,6066|false|false|false|C0013687|effusion|effusions
Anatomy|Body Part, Organ, or Organ Component|General Exam|6070,6076|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|Pelvis
Anatomy|Body Space or Junction|General Exam|6070,6076|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|Pelvis
Disorder|Neoplastic Process|General Exam|6070,6076|false|false|false|C0153663|Malignant neoplasm of pelvis|Pelvis
Finding|Finding|General Exam|6070,6076|false|false|false|C0812455|Pelvis problem|Pelvis
Phenomenon|Natural Phenomenon or Process|General Exam|6077,6081|false|false|false|C0043309|Roentgen Rays|Xray
Procedure|Diagnostic Procedure|General Exam|6077,6081|false|false|false|C0043299|Diagnostic radiologic examination|Xray
Finding|Intellectual Product|General Exam|6095,6100|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Disorder|Injury or Poisoning|General Exam|6101,6109|true|false|false|C0016658|Fracture|fracture
Disorder|Injury or Poisoning|General Exam|6113,6124|true|false|false|C0012691|Dislocations|dislocation
Finding|Pathologic Function|General Exam|6136,6141|true|false|false|C0024348|Lysis|lytic
Finding|Functional Concept|General Exam|6146,6155|false|false|false|C0036429;C0334135|Sclerosis;Sclerotic (qualifier value)|sclerotic
Finding|Pathologic Function|General Exam|6146,6155|false|false|false|C0036429;C0334135|Sclerosis;Sclerotic (qualifier value)|sclerotic
Anatomy|Body Part, Organ, or Organ Component|General Exam|6157,6164|false|false|false|C0262950;C4520924|Bone Tissue, Human;Skeletal bone|osseous
Anatomy|Tissue|General Exam|6157,6164|false|false|false|C0262950;C4520924|Bone Tissue, Human;Skeletal bone|osseous
Finding|Finding|General Exam|6165,6171|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|General Exam|6165,6171|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Idea or Concept|General Exam|6205,6212|false|false|false|C0376327|International Aspects|foreign
Disorder|Injury or Poisoning|General Exam|6205,6217|true|false|false|C0016542|Foreign Bodies|foreign body
Anatomy|Anatomical Structure|General Exam|6213,6217|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Anatomy|Body Part, Organ, or Organ Component|General Exam|6213,6217|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Finding|Intellectual Product|General Exam|6213,6217|true|false|false|C1551342|Document Body|body
Anatomy|Body Part, Organ, or Organ Component|General Exam|6221,6229|false|false|false|C0005847|Blood Vessel|Vascular
Finding|Finding|General Exam|6231,6245|false|false|false|C0006660;C2242558|Pathologic calcification, calcified structure;Physiologic calcification|calcifications
Finding|Organ or Tissue Function|General Exam|6231,6245|false|false|false|C0006660;C2242558|Pathologic calcification, calcified structure;Physiologic calcification|calcifications
Anatomy|Body Part, Organ, or Organ Component|General Exam|6273,6278|false|false|false|C0021853|Intestines|bowel
Drug|Biomedical or Dental Material|General Exam|6279,6282|false|false|false|C0017110;C1550641;C1704673|Gas - SpecimenType;Gas Dosage Form;Gases|gas
Drug|Chemical Viewed Structurally|General Exam|6279,6282|false|false|false|C0017110;C1550641;C1704673|Gas - SpecimenType;Gas Dosage Form;Gases|gas
Drug|Substance|General Exam|6279,6282|false|false|false|C0017110;C1550641;C1704673|Gas - SpecimenType;Gas Dosage Form;Gases|gas
Finding|Gene or Genome|General Exam|6279,6282|false|false|false|C0596601;C1414950;C1439341;C1540252;C1546643;C2266618;C2986619;C3812826;C5890923|GALNS gene;GALNS wt Allele;GAST gene;GAST wt Allele;Gas - Specimen Source Codes;PAGR1 gene;PAGR1 wt Allele;gastrointestinal gas;germacrene-A synthase activity|gas
Finding|Intellectual Product|General Exam|6279,6282|false|false|false|C0596601;C1414950;C1439341;C1540252;C1546643;C2266618;C2986619;C3812826;C5890923|GALNS gene;GALNS wt Allele;GAST gene;GAST wt Allele;Gas - Specimen Source Codes;PAGR1 gene;PAGR1 wt Allele;gastrointestinal gas;germacrene-A synthase activity|gas
Finding|Molecular Function|General Exam|6279,6282|false|false|false|C0596601;C1414950;C1439341;C1540252;C1546643;C2266618;C2986619;C3812826;C5890923|GALNS gene;GALNS wt Allele;GAST gene;GAST wt Allele;Gas - Specimen Source Codes;PAGR1 gene;PAGR1 wt Allele;gastrointestinal gas;germacrene-A synthase activity|gas
Finding|Sign or Symptom|General Exam|6279,6282|false|false|false|C0596601;C1414950;C1439341;C1540252;C1546643;C2266618;C2986619;C3812826;C5890923|GALNS gene;GALNS wt Allele;GAST gene;GAST wt Allele;Gas - Specimen Source Codes;PAGR1 gene;PAGR1 wt Allele;gastrointestinal gas;germacrene-A synthase activity|gas
Finding|Intellectual Product|General Exam|6315,6325|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|General Exam|6315,6325|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Intellectual Product|General Exam|6331,6336|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Disorder|Injury or Poisoning|General Exam|6337,6345|true|false|false|C0016658|Fracture|fracture
Disorder|Injury or Poisoning|General Exam|6349,6360|true|false|false|C0012691|Dislocations|dislocation
Anatomy|Body Location or Region|General Exam|6364,6369|false|false|false|C1548802|Body Site Modifier - Lower|Lower
Event|Activity|General Exam|6364,6369|false|false|false|C2003888|Lower (action)|Lower
Anatomy|Body Part, Organ, or Organ Component|General Exam|6364,6379|false|false|false|C0023216|Lower Extremity|Lower extremity
Anatomy|Body Part, Organ, or Organ Component|General Exam|6370,6379|false|false|false|C0015385|Limb structure|extremity
Finding|Functional Concept|General Exam|6380,6390|false|false|false|C0220934|Ultrasonic|ultrasound
Phenomenon|Natural Phenomenon or Process|General Exam|6380,6390|false|false|false|C0041621;C1456803|Ultrasonic Shockwave;Ultrasonics (sound)|ultrasound
Procedure|Diagnostic Procedure|General Exam|6380,6390|false|false|false|C0041618;C1315081|Ultrasonography;Urological ultrasound|ultrasound
Attribute|Clinical Attribute|General Exam|6395,6399|false|false|false|C4318566|Deep Resection Margin|Deep
Anatomy|Body Part, Organ, or Organ Component|General Exam|6395,6404|false|false|false|C0226514|Structure of deep vein|Deep vein
Disorder|Disease or Syndrome|General Exam|6395,6415|false|false|false|C0149871;C0340708|Deep Vein Thrombosis;Deep vein thrombosis of lower limb|Deep vein thrombosis
Anatomy|Body Part, Organ, or Organ Component|General Exam|6400,6404|false|false|false|C0042449|Veins|vein
Finding|Pathologic Function|General Exam|6400,6415|false|false|false|C0042487|Venous Thrombosis|vein thrombosis
Finding|Pathologic Function|General Exam|6405,6415|false|false|false|C0040053|Thrombosis|thrombosis
Finding|Functional Concept|General Exam|6423,6427|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Finding|Functional Concept|General Exam|6428,6434|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Finding|Intellectual Product|General Exam|6428,6434|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Anatomy|Body Part, Organ, or Organ Component|General Exam|6428,6447|false|false|false|C1275667|Common femoral vein|common femoral vein
Anatomy|Body Part, Organ, or Organ Component|General Exam|6435,6442|false|false|false|C0015811|Femur|femoral
Anatomy|Body Part, Organ, or Organ Component|General Exam|6435,6447|false|false|false|C0015809|Femoral vein|femoral vein
Anatomy|Body Part, Organ, or Organ Component|General Exam|6443,6447|false|false|false|C0042449|Veins|vein
Anatomy|Body Location or Region|General Exam|6478,6487|false|false|false|C0442037|popliteal|popliteal
Anatomy|Body Part, Organ, or Organ Component|General Exam|6478,6492|false|false|false|C0032652|Structure of popliteal vein|popliteal vein
Anatomy|Body Part, Organ, or Organ Component|General Exam|6488,6492|false|false|false|C0042449|Veins|vein
Finding|Functional Concept|General Exam|6495,6499|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Location or Region|General Exam|6495,6504|false|false|false|C0489800|Posterior part of left leg|Left calf
Anatomy|Body Location or Region|General Exam|6500,6504|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Part, Organ, or Organ Component|General Exam|6500,6504|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Part, Organ, or Organ Component|General Exam|6505,6510|false|false|false|C0042449|Veins|veins
Procedure|Therapeutic or Preventive Procedure|General Exam|6505,6510|false|false|false|C0398102|Procedure on vein|veins
Finding|Finding|General Exam|6542,6550|false|false|false|C0332149|Possible|possibly
Finding|Finding|General Exam|6556,6564|false|false|false|C0028778;C1947917|Obstruction;Occluded|occluded
Finding|Functional Concept|General Exam|6556,6564|false|false|false|C0028778;C1947917|Obstruction;Occluded|occluded
Finding|Functional Concept|General Exam|6574,6579|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|General Exam|6580,6583|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|General Exam|6580,6583|true|false|false|C2926618||DVT
Disorder|Disease or Syndrome|General Exam|6580,6583|true|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Lab|Laboratory or Test Result|General Exam|6592,6596|false|false|false|C0587081|Laboratory test finding|LABS
Finding|Body Substance|General Exam|6604,6613|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|General Exam|6604,6613|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|General Exam|6604,6613|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|General Exam|6604,6613|false|false|false|C0030685|Patient Discharge|DISCHARGE
Disorder|Disease or Syndrome|General Exam|6659,6664|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|6659,6664|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|6665,6668|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|6675,6678|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|6675,6678|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|6675,6678|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|6685,6688|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|6685,6688|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|6685,6688|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|6685,6688|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|6694,6697|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|6694,6697|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|6704,6707|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|General Exam|6704,6707|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|6704,6707|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|6704,6707|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|6713,6716|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|6713,6716|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|General Exam|6713,6716|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|6713,6716|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|6713,6716|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|General Exam|6723,6727|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|6755,6758|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|6775,6780|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|6775,6780|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|6775,6788|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|6775,6788|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|6775,6788|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|6781,6788|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|6781,6788|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|6781,6788|false|false|false|C0017725|glucose|Glucose
Lab|Laboratory or Test Result|General Exam|6781,6788|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|6781,6788|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|General Exam|6834,6838|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|6834,6838|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|General Exam|6834,6838|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|General Exam|6864,6869|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|6864,6869|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|6864,6877|false|false|false|C0853248|Blood albumin|BLOOD Albumin
Drug|Amino Acid, Peptide, or Protein|General Exam|6870,6877|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Biologically Active Substance|General Exam|6870,6877|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Pharmacologic Substance|General Exam|6870,6877|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Finding|Gene or Genome|General Exam|6870,6877|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Finding|Physiologic Function|General Exam|6870,6877|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Procedure|Laboratory Procedure|General Exam|6870,6877|false|false|false|C0201838|Albumin measurement|Albumin
Drug|Biologically Active Substance|General Exam|6883,6890|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|General Exam|6883,6890|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|General Exam|6883,6890|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|General Exam|6883,6890|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|General Exam|6883,6890|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Finding|Physiologic Function|General Exam|6883,6890|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|General Exam|6883,6890|false|false|false|C0201925|Calcium measurement|Calcium
Anatomy|Body Space or Junction|Hospital Course|6968,6971|false|false|false|C0262212|Choroidal fissure|CHF
Disorder|Disease or Syndrome|Hospital Course|6968,6971|false|false|false|C0018802|Congestive heart failure|CHF
Disorder|Disease or Syndrome|Hospital Course|6973,6977|false|false|false|C0004238|Atrial Fibrillation|Afib
Lab|Laboratory or Test Result|Hospital Course|6973,6977|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Afib
Finding|Finding|Hospital Course|6986,7001|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Finding|Physiologic Function|Hospital Course|6986,7001|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6986,7001|false|false|false|C0003281|Anticoagulation Therapy|anticoagulation
Finding|Finding|Hospital Course|7003,7009|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|Hospital Course|7003,7009|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Disorder|Disease or Syndrome|Hospital Course|7019,7028|false|false|false|C0002395|Alzheimer's Disease|Alzheimer
Disorder|Disease or Syndrome|Hospital Course|7019,7039|false|false|false|C0002395|Alzheimer's Disease|Alzheimer's dementia
Disorder|Mental or Behavioral Dysfunction|Hospital Course|7031,7039|false|false|false|C0011265;C0497327|Dementia;Presenile dementia|dementia
Disorder|Disease or Syndrome|Hospital Course|7042,7054|false|false|false|C0029456|Osteoporosis|osteoporosis
Finding|Finding|Hospital Course|7042,7054|false|false|false|C2911643|Encounter due to family history of osteoporosis|osteoporosis
Disorder|Disease or Syndrome|Hospital Course|7056,7059|false|false|false|C0020538|Hypertensive disease|HTN
Procedure|Health Care Activity|Hospital Course|7079,7094|false|false|false|C1456630|Assisted Living|assisted living
Finding|Conceptual Entity|Hospital Course|7088,7094|false|false|false|C0595998;C4520849;C4551704|Alive;Household composition;Living|living
Finding|Finding|Hospital Course|7088,7094|false|false|false|C0595998;C4520849;C4551704|Alive;Household composition;Living|living
Finding|Intellectual Product|Hospital Course|7095,7103|false|false|false|C4695111|ADMIN.FACILITY|facility
Anatomy|Body Location or Region|Hospital Course|7110,7115|false|false|false|C0524470|Right hip region structure|R hip
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7112,7115|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|hip
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7112,7115|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Biologically Active Substance|Hospital Course|7112,7115|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Pharmacologic Substance|Hospital Course|7112,7115|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Finding|Gene or Genome|Hospital Course|7112,7115|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|hip
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7112,7115|false|false|false|C1292890|Procedure on hip|hip
Attribute|Clinical Attribute|Hospital Course|7112,7120|false|false|false|C1716793||hip pain
Finding|Sign or Symptom|Hospital Course|7112,7120|false|false|false|C0019559;C4551516|Hip joint pain;Hip pain|hip pain
Attribute|Clinical Attribute|Hospital Course|7116,7120|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|7116,7120|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|7116,7120|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Anatomy|Body Location or Region|Hospital Course|7136,7139|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|Hospital Course|7136,7139|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|Hospital Course|7136,7139|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Finding|Functional Concept|Hospital Course|7140,7144|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Finding|Functional Concept|Hospital Course|7145,7151|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Finding|Intellectual Product|Hospital Course|7145,7151|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7145,7164|false|false|false|C1275667|Common femoral vein|common femoral vein
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7152,7159|false|false|false|C0015811|Femur|femoral
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7152,7164|false|false|false|C0015809|Femoral vein|femoral vein
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7160,7164|false|false|false|C0042449|Veins|vein
Finding|Intellectual Product|Hospital Course|7171,7177|false|false|false|C1705102|Volume (publication)|volume
Finding|Pathologic Function|Hospital Course|7171,7186|false|false|false|C0546817|Hypervolemia (finding)|volume overload
Event|Activity|Hospital Course|7197,7204|false|false|false|C0556656|Meetings|meeting
Finding|Body Substance|Hospital Course|7210,7217|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|7210,7217|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|7210,7217|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7222,7232|false|false|false|C3812393|ErbB Receptors|her family
Drug|Enzyme|Hospital Course|7222,7232|false|false|false|C3812393|ErbB Receptors|her family
Finding|Receptor|Hospital Course|7222,7232|false|false|false|C3812393|ErbB Receptors|her family
Finding|Classification|Hospital Course|7226,7232|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|Hospital Course|7226,7232|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|Hospital Course|7226,7232|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|Hospital Course|7226,7232|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Mental Process|Hospital Course|7235,7243|false|false|false|C0679006|Decision|decision
Disorder|Cell or Molecular Dysfunction|Hospital Course|7256,7266|false|false|false|C0599156|Transition Mutation|transition
Event|Activity|Hospital Course|7256,7266|false|false|false|C2700061|Transition (action)|transition
Procedure|Health Care Activity|Hospital Course|7256,7271|false|false|false|C4019071|Transitional Care|transition care
Event|Activity|Hospital Course|7267,7271|false|false|false|C1947933|care activity|care
Finding|Finding|Hospital Course|7267,7271|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Hospital Course|7267,7271|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Drug|Organic Chemical|Hospital Course|7275,7282|false|false|false|C1310585|Comfort brand of hydroxyethyl cellulose|comfort
Drug|Pharmacologic Substance|Hospital Course|7275,7282|false|false|false|C1310585|Comfort brand of hydroxyethyl cellulose|comfort
Finding|Mental Process|Hospital Course|7275,7282|false|false|false|C1331418|Comfort|comfort
Procedure|Health Care Activity|Hospital Course|7321,7328|false|false|false|C0085555|Hospice Care|hospice
Event|Occupational Activity|Hospital Course|7321,7337|false|false|false|C5423046|Purchased Services, Clinical and Biomedical, Home Healthcare, Hospice|hospice services
Event|Occupational Activity|Hospital Course|7329,7337|false|false|false|C0557854|Services|services
Procedure|Health Care Activity|Hospital Course|7329,7337|false|false|false|C1704289|Clinical Service|services
Finding|Body Substance|Hospital Course|7341,7350|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|7341,7350|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|7341,7350|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|7341,7350|false|false|false|C0030685|Patient Discharge|discharge
Disorder|Disease or Syndrome|Hospital Course|7385,7388|false|false|false|C0410422|Chronic multifocal osteomyelitis|CMO
Finding|Classification|Hospital Course|7405,7411|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|Hospital Course|7405,7411|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|Hospital Course|7405,7411|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|Hospital Course|7405,7411|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Event|Activity|Hospital Course|7412,7419|false|false|false|C0556656|Meetings|meeting
Finding|Mental Process|Hospital Course|7431,7439|false|false|false|C0679006|Decision|decision
Disorder|Cell or Molecular Dysfunction|Hospital Course|7453,7463|false|false|false|C0599156|Transition Mutation|transition
Event|Activity|Hospital Course|7453,7463|false|false|false|C2700061|Transition (action)|transition
Procedure|Health Care Activity|Hospital Course|7453,7468|false|false|false|C4019071|Transitional Care|transition care
Event|Activity|Hospital Course|7464,7468|false|false|false|C1947933|care activity|care
Finding|Finding|Hospital Course|7464,7468|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Hospital Course|7464,7468|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Disorder|Disease or Syndrome|Hospital Course|7472,7475|false|false|false|C0410422|Chronic multifocal osteomyelitis|CMO
Procedure|Health Care Activity|Hospital Course|7495,7502|false|false|false|C0085555|Hospice Care|hospice
Event|Occupational Activity|Hospital Course|7504,7512|false|false|false|C0557854|Services|services
Procedure|Health Care Activity|Hospital Course|7504,7512|false|false|false|C1704289|Clinical Service|services
Finding|Body Substance|Hospital Course|7516,7525|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|7516,7525|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|7516,7525|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|7516,7525|false|false|false|C0030685|Patient Discharge|discharge
Finding|Classification|Hospital Course|7527,7533|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|Hospital Course|7527,7533|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|Hospital Course|7527,7533|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|Hospital Course|7527,7533|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7565,7575|false|false|false|C0087111|Therapeutic procedure|treatments
Drug|Organic Chemical|Hospital Course|7584,7589|false|false|false|C0699992|Lasix|Lasix
Drug|Pharmacologic Substance|Hospital Course|7584,7589|false|false|false|C0699992|Lasix|Lasix
Disorder|Disease or Syndrome|Hospital Course|7633,7645|false|false|false|C0021167|Incontinence|incontinence
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7649,7654|false|false|false|C1456647|Childhood Vaccines|shots
Drug|Immunologic Factor|Hospital Course|7649,7654|false|false|false|C1456647|Childhood Vaccines|shots
Drug|Pharmacologic Substance|Hospital Course|7649,7654|false|false|false|C1456647|Childhood Vaccines|shots
Drug|Organic Chemical|Hospital Course|7663,7670|false|false|false|C0728963|Lovenox|lovenox
Drug|Pharmacologic Substance|Hospital Course|7663,7670|false|false|false|C0728963|Lovenox|lovenox
Finding|Conceptual Entity|Hospital Course|7675,7684|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|Hospital Course|7675,7684|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|Hospital Course|7675,7684|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7675,7684|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Anatomy|Body Location or Region|Hospital Course|7689,7692|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|Hospital Course|7689,7692|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|Hospital Course|7689,7692|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Finding|Idea or Concept|Hospital Course|7694,7698|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|7694,7698|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|7694,7698|false|false|false|C1553498|home health encounter|Home
Attribute|Clinical Attribute|Hospital Course|7699,7710|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Hospital Course|7699,7710|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|Hospital Course|7699,7710|false|false|false|C4284232|Medications|medications
Drug|Organic Chemical|Hospital Course|7711,7721|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|Hospital Course|7711,7721|false|false|false|C0025859|metoprolol|metoprolol
Drug|Organic Chemical|Hospital Course|7723,7732|false|false|false|C0527316|donepezil|donepezil
Drug|Pharmacologic Substance|Hospital Course|7723,7732|false|false|false|C0527316|donepezil|donepezil
Drug|Pharmacologic Substance|Hospital Course|7723,7746|false|false|false|C3652776|donepezil / memantine|donepezil and Memantine
Drug|Organic Chemical|Hospital Course|7737,7746|false|false|false|C0025242|memantine|Memantine
Drug|Pharmacologic Substance|Hospital Course|7737,7746|false|false|false|C0025242|memantine|Memantine
Drug|Organic Chemical|Hospital Course|7767,7774|false|false|false|C1310585|Comfort brand of hydroxyethyl cellulose|comfort
Drug|Pharmacologic Substance|Hospital Course|7767,7774|false|false|false|C1310585|Comfort brand of hydroxyethyl cellulose|comfort
Finding|Mental Process|Hospital Course|7767,7774|false|false|false|C1331418|Comfort|comfort
Finding|Intellectual Product|Hospital Course|7810,7818|false|false|false|C4695111|ADMIN.FACILITY|facility
Finding|Idea or Concept|Hospital Course|7828,7836|false|false|false|C1547192|Organization unit type - Hospital|HOSPITAL
Anatomy|Body Location or Region|Hospital Course|7870,7873|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|Hospital Course|7870,7873|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|Hospital Course|7870,7873|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Attribute|Clinical Attribute|Hospital Course|7875,7879|false|false|false|C4318566|Deep Resection Margin|Deep
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7875,7884|false|false|false|C0226514|Structure of deep vein|Deep vein
Disorder|Disease or Syndrome|Hospital Course|7875,7895|false|false|false|C0149871;C0340708|Deep Vein Thrombosis;Deep vein thrombosis of lower limb|Deep vein thrombosis
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7880,7884|false|false|false|C0042449|Veins|vein
Finding|Pathologic Function|Hospital Course|7880,7895|false|false|false|C0042487|Venous Thrombosis|vein thrombosis
Finding|Pathologic Function|Hospital Course|7885,7895|false|false|false|C0040053|Thrombosis|thrombosis
Finding|Functional Concept|Hospital Course|7903,7907|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Finding|Functional Concept|Hospital Course|7908,7914|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Finding|Intellectual Product|Hospital Course|7908,7914|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7908,7927|false|false|false|C1275667|Common femoral vein|common femoral vein
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7915,7922|false|false|false|C0015811|Femur|femoral
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7915,7927|false|false|false|C0015809|Femoral vein|femoral vein
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7923,7927|false|false|false|C0042449|Veins|vein
Anatomy|Body Location or Region|Hospital Course|7957,7966|false|false|false|C0442037|popliteal|popliteal
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7957,7971|false|false|false|C0032652|Structure of popliteal vein|popliteal vein
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7967,7971|false|false|false|C0042449|Veins|vein
Finding|Functional Concept|Hospital Course|7986,7996|false|false|false|C0220934|Ultrasonic|ultrasound
Phenomenon|Natural Phenomenon or Process|Hospital Course|7986,7996|false|false|false|C0041621;C1456803|Ultrasonic Shockwave;Ultrasonics (sound)|ultrasound
Procedure|Diagnostic Procedure|Hospital Course|7986,7996|false|false|false|C0041618;C1315081|Ultrasonography;Urological ultrasound|ultrasound
Procedure|Health Care Activity|Hospital Course|8000,8009|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Finding|Hospital Course|8020,8026|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Hospital Course|8020,8026|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Mental Process|Hospital Course|8043,8050|false|false|false|C0542559|contextual factors|setting
Finding|Finding|Hospital Course|8055,8065|false|false|false|C0231441|Immobile|immobility
Finding|Body Substance|Hospital Course|8074,8081|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|8074,8081|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|8074,8081|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Finding|Hospital Course|8110,8120|false|false|false|C2135586;C4321408|Wheelchair Usually Used;has wheelchair at home (history)|wheelchair
Procedure|Health Care Activity|Hospital Course|8128,8143|false|false|false|C1456630|Assisted Living|assisted living
Finding|Conceptual Entity|Hospital Course|8137,8143|false|false|false|C0595998;C4520849;C4551704|Alive;Household composition;Living|living
Finding|Finding|Hospital Course|8137,8143|false|false|false|C0595998;C4520849;C4551704|Alive;Household composition;Living|living
Finding|Idea or Concept|Hospital Course|8163,8168|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Intellectual Product|Hospital Course|8163,8168|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Functional Concept|Hospital Course|8169,8172|false|false|false|C0678226;C3146286|Due;Due to|due
Finding|Idea or Concept|Hospital Course|8169,8172|false|false|false|C0678226;C3146286|Due;Due to|due
Drug|Organic Chemical|Hospital Course|8222,8229|false|false|false|C0728963|Lovenox|Lovenox
Drug|Pharmacologic Substance|Hospital Course|8222,8229|false|false|false|C0728963|Lovenox|Lovenox
Finding|Conceptual Entity|Hospital Course|8235,8244|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|Hospital Course|8235,8244|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|Hospital Course|8235,8244|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8235,8244|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Finding|Mental Process|Hospital Course|8278,8285|false|false|false|C0542559|contextual factors|setting
Disorder|Cell or Molecular Dysfunction|Hospital Course|8289,8299|false|false|false|C0599156|Transition Mutation|transition
Event|Activity|Hospital Course|8289,8299|false|false|false|C2700061|Transition (action)|transition
Event|Activity|Hospital Course|8304,8308|false|false|false|C1947933|care activity|care
Finding|Finding|Hospital Course|8304,8308|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Hospital Course|8304,8308|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Disorder|Disease or Syndrome|Hospital Course|8312,8315|false|false|false|C0410422|Chronic multifocal osteomyelitis|CMO
Finding|Idea or Concept|Hospital Course|8319,8324|false|false|false|C1552828|Table Frame - above|above
Finding|Intellectual Product|Hospital Course|8330,8335|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|Acute
Anatomy|Body Space or Junction|Hospital Course|8336,8339|false|false|false|C0262212|Choroidal fissure|CHF
Disorder|Disease or Syndrome|Hospital Course|8336,8339|false|false|false|C0018802|Congestive heart failure|CHF
Finding|Body Substance|Hospital Course|8341,8348|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|8341,8348|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|8341,8348|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|8353,8359|false|false|false|C1705102|Volume (publication)|volume
Finding|Idea or Concept|Hospital Course|8374,8386|false|false|false|C0449450|Presentation|presentation
Anatomy|Tissue|Hospital Course|8393,8400|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|Hospital Course|8393,8400|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Pathologic Function|Hospital Course|8393,8410|false|false|false|C0032227|Pleural effusion (disorder)|pleural effusions
Finding|Pathologic Function|Hospital Course|8401,8410|false|false|false|C0013687|effusion|effusions
Drug|Organic Chemical|Hospital Course|8437,8442|false|false|false|C0699992|Lasix|Lasix
Drug|Pharmacologic Substance|Hospital Course|8437,8442|false|false|false|C0699992|Lasix|Lasix
Finding|Idea or Concept|Hospital Course|8444,8448|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|8444,8448|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|8444,8448|false|false|false|C1553498|home health encounter|Home
Drug|Organic Chemical|Hospital Course|8450,8460|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|Hospital Course|8450,8460|false|false|false|C0025859|metoprolol|metoprolol
Finding|Finding|Hospital Course|8480,8489|false|false|false|C0392756;C0442797|Decreasing;Reduced|decreased
Finding|Mental Process|Hospital Course|8503,8510|false|false|false|C0542559|contextual factors|setting
Disorder|Cell or Molecular Dysfunction|Hospital Course|8515,8525|false|false|false|C0599156|Transition Mutation|transition
Event|Activity|Hospital Course|8515,8525|false|false|false|C2700061|Transition (action)|transition
Event|Activity|Hospital Course|8529,8533|false|false|false|C1947933|care activity|care
Finding|Finding|Hospital Course|8529,8533|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Hospital Course|8529,8533|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Disorder|Disease or Syndrome|Hospital Course|8537,8540|false|false|false|C0410422|Chronic multifocal osteomyelitis|CMO
Drug|Organic Chemical|Hospital Course|8542,8547|false|false|false|C0699992|Lasix|Lasix
Drug|Pharmacologic Substance|Hospital Course|8542,8547|false|false|false|C0699992|Lasix|Lasix
Finding|Idea or Concept|Hospital Course|8575,8584|false|false|false|C0549178|Continuous|continued
Drug|Organic Chemical|Hospital Course|8588,8598|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|Hospital Course|8588,8598|false|false|false|C0025859|metoprolol|metoprolol
Drug|Organic Chemical|Hospital Course|8603,8610|false|false|false|C1310585|Comfort brand of hydroxyethyl cellulose|comfort
Drug|Pharmacologic Substance|Hospital Course|8603,8610|false|false|false|C1310585|Comfort brand of hydroxyethyl cellulose|comfort
Finding|Mental Process|Hospital Course|8603,8610|false|false|false|C1331418|Comfort|comfort
Finding|Finding|Hospital Course|8625,8636|false|false|false|C2709070|on room air|on room air
Drug|Inorganic Chemical|Hospital Course|8628,8636|false|false|false|C3846005|Room Air|room air
Drug|Inorganic Chemical|Hospital Course|8633,8636|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|Hospital Course|8633,8636|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|Hospital Course|8633,8636|false|false|false|C0001861;C3536832|Air (substance);air|air
Finding|Finding|Hospital Course|8633,8636|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|Hospital Course|8633,8636|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|Hospital Course|8633,8636|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Attribute|Clinical Attribute|Hospital Course|8646,8657|false|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|Hospital Course|8646,8657|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|Hospital Course|8646,8657|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|Hospital Course|8646,8657|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Sign or Symptom|Hospital Course|8646,8666|true|false|false|C0476273|Respiratory distress|respiratory distress
Finding|Finding|Hospital Course|8658,8666|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|Hospital Course|8658,8666|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Anatomy|Body Space or Junction|Hospital Course|8696,8701|false|false|false|C0030471;C1305231|Nasal sinus;Sinus - general anatomical term|sinus
Disorder|Anatomical Abnormality|Hospital Course|8696,8701|false|false|false|C0016169|pathologic fistula|sinus
Drug|Organic Chemical|Hospital Course|8696,8701|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Drug|Pharmacologic Substance|Hospital Course|8696,8701|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Finding|Finding|Hospital Course|8696,8708|false|false|false|C0232201;C2041122|Sinus rhythm|sinus rhythm
Finding|Finding|Hospital Course|8702,8708|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|Hospital Course|8702,8708|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Event|Activity|Hospital Course|8710,8714|false|false|false|C0871208|Rating (action)|rate
Finding|Idea or Concept|Hospital Course|8710,8714|false|false|false|C1549480|Amount type - Rate|rate
Drug|Organic Chemical|Hospital Course|8730,8740|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|Hospital Course|8730,8740|false|false|false|C0025859|metoprolol|metoprolol
Drug|Organic Chemical|Hospital Course|8742,8752|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|Hospital Course|8742,8752|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Organic Chemical|Hospital Course|8792,8799|false|false|false|C1310585|Comfort brand of hydroxyethyl cellulose|comfort
Drug|Pharmacologic Substance|Hospital Course|8792,8799|false|false|false|C1310585|Comfort brand of hydroxyethyl cellulose|comfort
Finding|Mental Process|Hospital Course|8792,8799|false|false|false|C1331418|Comfort|comfort
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8805,8808|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|Hip
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8805,8808|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|Hip
Drug|Biologically Active Substance|Hospital Course|8805,8808|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|Hip
Drug|Pharmacologic Substance|Hospital Course|8805,8808|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|Hip
Finding|Gene or Genome|Hospital Course|8805,8808|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|Hip
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8805,8808|false|false|false|C1292890|Procedure on hip|Hip
Attribute|Clinical Attribute|Hospital Course|8805,8813|false|false|false|C1716793||Hip pain
Finding|Sign or Symptom|Hospital Course|8805,8813|false|false|false|C0019559;C4551516|Hip joint pain;Hip pain|Hip pain
Attribute|Clinical Attribute|Hospital Course|8809,8813|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|8809,8813|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|8809,8813|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Functional Concept|Hospital Course|8819,8824|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|Hospital Course|8819,8828|false|false|false|C0524470|Right hip region structure|right hip
Finding|Sign or Symptom|Hospital Course|8819,8833|false|false|false|C2202100|Pain of right hip joint|right hip pain
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8825,8828|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|hip
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8825,8828|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Biologically Active Substance|Hospital Course|8825,8828|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Pharmacologic Substance|Hospital Course|8825,8828|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Finding|Gene or Genome|Hospital Course|8825,8828|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|hip
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8825,8828|false|false|false|C1292890|Procedure on hip|hip
Attribute|Clinical Attribute|Hospital Course|8825,8833|false|false|false|C1716793||hip pain
Finding|Sign or Symptom|Hospital Course|8825,8833|false|false|false|C0019559;C4551516|Hip joint pain;Hip pain|hip pain
Attribute|Clinical Attribute|Hospital Course|8829,8833|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|8829,8833|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|8829,8833|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|Hospital Course|8879,8883|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Hospital Course|8879,8883|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Hospital Course|8879,8883|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Procedure|Health Care Activity|Hospital Course|8887,8896|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8898,8904|false|false|false|C0030797|Pelvis|Pelvic
Phenomenon|Natural Phenomenon or Process|Hospital Course|8905,8909|false|false|false|C0043309|Roentgen Rays|xray
Procedure|Diagnostic Procedure|Hospital Course|8905,8909|false|false|false|C0043299|Diagnostic radiologic examination|xray
Disorder|Injury or Poisoning|Hospital Course|8923,8931|false|false|false|C0016658|Fracture|fracture
Drug|Organic Chemical|Hospital Course|8954,8961|false|false|false|C0699142|Tylenol|Tylenol
Drug|Pharmacologic Substance|Hospital Course|8954,8961|false|false|false|C0699142|Tylenol|Tylenol
Attribute|Clinical Attribute|Hospital Course|8976,8980|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|8976,8980|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|8976,8980|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|Hospital Course|8982,8989|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Pharmacologic Substance|Hospital Course|8982,8989|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Substance|Hospital Course|8982,8989|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Finding|Conceptual Entity|Hospital Course|8982,8989|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Functional Concept|Hospital Course|8982,8989|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Idea or Concept|Hospital Course|8982,8989|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9001,9009|false|false|false|C0011265;C0497327|Dementia;Presenile dementia|Dementia
Finding|Gene or Genome|Hospital Course|9019,9023|false|false|false|C1412433|AOX1 gene|AOx1
Drug|Biomedical or Dental Material|Hospital Course|9031,9039|false|false|false|C0168634|BaseLine dental cement|baseline
Finding|Idea or Concept|Hospital Course|9031,9039|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Finding|Classification|Hospital Course|9044,9050|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|Hospital Course|9044,9050|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|Hospital Course|9044,9050|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|Hospital Course|9044,9050|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Drug|Organic Chemical|Hospital Course|9082,9089|false|false|false|C0527315|Aricept|Aricept
Drug|Pharmacologic Substance|Hospital Course|9082,9089|false|false|false|C0527315|Aricept|Aricept
Drug|Organic Chemical|Hospital Course|9090,9097|false|false|false|C1330412|Namenda|Namenda
Drug|Pharmacologic Substance|Hospital Course|9090,9097|false|false|false|C1330412|Namenda|Namenda
Finding|Idea or Concept|Hospital Course|9102,9114|false|false|false|C1548597|Marketing basis - Transitional|TRANSITIONAL
Finding|Intellectual Product|Hospital Course|9150,9158|false|false|false|C4695111|ADMIN.FACILITY|facility
Finding|Intellectual Product|Hospital Course|9179,9185|false|false|false|C3244315|orders - HL7PublishingDomain|orders
Attribute|Clinical Attribute|Hospital Course|9191,9195|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|9191,9195|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|9191,9195|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9196,9203|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Finding|Sign or Symptom|Hospital Course|9196,9203|false|false|false|C0860603|Anxiety symptoms|anxiety
Finding|Body Substance|Hospital Course|9204,9214|false|false|false|C0036537|Bodily secretions|secretions
Finding|Functional Concept|Hospital Course|9225,9233|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Hospital Course|9225,9233|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Drug|Organic Chemical|Hospital Course|9248,9258|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|Hospital Course|9248,9258|false|false|false|C0025859|metoprolol|metoprolol
Drug|Organic Chemical|Hospital Course|9248,9268|false|false|false|C0724633|metoprolol succinate|metoprolol succinate
Drug|Pharmacologic Substance|Hospital Course|9248,9268|false|false|false|C0724633|metoprolol succinate|metoprolol succinate
Drug|Organic Chemical|Hospital Course|9259,9268|false|false|false|C0038617;C0220918|Succinates;succinate|succinate
Drug|Organic Chemical|Hospital Course|9273,9282|false|false|false|C0025242|memantine|Memantine
Drug|Pharmacologic Substance|Hospital Course|9273,9282|false|false|false|C0025242|memantine|Memantine
Drug|Organic Chemical|Hospital Course|9287,9296|false|false|false|C0527316|donepezil|donepezil
Drug|Pharmacologic Substance|Hospital Course|9287,9296|false|false|false|C0527316|donepezil|donepezil
Finding|Body Substance|Hospital Course|9301,9310|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|9301,9310|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|9301,9310|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|9301,9310|false|false|false|C0030685|Patient Discharge|discharge
Drug|Organic Chemical|Hospital Course|9315,9322|false|false|false|C1310585|Comfort brand of hydroxyethyl cellulose|comfort
Drug|Pharmacologic Substance|Hospital Course|9315,9322|false|false|false|C1310585|Comfort brand of hydroxyethyl cellulose|comfort
Finding|Mental Process|Hospital Course|9315,9322|false|false|false|C1331418|Comfort|comfort
Attribute|Clinical Attribute|Hospital Course|9346,9357|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Hospital Course|9346,9357|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|Hospital Course|9346,9357|false|false|false|C4284232|Medications|medications
Finding|Idea or Concept|Hospital Course|9385,9394|false|false|false|C1548438;C1549404|Patient Class - Inpatient;Referral category - Inpatient|inpatient
Procedure|Health Care Activity|Hospital Course|9385,9394|false|false|false|C1555324|inpatient encounter|inpatient
Procedure|Health Care Activity|Hospital Course|9395,9402|false|false|false|C0085555|Hospice Care|hospice
Attribute|Clinical Attribute|Hospital Course|9413,9417|false|false|false|C4255237||form
Finding|Functional Concept|Hospital Course|9413,9417|false|false|false|C1522492|Formation|form
Attribute|Clinical Attribute|Hospital Course|9419,9422|false|false|false|C4285234||DNR
Drug|Antibiotic|Hospital Course|9419,9422|false|false|false|C0011015|daunorubicin|DNR
Drug|Organic Chemical|Hospital Course|9419,9422|false|false|false|C0011015|daunorubicin|DNR
Finding|Finding|Hospital Course|9419,9422|false|false|false|C0079252;C0582114|Do not resuscitate status;Do-Not-Resuscitate Orders|DNR
Finding|Intellectual Product|Hospital Course|9419,9422|false|false|false|C0079252;C0582114|Do not resuscitate status;Do-Not-Resuscitate Orders|DNR
Event|Occupational Activity|Hospital Course|9454,9458|false|false|false|C0009219|Coding|CODE
Finding|Intellectual Product|Hospital Course|9454,9458|false|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|CODE
Attribute|Clinical Attribute|Hospital Course|9460,9463|false|false|false|C4285234||DNR
Drug|Antibiotic|Hospital Course|9460,9463|false|false|false|C0011015|daunorubicin|DNR
Drug|Organic Chemical|Hospital Course|9460,9463|false|false|false|C0011015|daunorubicin|DNR
Finding|Finding|Hospital Course|9460,9463|false|false|false|C0079252;C0582114|Do not resuscitate status;Do-Not-Resuscitate Orders|DNR
Finding|Intellectual Product|Hospital Course|9460,9463|false|false|false|C0079252;C0582114|Do not resuscitate status;Do-Not-Resuscitate Orders|DNR
Disorder|Disease or Syndrome|Hospital Course|9469,9472|false|false|false|C0410422|Chronic multifocal osteomyelitis|CMO
Event|Activity|Hospital Course|9476,9483|false|false|false|C3812666|Personal Contact|CONTACT
Finding|Functional Concept|Hospital Course|9476,9483|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Finding|Idea or Concept|Hospital Course|9476,9483|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Finding|Intellectual Product|Hospital Course|9476,9483|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Phenomenon|Phenomenon or Process|Hospital Course|9476,9483|false|false|false|C0392367|Physical contact|CONTACT
Disorder|Disease or Syndrome|Hospital Course|9485,9488|false|false|false|C0162531|Hereditary Coproporphyria|HCP
Finding|Gene or Genome|Hospital Course|9485,9488|false|false|false|C1335283;C1412376;C1413681;C1705637;C5780748|AMBP gene;AMBP wt Allele;CPOX gene;PTPN6 gene;PTPN6 wt Allele|HCP
Disorder|Neoplastic Process|Hospital Course|9518,9527|false|false|false|C0027627|Neoplasm Metastasis|secondary
Finding|Functional Concept|Hospital Course|9518,9527|false|false|false|C1522484|metastatic qualifier|secondary
Finding|Gene or Genome|Hospital Course|9533,9536|false|false|false|C1420310|SON gene|son
Attribute|Clinical Attribute|Hospital Course|9544,9555|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|9544,9555|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|Hospital Course|9544,9555|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|9544,9568|false|false|false|C1627937|Medications on admission|Medications on Admission
Procedure|Health Care Activity|Hospital Course|9559,9568|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|Hospital Course|9587,9597|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|Hospital Course|9587,9597|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|Hospital Course|9587,9602|false|false|false|C0746470|MEDICATION LIST|Medication list
Finding|Intellectual Product|Hospital Course|9598,9602|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Drug|Organic Chemical|Hospital Course|9619,9627|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|Hospital Course|9619,9627|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|Hospital Course|9619,9627|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Finding|Functional Concept|Hospital Course|9619,9627|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|Hospital Course|9619,9627|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Organic Chemical|Hospital Course|9632,9642|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|Hospital Course|9632,9642|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Organic Chemical|Hospital Course|9632,9652|false|false|false|C0724633|metoprolol succinate|Metoprolol Succinate
Drug|Pharmacologic Substance|Hospital Course|9632,9652|false|false|false|C0724633|metoprolol succinate|Metoprolol Succinate
Drug|Organic Chemical|Hospital Course|9643,9652|false|false|false|C0038617;C0220918|Succinates;succinate|Succinate
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9666,9669|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9666,9669|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|9666,9669|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|9666,9669|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|9674,9683|false|false|false|C0076840|torsemide|Torsemide
Drug|Pharmacologic Substance|Hospital Course|9674,9683|false|false|false|C0076840|torsemide|Torsemide
Drug|Organic Chemical|Hospital Course|9703,9710|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|Hospital Course|9703,9710|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|Hospital Course|9730,9739|false|false|false|C0527316|donepezil|Donepezil
Drug|Pharmacologic Substance|Hospital Course|9730,9739|false|false|false|C0527316|donepezil|Donepezil
Drug|Organic Chemical|Hospital Course|9757,9767|false|false|false|C0244404|raloxifene|raloxifene
Drug|Pharmacologic Substance|Hospital Course|9757,9767|false|false|false|C0244404|raloxifene|raloxifene
Anatomy|Body Space or Junction|Hospital Course|9774,9778|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|9774,9778|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|9774,9778|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|9774,9778|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Drug|Organic Chemical|Hospital Course|9789,9802|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|Hospital Course|9789,9802|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|Hospital Course|9789,9802|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Biomedical or Dental Material|Hospital Course|9805,9808|false|false|false|C0039225|Tablet Dosage Form|TAB
Drug|Organic Chemical|Hospital Course|9822,9829|false|false|false|C1330412|Namenda|Namenda
Drug|Pharmacologic Substance|Hospital Course|9822,9829|false|false|false|C1330412|Namenda|Namenda
Drug|Organic Chemical|Hospital Course|9822,9832|false|false|false|C1330412|Namenda|Namenda XR
Drug|Pharmacologic Substance|Hospital Course|9822,9832|false|false|false|C1330412|Namenda|Namenda XR
Drug|Organic Chemical|Hospital Course|9834,9843|false|false|false|C0025242|memantine|MEMAntine
Drug|Pharmacologic Substance|Hospital Course|9834,9843|false|false|false|C0025242|memantine|MEMAntine
Anatomy|Body Space or Junction|Hospital Course|9851,9855|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|9851,9855|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|9851,9855|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|9851,9855|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Drug|Organic Chemical|Hospital Course|9866,9879|false|false|false|C0003968|ascorbic acid|Ascorbic Acid
Drug|Pharmacologic Substance|Hospital Course|9866,9879|false|false|false|C0003968|ascorbic acid|Ascorbic Acid
Drug|Vitamin|Hospital Course|9866,9879|false|false|false|C0003968|ascorbic acid|Ascorbic Acid
Procedure|Laboratory Procedure|Hospital Course|9866,9879|false|false|false|C0201898|Ascorbic acid measurement|Ascorbic Acid
Drug|Biologically Active Substance|Hospital Course|9900,9907|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|Hospital Course|9900,9907|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|Hospital Course|9900,9907|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|Hospital Course|9900,9907|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|Hospital Course|9900,9907|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Finding|Physiologic Function|Hospital Course|9900,9907|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|Hospital Course|9900,9907|false|false|false|C0201925|Calcium measurement|Calcium
Drug|Inorganic Chemical|Hospital Course|9900,9917|false|false|false|C0006681|calcium carbonate|Calcium Carbonate
Drug|Pharmacologic Substance|Hospital Course|9900,9917|false|false|false|C0006681|calcium carbonate|Calcium Carbonate
Drug|Element, Ion, or Isotope|Hospital Course|9908,9917|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|Carbonate
Drug|Organic Chemical|Hospital Course|9908,9917|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|Carbonate
Drug|Pharmacologic Substance|Hospital Course|9908,9917|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|Carbonate
Drug|Organic Chemical|Hospital Course|9940,9947|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|Hospital Course|9940,9947|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|Hospital Course|9940,9947|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|Hospital Course|9940,9949|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|Hospital Course|9940,9949|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|Hospital Course|9940,9949|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|Hospital Course|9940,9949|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|Hospital Course|9940,9949|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Drug|Food|Hospital Course|9974,9978|false|false|false|C3257082;C4521129|Fish (substance);Fish extract|Fish
Drug|Organic Chemical|Hospital Course|9974,9978|false|false|false|C3257082;C4521129|Fish (substance);Fish extract|Fish
Finding|Gene or Genome|Hospital Course|9974,9978|false|false|false|C1822711;C3274826|SH3PXD2A gene;SH3PXD2A wt Allele|Fish
Procedure|Molecular Biology Research Technique|Hospital Course|9974,9978|false|false|false|C0162789|Fluorescent in Situ Hybridization|Fish
Drug|Organic Chemical|Hospital Course|9974,9982|false|false|false|C0016157|fish oils|Fish Oil
Drug|Pharmacologic Substance|Hospital Course|9974,9982|false|false|false|C0016157|fish oils|Fish Oil
Drug|Biomedical or Dental Material|Hospital Course|9979,9982|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|Oil
Drug|Food|Hospital Course|9979,9982|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|Oil
Drug|Organic Chemical|Hospital Course|9979,9982|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|Oil
Drug|Pharmacologic Substance|Hospital Course|9979,9982|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|Oil
Finding|Intellectual Product|Hospital Course|9984,9989|false|false|false|C1719844|Omega|Omega
Drug|Biologically Active Substance|Hospital Course|9984,9991|false|false|false|C0015689|omega-3 fatty acids|Omega 3
Drug|Organic Chemical|Hospital Course|9984,9991|false|false|false|C0015689|omega-3 fatty acids|Omega 3
Drug|Pharmacologic Substance|Hospital Course|9984,9991|false|false|false|C0015689|omega-3 fatty acids|Omega 3
Finding|Body Substance|Hospital Course|10014,10023|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|10014,10023|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|10014,10023|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|10014,10023|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|10014,10035|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|10024,10035|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|10024,10035|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|Hospital Course|10024,10035|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Hospital Course|10040,10049|false|false|false|C0527316|donepezil|Donepezil
Drug|Pharmacologic Substance|Hospital Course|10040,10049|false|false|false|C0527316|donepezil|Donepezil
Drug|Organic Chemical|Hospital Course|10067,10077|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|Hospital Course|10067,10077|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Organic Chemical|Hospital Course|10067,10087|false|false|false|C0724633|metoprolol succinate|Metoprolol Succinate
Drug|Pharmacologic Substance|Hospital Course|10067,10087|false|false|false|C0724633|metoprolol succinate|Metoprolol Succinate
Drug|Organic Chemical|Hospital Course|10078,10087|false|false|false|C0038617;C0220918|Succinates;succinate|Succinate
Drug|Organic Chemical|Hospital Course|10111,10118|false|false|false|C1330412|Namenda|Namenda
Drug|Pharmacologic Substance|Hospital Course|10111,10118|false|false|false|C1330412|Namenda|Namenda
Drug|Organic Chemical|Hospital Course|10111,10121|false|false|false|C1330412|Namenda|Namenda XR
Drug|Pharmacologic Substance|Hospital Course|10111,10121|false|false|false|C1330412|Namenda|Namenda XR
Drug|Organic Chemical|Hospital Course|10123,10132|false|false|false|C0025242|memantine|MEMAntine
Drug|Pharmacologic Substance|Hospital Course|10123,10132|false|false|false|C0025242|memantine|MEMAntine
Anatomy|Body Space or Junction|Hospital Course|10140,10144|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|10140,10144|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|10140,10144|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|10140,10144|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Drug|Organic Chemical|Hospital Course|10155,10168|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Hospital Course|10155,10168|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Procedure|Laboratory Procedure|Hospital Course|10155,10168|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Drug|Organic Chemical|Hospital Course|10188,10202|true|false|false|C0017970|glycopyrrolate|Glycopyrrolate
Drug|Pharmacologic Substance|Hospital Course|10188,10202|true|false|false|C0017970|glycopyrrolate|Glycopyrrolate
Finding|Gene or Genome|Hospital Course|10217,10220|false|false|false|C1422467|CIAO3 gene|PRN
Finding|Body Substance|Hospital Course|10228,10238|false|false|false|C0036537|Bodily secretions|secretions
Drug|Organic Chemical|Hospital Course|10243,10254|false|false|false|C0596004|hyoscyamine|Hyoscyamine
Drug|Pharmacologic Substance|Hospital Course|10243,10254|false|false|false|C0596004|hyoscyamine|Hyoscyamine
Finding|Gene or Genome|Hospital Course|10271,10274|false|false|false|C1422467|CIAO3 gene|PRN
Finding|Body Substance|Hospital Course|10282,10292|false|false|false|C0036537|Bodily secretions|secretions
Finding|Body Substance|Hospital Course|10298,10307|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|10298,10307|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|10298,10307|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|10298,10307|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|10298,10319|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|10298,10319|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|10308,10319|false|false|false|C2926604||Disposition
Procedure|Health Care Activity|Hospital Course|10308,10319|false|false|false|C0184758|Patient disposition|Disposition
Finding|Finding|Hospital Course|10321,10329|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|10321,10329|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Procedure|Health Care Activity|Hospital Course|10321,10334|false|false|false|C0023977|long-term care|Extended Care
Event|Activity|Hospital Course|10330,10334|false|false|false|C1947933|care activity|Care
Finding|Finding|Hospital Course|10330,10334|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|Hospital Course|10330,10334|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|Hospital Course|10337,10345|false|false|false|C4695111|ADMIN.FACILITY|Facility
Finding|Body Substance|Hospital Course|10353,10362|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|10353,10362|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|10353,10362|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|10353,10362|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|10353,10372|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|10363,10372|false|false|false|C0945731||Diagnosis
Finding|Classification|Hospital Course|10363,10372|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|10363,10372|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|10363,10372|false|false|false|C0011900|Diagnosis|Diagnosis
Attribute|Clinical Attribute|Principle Diagnosis|10411,10415|false|false|false|C4318566|Deep Resection Margin|Deep
Anatomy|Body Part, Organ, or Organ Component|Principle Diagnosis|10411,10420|false|false|false|C0226514|Structure of deep vein|Deep Vein
Disorder|Disease or Syndrome|Principle Diagnosis|10411,10431|false|false|false|C0149871;C0340708|Deep Vein Thrombosis;Deep vein thrombosis of lower limb|Deep Vein Thrombosis
Anatomy|Body Part, Organ, or Organ Component|Principle Diagnosis|10416,10420|false|false|false|C0042449|Veins|Vein
Finding|Pathologic Function|Principle Diagnosis|10416,10431|false|false|false|C0042487|Venous Thrombosis|Vein Thrombosis
Finding|Pathologic Function|Principle Diagnosis|10421,10431|false|false|false|C0040053|Thrombosis|Thrombosis
Disorder|Neoplastic Process|Principle Diagnosis|10436,10445|false|false|false|C0027627|Neoplasm Metastasis|Secondary
Finding|Functional Concept|Principle Diagnosis|10436,10445|false|false|false|C1522484|metastatic qualifier|Secondary
Attribute|Clinical Attribute|Principle Diagnosis|10436,10455|false|false|false|C4255018||Secondary Diagnosis
Finding|Finding|Principle Diagnosis|10436,10455|false|false|false|C0332138|Secondary diagnosis|Secondary Diagnosis
Attribute|Clinical Attribute|Principle Diagnosis|10446,10455|false|false|false|C0945731||Diagnosis
Finding|Classification|Principle Diagnosis|10446,10455|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Principle Diagnosis|10446,10455|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Principle Diagnosis|10446,10455|false|false|false|C0011900|Diagnosis|Diagnosis
Disorder|Disease or Syndrome|Principle Diagnosis|10478,10502|false|false|false|C0018802|Congestive heart failure|Congestive heart failure
Anatomy|Body Part, Organ, or Organ Component|Principle Diagnosis|10489,10494|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Principle Diagnosis|10489,10494|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Principle Diagnosis|10489,10494|false|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|Principle Diagnosis|10489,10502|false|false|false|C0018801;C0018802|Congestive heart failure;Heart failure|heart failure
Finding|Functional Concept|Principle Diagnosis|10495,10502|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|Principle Diagnosis|10495,10502|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|Principle Diagnosis|10495,10502|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Anatomy|Body Part, Organ, or Organ Component|Principle Diagnosis|10504,10510|false|false|false|C0018792|Heart Atrium|Atrial
Attribute|Clinical Attribute|Principle Diagnosis|10504,10523|false|false|false|C2926591||Atrial fibrillation
Disorder|Disease or Syndrome|Principle Diagnosis|10504,10523|false|false|false|C0004238|Atrial Fibrillation|Atrial fibrillation
Lab|Laboratory or Test Result|Principle Diagnosis|10504,10523|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Atrial fibrillation
Disorder|Disease or Syndrome|Principle Diagnosis|10511,10523|false|false|false|C0232197|Fibrillation|fibrillation
Finding|Sign or Symptom|Principle Diagnosis|10526,10538|false|false|false|C0009806|Constipation|Constipation
Disorder|Disease or Syndrome|Principle Diagnosis|10541,10553|false|false|false|C0162429|Malnutrition|Malnutrition
Disorder|Disease or Syndrome|Principle Diagnosis|10556,10568|false|false|false|C0020538|Hypertensive disease|Hypertension
Disorder|Disease or Syndrome|Principle Diagnosis|10571,10580|false|false|false|C0002395|Alzheimer's Disease|Alzheimer
Disorder|Disease or Syndrome|Principle Diagnosis|10571,10591|false|false|false|C0002395|Alzheimer's Disease|Alzheimer's dementia
Disorder|Mental or Behavioral Dysfunction|Principle Diagnosis|10583,10591|false|false|false|C0011265;C0497327|Dementia;Presenile dementia|dementia
Finding|Mental Process|Discharge Condition|10618,10624|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|10618,10631|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|10618,10631|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|10625,10631|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|10625,10631|false|false|false|C1546481|What subject filter - Status|Status
Disorder|Mental or Behavioral Dysfunction|Discharge Condition|10633,10641|false|false|false|C0009676|Confusion|Confused
Finding|Finding|Discharge Condition|10633,10641|false|false|false|C0683369;C1547301|Clouded consciousness;Precaution Code - Confused|Confused
Finding|Intellectual Product|Discharge Condition|10633,10641|false|false|false|C0683369;C1547301|Clouded consciousness;Precaution Code - Confused|Confused
Finding|Finding|Discharge Condition|10644,10650|false|false|false|C1549493;C3812891|All of the Time;Always - AcknowledgementCondition|always
Finding|Idea or Concept|Discharge Condition|10644,10650|false|false|false|C1549493;C3812891|All of the Time;Always - AcknowledgementCondition|always
Attribute|Clinical Attribute|Discharge Condition|10652,10674|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|10652,10674|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Finding|Finding|Discharge Condition|10661,10674|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|10661,10674|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|10676,10681|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|10676,10681|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|10676,10681|false|false|false|C0718338|Alert brand of caffeine|Alert
Finding|Finding|Discharge Condition|10676,10681|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|10676,10681|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|10676,10681|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|10686,10697|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|10699,10707|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|10699,10707|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|10699,10707|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|10708,10714|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|10708,10714|false|false|false|C1546481|What subject filter - Status|Status
Disorder|Disease or Syndrome|Discharge Condition|10723,10726|false|false|false|C3159311|BORNHOLM EYE DISEASE|Bed
Finding|Intellectual Product|Discharge Condition|10723,10726|false|false|false|C2346952|Bachelor of Education|Bed
Finding|Social Behavior|Discharge Condition|10732,10742|false|false|false|C0018896|Helping Behavior|assistance
Finding|Finding|Discharge Condition|10756,10766|false|false|false|C2135586;C4321408|Wheelchair Usually Used;has wheelchair at home (history)|wheelchair
Finding|Gene or Genome|Discharge Instructions|10795,10799|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Finding|Intellectual Product|Discharge Instructions|10816,10824|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|Discharge Instructions|10816,10824|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|Discharge Instructions|10832,10836|false|false|false|C1947933|care activity|care
Finding|Finding|Discharge Instructions|10832,10836|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|10832,10836|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|10832,10839|false|false|false|C1555558|care of - AddressPartType|care of
Procedure|Health Care Activity|Discharge Instructions|10857,10872|false|false|false|C0019993|Hospitalization|hospitalization
Finding|Functional Concept|Discharge Instructions|10910,10915|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|Discharge Instructions|10910,10919|false|false|false|C0524470|Right hip region structure|right hip
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|10916,10919|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|hip
Drug|Amino Acid, Peptide, or Protein|Discharge Instructions|10916,10919|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Biologically Active Substance|Discharge Instructions|10916,10919|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Pharmacologic Substance|Discharge Instructions|10916,10919|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Finding|Gene or Genome|Discharge Instructions|10916,10919|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|hip
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|10916,10919|false|false|false|C1292890|Procedure on hip|hip
Attribute|Clinical Attribute|Discharge Instructions|10921,10925|false|false|false|C2598155||pain
Finding|Functional Concept|Discharge Instructions|10921,10925|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|10921,10925|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Phenomenon|Natural Phenomenon or Process|Discharge Instructions|10934,10939|false|false|false|C0043309|Roentgen Rays|Xrays
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|10948,10951|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|hip
Drug|Amino Acid, Peptide, or Protein|Discharge Instructions|10948,10951|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Biologically Active Substance|Discharge Instructions|10948,10951|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Pharmacologic Substance|Discharge Instructions|10948,10951|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Finding|Gene or Genome|Discharge Instructions|10948,10951|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|hip
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|10948,10951|false|false|false|C1292890|Procedure on hip|hip
Disorder|Injury or Poisoning|Discharge Instructions|10975,10984|true|false|false|C0016658|Fracture|fractures
Finding|Finding|Discharge Instructions|10975,10984|true|false|false|C4554413|Fractured|fractures
Disorder|Disease or Syndrome|Discharge Instructions|11003,11008|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|Discharge Instructions|11003,11008|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Pathologic Function|Discharge Instructions|11003,11013|false|false|false|C0087086;C0302148|Blood Clot;Thrombus|blood clot
Drug|Organic Chemical|Discharge Instructions|11009,11013|false|false|false|C0009074|clotrimazole|clot
Drug|Pharmacologic Substance|Discharge Instructions|11009,11013|false|false|false|C0009074|clotrimazole|clot
Finding|Pathologic Function|Discharge Instructions|11009,11013|false|false|false|C0302148|Blood Clot|clot
Finding|Functional Concept|Discharge Instructions|11022,11026|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|11022,11030|false|false|false|C0230416;C0230443|Left lower extremity;Structure of left lower leg|left leg
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|11027,11030|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|11054,11059|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Discharge Instructions|11054,11059|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Discharge Instructions|11054,11059|false|false|false|C0795691|HEART PROBLEM|heart
Finding|Classification|Discharge Instructions|11122,11128|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|Discharge Instructions|11122,11128|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|Discharge Instructions|11122,11128|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|Discharge Instructions|11122,11128|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Gene or Genome|Discharge Instructions|11203,11207|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Finding|Intellectual Product|Discharge Instructions|11203,11207|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Event|Activity|Discharge Instructions|11211,11215|false|false|false|C1947933|care activity|care
Finding|Finding|Discharge Instructions|11211,11215|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|11211,11215|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Drug|Organic Chemical|Discharge Instructions|11272,11279|false|false|false|C1310585|Comfort brand of hydroxyethyl cellulose|comfort
Drug|Pharmacologic Substance|Discharge Instructions|11272,11279|false|false|false|C1310585|Comfort brand of hydroxyethyl cellulose|comfort
Finding|Mental Process|Discharge Instructions|11272,11279|false|false|false|C1331418|Comfort|comfort
Procedure|Health Care Activity|Discharge Instructions|11335,11342|false|false|false|C0085555|Hospice Care|hospice
Finding|Finding|Discharge Instructions|11335,11347|false|false|false|C0869461|Encounter for Hospice Care|hospice care
Procedure|Health Care Activity|Discharge Instructions|11335,11347|false|false|false|C0085555|Hospice Care|hospice care
Event|Activity|Discharge Instructions|11343,11347|false|false|false|C1947933|care activity|care
Finding|Finding|Discharge Instructions|11343,11347|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|11343,11347|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Classification|Discharge Instructions|11374,11380|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|Discharge Instructions|11374,11380|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|Discharge Instructions|11374,11380|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|Discharge Instructions|11374,11380|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|Discharge Instructions|11401,11410|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|Treatment
Finding|Functional Concept|Discharge Instructions|11401,11410|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|Treatment
Procedure|Health Care Activity|Discharge Instructions|11401,11410|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|Treatment
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|11401,11410|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|Treatment
Procedure|Health Care Activity|Discharge Instructions|11419,11427|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|11428,11440|false|false|false|C3263700||Instructions
Finding|Intellectual Product|Discharge Instructions|11428,11440|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

