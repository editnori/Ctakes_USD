 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|46,55|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|46,55|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|46,60|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|80,89|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|80,89|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|80,94|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|136,139|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|147,154|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|147,154|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|156,164|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|SIMPLE_SEGMENT|167,176|false|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|167,176|false|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|167,176|false|false|false|C0020517|Hypersensitivity|Allergies
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|179,189|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|179,189|false|false|false|C0065374|lisinopril|lisinopril
Event|Event|SIMPLE_SEGMENT|179,189|false|false|false|||lisinopril
Event|Event|SIMPLE_SEGMENT|192,201|false|false|false|||Attending
Finding|Functional Concept|SIMPLE_SEGMENT|192,201|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|SIMPLE_SEGMENT|209,224|false|false|false|C0277786|Chief complaint (finding)|Chief Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|215,224|false|false|false|C3864418||Complaint
Event|Event|SIMPLE_SEGMENT|215,224|false|false|false|||Complaint
Finding|Finding|SIMPLE_SEGMENT|215,224|false|false|false|C5441521|Complaint (finding)|Complaint
Anatomy|Body Location or Region|SIMPLE_SEGMENT|226,231|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|SIMPLE_SEGMENT|226,231|false|false|false|C0741025|Chest problem|Chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|226,236|false|false|false|C2926613||Chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|226,236|false|false|false|C0008031|Chest Pain|Chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|232,236|false|true|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|232,236|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|232,236|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|232,236|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Classification|SIMPLE_SEGMENT|239,244|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|SIMPLE_SEGMENT|245,253|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|245,253|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|257,275|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|266,275|false|false|false|C0945766||Procedure
Event|Event|SIMPLE_SEGMENT|266,275|false|false|false|||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|266,275|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|266,275|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|266,275|false|false|false|C0184661|Interventional procedure|Procedure
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|277,284|false|false|false|C0018787|Heart|Cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|277,284|false|false|false|C1314974|Cardiac attachment|Cardiac
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|277,289|false|false|false|C0018795|Cardiac Catheterization Procedures|Cardiac cath
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|285,289|false|false|false|C0007430|Catheterization|cath
Finding|Finding|SIMPLE_SEGMENT|299,319|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Event|Event|SIMPLE_SEGMENT|304,311|false|false|false|||Medical
Finding|Functional Concept|SIMPLE_SEGMENT|304,311|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|304,311|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|304,311|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|304,311|false|false|false|C0199168|Medical service|Medical
Finding|Finding|SIMPLE_SEGMENT|304,319|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|312,319|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|312,319|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|312,319|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|322,326|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|322,326|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|SIMPLE_SEGMENT|322,326|false|false|false|||COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|322,326|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|328,331|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|328,331|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|328,331|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|328,331|false|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|328,331|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|328,331|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|328,331|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|328,331|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|336,339|false|false|false|C0006430|Burning Mouth Syndrome|BMS
Event|Event|SIMPLE_SEGMENT|336,339|false|false|false|||BMS
Attribute|Clinical Attribute|SIMPLE_SEGMENT|340,348|false|false|false|C4489236|Proximal Resection Margin|proximal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|349,352|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|349,352|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|349,352|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|358,361|false|false|false|C4551552|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|DES
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|358,361|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Biologically Active Substance|SIMPLE_SEGMENT|358,361|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Hormone|SIMPLE_SEGMENT|358,361|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Organic Chemical|SIMPLE_SEGMENT|358,361|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|358,361|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Event|Event|SIMPLE_SEGMENT|358,361|false|false|false|||DES
Finding|Gene or Genome|SIMPLE_SEGMENT|358,361|false|false|false|C1413980|DES gene|DES
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|369,372|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|369,372|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|SIMPLE_SEGMENT|369,372|false|false|false|||LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|369,372|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|378,381|false|false|false|C4551552|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|DES
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|378,381|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Biologically Active Substance|SIMPLE_SEGMENT|378,381|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Hormone|SIMPLE_SEGMENT|378,381|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Organic Chemical|SIMPLE_SEGMENT|378,381|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|378,381|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Event|Event|SIMPLE_SEGMENT|378,381|false|false|false|||DES
Finding|Gene or Genome|SIMPLE_SEGMENT|378,381|false|false|false|C1413980|DES gene|DES
Event|Event|SIMPLE_SEGMENT|385,389|false|false|false|||edge
Finding|Conceptual Entity|SIMPLE_SEGMENT|385,389|false|false|false|C2697523|Graph Edge|edge
Event|Event|SIMPLE_SEGMENT|391,394|false|false|false|||ISR
Finding|Cell Function|SIMPLE_SEGMENT|391,394|false|false|false|C5445058|integrated stress response signaling|ISR
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|402,405|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|402,405|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|402,405|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|406,409|false|false|false|C4551552|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|DES
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|406,409|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Biologically Active Substance|SIMPLE_SEGMENT|406,409|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Hormone|SIMPLE_SEGMENT|406,409|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Organic Chemical|SIMPLE_SEGMENT|406,409|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|406,409|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Event|Event|SIMPLE_SEGMENT|406,409|false|false|false|||DES
Finding|Gene or Genome|SIMPLE_SEGMENT|406,409|false|false|false|C1413980|DES gene|DES
Event|Event|SIMPLE_SEGMENT|414,422|false|false|false|||stenosis
Finding|Pathologic Function|SIMPLE_SEGMENT|414,422|false|false|false|C1261287|Stenosis|stenosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|423,429|false|false|false|C4522154|Distal Resection Margin|distal
Event|Event|SIMPLE_SEGMENT|433,438|false|false|false|||stent
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|444,447|false|false|false|C4551552|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|DES
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|444,447|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Biologically Active Substance|SIMPLE_SEGMENT|444,447|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Hormone|SIMPLE_SEGMENT|444,447|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Organic Chemical|SIMPLE_SEGMENT|444,447|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|444,447|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Event|Event|SIMPLE_SEGMENT|444,447|false|false|false|||DES
Finding|Gene or Genome|SIMPLE_SEGMENT|444,447|false|false|false|C1413980|DES gene|DES
Event|Event|SIMPLE_SEGMENT|469,473|false|false|false|||CABG
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|469,473|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|479,482|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|479,482|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|SIMPLE_SEGMENT|479,482|false|false|false|||LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|479,482|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|507,517|false|false|false|C0011570;C0011581;C0344315;C0812393|Cancer patients and suicide and depression;Depressed mood;Depressive disorder;Mental Depression|Depression
Event|Event|SIMPLE_SEGMENT|507,517|false|false|false|||Depression
Finding|Functional Concept|SIMPLE_SEGMENT|507,517|false|false|false|C0460137;C1579931|Depression - motion|Depression
Finding|Sign or Symptom|SIMPLE_SEGMENT|507,517|false|false|false|C0460137;C1579931|Depression - motion|Depression
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|527,531|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Event|Event|SIMPLE_SEGMENT|527,531|false|false|false|||GERD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|535,547|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|SIMPLE_SEGMENT|535,547|false|false|false|||Hypertension
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|549,558|false|false|false|C0149931|Migraine Disorders|Migraines
Event|Event|SIMPLE_SEGMENT|549,558|false|false|false|||Migraines
Finding|Intellectual Product|SIMPLE_SEGMENT|560,567|false|false|false|C1547296|Chronic - Admission Level of Care Code|Chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|560,567|false|false|false|C1555457|Provision of recurring care for chronic illness|Chronic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|560,581|false|false|false|C0748678|shoulder pain chronic|Chronic shoulder pain
Anatomy|Body Location or Region|SIMPLE_SEGMENT|568,576|false|false|false|C0037004;C4299050|Shoulder;Upper extremity>Shoulder|shoulder
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|568,576|false|false|false|C0221590;C0869975|Examination of shoulder(s);Procedures on Shoulder|shoulder
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|568,576|false|false|false|C0221590;C0869975|Examination of shoulder(s);Procedures on Shoulder|shoulder
Finding|Sign or Symptom|SIMPLE_SEGMENT|568,581|false|false|false|C0037011|Shoulder Pain|shoulder pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|577,581|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|577,581|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|577,581|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|577,581|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|585,594|false|false|false|C0027415|Narcotics|narcotics
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|585,594|false|false|false|C0027415|Narcotics|narcotics
Event|Event|SIMPLE_SEGMENT|585,594|false|false|false|||narcotics
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|596,599|false|false|false|C0520679|Sleep Apnea, Obstructive|OSA
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|596,599|false|false|false|C0764906|OSA protein, Drosophila|OSA
Drug|Biologically Active Substance|SIMPLE_SEGMENT|596,599|false|false|false|C0764906|OSA protein, Drosophila|OSA
Event|Event|SIMPLE_SEGMENT|596,599|false|false|false|||OSA
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|601,622|false|false|false|C0031117;C4721453|Peripheral Nervous System Diseases;Peripheral Neuropathy|Peripheral neuropathy
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|612,622|false|false|false|C0442874|Neuropathy|neuropathy
Event|Event|SIMPLE_SEGMENT|612,622|false|false|false|||neuropathy
Finding|Sign or Symptom|SIMPLE_SEGMENT|624,632|false|false|false|C0085631;C3887611|Agitation;Restlessness|Restless
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|624,636|false|false|false|C0035258|Restless Legs Syndrome|Restless leg
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|633,636|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Finding|Functional Concept|SIMPLE_SEGMENT|639,645|false|false|false|C0728831|Social|Social
Finding|Finding|SIMPLE_SEGMENT|639,653|false|false|false|C0424945;C3714536|Social History;Social and personal history|Social History
Event|Event|SIMPLE_SEGMENT|646,653|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|646,653|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|646,653|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|646,653|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Classification|SIMPLE_SEGMENT|659,665|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|SIMPLE_SEGMENT|659,665|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|SIMPLE_SEGMENT|659,665|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|SIMPLE_SEGMENT|659,665|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Finding|SIMPLE_SEGMENT|659,673|false|false|false|C0241889|Family Medical History|Family History
Event|Event|SIMPLE_SEGMENT|666,673|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|666,673|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|666,673|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|666,673|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Body Substance|SIMPLE_SEGMENT|675,682|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|675,682|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|675,682|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|687,691|true|false|false|||ward
Finding|Functional Concept|SIMPLE_SEGMENT|699,704|true|false|false|C1442792|State|state
Event|Event|SIMPLE_SEGMENT|714,718|true|false|false|||know
Event|Event|SIMPLE_SEGMENT|724,731|true|false|false|||details
Finding|Classification|SIMPLE_SEGMENT|736,742|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|736,742|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|736,742|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|736,742|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Finding|SIMPLE_SEGMENT|736,750|true|false|false|C0241889|Family Medical History|family history
Event|Event|SIMPLE_SEGMENT|743,750|true|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|743,750|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|743,750|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|743,750|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Event|Event|SIMPLE_SEGMENT|752,758|false|false|false|||Mother
Finding|Idea or Concept|SIMPLE_SEGMENT|752,758|false|false|false|C1546508|Relationship - Mother|Mother
Finding|Finding|SIMPLE_SEGMENT|764,772|false|false|false|C0332149|Possible|possible
Drug|Organic Chemical|SIMPLE_SEGMENT|773,780|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|773,780|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Event|Event|SIMPLE_SEGMENT|773,780|false|false|false|||alcohol
Finding|Intellectual Product|SIMPLE_SEGMENT|773,780|false|false|false|C1547288|Alcohol - Recreational Drug Use Code|alcohol
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|773,786|false|true|false|C0085762|Alcohol abuse|alcohol abuse
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|781,786|false|false|false|C0013146|Drug abuse|abuse
Event|Event|SIMPLE_SEGMENT|781,786|false|false|false|||abuse
Event|Event|SIMPLE_SEGMENT|781,786|false|false|false|C1546935|Abuse|abuse
Finding|Finding|SIMPLE_SEGMENT|781,786|false|false|false|C0562381|Victim of abuse (finding)|abuse
Finding|Conceptual Entity|SIMPLE_SEGMENT|788,794|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Idea or Concept|SIMPLE_SEGMENT|788,794|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Event|Event|SIMPLE_SEGMENT|796,804|false|false|false|||deceased
Finding|Finding|SIMPLE_SEGMENT|796,804|false|false|false|C0011065;C1549464;C1704456|Cessation of life;Deceased - ActIneligibilityReason;Deceased - Military Status|deceased
Finding|Organism Function|SIMPLE_SEGMENT|796,804|false|false|false|C0011065;C1549464;C1704456|Cessation of life;Deceased - ActIneligibilityReason;Deceased - Military Status|deceased
Disorder|Neoplastic Process|SIMPLE_SEGMENT|817,824|false|false|false|C0019829|Hodgkin Disease|Hodgkin
Disorder|Neoplastic Process|SIMPLE_SEGMENT|817,834|false|false|false|C0019829|Hodgkin Disease|Hodgkin's Disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|827,834|false|false|false|C0012634|Disease|Disease
Event|Event|SIMPLE_SEGMENT|827,834|false|false|false|||Disease
Event|Event|SIMPLE_SEGMENT|843,850|false|false|false|||records
Finding|Idea or Concept|SIMPLE_SEGMENT|843,850|false|false|false|C0034869;C1548330|Quantity limited request - Records;Records|records
Finding|Intellectual Product|SIMPLE_SEGMENT|843,850|false|false|false|C0034869;C1548330|Quantity limited request - Records;Records|records
Event|Event|SIMPLE_SEGMENT|854,862|false|false|false|||Physical
Finding|Finding|SIMPLE_SEGMENT|854,862|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|854,862|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|854,862|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|854,867|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|854,867|false|false|false|C0031809|Physical Examination|Physical Exam
Event|Event|SIMPLE_SEGMENT|863,867|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|863,867|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|863,867|false|false|false|C0582103|Medical Examination|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|869,878|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|SIMPLE_SEGMENT|879,883|false|false|false|||EXAM
Finding|Functional Concept|SIMPLE_SEGMENT|879,883|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|SIMPLE_SEGMENT|879,883|false|false|false|C0582103|Medical Examination|EXAM
Event|Event|SIMPLE_SEGMENT|899,906|false|false|false|||GENERAL
Finding|Classification|SIMPLE_SEGMENT|899,906|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|899,906|false|false|false|C3812897|General medical service|GENERAL
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|907,910|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|907,910|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|907,910|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|907,910|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|907,910|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|SIMPLE_SEGMENT|907,910|false|false|false|||NAD
Finding|Finding|SIMPLE_SEGMENT|907,910|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Event|Event|SIMPLE_SEGMENT|916,924|false|false|false|||Pleasant
Finding|Mental Process|SIMPLE_SEGMENT|916,924|false|false|false|C2987187|Pleasant|Pleasant
Anatomy|Body Location or Region|SIMPLE_SEGMENT|933,938|false|false|false|C1512338|HEENT|HEENT
Event|Event|SIMPLE_SEGMENT|940,944|false|false|false|||NCAT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|946,952|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|946,952|false|false|false|C0036412|Scleral Diseases|Sclera
Event|Event|SIMPLE_SEGMENT|946,952|false|false|false|||Sclera
Procedure|Health Care Activity|SIMPLE_SEGMENT|946,952|false|false|false|C2228481|examination of sclera|Sclera
Event|Event|SIMPLE_SEGMENT|953,962|false|false|false|||anicteric
Finding|Finding|SIMPLE_SEGMENT|953,962|false|false|false|C0205180|Anicteric|anicteric
Event|Event|SIMPLE_SEGMENT|964,969|false|false|false|||PERRL
Finding|Finding|SIMPLE_SEGMENT|964,969|false|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Event|Event|SIMPLE_SEGMENT|971,975|false|false|false|||EOMI
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|977,988|true|false|false|C0009758;C0229274|Structure of palpebral conjunctiva;conjunctiva|Conjunctiva
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|977,988|true|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|Conjunctiva
Disorder|Neoplastic Process|SIMPLE_SEGMENT|977,988|true|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|Conjunctiva
Event|Event|SIMPLE_SEGMENT|977,988|true|false|false|||Conjunctiva
Finding|Body Substance|SIMPLE_SEGMENT|977,988|true|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|Conjunctiva
Finding|Intellectual Product|SIMPLE_SEGMENT|977,988|true|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|Conjunctiva
Procedure|Health Care Activity|SIMPLE_SEGMENT|977,988|true|false|false|C0872390;C2228431|Procedure on conjunctiva;examination of conjunctiva|Conjunctiva
Event|Event|SIMPLE_SEGMENT|999,1005|true|false|false|||pallor
Finding|Finding|SIMPLE_SEGMENT|999,1005|true|false|false|C0241137|Pallor of skin|pallor
Event|Event|SIMPLE_SEGMENT|1009,1017|true|false|false|||cyanosis
Finding|Sign or Symptom|SIMPLE_SEGMENT|1009,1017|true|false|false|C0010520|Cyanosis|cyanosis
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|1025,1029|true|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|1025,1029|true|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|1025,1029|true|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|1025,1029|true|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1025,1036|true|false|false|C0026639|Oral mucous membrane structure|oral mucosa
Anatomy|Tissue|SIMPLE_SEGMENT|1030,1036|false|false|false|C0026724|Mucous Membrane|mucosa
Finding|Intellectual Product|SIMPLE_SEGMENT|1030,1036|false|false|false|C1561514||mucosa
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1037,1041|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|SIMPLE_SEGMENT|1037,1041|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|SIMPLE_SEGMENT|1037,1041|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Event|Event|SIMPLE_SEGMENT|1043,1049|true|false|false|||Supple
Finding|Functional Concept|SIMPLE_SEGMENT|1043,1049|true|false|false|C0332254|Supple|Supple
Event|Event|SIMPLE_SEGMENT|1058,1061|true|false|false|||JVD
Finding|Finding|SIMPLE_SEGMENT|1058,1061|true|false|false|C0425687|Jugular venous engorgement|JVD
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1062,1069|true|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|SIMPLE_SEGMENT|1062,1069|true|false|false|C1314974|Cardiac attachment|CARDIAC
Event|Event|SIMPLE_SEGMENT|1071,1074|false|false|false|||RRR
Event|Event|SIMPLE_SEGMENT|1092,1099|true|false|false|||thrills
Finding|Finding|SIMPLE_SEGMENT|1092,1099|true|false|false|C0232269|Cardiac thrill (finding)|thrills
Event|Event|SIMPLE_SEGMENT|1101,1106|true|false|false|||lifts
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1110,1115|false|false|false|C0024109|Lung|LUNGS
Drug|Organic Chemical|SIMPLE_SEGMENT|1117,1121|false|false|false|C0951233|cetrimonium bromide|CTAB
Event|Event|SIMPLE_SEGMENT|1117,1121|false|false|false|||CTAB
Event|Event|SIMPLE_SEGMENT|1126,1134|true|false|false|||crackles
Finding|Finding|SIMPLE_SEGMENT|1126,1134|true|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Event|Event|SIMPLE_SEGMENT|1136,1143|true|false|false|||wheezes
Finding|Sign or Symptom|SIMPLE_SEGMENT|1136,1143|true|false|false|C0043144|Wheezing|wheezes
Event|Event|SIMPLE_SEGMENT|1147,1154|true|false|false|||rhonchi
Finding|Finding|SIMPLE_SEGMENT|1147,1154|true|false|false|C0035508|Rhonchi|rhonchi
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1158,1165|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1158,1165|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Event|Event|SIMPLE_SEGMENT|1158,1165|false|false|false|||ABDOMEN
Finding|Finding|SIMPLE_SEGMENT|1158,1165|false|false|false|C0941288|Abdomen problem|ABDOMEN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1167,1171|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Event|Event|SIMPLE_SEGMENT|1167,1171|false|false|false|||Soft
Event|Event|SIMPLE_SEGMENT|1173,1177|false|false|false|||NTND
Event|Event|SIMPLE_SEGMENT|1182,1185|true|false|false|||HSM
Finding|Gene or Genome|SIMPLE_SEGMENT|1182,1185|true|false|false|C1537594|LRRC4B gene|HSM
Event|Event|SIMPLE_SEGMENT|1189,1199|true|false|false|||tenderness
Finding|Mental Process|SIMPLE_SEGMENT|1189,1199|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|SIMPLE_SEGMENT|1189,1199|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1203,1214|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1223,1228|true|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|1223,1228|true|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|1223,1228|true|false|false|C0013604|Edema|edema
Drug|Food|SIMPLE_SEGMENT|1229,1235|true|false|false|C5890763||PULSES
Event|Event|SIMPLE_SEGMENT|1229,1235|true|false|false|||PULSES
Finding|Physiologic Function|SIMPLE_SEGMENT|1229,1235|true|false|false|C0391850|Physiologic pulse|PULSES
Procedure|Health Care Activity|SIMPLE_SEGMENT|1229,1235|true|false|false|C0034107|Pulse taking|PULSES
Finding|Functional Concept|SIMPLE_SEGMENT|1264,1269|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Event|Event|SIMPLE_SEGMENT|1284,1288|true|false|false|||take
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|1290,1297|true|false|false|C2346961|Bandage Dosage Form|bandage
Event|Event|SIMPLE_SEGMENT|1290,1297|true|false|false|||bandage
Event|Event|SIMPLE_SEGMENT|1307,1311|true|false|false|||exam
Finding|Functional Concept|SIMPLE_SEGMENT|1307,1311|true|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|1307,1311|true|false|false|C0582103|Medical Examination|exam
Event|Event|SIMPLE_SEGMENT|1333,1340|false|false|false|||dressed
Finding|Body Substance|SIMPLE_SEGMENT|1346,1355|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|1346,1355|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|1346,1355|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|1346,1355|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|SIMPLE_SEGMENT|1356,1360|false|false|false|||EXAM
Finding|Functional Concept|SIMPLE_SEGMENT|1356,1360|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|SIMPLE_SEGMENT|1356,1360|false|false|false|C0582103|Medical Examination|EXAM
Event|Event|SIMPLE_SEGMENT|1376,1382|false|false|false|||VITALS
Event|Event|SIMPLE_SEGMENT|1394,1398|false|false|false|||Temp
Finding|Gene or Genome|SIMPLE_SEGMENT|1394,1398|false|false|false|C1823816|C1orf210 gene|Temp
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1394,1398|false|false|false|C0279848|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Temp
Finding|Individual Behavior|SIMPLE_SEGMENT|1421,1426|false|false|false|C0600261|Telling untruths|Lying
Event|Event|SIMPLE_SEGMENT|1427,1429|false|false|false|||HR
Event|Event|SIMPLE_SEGMENT|1456,1464|false|false|false|||delivery
Finding|Finding|SIMPLE_SEGMENT|1456,1464|false|false|false|C1314680;C1705822;C2053584|Transfer Technique;delivery (history)|delivery
Finding|Functional Concept|SIMPLE_SEGMENT|1456,1464|false|false|false|C1314680;C1705822;C2053584|Transfer Technique;delivery (history)|delivery
Finding|Organism Function|SIMPLE_SEGMENT|1456,1464|false|false|false|C1314680;C1705822;C2053584|Transfer Technique;delivery (history)|delivery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1456,1464|false|false|false|C0011209|Obstetric Delivery|delivery
Event|Event|SIMPLE_SEGMENT|1470,1477|false|false|false|||GENERAL
Finding|Classification|SIMPLE_SEGMENT|1470,1477|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|1470,1477|false|false|false|C3812897|General medical service|GENERAL
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1478,1481|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1478,1481|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1478,1481|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|1478,1481|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1478,1481|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|SIMPLE_SEGMENT|1478,1481|false|false|false|||NAD
Finding|Finding|SIMPLE_SEGMENT|1478,1481|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Event|Event|SIMPLE_SEGMENT|1487,1495|false|false|false|||Pleasant
Finding|Mental Process|SIMPLE_SEGMENT|1487,1495|false|false|false|C2987187|Pleasant|Pleasant
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1504,1509|false|false|false|C1512338|HEENT|HEENT
Event|Event|SIMPLE_SEGMENT|1511,1515|false|false|false|||NCAT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1517,1523|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1517,1523|false|false|false|C0036412|Scleral Diseases|Sclera
Event|Event|SIMPLE_SEGMENT|1517,1523|false|false|false|||Sclera
Procedure|Health Care Activity|SIMPLE_SEGMENT|1517,1523|false|false|false|C2228481|examination of sclera|Sclera
Event|Event|SIMPLE_SEGMENT|1524,1533|false|false|false|||anicteric
Finding|Finding|SIMPLE_SEGMENT|1524,1533|false|false|false|C0205180|Anicteric|anicteric
Event|Event|SIMPLE_SEGMENT|1535,1540|false|false|false|||PERRL
Finding|Finding|SIMPLE_SEGMENT|1535,1540|false|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Event|Event|SIMPLE_SEGMENT|1542,1546|false|false|false|||EOMI
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1548,1559|true|false|false|C0009758;C0229274|Structure of palpebral conjunctiva;conjunctiva|Conjunctiva
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1548,1559|true|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|Conjunctiva
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1548,1559|true|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|Conjunctiva
Event|Event|SIMPLE_SEGMENT|1548,1559|true|false|false|||Conjunctiva
Finding|Body Substance|SIMPLE_SEGMENT|1548,1559|true|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|Conjunctiva
Finding|Intellectual Product|SIMPLE_SEGMENT|1548,1559|true|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|Conjunctiva
Procedure|Health Care Activity|SIMPLE_SEGMENT|1548,1559|true|false|false|C0872390;C2228431|Procedure on conjunctiva;examination of conjunctiva|Conjunctiva
Event|Event|SIMPLE_SEGMENT|1569,1575|true|false|false|||pallor
Finding|Finding|SIMPLE_SEGMENT|1569,1575|true|false|false|C0241137|Pallor of skin|pallor
Event|Event|SIMPLE_SEGMENT|1579,1587|true|false|false|||cyanosis
Finding|Sign or Symptom|SIMPLE_SEGMENT|1579,1587|true|false|false|C0010520|Cyanosis|cyanosis
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|1595,1599|true|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|1595,1599|true|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|1595,1599|true|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|1595,1599|true|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1595,1606|true|false|false|C0026639|Oral mucous membrane structure|oral mucosa
Anatomy|Tissue|SIMPLE_SEGMENT|1600,1606|false|false|false|C0026724|Mucous Membrane|mucosa
Finding|Intellectual Product|SIMPLE_SEGMENT|1600,1606|false|false|false|C1561514||mucosa
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1607,1611|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|SIMPLE_SEGMENT|1607,1611|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|SIMPLE_SEGMENT|1607,1611|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Event|Event|SIMPLE_SEGMENT|1613,1619|true|false|false|||Supple
Finding|Functional Concept|SIMPLE_SEGMENT|1613,1619|true|false|false|C0332254|Supple|Supple
Event|Event|SIMPLE_SEGMENT|1628,1631|true|false|false|||JVD
Finding|Finding|SIMPLE_SEGMENT|1628,1631|true|false|false|C0425687|Jugular venous engorgement|JVD
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1632,1639|true|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|SIMPLE_SEGMENT|1632,1639|true|false|false|C1314974|Cardiac attachment|CARDIAC
Event|Event|SIMPLE_SEGMENT|1641,1644|false|false|false|||RRR
Event|Event|SIMPLE_SEGMENT|1662,1669|true|false|false|||thrills
Finding|Finding|SIMPLE_SEGMENT|1662,1669|true|false|false|C0232269|Cardiac thrill (finding)|thrills
Event|Event|SIMPLE_SEGMENT|1671,1676|true|false|false|||lifts
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1680,1685|false|false|false|C0024109|Lung|LUNGS
Drug|Organic Chemical|SIMPLE_SEGMENT|1687,1691|false|false|false|C0951233|cetrimonium bromide|CTAB
Event|Event|SIMPLE_SEGMENT|1687,1691|false|false|false|||CTAB
Event|Event|SIMPLE_SEGMENT|1696,1704|true|false|false|||crackles
Finding|Finding|SIMPLE_SEGMENT|1696,1704|true|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Event|Event|SIMPLE_SEGMENT|1706,1713|true|false|false|||wheezes
Finding|Sign or Symptom|SIMPLE_SEGMENT|1706,1713|true|false|false|C0043144|Wheezing|wheezes
Event|Event|SIMPLE_SEGMENT|1717,1724|true|false|false|||rhonchi
Finding|Finding|SIMPLE_SEGMENT|1717,1724|true|false|false|C0035508|Rhonchi|rhonchi
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1728,1735|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1728,1735|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Event|Event|SIMPLE_SEGMENT|1728,1735|false|false|false|||ABDOMEN
Finding|Finding|SIMPLE_SEGMENT|1728,1735|false|false|false|C0941288|Abdomen problem|ABDOMEN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1737,1741|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Event|Event|SIMPLE_SEGMENT|1737,1741|false|false|false|||Soft
Event|Event|SIMPLE_SEGMENT|1743,1747|false|false|false|||NTND
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1750,1761|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1770,1775|true|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|1770,1775|true|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|1770,1775|true|false|false|C0013604|Edema|edema
Drug|Food|SIMPLE_SEGMENT|1776,1782|true|false|false|C5890763||PULSES
Event|Event|SIMPLE_SEGMENT|1776,1782|true|false|false|||PULSES
Finding|Physiologic Function|SIMPLE_SEGMENT|1776,1782|true|false|false|C0391850|Physiologic pulse|PULSES
Procedure|Health Care Activity|SIMPLE_SEGMENT|1776,1782|true|false|false|C0034107|Pulse taking|PULSES
Finding|Functional Concept|SIMPLE_SEGMENT|1811,1816|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Event|Event|SIMPLE_SEGMENT|1831,1835|true|false|false|||take
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|1836,1843|true|false|false|C2346961|Bandage Dosage Form|bandage
Event|Event|SIMPLE_SEGMENT|1836,1843|true|false|false|||bandage
Event|Event|SIMPLE_SEGMENT|1853,1857|true|false|false|||exam
Finding|Functional Concept|SIMPLE_SEGMENT|1853,1857|true|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|1853,1857|true|false|false|C0582103|Medical Examination|exam
Event|Event|SIMPLE_SEGMENT|1879,1886|false|false|false|||dressed
Event|Event|SIMPLE_SEGMENT|1902,1906|false|false|false|||exam
Finding|Functional Concept|SIMPLE_SEGMENT|1902,1906|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|1902,1906|false|false|false|C0582103|Medical Examination|exam
Event|Event|SIMPLE_SEGMENT|1927,1934|false|false|false|||picture
Event|Event|SIMPLE_SEGMENT|1938,1941|false|false|false|||OMR
Finding|Gene or Genome|SIMPLE_SEGMENT|1938,1941|false|false|false|C1412647|ATP5F1A gene|OMR
Drug|Food|SIMPLE_SEGMENT|1947,1953|false|false|false|C5890763||pulses
Event|Event|SIMPLE_SEGMENT|1947,1953|false|false|false|||pulses
Finding|Physiologic Function|SIMPLE_SEGMENT|1947,1953|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|SIMPLE_SEGMENT|1947,1953|false|false|false|C0034107|Pulse taking|pulses
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1968,1971|false|false|false|C1332833|Calcifying Fibrous Pseudotumor|CFT
Event|Event|SIMPLE_SEGMENT|1968,1971|false|false|false|||CFT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1968,1971|false|false|false|C0280462;C4552804|Cisplatin/Fluorouracil/Trastuzumab Regimen;Cyclophosphamide/Fluorouracil/Tamoxifen|CFT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1975,1978|false|false|false|C0059387;C0074289|selenocysteine;staphylococcal enterotoxin C|sec
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1975,1978|false|false|false|C0059387;C0074289|selenocysteine;staphylococcal enterotoxin C|sec
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|1975,1978|false|false|false|C0059387;C0074289|selenocysteine;staphylococcal enterotoxin C|sec
Drug|Immunologic Factor|SIMPLE_SEGMENT|1975,1978|false|false|false|C0059387;C0074289|selenocysteine;staphylococcal enterotoxin C|sec
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1982,1988|false|false|false|C0582802|Digit structure|digits
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2015,2021|false|false|false|C0018534|Hallux structure|hallux
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|2022,2027|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|wound
Event|Event|SIMPLE_SEGMENT|2022,2027|false|false|false|||wound
Finding|Body Substance|SIMPLE_SEGMENT|2022,2027|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Functional Concept|SIMPLE_SEGMENT|2022,2027|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Intellectual Product|SIMPLE_SEGMENT|2022,2027|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Event|Event|SIMPLE_SEGMENT|2028,2035|false|false|false|||present
Finding|Finding|SIMPLE_SEGMENT|2028,2035|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|SIMPLE_SEGMENT|2028,2035|false|false|false|C0150312;C0449450|Present;Presentation|present
Event|Event|SIMPLE_SEGMENT|2050,2056|false|false|false|||aspect
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2064,2067|false|false|false|C0040357;C4299090|Lower extremity>Toes;Toes|toe
Event|Event|SIMPLE_SEGMENT|2088,2091|false|false|false|||IPJ
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|2093,2098|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|Wound
Event|Event|SIMPLE_SEGMENT|2093,2098|false|false|false|||Wound
Finding|Body Substance|SIMPLE_SEGMENT|2093,2098|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|Wound
Finding|Functional Concept|SIMPLE_SEGMENT|2093,2098|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|Wound
Finding|Intellectual Product|SIMPLE_SEGMENT|2093,2098|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|Wound
Finding|Pathologic Function|SIMPLE_SEGMENT|2103,2109|false|false|false|C0521172|Eschar|eschar
Event|Event|SIMPLE_SEGMENT|2110,2114|false|false|false|||over
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2126,2130|false|false|false|C2987514|Anatomical base|base
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|2126,2130|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Chemical Viewed Functionally|SIMPLE_SEGMENT|2126,2130|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|2126,2130|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Finding|Gene or Genome|SIMPLE_SEGMENT|2126,2130|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Finding|Idea or Concept|SIMPLE_SEGMENT|2126,2130|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Finding|Functional Concept|SIMPLE_SEGMENT|2146,2160|false|false|false|C0334012|Hyperkeratotic|hyperkeratotic
Anatomy|Body System|SIMPLE_SEGMENT|2161,2165|false|false|false|C1123023;C4520765|Skin;Skin, Human|skin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2161,2165|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2161,2165|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Event|Event|SIMPLE_SEGMENT|2161,2165|false|false|false|||skin
Finding|Body Substance|SIMPLE_SEGMENT|2161,2165|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Finding|Intellectual Product|SIMPLE_SEGMENT|2161,2165|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2182,2190|false|false|false|C0041834|Erythema|erythema
Event|Event|SIMPLE_SEGMENT|2182,2190|false|false|false|||erythema
Event|Event|SIMPLE_SEGMENT|2204,2211|true|false|false|||malodor
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2215,2223|true|false|false|C4489236|Proximal Resection Margin|proximal
Event|Event|SIMPLE_SEGMENT|2224,2233|true|false|false|||streaking
Event|Event|SIMPLE_SEGMENT|2234,2241|true|false|false|||present
Finding|Finding|SIMPLE_SEGMENT|2234,2241|true|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|SIMPLE_SEGMENT|2234,2241|true|false|false|C0150312;C0449450|Present;Presentation|present
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|2252,2257|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|wound
Event|Event|SIMPLE_SEGMENT|2252,2257|false|false|false|||wound
Finding|Body Substance|SIMPLE_SEGMENT|2252,2257|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Functional Concept|SIMPLE_SEGMENT|2252,2257|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Intellectual Product|SIMPLE_SEGMENT|2252,2257|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Event|Event|SIMPLE_SEGMENT|2262,2270|false|false|false|||debrided
Event|Event|SIMPLE_SEGMENT|2279,2285|false|false|false|||eschar
Finding|Pathologic Function|SIMPLE_SEGMENT|2279,2285|false|false|false|C0521172|Eschar|eschar
Anatomy|Body System|SIMPLE_SEGMENT|2319,2323|false|false|false|C1123023;C4520765|Skin;Skin, Human|skin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2319,2323|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2319,2323|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Event|Event|SIMPLE_SEGMENT|2319,2323|false|false|false|||skin
Finding|Body Substance|SIMPLE_SEGMENT|2319,2323|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Finding|Intellectual Product|SIMPLE_SEGMENT|2319,2323|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2331,2335|false|false|false|C2987514|Anatomical base|base
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|2331,2335|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Chemical Viewed Functionally|SIMPLE_SEGMENT|2331,2335|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|2331,2335|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Finding|Gene or Genome|SIMPLE_SEGMENT|2331,2335|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Finding|Idea or Concept|SIMPLE_SEGMENT|2331,2335|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|2343,2348|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|wound
Event|Event|SIMPLE_SEGMENT|2343,2348|false|false|false|||wound
Finding|Body Substance|SIMPLE_SEGMENT|2343,2348|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Functional Concept|SIMPLE_SEGMENT|2343,2348|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Intellectual Product|SIMPLE_SEGMENT|2343,2348|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Drug|Chemical Viewed Functionally|SIMPLE_SEGMENT|2362,2367|true|false|false|C0728863;C2347609|Chemical Probe;Probe brand of methazole herbicide|probe
Drug|Organic Chemical|SIMPLE_SEGMENT|2362,2367|true|false|false|C0728863;C2347609|Chemical Probe;Probe brand of methazole herbicide|probe
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2362,2367|true|false|false|C0728863;C2347609|Chemical Probe;Probe brand of methazole herbicide|probe
Event|Event|SIMPLE_SEGMENT|2362,2367|true|false|false|||probe
Finding|Gene or Genome|SIMPLE_SEGMENT|2362,2367|true|false|false|C1704681|probe gene fragment|probe
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2362,2367|true|false|false|C1442917|DNA probe method|probe
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2368,2372|true|false|false|C4318566|Deep Resection Margin|deep
Event|Event|SIMPLE_SEGMENT|2368,2372|true|false|false|||deep
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2376,2380|true|false|false|C0262950;C1442209|Skeletal bone;XXX bone|bone
Finding|Body Substance|SIMPLE_SEGMENT|2376,2380|true|false|false|C1546560;C1550616|Specimen Type - Bone|bone
Finding|Intellectual Product|SIMPLE_SEGMENT|2376,2380|true|false|false|C1546560;C1550616|Specimen Type - Bone|bone
Finding|Finding|SIMPLE_SEGMENT|2389,2406|false|false|false|C0517630|Purulent drainage|purulent drainage
Event|Event|SIMPLE_SEGMENT|2398,2406|false|false|false|||drainage
Finding|Body Substance|SIMPLE_SEGMENT|2398,2406|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Finding|Sign or Symptom|SIMPLE_SEGMENT|2398,2406|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2398,2406|false|false|false|C0013103|Drainage procedure|drainage
Event|Event|SIMPLE_SEGMENT|2411,2420|false|false|false|||expressed
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|2433,2438|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|Wound
Event|Event|SIMPLE_SEGMENT|2433,2438|false|false|false|||Wound
Finding|Body Substance|SIMPLE_SEGMENT|2433,2438|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|Wound
Finding|Functional Concept|SIMPLE_SEGMENT|2433,2438|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|Wound
Finding|Intellectual Product|SIMPLE_SEGMENT|2433,2438|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|Wound
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2452,2455|false|false|false|C0034155;C1268935|Congenital Thrombotic Thrombocytopenic Purpura;Purpura, Thrombotic Thrombocytopenic|TTP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2452,2455|false|false|false|C1506603;C4723973|ZFP36 protein, human;thiamine triphosphorate|TTP
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2452,2455|false|false|false|C1506603;C4723973|ZFP36 protein, human;thiamine triphosphorate|TTP
Drug|Organic Chemical|SIMPLE_SEGMENT|2452,2455|false|false|false|C1506603;C4723973|ZFP36 protein, human;thiamine triphosphorate|TTP
Drug|Vitamin|SIMPLE_SEGMENT|2452,2455|false|false|false|C1506603;C4723973|ZFP36 protein, human;thiamine triphosphorate|TTP
Event|Event|SIMPLE_SEGMENT|2452,2455|false|false|false|||TTP
Finding|Gene or Genome|SIMPLE_SEGMENT|2452,2455|false|false|false|C1413036;C1421571;C3539814|ADAMTS13 gene;ZFP36 gene;ZFP36 wt Allele|TTP
Event|Event|SIMPLE_SEGMENT|2463,2472|false|false|false|||sensation
Finding|Finding|SIMPLE_SEGMENT|2463,2472|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|2463,2472|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|SIMPLE_SEGMENT|2463,2472|false|false|false|C2229507|sensory exam|sensation
Event|Event|SIMPLE_SEGMENT|2476,2482|false|false|false|||intact
Finding|Finding|SIMPLE_SEGMENT|2476,2482|false|false|false|C1554187|Gender Status - Intact|intact
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2490,2495|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|2490,2495|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2490,2507|false|false|false|C0023216|Lower Extremity|lower extremities
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2496,2507|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2509,2512|false|false|false|C0796068|Oculodigitoesophagoduodenal syndrome|MMT
Drug|Organic Chemical|SIMPLE_SEGMENT|2509,2512|false|false|false|C0046370|2-methylcyclopentadienyl manganese tricarbonyl|MMT
Event|Event|SIMPLE_SEGMENT|2509,2512|false|false|false|||MMT
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2509,2512|false|false|false|C0699782|Manual muscle testing|MMT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2528,2534|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Anatomy|Tissue|SIMPLE_SEGMENT|2528,2534|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Event|Event|SIMPLE_SEGMENT|2535,2541|false|false|false|||groups
Finding|Idea or Concept|SIMPLE_SEGMENT|2535,2541|false|false|false|C0441833;C1552839|Groups;Table Rules - groups|groups
Finding|Intellectual Product|SIMPLE_SEGMENT|2535,2541|false|false|false|C0441833;C1552839|Groups;Table Rules - groups|groups
Event|Event|SIMPLE_SEGMENT|2542,2550|false|false|false|||crossing
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2555,2560|false|false|false|C0003086;C0003087;C4284979|Ankle;Ankle joint structure;Lower extremity>Ankle|ankle
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|2555,2560|false|false|false|C0003086;C0003087;C4284979|Ankle;Ankle joint structure;Lower extremity>Ankle|ankle
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|2574,2585|true|false|false|C0000768|Congenital Abnormality|deformities
Event|Event|SIMPLE_SEGMENT|2574,2585|true|false|false|||deformities
Event|Event|SIMPLE_SEGMENT|2586,2591|true|false|false|||noted
Procedure|Health Care Activity|SIMPLE_SEGMENT|2615,2624|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|SIMPLE_SEGMENT|2625,2629|false|false|false|||LABS
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2625,2629|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2657,2662|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|2657,2662|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|2657,2662|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|2663,2666|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|2673,2676|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2673,2676|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2673,2676|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2682,2685|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2682,2685|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|2682,2685|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2682,2685|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2691,2694|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2691,2694|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|2701,2704|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|2701,2704|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2701,2704|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2701,2704|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2701,2704|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|2708,2711|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2708,2711|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|2708,2711|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|2708,2711|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|2708,2711|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2708,2711|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2718,2722|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2748,2751|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2768,2773|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|2768,2773|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|2768,2773|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|2768,2781|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2768,2781|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2768,2781|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2774,2781|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|2774,2781|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2774,2781|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|2774,2781|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2774,2781|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2774,2781|false|false|false|C0337438|Glucose measurement|Glucose
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2860,2865|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|2860,2865|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|2860,2865|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2892,2897|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|2892,2897|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|2892,2897|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2924,2929|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|2924,2929|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|2924,2929|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2956,2961|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|2956,2961|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|2956,2961|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2962,2967|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|SIMPLE_SEGMENT|2962,2967|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|SIMPLE_SEGMENT|2962,2967|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2962,2967|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Event|Event|SIMPLE_SEGMENT|2965,2967|false|false|false|||MB
Finding|Gene or Genome|SIMPLE_SEGMENT|2965,2969|false|false|false|C1413238;C3273407|CD79A gene;CD79A wt Allele|MB-1
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2996,3001|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|2996,3001|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|2996,3001|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2996,3009|false|false|false|C0853248|Blood albumin|BLOOD Albumin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3002,3009|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3002,3009|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3002,3009|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Event|Event|SIMPLE_SEGMENT|3002,3009|false|false|false|||Albumin
Finding|Gene or Genome|SIMPLE_SEGMENT|3002,3009|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Finding|Physiologic Function|SIMPLE_SEGMENT|3002,3009|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3002,3009|false|false|false|C0201838|Albumin measurement|Albumin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3014,3021|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|3014,3021|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|3014,3021|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3014,3021|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|3014,3021|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|SIMPLE_SEGMENT|3014,3021|false|false|false|||Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|3014,3021|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3014,3021|false|false|false|C0201925|Calcium measurement|Calcium
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3054,3059|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3054,3059|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3054,3059|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3061,3066|false|false|false|C0019018|Glycosylated hemoglobin A|HbA1c
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3061,3066|false|false|false|C0019018|Glycosylated hemoglobin A|HbA1c
Event|Event|SIMPLE_SEGMENT|3061,3066|false|false|false|||HbA1c
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3061,3066|false|false|false|C0202054|Glucohemoglobin measurement|HbA1c
Finding|Gene or Genome|SIMPLE_SEGMENT|3073,3076|false|false|false|C1416571|KCNH1 gene|eAG
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3094,3099|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3094,3099|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3094,3099|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3100,3103|false|false|false|C0006560;C4048285|C-Reactive Protein, human;C-reactive protein|CRP
Drug|Immunologic Factor|SIMPLE_SEGMENT|3100,3103|false|false|false|C0006560;C4048285|C-Reactive Protein, human;C-reactive protein|CRP
Event|Event|SIMPLE_SEGMENT|3100,3103|false|false|false|||CRP
Finding|Gene or Genome|SIMPLE_SEGMENT|3100,3103|false|false|false|C1413716;C1413766;C1826658;C1879974|CRP gene;CRP wt Allele;CSRP1 gene;PPIAP10 gene|CRP
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3122,3127|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3122,3127|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3122,3127|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3128,3131|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Enzyme|SIMPLE_SEGMENT|3128,3131|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Organic Chemical|SIMPLE_SEGMENT|3128,3131|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3128,3131|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Event|Event|SIMPLE_SEGMENT|3128,3131|false|false|false|||ASA
Finding|Gene or Genome|SIMPLE_SEGMENT|3128,3131|false|false|false|C1412553|ARSA gene|ASA
Event|Event|SIMPLE_SEGMENT|3132,3135|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|3132,3135|false|false|false|C5848551|Neg - answer|NEG
Finding|Finding|SIMPLE_SEGMENT|3144,3147|false|false|false|C5848551|Neg - answer|NEG
Event|Event|SIMPLE_SEGMENT|3156,3159|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|3156,3159|false|false|false|C5848551|Neg - answer|NEG
Event|Event|SIMPLE_SEGMENT|3161,3168|false|false|false|||STUDIES
Procedure|Research Activity|SIMPLE_SEGMENT|3161,3168|false|false|false|C0947630|Scientific Study|STUDIES
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3181,3189|false|false|false|C0018787|Heart|Coronary
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3181,3199|false|false|false|C0085532|Coronary angiography|Coronary Angiogram
Event|Event|SIMPLE_SEGMENT|3190,3199|false|false|false|||Angiogram
Finding|Finding|SIMPLE_SEGMENT|3190,3199|false|false|false|C4255126;C5551379|Angiogram (image);Angiogram - result|Angiogram
Finding|Intellectual Product|SIMPLE_SEGMENT|3190,3199|false|false|false|C4255126;C5551379|Angiogram (image);Angiogram - result|Angiogram
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3190,3199|false|false|false|C0002978;C1548816|Angiogram - Consent Type;angiogram|Angiogram
Procedure|Health Care Activity|SIMPLE_SEGMENT|3190,3199|false|false|false|C0002978;C1548816|Angiogram - Consent Type;angiogram|Angiogram
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3200,3208|false|false|false|C0018787|Heart|Coronary
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|3209,3216|false|false|false|C0700276|Anatomical structure|Anatomy
Event|Event|SIMPLE_SEGMENT|3217,3226|false|false|false|||Dominance
Finding|Finding|SIMPLE_SEGMENT|3217,3226|false|false|false|C0870441;C1287621|Dominance;Finding of eye dominance|Dominance
Finding|Idea or Concept|SIMPLE_SEGMENT|3217,3226|false|false|false|C0870441;C1287621|Dominance;Finding of eye dominance|Dominance
Finding|Functional Concept|SIMPLE_SEGMENT|3228,3233|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Finding|Functional Concept|SIMPLE_SEGMENT|3236,3240|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3236,3261|false|false|false|C1261082|Left coronary artery structure|Left Main Coronary Artery
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3246,3254|false|false|false|C0018787|Heart|Coronary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3246,3261|false|false|false|C0205042|Coronary artery|Coronary Artery
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3255,3261|false|false|false|C0003842;C0226004|Arterial system;Arteries|Artery
Anatomy|Body System|SIMPLE_SEGMENT|3255,3261|false|false|false|C0003842;C0226004|Arterial system;Arteries|Artery
Drug|Organic Chemical|SIMPLE_SEGMENT|3266,3270|false|false|false|C2828271|levomefolate calcium|LMCA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3266,3270|false|false|false|C2828271|levomefolate calcium|LMCA
Drug|Vitamin|SIMPLE_SEGMENT|3266,3270|false|false|false|C2828271|levomefolate calcium|LMCA
Event|Event|SIMPLE_SEGMENT|3266,3270|false|false|false|||LMCA
Finding|Functional Concept|SIMPLE_SEGMENT|3277,3281|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3282,3290|false|false|false|C0751437|Adenohypophyseal Diseases|Anterior
Event|Event|SIMPLE_SEGMENT|3291,3301|false|false|false|||Descending
Finding|Functional Concept|SIMPLE_SEGMENT|3291,3301|false|false|false|C1547177|Sequencing - Descending|Descending
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3306,3309|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3306,3309|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|SIMPLE_SEGMENT|3306,3309|false|false|false|||LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|3306,3309|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Finding|Pathologic Function|SIMPLE_SEGMENT|3329,3345|false|false|false|C3272317|Stent restenosis|stent restenosis
Event|Event|SIMPLE_SEGMENT|3335,3345|false|false|false|||restenosis
Finding|Pathologic Function|SIMPLE_SEGMENT|3335,3345|false|false|false|C0333186|Restenosis|restenosis
Finding|Intellectual Product|SIMPLE_SEGMENT|3351,3357|false|false|false|C0030650|Legal patent|patent
Event|Event|SIMPLE_SEGMENT|3358,3362|false|false|false|||LIMA
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3367,3373|false|false|false|C4522154|Distal Resection Margin|distal
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3374,3380|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3374,3380|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Event|Event|SIMPLE_SEGMENT|3463,3471|false|false|false|||occluded
Finding|Finding|SIMPLE_SEGMENT|3463,3471|false|false|false|C0028778;C1947917|Obstruction;Occluded|occluded
Finding|Functional Concept|SIMPLE_SEGMENT|3463,3471|false|false|false|C0028778;C1947917|Obstruction;Occluded|occluded
Event|Event|SIMPLE_SEGMENT|3502,3508|false|false|false|||patent
Finding|Intellectual Product|SIMPLE_SEGMENT|3502,3508|false|false|false|C0030650|Legal patent|patent
Event|Event|SIMPLE_SEGMENT|3510,3513|false|false|false|||SVG
Finding|Functional Concept|SIMPLE_SEGMENT|3524,3529|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3524,3545|false|false|false|C0226042;C1261316|Right coronary artery structure|Right Coronary Artery
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3530,3538|false|false|false|C0018787|Heart|Coronary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3530,3545|false|false|false|C0205042|Coronary artery|Coronary Artery
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3539,3545|false|false|false|C0003842;C0226004|Arterial system;Arteries|Artery
Anatomy|Body System|SIMPLE_SEGMENT|3539,3545|false|false|false|C0003842;C0226004|Arterial system;Arteries|Artery
Event|Event|SIMPLE_SEGMENT|3558,3563|false|false|false|||focal
Event|Event|SIMPLE_SEGMENT|3572,3580|false|false|false|||stenosis
Finding|Pathologic Function|SIMPLE_SEGMENT|3572,3580|false|false|false|C1261287|Stenosis|stenosis
Event|Event|SIMPLE_SEGMENT|3582,3585|false|false|false|||SVG
Event|Event|SIMPLE_SEGMENT|3592,3598|false|false|false|||patent
Finding|Intellectual Product|SIMPLE_SEGMENT|3592,3598|false|false|false|C0030650|Legal patent|patent
Event|Event|SIMPLE_SEGMENT|3600,3604|false|false|false|||LIMA
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3608,3611|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3608,3611|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|3608,3611|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Event|Event|SIMPLE_SEGMENT|3612,3618|false|false|false|||patent
Finding|Intellectual Product|SIMPLE_SEGMENT|3612,3618|false|false|false|C0030650|Legal patent|patent
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3637,3650|true|false|false|C0802632||Complications
Event|Event|SIMPLE_SEGMENT|3637,3650|false|false|false|||Complications
Finding|Functional Concept|SIMPLE_SEGMENT|3637,3650|true|false|false|C0009566;C1171258|Complication;complication aspects|Complications
Finding|Pathologic Function|SIMPLE_SEGMENT|3637,3650|true|false|false|C0009566;C1171258|Complication;complication aspects|Complications
Event|Event|SIMPLE_SEGMENT|3657,3668|true|false|false|||Impressions
Finding|Mental Process|SIMPLE_SEGMENT|3657,3668|true|false|false|C0596764|impression (attitude)|Impressions
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3679,3685|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3679,3685|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3686,3689|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3686,3689|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|3686,3689|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|3686,3689|false|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|3686,3689|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3686,3689|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|3686,3689|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3686,3689|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Finding|Intellectual Product|SIMPLE_SEGMENT|3694,3700|false|false|false|C0030650|Legal patent|Patent
Event|Event|SIMPLE_SEGMENT|3701,3704|false|false|false|||SVG
Event|Event|SIMPLE_SEGMENT|3715,3719|false|false|false|||LIMA
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3723,3726|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3723,3726|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|SIMPLE_SEGMENT|3723,3726|false|false|false|||LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|3723,3726|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Event|Event|SIMPLE_SEGMENT|3728,3743|false|false|false|||Recommendations
Finding|Idea or Concept|SIMPLE_SEGMENT|3728,3743|false|false|false|C0034866|Recommendation|Recommendations
Finding|Functional Concept|SIMPLE_SEGMENT|3747,3754|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|3747,3754|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|3747,3754|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|3747,3754|false|false|false|C0199168|Medical service|Medical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3747,3762|false|false|false|C0418981;C2069680|Medical therapy;disposition medical therapy|Medical therapy
Event|Event|SIMPLE_SEGMENT|3755,3762|false|false|false|||therapy
Finding|Finding|SIMPLE_SEGMENT|3755,3762|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|SIMPLE_SEGMENT|3755,3762|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3755,3762|false|false|false|C0087111|Therapeutic procedure|therapy
Finding|Functional Concept|SIMPLE_SEGMENT|3765,3780|false|false|false|C0205464|pharmacological|Pharmacological
Event|Event|SIMPLE_SEGMENT|3781,3785|false|false|false|||MIBI
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3781,3785|false|false|false|C5557372|Multiplexed Ion Beam Imaging|MIBI
Event|Event|SIMPLE_SEGMENT|3790,3800|false|false|false|||IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|3790,3800|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|3790,3800|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Event|Event|SIMPLE_SEGMENT|3809,3819|false|false|false|||Reversible
Finding|Functional Concept|SIMPLE_SEGMENT|3809,3819|false|false|false|C0205343|Reversible|Reversible
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|3821,3827|false|false|false|C0010454;C1705217|Culture Media;Medium (Substance)|medium
Drug|Substance|SIMPLE_SEGMENT|3821,3827|false|false|false|C0010454;C1705217|Culture Media;Medium (Substance)|medium
Event|Event|SIMPLE_SEGMENT|3821,3827|false|false|false|||medium
Finding|Finding|SIMPLE_SEGMENT|3821,3827|false|false|false|C0009458;C4522282;C4522283|A Medium Amount;A Medium Amount of Time;Communications Media|medium
Finding|Intellectual Product|SIMPLE_SEGMENT|3821,3827|false|false|false|C0009458;C4522282;C4522283|A Medium Amount;A Medium Amount of Time;Communications Media|medium
Finding|Finding|SIMPLE_SEGMENT|3835,3843|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|SIMPLE_SEGMENT|3835,3843|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Event|Event|SIMPLE_SEGMENT|3853,3862|false|false|false|||perfusion
Finding|Functional Concept|SIMPLE_SEGMENT|3853,3862|false|false|false|C4281794;C4723760|Perfusion (biological);Perfusion route|perfusion
Finding|Organism Function|SIMPLE_SEGMENT|3853,3862|false|false|false|C4281794;C4723760|Perfusion (biological);Perfusion route|perfusion
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3853,3862|false|false|false|C0031001;C4721534|Chemotherapeutic Perfusion;Perfusion (procedure)|perfusion
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3863,3869|false|false|false|C1861101|THYROID HORMONE PLASMA MEMBRANE TRANSPORT DEFECT|defect
Event|Event|SIMPLE_SEGMENT|3863,3869|false|false|false|||defect
Finding|Functional Concept|SIMPLE_SEGMENT|3863,3869|false|false|false|C1457869|Defect|defect
Event|Event|SIMPLE_SEGMENT|3871,3880|false|false|false|||involving
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3886,3889|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3886,3889|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|SIMPLE_SEGMENT|3886,3889|false|false|false|||LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|3886,3889|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Event|Event|SIMPLE_SEGMENT|3890,3899|false|false|false|||territory
Finding|Functional Concept|SIMPLE_SEGMENT|3915,3919|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|3915,3938|false|false|false|C0503990|Cavity of left ventricle|left ventricular cavity
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3915,3943|false|false|false|C0455830|Left ventricular cavity size|left ventricular cavity size
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3920,3931|false|false|false|C0018827|Heart Ventricle|ventricular
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|3920,3938|false|false|false|C0507083|Cavity of ventricle|ventricular cavity
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|3932,3938|false|false|false|C0333343|Body cavities|cavity
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|3932,3938|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3932,3938|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|3948,3956|false|false|false|C0039155|Systole|systolic
Event|Event|SIMPLE_SEGMENT|3957,3965|false|false|false|||function
Finding|Finding|SIMPLE_SEGMENT|3957,3965|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|SIMPLE_SEGMENT|3957,3965|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|SIMPLE_SEGMENT|3957,3965|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|SIMPLE_SEGMENT|3957,3965|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Event|Event|SIMPLE_SEGMENT|3973,3981|false|false|false|||Compared
Event|Event|SIMPLE_SEGMENT|3995,4000|false|false|false|||study
Finding|Intellectual Product|SIMPLE_SEGMENT|3995,4000|false|false|false|C1705923|Study Object|study
Procedure|Research Activity|SIMPLE_SEGMENT|3995,4000|false|false|false|C0008972;C0947630;C2603343|Clinical Research;Scientific Study;Study|study
Finding|Functional Concept|SIMPLE_SEGMENT|4013,4022|false|false|false|C4281794;C4723760|Perfusion (biological);Perfusion route|perfusion
Finding|Organism Function|SIMPLE_SEGMENT|4013,4022|false|false|false|C4281794;C4723760|Perfusion (biological);Perfusion route|perfusion
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4013,4022|false|false|false|C0031001;C4721534|Chemotherapeutic Perfusion;Perfusion (procedure)|perfusion
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4023,4029|false|false|false|C1861101|THYROID HORMONE PLASMA MEMBRANE TRANSPORT DEFECT|defect
Event|Event|SIMPLE_SEGMENT|4023,4029|false|false|false|||defect
Finding|Functional Concept|SIMPLE_SEGMENT|4023,4029|false|false|false|C1457869|Defect|defect
Event|Event|SIMPLE_SEGMENT|4034,4037|false|false|false|||new
Finding|Finding|SIMPLE_SEGMENT|4034,4037|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|4034,4037|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Event|Event|SIMPLE_SEGMENT|4044,4048|false|false|false|||ECHO
Procedure|Health Care Activity|SIMPLE_SEGMENT|4044,4048|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4044,4048|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Event|Event|SIMPLE_SEGMENT|4053,4057|false|false|false|||LEFT
Finding|Functional Concept|SIMPLE_SEGMENT|4053,4057|false|false|false|C1552822|Table Cell Horizontal Align - left|LEFT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4053,4064|false|false|false|C0225860|Left atrial structure|LEFT ATRIUM
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4058,4064|false|false|false|C0018792|Heart Atrium|ATRIUM
Finding|Intellectual Product|SIMPLE_SEGMENT|4076,4082|false|false|false|C1705102|Volume (publication)|volume
Event|Event|SIMPLE_SEGMENT|4083,4088|false|false|false|||index
Finding|Idea or Concept|SIMPLE_SEGMENT|4083,4088|false|false|false|C0600653;C0918012;C1552854|Html Link Type - index;Index;Indexes|index
Finding|Intellectual Product|SIMPLE_SEGMENT|4083,4088|false|false|false|C0600653;C0918012;C1552854|Html Link Type - index;Index;Indexes|index
Event|Event|SIMPLE_SEGMENT|4092,4096|false|false|false|||LEFT
Finding|Functional Concept|SIMPLE_SEGMENT|4092,4096|false|false|false|C1552822|Table Cell Horizontal Align - left|LEFT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4092,4106|false|false|false|C0225897;C4266612|Chest>Heart.ventricle.left;Left ventricular structure|LEFT VENTRICLE
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4097,4106|false|false|false|C0007799;C0018827;C2355627|Cerebral Ventricles;Heart Ventricle;Ventricle|VENTRICLE
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4097,4106|false|false|false|C0007799;C0018827;C2355627|Cerebral Ventricles;Heart Ventricle;Ventricle|VENTRICLE
Event|Event|SIMPLE_SEGMENT|4108,4114|false|false|false|||Normal
Event|Event|SIMPLE_SEGMENT|4123,4132|false|false|false|||thickness
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4134,4140|false|false|false|C0333343|Body cavities|cavity
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|4134,4140|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4134,4140|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|4168,4176|false|false|false|C0039155|Systole|systolic
Event|Event|SIMPLE_SEGMENT|4177,4185|false|false|false|||function
Finding|Finding|SIMPLE_SEGMENT|4177,4185|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|SIMPLE_SEGMENT|4177,4185|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|SIMPLE_SEGMENT|4177,4185|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|SIMPLE_SEGMENT|4177,4185|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4195,4199|false|false|false|C0428772|Left ventricular ejection fraction|LVEF
Event|Event|SIMPLE_SEGMENT|4195,4199|false|false|false|||LVEF
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4195,4199|false|false|false|C3837267|LVEF (procedure)|LVEF
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4206,4213|false|false|false|C0554756|Doppler studies|Doppler
Event|Event|SIMPLE_SEGMENT|4215,4225|false|false|false|||parameters
Finding|Finding|SIMPLE_SEGMENT|4215,4225|false|false|false|C0449381|Observation parameter|parameters
Event|Event|SIMPLE_SEGMENT|4235,4245|false|false|false|||consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|4235,4245|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|4235,4250|false|false|false|C0332290|Consistent with|consistent with
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4261,4270|false|false|false|C0012000|Diastole|diastolic
Event|Event|SIMPLE_SEGMENT|4261,4270|false|false|false|||diastolic
Event|Event|SIMPLE_SEGMENT|4272,4280|false|false|false|||function
Finding|Finding|SIMPLE_SEGMENT|4272,4280|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|SIMPLE_SEGMENT|4272,4280|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|SIMPLE_SEGMENT|4272,4280|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|SIMPLE_SEGMENT|4272,4280|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|SIMPLE_SEGMENT|4284,4289|false|false|false|C1552823|Table Cell Horizontal Align - right|RIGHT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4284,4299|false|false|false|C0225883|Right ventricular structure|RIGHT VENTRICLE
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4290,4299|false|false|false|C0007799;C0018827;C2355627|Cerebral Ventricles;Heart Ventricle;Ventricle|VENTRICLE
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4290,4299|false|false|false|C0007799;C0018827;C2355627|Cerebral Ventricles;Heart Ventricle;Ventricle|VENTRICLE
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4311,4318|false|false|false|C0935616|chamber [body part]|chamber
Event|Event|SIMPLE_SEGMENT|4328,4332|false|false|false|||free
Finding|Functional Concept|SIMPLE_SEGMENT|4328,4332|false|false|false|C0332296|Free of (attribute)|free
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4333,4344|false|false|false|C1980023|Wall motion|wall motion
Event|Event|SIMPLE_SEGMENT|4338,4344|false|false|false|||motion
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|4338,4344|false|false|false|C0026597|Motion|motion
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|4364,4370|false|false|false|C0026597|Motion|motion
Event|Event|SIMPLE_SEGMENT|4371,4381|false|false|false|||consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|4371,4381|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|4371,4386|false|false|false|C0332290|Consistent with|consistent with
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4393,4400|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|4393,4400|false|false|false|C1314974|Cardiac attachment|cardiac
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4393,4408|false|false|false|C0018821|Cardiac Surgery procedures|cardiac surgery
Event|Event|SIMPLE_SEGMENT|4401,4408|false|false|false|||surgery
Finding|Finding|SIMPLE_SEGMENT|4401,4408|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|SIMPLE_SEGMENT|4401,4408|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|SIMPLE_SEGMENT|4401,4408|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4401,4408|false|false|false|C0543467|Operative Surgical Procedures|surgery
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4412,4417|false|false|false|C0003483;C4037978|Aorta;Chest+Abdomen>Aorta|AORTA
Procedure|Health Care Activity|SIMPLE_SEGMENT|4412,4417|false|false|false|C0869784|Procedure on aorta|AORTA
Finding|Finding|SIMPLE_SEGMENT|4426,4443|false|false|false|C0579133|Aortic diameter|diameter of aorta
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4438,4443|false|false|false|C0003483;C4037978|Aorta;Chest+Abdomen>Aorta|aorta
Procedure|Health Care Activity|SIMPLE_SEGMENT|4438,4443|false|false|false|C0869784|Procedure on aorta|aorta
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4451,4456|false|false|false|C0030471;C1305231|Nasal sinus;Sinus - general anatomical term|sinus
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|4451,4456|false|false|false|C0016169|pathologic fistula|sinus
Drug|Organic Chemical|SIMPLE_SEGMENT|4451,4456|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4451,4456|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Event|Event|SIMPLE_SEGMENT|4458,4467|false|false|false|||ascending
Finding|Functional Concept|SIMPLE_SEGMENT|4458,4467|false|false|false|C1547175;C1962987|Ascend (action);Sequencing - Ascending|ascending
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4472,4476|false|false|false|C0003741;C0230467;C0741204|ARCH;Arch of foot;Structure of nucleus infundibularis hypothalami|arch
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4472,4476|false|false|false|C0003741;C0230467;C0741204|ARCH;Arch of foot;Structure of nucleus infundibularis hypothalami|arch
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4472,4476|false|false|false|C0003741;C0230467;C0741204|ARCH;Arch of foot;Structure of nucleus infundibularis hypothalami|arch
Finding|Finding|SIMPLE_SEGMENT|4472,4476|false|false|false|C1538146;C4722404|Age-Related Clonal Hematopoiesis;ZBTB8OS gene|arch
Finding|Gene or Genome|SIMPLE_SEGMENT|4472,4476|false|false|false|C1538146;C4722404|Age-Related Clonal Hematopoiesis;ZBTB8OS gene|arch
Event|Event|SIMPLE_SEGMENT|4478,4484|false|false|false|||levels
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4488,4494|false|false|false|C0003483|Aorta|AORTIC
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4488,4500|false|false|false|C0003501;C4533215|Aortic valve structure;Chest>Aortic valve|AORTIC VALVE
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4495,4500|false|false|false|C1186983|Anatomical valve|VALVE
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4509,4515|false|false|false|C0003483|Aorta|aortic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4509,4521|false|false|false|C0003501;C4533215|Aortic valve structure;Chest>Aortic valve|aortic valve
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4516,4521|false|false|false|C1186983|Anatomical valve|valve
Event|Event|SIMPLE_SEGMENT|4522,4530|false|false|false|||leaflets
Event|Event|SIMPLE_SEGMENT|4539,4541|true|false|false|||AS
Event|Event|SIMPLE_SEGMENT|4546,4548|true|false|false|||AR
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4552,4564|false|false|false|C0026264|Mitral Valve|MITRAL VALVE
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4559,4564|false|false|false|C1186983|Anatomical valve|VALVE
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4573,4585|false|false|false|C0026264|Mitral Valve|mitral valve
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4580,4585|false|false|false|C1186983|Anatomical valve|valve
Event|Event|SIMPLE_SEGMENT|4586,4594|false|false|false|||leaflets
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4617,4629|false|false|false|C0026264|Mitral Valve|mitral valve
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4624,4629|false|false|false|C1186983|Anatomical valve|valve
Event|Event|SIMPLE_SEGMENT|4641,4651|false|false|false|||structures
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4666,4671|false|false|false|C1186983|Anatomical valve|VALVE
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4680,4695|false|false|false|C0040960|Tricuspid valve structure|tricuspid valve
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4690,4695|false|false|false|C1186983|Anatomical valve|valve
Event|Event|SIMPLE_SEGMENT|4696,4704|false|false|false|||leaflets
Event|Event|SIMPLE_SEGMENT|4723,4729|false|false|false|||Normal
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|4733,4741|false|false|false|C0039155|Systole|systolic
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4733,4750|false|false|false|C0871470|Systolic Pressure|systolic pressure
Event|Event|SIMPLE_SEGMENT|4742,4750|false|false|false|||pressure
Finding|Finding|SIMPLE_SEGMENT|4742,4750|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|SIMPLE_SEGMENT|4742,4750|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|4742,4750|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|4742,4750|false|false|false|C0033095||pressure
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4754,4768|false|false|false|C0034086|Pulmonary valve structure|PULMONIC VALVE
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4763,4768|false|false|false|C1186983|Anatomical valve|VALVE
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4769,4778|false|false|false|C0024109|Lung|PULMONARY
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4769,4778|false|false|false|C2707265||PULMONARY
Finding|Finding|SIMPLE_SEGMENT|4769,4778|false|false|false|C4522268|Pulmonary (intended site)|PULMONARY
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4769,4785|false|false|false|C0034052|Pulmonary artery structure|PULMONARY ARTERY
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4779,4785|false|false|false|C0003842;C0226004|Arterial system;Arteries|ARTERY
Anatomy|Body System|SIMPLE_SEGMENT|4779,4785|false|false|false|C0003842;C0226004|Arterial system;Arteries|ARTERY
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4787,4801|true|false|false|C0034086|Pulmonary valve structure|Pulmonic valve
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4796,4801|true|false|false|C1186983|Anatomical valve|valve
Event|Event|SIMPLE_SEGMENT|4806,4816|true|false|false|||visualized
Event|Event|SIMPLE_SEGMENT|4822,4824|true|false|false|||PS
Finding|Functional Concept|SIMPLE_SEGMENT|4826,4837|false|false|false|C0205463|Physiological|Physiologic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4844,4855|false|false|false|C0031050|Pericardial sac structure|PERICARDIUM
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4860,4871|true|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4860,4871|true|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4860,4880|true|false|false|C0031039|Pericardial effusion|pericardial effusion
Finding|Body Substance|SIMPLE_SEGMENT|4860,4880|true|false|false|C1253937|Pericardial effusion body substance|pericardial effusion
Event|Event|SIMPLE_SEGMENT|4872,4880|true|false|false|||effusion
Finding|Body Substance|SIMPLE_SEGMENT|4872,4880|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|SIMPLE_SEGMENT|4872,4880|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|4872,4880|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Event|Event|SIMPLE_SEGMENT|4885,4896|false|false|false|||Conclusions
Finding|Idea or Concept|SIMPLE_SEGMENT|4885,4896|false|false|false|C1707478|Conclusion|Conclusions
Finding|Functional Concept|SIMPLE_SEGMENT|4905,4909|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Finding|Finding|SIMPLE_SEGMENT|4905,4923|false|false|false|C2059558||left atrial volume
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4910,4916|false|false|false|C0018792|Heart Atrium|atrial
Finding|Intellectual Product|SIMPLE_SEGMENT|4917,4923|false|false|false|C1705102|Volume (publication)|volume
Event|Event|SIMPLE_SEGMENT|4924,4929|false|false|false|||index
Finding|Idea or Concept|SIMPLE_SEGMENT|4924,4929|false|false|false|C0600653;C0918012;C1552854|Html Link Type - index;Index;Indexes|index
Finding|Intellectual Product|SIMPLE_SEGMENT|4924,4929|false|false|false|C0600653;C0918012;C1552854|Html Link Type - index;Index;Indexes|index
Event|Event|SIMPLE_SEGMENT|4933,4939|false|false|false|||normal
Finding|Functional Concept|SIMPLE_SEGMENT|4948,4952|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4953,4964|false|false|false|C0018827|Heart Ventricle|ventricular
Event|Event|SIMPLE_SEGMENT|4971,4980|false|false|false|||thickness
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4982,4988|false|false|false|C0333343|Body cavities|cavity
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|4982,4988|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4982,4988|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Event|Event|SIMPLE_SEGMENT|5015,5023|false|false|false|||systolic
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|5015,5023|false|false|false|C0039155|Systole|systolic
Event|Event|SIMPLE_SEGMENT|5025,5033|false|false|false|||function
Finding|Finding|SIMPLE_SEGMENT|5025,5033|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|SIMPLE_SEGMENT|5025,5033|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|SIMPLE_SEGMENT|5025,5033|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|SIMPLE_SEGMENT|5025,5033|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5043,5047|false|false|false|C0428772|Left ventricular ejection fraction|LVEF
Event|Event|SIMPLE_SEGMENT|5043,5047|false|false|false|||LVEF
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5043,5047|false|false|false|C3837267|LVEF (procedure)|LVEF
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5057,5064|false|false|false|C0554756|Doppler studies|Doppler
Event|Event|SIMPLE_SEGMENT|5065,5075|false|false|false|||parameters
Finding|Finding|SIMPLE_SEGMENT|5065,5075|false|false|false|C0449381|Observation parameter|parameters
Event|Event|SIMPLE_SEGMENT|5086,5096|false|false|false|||consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|5086,5096|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|5086,5101|false|false|false|C0332290|Consistent with|consistent with
Finding|Functional Concept|SIMPLE_SEGMENT|5109,5113|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5114,5125|false|false|false|C0018827|Heart Ventricle|ventricular
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5126,5135|false|false|false|C0012000|Diastole|diastolic
Event|Event|SIMPLE_SEGMENT|5136,5144|false|false|false|||function
Finding|Finding|SIMPLE_SEGMENT|5136,5144|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|SIMPLE_SEGMENT|5136,5144|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|SIMPLE_SEGMENT|5136,5144|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|SIMPLE_SEGMENT|5136,5144|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|SIMPLE_SEGMENT|5147,5152|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5153,5164|false|false|false|C0018827|Heart Ventricle|ventricular
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5165,5172|false|false|false|C0935616|chamber [body part]|chamber
Event|Event|SIMPLE_SEGMENT|5182,5186|false|false|false|||free
Finding|Functional Concept|SIMPLE_SEGMENT|5182,5186|false|false|false|C0332296|Free of (attribute)|free
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5187,5198|false|false|false|C1980023|Wall motion|wall motion
Event|Event|SIMPLE_SEGMENT|5192,5198|false|false|false|||motion
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|5192,5198|false|false|false|C0026597|Motion|motion
Event|Event|SIMPLE_SEGMENT|5203,5209|false|false|false|||normal
Event|Event|SIMPLE_SEGMENT|5216,5225|false|false|false|||diameters
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5229,5234|false|false|false|C0003483;C4037978|Aorta;Chest+Abdomen>Aorta|aorta
Procedure|Health Care Activity|SIMPLE_SEGMENT|5229,5234|false|false|false|C0869784|Procedure on aorta|aorta
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5242,5247|false|false|false|C0030471;C1305231|Nasal sinus;Sinus - general anatomical term|sinus
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|5242,5247|false|false|false|C0016169|pathologic fistula|sinus
Drug|Organic Chemical|SIMPLE_SEGMENT|5242,5247|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5242,5247|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Event|Event|SIMPLE_SEGMENT|5249,5258|false|false|false|||ascending
Finding|Functional Concept|SIMPLE_SEGMENT|5249,5258|false|false|false|C1547175;C1962987|Ascend (action);Sequencing - Ascending|ascending
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5263,5267|false|false|false|C0003741;C0230467;C0741204|ARCH;Arch of foot;Structure of nucleus infundibularis hypothalami|arch
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5263,5267|false|false|false|C0003741;C0230467;C0741204|ARCH;Arch of foot;Structure of nucleus infundibularis hypothalami|arch
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5263,5267|false|false|false|C0003741;C0230467;C0741204|ARCH;Arch of foot;Structure of nucleus infundibularis hypothalami|arch
Finding|Finding|SIMPLE_SEGMENT|5263,5267|false|false|false|C1538146;C4722404|Age-Related Clonal Hematopoiesis;ZBTB8OS gene|arch
Finding|Gene or Genome|SIMPLE_SEGMENT|5263,5267|false|false|false|C1538146;C4722404|Age-Related Clonal Hematopoiesis;ZBTB8OS gene|arch
Event|Event|SIMPLE_SEGMENT|5268,5274|false|false|false|||levels
Event|Event|SIMPLE_SEGMENT|5280,5286|false|false|false|||normal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5292,5298|false|false|false|C0003483|Aorta|aortic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5292,5304|false|false|false|C0003501;C4533215|Aortic valve structure;Chest>Aortic valve|aortic valve
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5299,5304|false|false|false|C1186983|Anatomical valve|valve
Event|Event|SIMPLE_SEGMENT|5305,5313|false|false|false|||leaflets
Event|Event|SIMPLE_SEGMENT|5339,5345|true|false|false|||normal
Finding|Idea or Concept|SIMPLE_SEGMENT|5351,5355|true|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Finding|Intellectual Product|SIMPLE_SEGMENT|5356,5363|true|false|false|C3273178|Leaflet|leaflet
Event|Event|SIMPLE_SEGMENT|5364,5373|true|false|false|||excursion
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5381,5387|true|false|false|C0003483|Aorta|aortic
Finding|Pathologic Function|SIMPLE_SEGMENT|5381,5396|true|false|false|C0003507|Aortic Valve Stenosis|aortic stenosis
Event|Event|SIMPLE_SEGMENT|5388,5396|true|false|false|||stenosis
Finding|Pathologic Function|SIMPLE_SEGMENT|5388,5396|true|false|false|C1261287|Stenosis|stenosis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5401,5407|true|false|false|C0003483|Aorta|aortic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5401,5421|true|false|false|C0003504|Aortic Valve Insufficiency|aortic regurgitation
Event|Event|SIMPLE_SEGMENT|5408,5421|true|false|false|||regurgitation
Finding|Finding|SIMPLE_SEGMENT|5408,5421|true|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|SIMPLE_SEGMENT|5408,5421|true|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|SIMPLE_SEGMENT|5408,5421|true|false|false|C0460152|Regurgitation - mechanism|regurgitation
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5427,5439|false|false|false|C0026264|Mitral Valve|mitral valve
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5434,5439|false|false|false|C1186983|Anatomical valve|valve
Event|Event|SIMPLE_SEGMENT|5462,5468|false|false|false|||normal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5482,5502|false|false|false|C0026266|Mitral Valve Insufficiency|mitral regurgitation
Event|Event|SIMPLE_SEGMENT|5489,5502|false|false|false|||regurgitation
Finding|Finding|SIMPLE_SEGMENT|5489,5502|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|SIMPLE_SEGMENT|5489,5502|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|SIMPLE_SEGMENT|5489,5502|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5519,5528|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5519,5528|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|5519,5528|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5519,5535|false|false|false|C0034052|Pulmonary artery structure|pulmonary artery
Finding|Finding|SIMPLE_SEGMENT|5519,5553|false|false|false|C0428643|Pulmonary artery systolic pressure|pulmonary artery systolic pressure
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5529,5535|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|SIMPLE_SEGMENT|5529,5535|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|5536,5544|false|false|false|C0039155|Systole|systolic
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5536,5553|false|false|false|C0871470|Systolic Pressure|systolic pressure
Event|Event|SIMPLE_SEGMENT|5545,5553|false|false|false|||pressure
Finding|Finding|SIMPLE_SEGMENT|5545,5553|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|SIMPLE_SEGMENT|5545,5553|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|5545,5553|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|5545,5553|false|false|false|C0033095||pressure
Event|Event|SIMPLE_SEGMENT|5557,5563|false|false|false|||normal
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5578,5589|true|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5578,5589|true|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5578,5598|true|false|false|C0031039|Pericardial effusion|pericardial effusion
Finding|Body Substance|SIMPLE_SEGMENT|5578,5598|true|false|false|C1253937|Pericardial effusion body substance|pericardial effusion
Event|Event|SIMPLE_SEGMENT|5590,5598|true|false|false|||effusion
Finding|Body Substance|SIMPLE_SEGMENT|5590,5598|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|SIMPLE_SEGMENT|5590,5598|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|5590,5598|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Event|Event|SIMPLE_SEGMENT|5603,5613|false|false|false|||IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|5603,5613|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|5603,5613|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|5657,5665|false|false|false|C0039155|Systole|systolic
Event|Event|SIMPLE_SEGMENT|5666,5674|false|false|false|||function
Finding|Finding|SIMPLE_SEGMENT|5666,5674|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|SIMPLE_SEGMENT|5666,5674|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|SIMPLE_SEGMENT|5666,5674|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|SIMPLE_SEGMENT|5666,5674|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Event|Event|SIMPLE_SEGMENT|5703,5708|false|false|false|||study
Finding|Intellectual Product|SIMPLE_SEGMENT|5703,5708|false|false|false|C1705923|Study Object|study
Procedure|Research Activity|SIMPLE_SEGMENT|5703,5708|false|false|false|C0008972;C0947630;C2603343|Clinical Research;Scientific Study;Study|study
Event|Event|SIMPLE_SEGMENT|5717,5725|false|false|false|||reviewed
Finding|Idea or Concept|SIMPLE_SEGMENT|5750,5761|true|false|false|C0750502|Significant|significant
Event|Event|SIMPLE_SEGMENT|5762,5768|true|false|false|||change
Finding|Functional Concept|SIMPLE_SEGMENT|5762,5768|true|false|false|C0392747|Changing|change
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5762,5768|true|false|false|C4319952|Change - procedure|change
Event|Event|SIMPLE_SEGMENT|5769,5774|true|false|false|||noted
Finding|Body Substance|SIMPLE_SEGMENT|5777,5786|true|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|5777,5786|true|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|5777,5786|true|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|5777,5786|true|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|SIMPLE_SEGMENT|5787,5791|false|false|false|||LABS
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5787,5791|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5819,5824|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5819,5824|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5819,5824|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|5825,5828|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|5833,5836|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5833,5836|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5833,5836|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5843,5846|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5843,5846|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|5843,5846|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5843,5846|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5852,5855|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5852,5855|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|5863,5866|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|5863,5866|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5863,5866|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5863,5866|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5863,5866|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|5870,5873|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5870,5873|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|5870,5873|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|5870,5873|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|5870,5873|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5870,5873|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|SIMPLE_SEGMENT|5880,5884|false|false|false|||MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5880,5884|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5910,5913|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5930,5935|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5930,5935|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5930,5935|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|5930,5943|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5930,5943|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5930,5943|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5936,5943|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|5936,5943|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5936,5943|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|5936,5943|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5936,5943|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5936,5943|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5989,5993|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5989,5993|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5989,5993|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6018,6023|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|6018,6023|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|6018,6023|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6024,6027|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6024,6027|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|SIMPLE_SEGMENT|6024,6027|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|SIMPLE_SEGMENT|6024,6027|false|false|false|||ALT
Finding|Gene or Genome|SIMPLE_SEGMENT|6024,6027|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|SIMPLE_SEGMENT|6024,6027|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|SIMPLE_SEGMENT|6024,6027|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6024,6027|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|6031,6034|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6031,6034|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6031,6034|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6031,6034|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|SIMPLE_SEGMENT|6031,6034|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|SIMPLE_SEGMENT|6031,6034|false|false|false|||AST
Finding|Gene or Genome|SIMPLE_SEGMENT|6031,6034|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6038,6045|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|SIMPLE_SEGMENT|6038,6045|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6073,6078|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|6073,6078|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|6073,6078|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6073,6086|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6079,6086|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|6079,6086|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|6079,6086|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6079,6086|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|6079,6086|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|SIMPLE_SEGMENT|6079,6086|false|false|false|||Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|6079,6086|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6079,6086|false|false|false|C0201925|Calcium measurement|Calcium
Finding|Idea or Concept|SIMPLE_SEGMENT|6111,6115|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|SIMPLE_SEGMENT|6111,6115|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Event|Event|SIMPLE_SEGMENT|6116,6119|false|false|false|||old
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6132,6135|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6132,6135|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|6132,6135|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|6132,6135|false|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|6132,6135|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6132,6135|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|6132,6135|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6132,6135|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6140,6143|false|false|false|C0006430|Burning Mouth Syndrome|BMS
Event|Event|SIMPLE_SEGMENT|6140,6143|false|false|false|||BMS
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6144,6152|false|false|false|C4489236|Proximal Resection Margin|proximal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6153,6156|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6153,6156|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|6153,6156|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6162,6165|false|false|false|C4551552|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|DES
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6162,6165|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6162,6165|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Hormone|SIMPLE_SEGMENT|6162,6165|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Organic Chemical|SIMPLE_SEGMENT|6162,6165|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6162,6165|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Event|Event|SIMPLE_SEGMENT|6162,6165|false|false|false|||DES
Finding|Gene or Genome|SIMPLE_SEGMENT|6162,6165|false|false|false|C1413980|DES gene|DES
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6174,6177|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6174,6177|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|SIMPLE_SEGMENT|6174,6177|false|false|false|||LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|6174,6177|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6183,6186|false|false|false|C4551552|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|DES
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6183,6186|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6183,6186|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Hormone|SIMPLE_SEGMENT|6183,6186|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Organic Chemical|SIMPLE_SEGMENT|6183,6186|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6183,6186|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Event|Event|SIMPLE_SEGMENT|6183,6186|false|false|false|||DES
Finding|Gene or Genome|SIMPLE_SEGMENT|6183,6186|false|false|false|C1413980|DES gene|DES
Event|Event|SIMPLE_SEGMENT|6190,6194|false|false|false|||edge
Finding|Conceptual Entity|SIMPLE_SEGMENT|6190,6194|false|false|false|C2697523|Graph Edge|edge
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6206,6209|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6206,6209|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|6206,6209|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6210,6213|false|false|false|C4551552|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|DES
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6210,6213|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6210,6213|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Hormone|SIMPLE_SEGMENT|6210,6213|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Organic Chemical|SIMPLE_SEGMENT|6210,6213|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6210,6213|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Event|Event|SIMPLE_SEGMENT|6210,6213|false|false|false|||DES
Finding|Gene or Genome|SIMPLE_SEGMENT|6210,6213|false|false|false|C1413980|DES gene|DES
Event|Event|SIMPLE_SEGMENT|6218,6226|false|false|false|||stenosis
Finding|Pathologic Function|SIMPLE_SEGMENT|6218,6226|false|false|false|C1261287|Stenosis|stenosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6227,6233|false|false|false|C4522154|Distal Resection Margin|distal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6249,6252|false|false|false|C4551552|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|DES
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6249,6252|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6249,6252|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Hormone|SIMPLE_SEGMENT|6249,6252|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Organic Chemical|SIMPLE_SEGMENT|6249,6252|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6249,6252|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Event|Event|SIMPLE_SEGMENT|6249,6252|false|false|false|||DES
Finding|Gene or Genome|SIMPLE_SEGMENT|6249,6252|false|false|false|C1413980|DES gene|DES
Event|Event|SIMPLE_SEGMENT|6269,6273|false|false|false|||CABG
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6269,6273|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6279,6282|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6279,6282|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|SIMPLE_SEGMENT|6279,6282|false|false|false|||LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|6279,6282|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Finding|Finding|SIMPLE_SEGMENT|6301,6309|false|false|false|C0028778;C1947917|Obstruction;Occluded|occluded
Finding|Functional Concept|SIMPLE_SEGMENT|6301,6309|false|false|false|C0028778;C1947917|Obstruction;Occluded|occluded
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6323,6327|false|false|false|C0011854|Diabetes Mellitus, Insulin-Dependent|IDDM
Event|Event|SIMPLE_SEGMENT|6323,6327|false|false|false|||IDDM
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6329,6332|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|SIMPLE_SEGMENT|6329,6332|false|false|false|||HTN
Event|Event|SIMPLE_SEGMENT|6338,6347|false|false|false|||presented
Finding|Finding|SIMPLE_SEGMENT|6353,6365|false|false|false|C3845714|Several days|several days
Finding|Finding|SIMPLE_SEGMENT|6366,6374|false|false|false|C0741302|atypia morphology|atypical
Finding|Sign or Symptom|SIMPLE_SEGMENT|6366,6385|false|false|false|C0262384|Atypical chest pain|atypical chest pain
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6375,6380|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|6375,6380|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6375,6385|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|6375,6385|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6381,6385|false|true|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|6381,6385|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|6381,6385|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|6381,6385|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|6397,6405|false|false|false|||exertion
Finding|Organism Function|SIMPLE_SEGMENT|6397,6405|false|false|false|C0015264|Exertion|exertion
Finding|Functional Concept|SIMPLE_SEGMENT|6410,6417|false|false|false|C0443144|At rest (qualifier value)|at rest
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6413,6417|false|false|false|C1742913|REST protein, human|rest
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6413,6417|false|false|false|C1742913|REST protein, human|rest
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|6413,6417|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Gene or Genome|SIMPLE_SEGMENT|6413,6417|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Molecular Function|SIMPLE_SEGMENT|6413,6417|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Intellectual Product|SIMPLE_SEGMENT|6424,6428|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Finding|SIMPLE_SEGMENT|6429,6435|false|false|false|C0429103|T wave feature|T wave
Finding|Gene or Genome|SIMPLE_SEGMENT|6431,6435|false|false|false|C1421479|WASF1 gene|wave
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|6431,6435|false|false|false|C0678544||wave
Event|Event|SIMPLE_SEGMENT|6436,6445|false|false|false|||deepening
Event|Event|SIMPLE_SEGMENT|6460,6463|true|false|false|||EKG
Finding|Intellectual Product|SIMPLE_SEGMENT|6460,6463|true|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6460,6463|true|false|false|C1623258|Electrocardiography|EKG
Event|Event|SIMPLE_SEGMENT|6464,6471|true|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|6464,6471|true|false|false|C0392747|Changing|changes
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6475,6483|true|false|false|C0041199|Troponin|troponin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6475,6483|true|false|false|C0041199|Troponin|troponin
Event|Event|SIMPLE_SEGMENT|6475,6483|true|false|false|||troponin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6475,6483|true|false|false|C0523952|Troponin measurement|troponin
Event|Event|SIMPLE_SEGMENT|6494,6503|false|false|false|||presented
Finding|Intellectual Product|SIMPLE_SEGMENT|6509,6513|false|false|false|C1547225|Mild Severity of Illness Code|mild
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6514,6517|false|false|false|C0011880|Diabetic Ketoacidosis|DKA
Event|Event|SIMPLE_SEGMENT|6514,6517|false|false|false|||DKA
Finding|Finding|SIMPLE_SEGMENT|6523,6531|false|false|false|C0241863|Diabetic|diabetic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6523,6536|false|false|false|C0206172|Diabetic Foot|diabetic foot
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6523,6542|false|false|false|C1456868|Diabetic foot ulcer|diabetic foot ulcer
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6532,6536|false|false|false|C0016504;C4299097|Foot;Lower extremity>Foot|foot
Finding|Finding|SIMPLE_SEGMENT|6532,6536|false|false|false|C0555980|Foot problem|foot
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6532,6542|false|false|false|C0085119|Foot Ulcer|foot ulcer
Event|Event|SIMPLE_SEGMENT|6537,6542|false|false|false|||ulcer
Finding|Body Substance|SIMPLE_SEGMENT|6537,6542|false|false|false|C0041582;C1547940;C1550672|Specimen Type - Ulcer;Ulcer|ulcer
Finding|Intellectual Product|SIMPLE_SEGMENT|6537,6542|false|false|false|C0041582;C1547940;C1550672|Specimen Type - Ulcer;Ulcer|ulcer
Finding|Pathologic Function|SIMPLE_SEGMENT|6537,6542|false|false|false|C0041582;C1547940;C1550672|Specimen Type - Ulcer;Ulcer|ulcer
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6554,6560|false|false|false|C1718621|W stress|stress
Drug|Organic Chemical|SIMPLE_SEGMENT|6554,6560|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6554,6560|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Finding|Finding|SIMPLE_SEGMENT|6554,6560|false|false|false|C0038435|Stress|stress
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6554,6565|false|false|false|C0015260;C3494508|Exercise stress test;Stress Test|stress test
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6561,6565|false|false|false|C4318744|Test - temporal region|test
Event|Event|SIMPLE_SEGMENT|6561,6565|false|false|false|||test
Finding|Functional Concept|SIMPLE_SEGMENT|6561,6565|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Finding|Intellectual Product|SIMPLE_SEGMENT|6561,6565|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6561,6565|false|false|false|C0456984|Test Result|test
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6561,6565|false|false|false|C0022885|Laboratory Procedures|test
Event|Event|SIMPLE_SEGMENT|6571,6581|false|false|false|||reversible
Finding|Functional Concept|SIMPLE_SEGMENT|6571,6581|false|false|false|C0205343|Reversible|reversible
Event|Event|SIMPLE_SEGMENT|6583,6591|false|false|false|||ischemia
Finding|Pathologic Function|SIMPLE_SEGMENT|6583,6591|false|false|false|C0022116|Ischemia|ischemia
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6583,6591|false|false|false|C4321499|Ischemia Procedure|ischemia
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6599,6602|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6599,6602|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|6599,6602|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Event|Event|SIMPLE_SEGMENT|6623,6627|false|false|false|||went
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6631,6638|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|6631,6638|false|false|false|C1314974|Cardiac attachment|cardiac
Event|Event|SIMPLE_SEGMENT|6640,6655|false|false|false|||catheterization
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6640,6655|false|false|false|C0007430|Catheterization|catheterization
Event|Event|SIMPLE_SEGMENT|6666,6672|true|false|false|||showed
Finding|Intellectual Product|SIMPLE_SEGMENT|6673,6679|true|false|false|C1547311|Patient Condition Code - Stable|stable
Finding|Classification|SIMPLE_SEGMENT|6673,6687|true|false|false|C0677946;C3538874;C4724041;C5203101;C5203102;C5203130;C5575532|Global Stable Disease in Skin;IMWG Stable Disease;ITMIG MRECIST Stable Disease;RECIL SD;Stable Disease;Stable chronic Graft vs Host Disease;irSD (Immune-Related Response Criteria)|stable disease
Finding|Finding|SIMPLE_SEGMENT|6673,6687|true|false|false|C0677946;C3538874;C4724041;C5203101;C5203102;C5203130;C5575532|Global Stable Disease in Skin;IMWG Stable Disease;ITMIG MRECIST Stable Disease;RECIL SD;Stable Disease;Stable chronic Graft vs Host Disease;irSD (Immune-Related Response Criteria)|stable disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6680,6687|true|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|6680,6687|true|false|false|||disease
Finding|Finding|SIMPLE_SEGMENT|6695,6698|true|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|6695,6698|true|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Functional Concept|SIMPLE_SEGMENT|6700,6711|true|false|false|C0549186|Obstructed|obstructive
Event|Event|SIMPLE_SEGMENT|6712,6719|true|false|false|||lesions
Finding|Finding|SIMPLE_SEGMENT|6712,6719|true|false|false|C0221198|Lesion|lesions
Finding|Intellectual Product|SIMPLE_SEGMENT|6721,6728|false|false|false|C0282416|Overall Publication Type|Overall
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6733,6738|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|6733,6738|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6733,6743|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|6733,6743|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6739,6743|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|6739,6743|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|6739,6743|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|6739,6743|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|6748,6752|false|false|false|||felt
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6774,6789|false|false|false|C2707260||musculoskeletal
Event|Event|SIMPLE_SEGMENT|6774,6789|false|false|false|||musculoskeletal
Finding|Functional Concept|SIMPLE_SEGMENT|6774,6789|false|false|false|C0497254|Musculoskeletal|musculoskeletal
Event|Event|SIMPLE_SEGMENT|6793,6799|false|false|false|||demand
Finding|Idea or Concept|SIMPLE_SEGMENT|6793,6799|false|false|false|C0699784|Economic demand|demand
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6793,6799|false|false|false|C0441516|Demand (clinical)|demand
Finding|Mental Process|SIMPLE_SEGMENT|6807,6814|false|false|false|C0542559|contextual factors|setting
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6818,6821|false|false|false|C0011880|Diabetic Ketoacidosis|DKA
Event|Event|SIMPLE_SEGMENT|6818,6821|false|false|false|||DKA
Finding|Finding|SIMPLE_SEGMENT|6827,6835|false|false|false|C0241863|Diabetic|diabetic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6827,6840|false|false|false|C0206172|Diabetic Foot|diabetic foot
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6827,6846|false|false|false|C1456868|Diabetic foot ulcer|diabetic foot ulcer
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6836,6840|false|false|false|C0016504;C4299097|Foot;Lower extremity>Foot|foot
Finding|Finding|SIMPLE_SEGMENT|6836,6840|false|false|false|C0555980|Foot problem|foot
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6836,6846|false|false|false|C0085119|Foot Ulcer|foot ulcer
Event|Event|SIMPLE_SEGMENT|6841,6846|false|false|false|||ulcer
Finding|Body Substance|SIMPLE_SEGMENT|6841,6846|false|false|false|C0041582;C1547940;C1550672|Specimen Type - Ulcer;Ulcer|ulcer
Finding|Intellectual Product|SIMPLE_SEGMENT|6841,6846|false|false|false|C0041582;C1547940;C1550672|Specimen Type - Ulcer;Ulcer|ulcer
Finding|Pathologic Function|SIMPLE_SEGMENT|6841,6846|false|false|false|C0041582;C1547940;C1550672|Specimen Type - Ulcer;Ulcer|ulcer
Event|Event|SIMPLE_SEGMENT|6856,6866|false|false|false|||discharged
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6870,6873|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Enzyme|SIMPLE_SEGMENT|6870,6873|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Organic Chemical|SIMPLE_SEGMENT|6870,6873|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6870,6873|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Event|Event|SIMPLE_SEGMENT|6870,6873|false|false|false|||ASA
Finding|Gene or Genome|SIMPLE_SEGMENT|6870,6873|false|false|false|C1412553|ARSA gene|ASA
Drug|Organic Chemical|SIMPLE_SEGMENT|6878,6890|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6878,6890|false|false|false|C0286651|atorvastatin|atorvastatin
Event|Event|SIMPLE_SEGMENT|6878,6890|false|false|false|||atorvastatin
Drug|Organic Chemical|SIMPLE_SEGMENT|6896,6906|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6896,6906|false|false|false|C0025859|metoprolol|Metoprolol
Event|Event|SIMPLE_SEGMENT|6910,6915|false|false|false|||100mg
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6926,6929|false|false|false|C0011880|Diabetic Ketoacidosis|DKA
Event|Event|SIMPLE_SEGMENT|6926,6929|false|false|false|||DKA
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6930,6934|false|false|false|C0011854|Diabetes Mellitus, Insulin-Dependent|IDDM
Finding|Body Substance|SIMPLE_SEGMENT|6936,6943|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|6936,6943|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|6936,6943|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|6944,6953|false|false|false|||presented
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|6959,6964|false|false|false|C0003075|Anions|anion
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6959,6968|false|false|false|C0003074|Anion Gap|anion gap
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6959,6968|false|false|false|C1509129|Anion gap result|anion gap
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6959,6968|false|false|false|C0201889;C2189246|Anion gap measurement;blood anion gap (lab test)|anion gap
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6965,6968|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|gap
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6965,6968|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|gap
Event|Event|SIMPLE_SEGMENT|6965,6968|false|false|false|||gap
Finding|Gene or Genome|SIMPLE_SEGMENT|6965,6968|false|false|false|C1419277;C2984552|RASA1 gene;RASA1 wt Allele|gap
Event|Event|SIMPLE_SEGMENT|6969,6978|false|false|false|||metabolic
Finding|Cell Function|SIMPLE_SEGMENT|6969,6978|false|false|false|C0311400;C1524026|Metabolic;Metabolic Process, Cellular|metabolic
Finding|Functional Concept|SIMPLE_SEGMENT|6969,6978|false|false|false|C0311400;C1524026|Metabolic;Metabolic Process, Cellular|metabolic
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6969,6978|false|false|false|C4263342|Multisection metabolic|metabolic
Finding|Pathologic Function|SIMPLE_SEGMENT|6969,6987|false|false|false|C0220981|Metabolic acidosis|metabolic acidosis
Event|Event|SIMPLE_SEGMENT|6979,6987|false|false|false|||acidosis
Finding|Pathologic Function|SIMPLE_SEGMENT|6979,6987|false|false|false|C0001122|Acidosis|acidosis
Event|Event|SIMPLE_SEGMENT|6993,6997|false|false|false|||felt
Finding|Intellectual Product|SIMPLE_SEGMENT|7007,7011|false|false|false|C1547225|Mild Severity of Illness Code|mild
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7012,7015|false|false|false|C0011880|Diabetic Ketoacidosis|DKA
Event|Event|SIMPLE_SEGMENT|7012,7015|false|false|false|||DKA
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7025,7032|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|SIMPLE_SEGMENT|7025,7032|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7025,7032|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|SIMPLE_SEGMENT|7025,7032|false|false|false|||insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|7025,7032|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7025,7032|false|false|false|C0202098|Insulin measurement|insulin
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7033,7036|false|false|false|C1135868|Gestational Trophoblastic Neoplasms|gtt
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7033,7036|false|false|false|C0991568|Drops - Drug Form|gtt
Event|Event|SIMPLE_SEGMENT|7033,7036|false|false|false|||gtt
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7033,7036|false|false|false|C0017741|Glucose tolerance test|gtt
Event|Event|SIMPLE_SEGMENT|7064,7072|false|false|false|||switched
Finding|Functional Concept|SIMPLE_SEGMENT|7076,7088|false|false|false|C1522438|Subcutaneous Route of Administration|subcutaneous
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7089,7096|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|SIMPLE_SEGMENT|7089,7096|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7089,7096|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|SIMPLE_SEGMENT|7089,7096|false|false|false|||insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|7089,7096|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7089,7096|false|false|false|C0202098|Insulin measurement|insulin
Event|Event|SIMPLE_SEGMENT|7102,7105|false|false|false|||A1c
Finding|Classification|SIMPLE_SEGMENT|7102,7105|false|false|false|C4521595|United States Military enlisted E3 (qualifier value)|A1c
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7102,7105|false|false|false|C0474680|Hemoglobin A1c measurement|A1c
Event|Event|SIMPLE_SEGMENT|7106,7114|false|false|false|||returned
Event|Event|SIMPLE_SEGMENT|7137,7144|false|false|false|||highest
Event|Event|SIMPLE_SEGMENT|7157,7165|false|false|false|||recorded
Event|Event|SIMPLE_SEGMENT|7182,7189|false|false|false|||records
Finding|Idea or Concept|SIMPLE_SEGMENT|7182,7189|false|false|false|C0034869;C1548330|Quantity limited request - Records;Records|records
Finding|Intellectual Product|SIMPLE_SEGMENT|7182,7189|false|false|false|C0034869;C1548330|Quantity limited request - Records;Records|records
Drug|Organic Chemical|SIMPLE_SEGMENT|7240,7253|false|false|false|C2974540|canagliflozin|canagliflozin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7240,7253|false|false|false|C2974540|canagliflozin|canagliflozin
Event|Event|SIMPLE_SEGMENT|7240,7253|false|false|false|||canagliflozin
Drug|Organic Chemical|SIMPLE_SEGMENT|7258,7267|false|false|false|C0017642|glipizide|glipizide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7258,7267|false|false|false|C0017642|glipizide|glipizide
Event|Event|SIMPLE_SEGMENT|7258,7267|false|false|false|||glipizide
Finding|Finding|SIMPLE_SEGMENT|7271,7275|false|false|false|C5575035|Well (answer to question)|well
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7282,7289|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|SIMPLE_SEGMENT|7282,7289|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7282,7289|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|SIMPLE_SEGMENT|7282,7289|false|false|false|||insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|7282,7289|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7282,7289|false|false|false|C0202098|Insulin measurement|insulin
Event|Event|SIMPLE_SEGMENT|7300,7309|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|7300,7309|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|SIMPLE_SEGMENT|7324,7332|false|false|false|||reported
Event|Event|SIMPLE_SEGMENT|7346,7355|false|false|false|||adherence
Finding|Functional Concept|SIMPLE_SEGMENT|7346,7355|false|false|false|C1510802|Adherence (attribute)|adherence
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7364,7375|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7364,7375|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|7364,7375|false|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|7364,7375|false|false|false|C4284232|Medications|medications
Finding|Finding|SIMPLE_SEGMENT|7393,7399|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|7393,7399|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|SIMPLE_SEGMENT|7400,7406|false|false|false|||reason
Finding|Idea or Concept|SIMPLE_SEGMENT|7400,7406|false|false|false|C0392360|Indication of (contextual qualifier)|reason
Finding|Idea or Concept|SIMPLE_SEGMENT|7400,7410|false|true|false|C0392360|Indication of (contextual qualifier)|reason for
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7415,7418|false|false|false|C0011880|Diabetic Ketoacidosis|DKA
Event|Event|SIMPLE_SEGMENT|7415,7418|false|false|false|||DKA
Event|Event|SIMPLE_SEGMENT|7475,7478|false|false|false|||met
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7487,7495|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|diabetes
Event|Event|SIMPLE_SEGMENT|7487,7495|false|false|false|||diabetes
Drug|Organic Chemical|SIMPLE_SEGMENT|7510,7523|false|false|false|C2974540|canagliflozin|canagliflozin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7510,7523|false|false|false|C2974540|canagliflozin|canagliflozin
Event|Event|SIMPLE_SEGMENT|7510,7523|false|false|false|||canagliflozin
Event|Event|SIMPLE_SEGMENT|7528,7535|false|false|false|||stopped
Event|Event|SIMPLE_SEGMENT|7540,7549|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|7540,7549|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|7540,7549|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|7540,7549|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|7540,7549|false|false|false|C0030685|Patient Discharge|discharge
Finding|Finding|SIMPLE_SEGMENT|7557,7571|false|false|false|C4699158|Increased risk|increased risk
Event|Event|SIMPLE_SEGMENT|7567,7571|false|false|false|||risk
Finding|Idea or Concept|SIMPLE_SEGMENT|7567,7571|false|false|false|C0035647|Risk|risk
Finding|Idea or Concept|SIMPLE_SEGMENT|7567,7574|false|false|false|C0035647|Risk|risk of
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|7575,7585|false|false|false|C0332840|Amputated structure (morphologic abnormality)|amputation
Event|Event|SIMPLE_SEGMENT|7575,7585|false|false|false|||amputation
Finding|Intellectual Product|SIMPLE_SEGMENT|7575,7585|false|false|false|C1546539|Amputation Specimen Code|amputation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7575,7585|false|false|false|C0002688|Amputation|amputation
Finding|Finding|SIMPLE_SEGMENT|7590,7598|false|false|false|C0241863|Diabetic|Diabetic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7590,7603|false|false|false|C0206172|Diabetic Foot|Diabetic foot
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7590,7609|false|false|false|C1456868|Diabetic foot ulcer|Diabetic foot ulcer
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7599,7603|false|false|false|C0016504;C4299097|Foot;Lower extremity>Foot|foot
Finding|Finding|SIMPLE_SEGMENT|7599,7603|false|false|false|C0555980|Foot problem|foot
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7599,7609|false|false|false|C0085119|Foot Ulcer|foot ulcer
Event|Event|SIMPLE_SEGMENT|7604,7609|false|false|false|||ulcer
Finding|Body Substance|SIMPLE_SEGMENT|7604,7609|false|false|false|C0041582;C1547940;C1550672|Specimen Type - Ulcer;Ulcer|ulcer
Finding|Intellectual Product|SIMPLE_SEGMENT|7604,7609|false|false|false|C0041582;C1547940;C1550672|Specimen Type - Ulcer;Ulcer|ulcer
Finding|Pathologic Function|SIMPLE_SEGMENT|7604,7609|false|false|false|C0041582;C1547940;C1550672|Specimen Type - Ulcer;Ulcer|ulcer
Finding|Finding|SIMPLE_SEGMENT|7611,7618|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Idea or Concept|SIMPLE_SEGMENT|7611,7618|false|false|false|C0150312;C0449450|Present;Presentation|Present
Event|Event|SIMPLE_SEGMENT|7650,7659|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|7650,7659|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|SIMPLE_SEGMENT|7683,7694|false|false|false|||debridement
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7683,7694|false|false|false|C0011079;C3245462|Debridement;Sterile maggot wound debridement|debridement
Event|Event|SIMPLE_SEGMENT|7718,7727|false|false|false|||suggested
Event|Event|SIMPLE_SEGMENT|7728,7736|false|false|false|||presence
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7728,7736|false|false|false|C0392148|Providing presence (regime/therapy)|presence
Finding|Finding|SIMPLE_SEGMENT|7728,7739|false|false|false|C0150312|Present|presence of
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7740,7753|false|false|false|C0029443|Osteomyelitis|osteomyelitis
Event|Event|SIMPLE_SEGMENT|7740,7753|false|false|false|||osteomyelitis
Event|Event|SIMPLE_SEGMENT|7764,7774|false|false|false|||maintained
Event|Event|SIMPLE_SEGMENT|7779,7783|false|false|false|||vanc
Drug|Antibiotic|SIMPLE_SEGMENT|7784,7792|false|false|false|C0055003|cefepime|cefepime
Drug|Organic Chemical|SIMPLE_SEGMENT|7784,7792|false|false|false|C0055003|cefepime|cefepime
Event|Event|SIMPLE_SEGMENT|7784,7792|false|false|false|||cefepime
Drug|Organic Chemical|SIMPLE_SEGMENT|7793,7799|false|false|false|C0699678|Flagyl|flagyl
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7793,7799|false|false|false|C0699678|Flagyl|flagyl
Event|Event|SIMPLE_SEGMENT|7793,7799|false|false|false|||flagyl
Event|Event|SIMPLE_SEGMENT|7818,7826|false|false|false|||switched
Drug|Organic Chemical|SIMPLE_SEGMENT|7830,7835|false|false|false|C0701042|Cipro|cipro
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7830,7835|false|false|false|C0701042|Cipro|cipro
Event|Event|SIMPLE_SEGMENT|7847,7856|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|7847,7856|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|7847,7856|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|7847,7856|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|7847,7856|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|SIMPLE_SEGMENT|7870,7874|false|false|false|||recs
Event|Event|SIMPLE_SEGMENT|7880,7885|false|false|false|||plans
Finding|Finding|SIMPLE_SEGMENT|7890,7895|false|false|false|C0587267;C3810854|Close;Closed|close
Finding|Functional Concept|SIMPLE_SEGMENT|7890,7895|false|false|false|C0587267;C3810854|Close;Closed|close
Event|Event|SIMPLE_SEGMENT|7896,7902|false|false|false|||follow
Finding|Functional Concept|SIMPLE_SEGMENT|7896,7902|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|SIMPLE_SEGMENT|7896,7902|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|SIMPLE_SEGMENT|7896,7905|false|false|false|C0589120|Follow-up status|follow up
Procedure|Health Care Activity|SIMPLE_SEGMENT|7896,7905|false|false|false|C1522577|follow-up|follow up
Event|Event|SIMPLE_SEGMENT|7903,7905|false|false|false|||up
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|7912,7917|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|wound
Event|Event|SIMPLE_SEGMENT|7912,7917|false|false|false|||wound
Finding|Body Substance|SIMPLE_SEGMENT|7912,7917|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Functional Concept|SIMPLE_SEGMENT|7912,7917|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Intellectual Product|SIMPLE_SEGMENT|7912,7917|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Body Substance|SIMPLE_SEGMENT|7912,7922|false|false|false|C0438733|Wound swab (specimen)|wound swab
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7912,7922|false|false|false|C2266642|wound swab (lab test)|wound swab
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7918,7922|false|false|false|C0183753;C1706069|Swab Dosage Form;Swab specimen|swab
Drug|Substance|SIMPLE_SEGMENT|7918,7922|false|false|false|C0183753;C1706069|Swab Dosage Form;Swab specimen|swab
Event|Event|SIMPLE_SEGMENT|7918,7922|false|false|false|||swab
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7918,7922|false|false|false|C0563454|Taking of swab|swab
Finding|Finding|SIMPLE_SEGMENT|7926,7930|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|7926,7930|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|7926,7930|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|SIMPLE_SEGMENT|7934,7943|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|7934,7943|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|7934,7943|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|7934,7943|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|7934,7943|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|SIMPLE_SEGMENT|7948,7961|false|false|false|||polymicrobial
Finding|Body Substance|SIMPLE_SEGMENT|7979,7984|false|false|false|C0441833;C1519504;C1561557;C1705428|Group Object;Group Specimen;Groups;Stage Grouping|Group
Finding|Conceptual Entity|SIMPLE_SEGMENT|7979,7984|false|false|false|C0441833;C1519504;C1561557;C1705428|Group Object;Group Specimen;Groups;Stage Grouping|Group
Finding|Functional Concept|SIMPLE_SEGMENT|7979,7984|false|false|false|C0441833;C1519504;C1561557;C1705428|Group Object;Group Specimen;Groups;Stage Grouping|Group
Finding|Idea or Concept|SIMPLE_SEGMENT|7979,7984|false|false|false|C0441833;C1519504;C1561557;C1705428|Group Object;Group Specimen;Groups;Stage Grouping|Group
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7979,7986|false|false|false|C0348801|Group B streptococcal pneumonia|Group B
Finding|Classification|SIMPLE_SEGMENT|7979,7986|false|false|false|C0441836;C4522078|Group B;Group B rank|Group B
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7987,7992|false|false|false|C0038395|Streptococcal Infections|strep
Event|Event|SIMPLE_SEGMENT|7994,8007|false|false|false|||sensitivities
Finding|Finding|SIMPLE_SEGMENT|7994,8007|false|false|false|C0427965|Antimicrobial susceptibility|sensitivities
Event|Event|SIMPLE_SEGMENT|8008,8015|false|false|false|||pending
Finding|Idea or Concept|SIMPLE_SEGMENT|8008,8015|false|false|false|C1691786;C1704475|Pending - Allergy Clinical Status;Pending - referral status|pending
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8021,8031|false|false|false|C0519030|Pneumonia due to Klebsiella pneumoniae|klebsiella
Event|Event|SIMPLE_SEGMENT|8021,8031|false|false|false|||klebsiella
Anatomy|Cell Component|SIMPLE_SEGMENT|8034,8037|false|false|false|C2244316|proteasome-activating nucleotidase complex|pan
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8034,8037|false|false|false|C0031036|Polyarteritis Nodosa|pan
Finding|Gene or Genome|SIMPLE_SEGMENT|8034,8037|false|false|false|C5401218|ADA2 wt Allele|pan
Event|Event|SIMPLE_SEGMENT|8038,8047|false|false|false|||sensitive
Finding|Functional Concept|SIMPLE_SEGMENT|8038,8047|false|false|false|C0332324|Sensitive|sensitive
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|8053,8056|false|false|false|C0026760|Multiple Epiphyseal Dysplasia|Med
Finding|Gene or Genome|SIMPLE_SEGMENT|8053,8056|false|false|false|C1413596;C1413597;C1419866;C1456376;C1549978;C4321267;C5781216|COL9A2 gene;COL9A3 gene;COMP gene;COMP wt Allele;Master of Education;SCN8A gene;SCN8A wt Allele|Med
Finding|Intellectual Product|SIMPLE_SEGMENT|8053,8056|false|false|false|C1413596;C1413597;C1419866;C1456376;C1549978;C4321267;C5781216|COL9A2 gene;COL9A3 gene;COMP gene;COMP wt Allele;Master of Education;SCN8A gene;SCN8A wt Allele|Med
Event|Event|SIMPLE_SEGMENT|8057,8070|false|false|false|||noncompliance
Event|Event|SIMPLE_SEGMENT|8076,8084|false|false|false|||reported
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8098,8108|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|8098,8108|false|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|8098,8108|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|SIMPLE_SEGMENT|8110,8120|false|false|false|||compliance
Finding|Finding|SIMPLE_SEGMENT|8110,8120|false|false|false|C1321605;C3244300;C4054143|Compliance behavior;Operational Compliance;Pulmonary compliance|compliance
Finding|Idea or Concept|SIMPLE_SEGMENT|8110,8120|false|false|false|C1321605;C3244300;C4054143|Compliance behavior;Operational Compliance;Pulmonary compliance|compliance
Finding|Individual Behavior|SIMPLE_SEGMENT|8110,8120|false|false|false|C1321605;C3244300;C4054143|Compliance behavior;Operational Compliance;Pulmonary compliance|compliance
Drug|Organic Chemical|SIMPLE_SEGMENT|8121,8128|false|false|false|C0163712|Relate - vinyl resin|related
Event|Event|SIMPLE_SEGMENT|8121,8128|false|false|false|||related
Finding|Finding|SIMPLE_SEGMENT|8121,8128|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Finding|Functional Concept|SIMPLE_SEGMENT|8121,8128|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Event|Event|SIMPLE_SEGMENT|8132,8142|false|false|false|||difficulty
Finding|Finding|SIMPLE_SEGMENT|8132,8142|false|false|false|C1299586|Has difficulty doing (qualifier value)|difficulty
Event|Event|SIMPLE_SEGMENT|8143,8154|false|false|false|||remembering
Event|Event|SIMPLE_SEGMENT|8158,8162|false|false|false|||take
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8168,8179|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8168,8179|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|8168,8179|false|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|8168,8179|false|false|false|C4284232|Medications|medications
Finding|Finding|SIMPLE_SEGMENT|8183,8187|false|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|8191,8198|false|false|false|||periods
Finding|Organism Function|SIMPLE_SEGMENT|8191,8198|false|false|false|C0025344|Menstruation|periods
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|8202,8212|false|false|false|C0011570;C0011581;C0344315;C0812393|Cancer patients and suicide and depression;Depressed mood;Depressive disorder;Mental Depression|depression
Event|Event|SIMPLE_SEGMENT|8202,8212|false|false|false|||depression
Finding|Functional Concept|SIMPLE_SEGMENT|8202,8212|false|false|false|C0460137;C1579931|Depression - motion|depression
Finding|Sign or Symptom|SIMPLE_SEGMENT|8202,8212|false|false|false|C0460137;C1579931|Depression - motion|depression
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8217,8223|true|false|false|C1718621|W stress|stress
Drug|Organic Chemical|SIMPLE_SEGMENT|8217,8223|true|false|false|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8217,8223|true|false|false|C0723460|Stress bismuth subsalicylate|stress
Event|Event|SIMPLE_SEGMENT|8217,8223|true|false|false|||stress
Finding|Finding|SIMPLE_SEGMENT|8217,8223|true|false|false|C0038435|Stress|stress
Event|Event|SIMPLE_SEGMENT|8231,8237|true|false|false|||taking
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8242,8252|true|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|8242,8252|true|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|8242,8252|true|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|SIMPLE_SEGMENT|8263,8271|true|false|false|||priority
Finding|Mental Process|SIMPLE_SEGMENT|8263,8271|true|false|false|C0699033|Personal priorities|priority
Event|Event|SIMPLE_SEGMENT|8302,8309|false|false|false|||pillbox
Event|Event|SIMPLE_SEGMENT|8335,8342|false|false|false|||helping
Event|Event|SIMPLE_SEGMENT|8353,8364|false|false|false|||remembering
Event|Event|SIMPLE_SEGMENT|8368,8372|false|false|false|||take
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8377,8388|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8377,8388|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|8377,8388|false|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|8377,8388|false|false|false|C4284232|Medications|medications
Drug|Organic Chemical|SIMPLE_SEGMENT|8400,8410|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8400,8410|false|false|false|C0025859|metoprolol|Metoprolol
Finding|Idea or Concept|SIMPLE_SEGMENT|8414,8419|false|false|false|C1552828|Table Frame - above|above
Event|Event|SIMPLE_SEGMENT|8421,8430|false|false|false|||continued
Drug|Organic Chemical|SIMPLE_SEGMENT|8431,8440|false|false|false|C0076840|torsemide|torsemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8431,8440|false|false|false|C0076840|torsemide|torsemide
Event|Event|SIMPLE_SEGMENT|8464,8473|false|false|false|||euvolemic
Event|Event|SIMPLE_SEGMENT|8485,8494|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|8485,8494|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Drug|Organic Chemical|SIMPLE_SEGMENT|8512,8524|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8512,8524|false|false|false|C0286651|atorvastatin|atorvastatin
Event|Event|SIMPLE_SEGMENT|8512,8524|false|false|false|||atorvastatin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8526,8529|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|SIMPLE_SEGMENT|8526,8529|false|false|false|||HTN
Drug|Organic Chemical|SIMPLE_SEGMENT|8531,8541|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8531,8541|false|false|false|C0025859|metoprolol|Metoprolol
Event|Event|SIMPLE_SEGMENT|8542,8549|false|false|false|||lowered
Drug|Organic Chemical|SIMPLE_SEGMENT|8569,8577|false|false|false|C0126174|losartan|losartan
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8569,8577|false|false|false|C0126174|losartan|losartan
Event|Event|SIMPLE_SEGMENT|8569,8577|false|false|false|||losartan
Event|Event|SIMPLE_SEGMENT|8578,8582|false|false|false|||kept
Drug|Organic Chemical|SIMPLE_SEGMENT|8599,8604|false|false|false|C0590690|Imdur|Imdur
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8599,8604|false|false|false|C0590690|Imdur|Imdur
Event|Event|SIMPLE_SEGMENT|8605,8612|false|false|false|||stopped
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8615,8619|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8615,8619|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|SIMPLE_SEGMENT|8615,8619|false|false|false|||COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|8615,8619|false|false|false|C1412502|ARCN1 gene|COPD
Event|Event|SIMPLE_SEGMENT|8643,8652|false|false|false|||continued
Finding|Idea or Concept|SIMPLE_SEGMENT|8653,8657|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|8653,8657|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|8653,8657|false|false|false|C1553498|home health encounter|home
Event|Event|SIMPLE_SEGMENT|8658,8666|false|false|false|||inhalers
Event|Event|SIMPLE_SEGMENT|8671,8680|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|8671,8680|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|8671,8680|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|8671,8680|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|8671,8680|false|false|false|C0030685|Patient Discharge|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|8684,8692|false|false|false|C0085631;C3887611|Agitation;Restlessness|Restless
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8684,8697|false|false|false|C0035258|Restless Legs Syndrome|Restless legs
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8693,8697|false|false|false|C1140621|Leg|legs
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8693,8697|false|false|false|C5781420||legs
Event|Event|SIMPLE_SEGMENT|8699,8708|false|false|false|||continued
Finding|Idea or Concept|SIMPLE_SEGMENT|8722,8734|false|false|false|C1548597|Marketing basis - Transitional|Transitional
Event|Event|SIMPLE_SEGMENT|8735,8741|false|false|false|||issues
Event|Event|SIMPLE_SEGMENT|8753,8759|false|false|false|||follow
Finding|Finding|SIMPLE_SEGMENT|8767,8775|false|false|false|C0241863|Diabetic|diabetic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8767,8780|false|false|false|C0206172|Diabetic Foot|diabetic foot
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8767,8786|false|false|false|C1456868|Diabetic foot ulcer|diabetic foot ulcer
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8776,8780|false|false|false|C0016504;C4299097|Foot;Lower extremity>Foot|foot
Finding|Finding|SIMPLE_SEGMENT|8776,8780|false|false|false|C0555980|Foot problem|foot
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8776,8786|false|false|false|C0085119|Foot Ulcer|foot ulcer
Event|Event|SIMPLE_SEGMENT|8781,8786|false|false|false|||ulcer
Finding|Body Substance|SIMPLE_SEGMENT|8781,8786|false|false|false|C0041582;C1547940;C1550672|Specimen Type - Ulcer;Ulcer|ulcer
Finding|Intellectual Product|SIMPLE_SEGMENT|8781,8786|false|false|false|C0041582;C1547940;C1550672|Specimen Type - Ulcer;Ulcer|ulcer
Finding|Pathologic Function|SIMPLE_SEGMENT|8781,8786|false|false|false|C0041582;C1547940;C1550672|Specimen Type - Ulcer;Ulcer|ulcer
Event|Event|SIMPLE_SEGMENT|8794,8800|false|false|false|||clinic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8803,8807|false|false|false|C0270724|Infantile Neuroaxonal Dystrophy|Plan
Event|Event|SIMPLE_SEGMENT|8803,8807|false|false|false|||Plan
Finding|Functional Concept|SIMPLE_SEGMENT|8803,8807|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|Plan
Finding|Intellectual Product|SIMPLE_SEGMENT|8803,8807|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|Plan
Finding|Mental Process|SIMPLE_SEGMENT|8803,8807|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|Plan
Finding|Finding|SIMPLE_SEGMENT|8811,8815|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|8811,8815|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|8811,8815|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|SIMPLE_SEGMENT|8819,8828|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|8819,8828|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|8819,8828|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|8819,8828|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|8819,8828|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|SIMPLE_SEGMENT|8836,8840|false|false|false|||take
Event|Event|SIMPLE_SEGMENT|8859,8867|false|false|false|||surgical
Procedure|Health Care Activity|SIMPLE_SEGMENT|8859,8867|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8859,8867|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Event|Event|SIMPLE_SEGMENT|8869,8880|false|false|false|||debridement
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8869,8880|false|false|false|C0011079;C3245462|Debridement;Sterile maggot wound debridement|debridement
Finding|Body Substance|SIMPLE_SEGMENT|8882,8889|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|8882,8889|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|8882,8889|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|8894,8904|false|false|false|||discharged
Drug|Organic Chemical|SIMPLE_SEGMENT|8910,8915|false|false|false|C0701042|Cipro|cipro
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8910,8915|false|false|false|C0701042|Cipro|cipro
Event|Event|SIMPLE_SEGMENT|8910,8915|false|false|false|||cipro
Finding|Functional Concept|SIMPLE_SEGMENT|8939,8945|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|SIMPLE_SEGMENT|8939,8945|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|SIMPLE_SEGMENT|8939,8948|false|false|false|C0589120|Follow-up status|follow up
Procedure|Health Care Activity|SIMPLE_SEGMENT|8939,8948|false|false|false|C1522577|follow-up|follow up
Event|Event|SIMPLE_SEGMENT|8946,8948|false|false|false|||up
Event|Event|SIMPLE_SEGMENT|8959,8965|false|false|false|||review
Finding|Idea or Concept|SIMPLE_SEGMENT|8959,8965|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Finding|Intellectual Product|SIMPLE_SEGMENT|8959,8965|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8970,8975|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|8970,8975|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|8970,8975|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Drug|Organic Chemical|SIMPLE_SEGMENT|8970,8982|false|false|false|C0005802|Blood Glucose|blood sugars
Drug|Organic Chemical|SIMPLE_SEGMENT|8976,8982|false|false|false|C0242209|Sugars|sugars
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8976,8982|false|false|false|C0242209|Sugars|sugars
Event|Event|SIMPLE_SEGMENT|8976,8982|false|false|false|||sugars
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8976,8982|false|false|false|C2239291|sugars (lab test)|sugars
Finding|Finding|SIMPLE_SEGMENT|8983,8990|false|false|false|C4534363|At home|at home
Event|Event|SIMPLE_SEGMENT|8986,8990|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|8986,8990|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|8986,8990|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|8986,8990|false|false|false|C1553498|home health encounter|home
Event|Event|SIMPLE_SEGMENT|8995,9003|false|false|false|||continue
Event|Event|SIMPLE_SEGMENT|9018,9028|false|false|false|||compliance
Finding|Finding|SIMPLE_SEGMENT|9018,9028|false|false|false|C1321605;C3244300;C4054143|Compliance behavior;Operational Compliance;Pulmonary compliance|compliance
Finding|Idea or Concept|SIMPLE_SEGMENT|9018,9028|false|false|false|C1321605;C3244300;C4054143|Compliance behavior;Operational Compliance;Pulmonary compliance|compliance
Finding|Individual Behavior|SIMPLE_SEGMENT|9018,9028|false|false|false|C1321605;C3244300;C4054143|Compliance behavior;Operational Compliance;Pulmonary compliance|compliance
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9034,9042|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|diabetes
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9043,9054|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9043,9054|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|9043,9054|false|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|9043,9054|false|false|false|C4284232|Medications|medications
Drug|Organic Chemical|SIMPLE_SEGMENT|9061,9074|false|false|false|C2974540|canagliflozin|Canagliflozin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9061,9074|false|false|false|C2974540|canagliflozin|Canagliflozin
Event|Event|SIMPLE_SEGMENT|9061,9074|false|false|false|||Canagliflozin
Event|Event|SIMPLE_SEGMENT|9079,9086|false|false|false|||stopped
Finding|Finding|SIMPLE_SEGMENT|9094,9108|false|false|false|C4699158|Increased risk|increased risk
Event|Event|SIMPLE_SEGMENT|9104,9108|false|false|false|||risk
Finding|Idea or Concept|SIMPLE_SEGMENT|9104,9108|false|false|false|C0035647|Risk|risk
Finding|Idea or Concept|SIMPLE_SEGMENT|9104,9111|false|false|false|C0035647|Risk|risk of
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|9112,9122|false|false|false|C0332840|Amputated structure (morphologic abnormality)|amputation
Event|Event|SIMPLE_SEGMENT|9112,9122|false|false|false|||amputation
Finding|Intellectual Product|SIMPLE_SEGMENT|9112,9122|false|false|false|C1546539|Amputation Specimen Code|amputation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9112,9122|false|false|false|C0002688|Amputation|amputation
Event|Event|SIMPLE_SEGMENT|9125,9133|false|false|false|||Consider
Drug|Organic Chemical|SIMPLE_SEGMENT|9148,9157|false|false|false|C0025598|metformin|metformin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9148,9157|false|false|false|C0025598|metformin|metformin
Event|Event|SIMPLE_SEGMENT|9148,9157|false|false|false|||metformin
Event|Event|SIMPLE_SEGMENT|9170,9177|false|false|false|||stopped
Finding|Gene or Genome|SIMPLE_SEGMENT|9188,9191|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Event|Event|SIMPLE_SEGMENT|9197,9205|false|false|false|||diarrhea
Finding|Finding|SIMPLE_SEGMENT|9197,9205|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|SIMPLE_SEGMENT|9197,9205|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Idea or Concept|SIMPLE_SEGMENT|9219,9225|false|true|false|C1550462|Observation Interpretation - better|better
Event|Event|SIMPLE_SEGMENT|9226,9232|false|false|false|||option
Finding|Functional Concept|SIMPLE_SEGMENT|9226,9232|false|true|false|C1518601;C1550456|Options;option - ActMoodPredicate|option
Finding|Idea or Concept|SIMPLE_SEGMENT|9226,9232|false|true|false|C1518601;C1550456|Options;option - ActMoodPredicate|option
Event|Event|SIMPLE_SEGMENT|9245,9251|false|false|false|||Follow
Finding|Functional Concept|SIMPLE_SEGMENT|9245,9251|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|Follow
Finding|Intellectual Product|SIMPLE_SEGMENT|9245,9251|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|Follow
Finding|Finding|SIMPLE_SEGMENT|9245,9254|false|false|false|C0589120|Follow-up status|Follow up
Procedure|Health Care Activity|SIMPLE_SEGMENT|9245,9254|false|false|false|C1522577|follow-up|Follow up
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9255,9260|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|9255,9260|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|9255,9260|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Finding|SIMPLE_SEGMENT|9255,9270|false|false|false|C1272641|Systemic arterial pressure|blood pressures
Event|Event|SIMPLE_SEGMENT|9261,9270|false|false|false|||pressures
Finding|Finding|SIMPLE_SEGMENT|9261,9270|false|false|false|C0460139|Pressure (finding)|pressures
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|9261,9270|false|false|false|C0033095||pressures
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9275,9280|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|9275,9280|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|9275,9280|false|false|false|C0795691|HEART PROBLEM|heart
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9275,9285|false|false|false|C0018810;C0488794|heart rate|heart rate
Finding|Finding|SIMPLE_SEGMENT|9275,9285|false|false|false|C2041121||heart rate
Procedure|Health Care Activity|SIMPLE_SEGMENT|9275,9285|false|false|false|C2197023|examination of heart rate|heart rate
Event|Activity|SIMPLE_SEGMENT|9281,9285|false|false|false|C0871208|Rating (action)|rate
Event|Event|SIMPLE_SEGMENT|9281,9285|false|false|false|||rate
Finding|Idea or Concept|SIMPLE_SEGMENT|9281,9285|false|false|false|C1549480|Amount type - Rate|rate
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|9293,9300|false|false|false|C1705970|Electrical Current|current
Event|Event|SIMPLE_SEGMENT|9302,9309|false|false|false|||regimen
Finding|Intellectual Product|SIMPLE_SEGMENT|9302,9309|false|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9302,9309|false|false|false|C0040808|Treatment Protocols|regimen
Event|Event|SIMPLE_SEGMENT|9331,9344|false|false|false|||noncompliance
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9349,9360|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9349,9360|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|9349,9360|false|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|9349,9360|false|false|false|C4284232|Medications|medications
Event|Event|SIMPLE_SEGMENT|9367,9377|false|false|false|||uptitrated
Event|Event|SIMPLE_SEGMENT|9388,9393|false|false|false|||doses
Event|Event|SIMPLE_SEGMENT|9412,9417|false|false|false|||needs
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9422,9425|false|false|false|C0228549|Cuneate tubercle structure|cut
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|9422,9425|false|false|false|C0000925|Incised wound|cut
Finding|Finding|SIMPLE_SEGMENT|9422,9425|false|false|false|C1413827;C2136694|CUX1 gene;reported cut of tissue (history)|cut
Finding|Gene or Genome|SIMPLE_SEGMENT|9422,9425|false|false|false|C1413827;C2136694|CUX1 gene;reported cut of tissue (history)|cut
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|9422,9430|false|false|false|C0561296|Cut of back|cut back
Drug|Organic Chemical|SIMPLE_SEGMENT|9436,9446|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9436,9446|false|false|false|C0025859|metoprolol|Metoprolol
Event|Event|SIMPLE_SEGMENT|9451,9457|false|false|false|||stoped
Drug|Organic Chemical|SIMPLE_SEGMENT|9462,9467|false|false|false|C0590690|Imdur|imdur
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9462,9467|false|false|false|C0590690|Imdur|imdur
Event|Event|SIMPLE_SEGMENT|9462,9467|false|false|false|||imdur
Event|Event|SIMPLE_SEGMENT|9474,9481|false|false|false|||restart
Drug|Organic Chemical|SIMPLE_SEGMENT|9482,9487|false|false|false|C0590690|Imdur|imdur
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9482,9487|false|false|false|C0590690|Imdur|imdur
Event|Event|SIMPLE_SEGMENT|9482,9487|false|false|false|||imdur
Event|Event|SIMPLE_SEGMENT|9491,9500|false|false|false|||requiring
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9505,9510|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|9505,9510|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9505,9515|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|9505,9515|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9511,9515|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|9511,9515|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|9511,9515|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|9511,9515|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|9519,9529|false|false|false|||outpatient
Finding|Classification|SIMPLE_SEGMENT|9519,9529|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|9519,9529|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9531,9536|false|false|false|C1874451|Basis|basis
Event|Event|SIMPLE_SEGMENT|9531,9536|false|false|false|||basis
Finding|Functional Concept|SIMPLE_SEGMENT|9531,9536|false|false|false|C1527178|Basis - conceptual entity|basis
Event|Event|SIMPLE_SEGMENT|9546,9554|false|false|false|||continue
Event|Event|SIMPLE_SEGMENT|9558,9562|false|false|false|||work
Finding|Body Substance|SIMPLE_SEGMENT|9568,9575|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|9568,9575|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|9568,9575|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|9579,9582|false|false|false|C0026760|Multiple Epiphyseal Dysplasia|med
Event|Event|SIMPLE_SEGMENT|9579,9582|false|false|false|||med
Finding|Gene or Genome|SIMPLE_SEGMENT|9579,9582|false|false|false|C1413596;C1413597;C1419866;C1456376;C1549978;C4321267;C5781216|COL9A2 gene;COL9A3 gene;COMP gene;COMP wt Allele;Master of Education;SCN8A gene;SCN8A wt Allele|med
Finding|Intellectual Product|SIMPLE_SEGMENT|9579,9582|false|false|false|C1413596;C1413597;C1419866;C1456376;C1549978;C4321267;C5781216|COL9A2 gene;COL9A3 gene;COMP gene;COMP wt Allele;Master of Education;SCN8A gene;SCN8A wt Allele|med
Event|Event|SIMPLE_SEGMENT|9583,9593|false|false|false|||compliance
Finding|Finding|SIMPLE_SEGMENT|9583,9593|false|false|false|C1321605;C3244300;C4054143|Compliance behavior;Operational Compliance;Pulmonary compliance|compliance
Finding|Idea or Concept|SIMPLE_SEGMENT|9583,9593|false|false|false|C1321605;C3244300;C4054143|Compliance behavior;Operational Compliance;Pulmonary compliance|compliance
Finding|Individual Behavior|SIMPLE_SEGMENT|9583,9593|false|false|false|C1321605;C3244300;C4054143|Compliance behavior;Operational Compliance;Pulmonary compliance|compliance
Finding|Finding|SIMPLE_SEGMENT|9599,9607|false|false|false|C0332149|Possible|possible
Event|Event|SIMPLE_SEGMENT|9608,9616|false|false|false|||barriers
Event|Event|SIMPLE_SEGMENT|9622,9628|false|false|false|||denied
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|9629,9639|true|false|false|C0011570;C0011581;C0344315;C0812393|Cancer patients and suicide and depression;Depressed mood;Depressive disorder;Mental Depression|depression
Event|Event|SIMPLE_SEGMENT|9629,9639|true|false|false|||depression
Finding|Functional Concept|SIMPLE_SEGMENT|9629,9639|true|false|false|C0460137;C1579931|Depression - motion|depression
Finding|Sign or Symptom|SIMPLE_SEGMENT|9629,9639|true|false|false|C0460137;C1579931|Depression - motion|depression
Finding|Functional Concept|SIMPLE_SEGMENT|9649,9655|true|false|false|C0728831|Social|social
Event|Event|SIMPLE_SEGMENT|9673,9680|false|false|false|||endorse
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9686,9692|false|false|false|C1718621|W stress|stress
Drug|Organic Chemical|SIMPLE_SEGMENT|9686,9692|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9686,9692|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Event|Event|SIMPLE_SEGMENT|9686,9692|false|false|false|||stress
Finding|Finding|SIMPLE_SEGMENT|9686,9692|false|false|false|C0038435|Stress|stress
Event|Event|SIMPLE_SEGMENT|9693,9698|false|false|false|||makes
Event|Event|SIMPLE_SEGMENT|9702,9706|false|false|false|||hard
Event|Event|SIMPLE_SEGMENT|9710,9714|false|false|false|||take
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9720,9731|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9720,9731|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|9720,9731|false|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|9720,9731|false|false|false|C4284232|Medications|medications
Finding|Idea or Concept|SIMPLE_SEGMENT|9740,9745|false|false|false|C1546485|Diagnosis Type - Final|final
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|9746,9751|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|wound
Event|Event|SIMPLE_SEGMENT|9746,9751|false|false|false|||wound
Finding|Body Substance|SIMPLE_SEGMENT|9746,9751|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Functional Concept|SIMPLE_SEGMENT|9746,9751|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Intellectual Product|SIMPLE_SEGMENT|9746,9751|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Body Substance|SIMPLE_SEGMENT|9746,9756|false|false|false|C0438733|Wound swab (specimen)|wound swab
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9746,9756|false|false|false|C2266642|wound swab (lab test)|wound swab
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9752,9756|false|false|false|C0183753;C1706069|Swab Dosage Form;Swab specimen|swab
Drug|Substance|SIMPLE_SEGMENT|9752,9756|false|false|false|C0183753;C1706069|Swab Dosage Form;Swab specimen|swab
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|9752,9756|false|false|false|C0563454|Taking of swab|swab
Event|Event|SIMPLE_SEGMENT|9757,9765|false|false|false|||cultures
Finding|Idea or Concept|SIMPLE_SEGMENT|9757,9765|false|true|false|C0010453|Culture (Anthropological)|cultures
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9770,9781|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9770,9781|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|9770,9781|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|9770,9781|false|false|false|C4284232|Medications|Medications
Finding|Finding|SIMPLE_SEGMENT|9770,9794|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|SIMPLE_SEGMENT|9785,9794|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|9785,9794|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9813,9823|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|9813,9823|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|9813,9828|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|SIMPLE_SEGMENT|9824,9828|false|false|false|||list
Finding|Intellectual Product|SIMPLE_SEGMENT|9824,9828|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|SIMPLE_SEGMENT|9832,9840|false|false|false|||accurate
Drug|Organic Chemical|SIMPLE_SEGMENT|9845,9853|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9845,9853|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|SIMPLE_SEGMENT|9845,9853|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|SIMPLE_SEGMENT|9845,9853|false|false|false|||complete
Finding|Functional Concept|SIMPLE_SEGMENT|9845,9853|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|SIMPLE_SEGMENT|9845,9853|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Organic Chemical|SIMPLE_SEGMENT|9858,9866|false|false|false|C0126174|losartan|Losartan
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9858,9866|false|false|false|C0126174|losartan|Losartan
Event|Event|SIMPLE_SEGMENT|9858,9866|false|false|false|||Losartan
Drug|Organic Chemical|SIMPLE_SEGMENT|9858,9876|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9858,9876|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9867,9876|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|9867,9876|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Food|SIMPLE_SEGMENT|9867,9876|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|9867,9876|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9867,9876|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Event|Event|SIMPLE_SEGMENT|9867,9876|false|false|false|||Potassium
Finding|Physiologic Function|SIMPLE_SEGMENT|9867,9876|false|false|false|C4553027|Potassium metabolic function|Potassium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9867,9876|false|false|false|C0202194|Potassium measurement|Potassium
Drug|Organic Chemical|SIMPLE_SEGMENT|9896,9909|false|false|false|C0025872|metronidazole|MetronidAZOLE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9896,9909|false|false|false|C0025872|metronidazole|MetronidAZOLE
Event|Event|SIMPLE_SEGMENT|9896,9909|false|false|false|||MetronidAZOLE
Drug|Clinical Drug|SIMPLE_SEGMENT|9896,9917|false|false|false|C0360349||MetronidAZOLE Topical
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9910,9917|false|false|false|C1710439|Topical Dosage Form|Topical
Finding|Functional Concept|SIMPLE_SEGMENT|9910,9917|false|false|false|C1522168|Topical Route of Administration|Topical
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9922,9925|false|false|false|C0017243;C0972569;C1382104;C1551386|Electrophoresis Gel;Gel;Gel - ContainerSeparator;Gel physical state|Gel
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|9922,9925|false|false|false|C0017243;C0972569;C1382104;C1551386|Electrophoresis Gel;Gel;Gel - ContainerSeparator;Gel physical state|Gel
Drug|Substance|SIMPLE_SEGMENT|9922,9925|false|false|false|C0017243;C0972569;C1382104;C1551386|Electrophoresis Gel;Gel;Gel - ContainerSeparator;Gel physical state|Gel
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9922,9925|false|false|false|C5977403|Blood group antibody screen.GEL|Gel
Finding|Gene or Genome|SIMPLE_SEGMENT|9928,9932|false|false|false|C1858559|APPL1 gene|Appl
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|9936,9939|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9936,9939|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9936,9939|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|9936,9939|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|9936,9939|false|false|false|C1332410|BID gene|BID
Event|Event|SIMPLE_SEGMENT|9940,9943|false|false|false|||PRN
Finding|Gene or Genome|SIMPLE_SEGMENT|9940,9943|false|false|false|C1422467|CIAO3 gene|PRN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9944,9951|false|false|false|C0035854|Rosacea|Rosacea
Event|Event|SIMPLE_SEGMENT|9944,9951|false|false|false|||Rosacea
Drug|Organic Chemical|SIMPLE_SEGMENT|9956,9966|false|false|false|C0060926|gabapentin|Gabapentin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9956,9966|false|false|false|C0060926|gabapentin|Gabapentin
Finding|Gene or Genome|SIMPLE_SEGMENT|9981,9984|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|SIMPLE_SEGMENT|9985,9993|false|false|false|||Headache
Finding|Sign or Symptom|SIMPLE_SEGMENT|9985,9993|false|false|false|C0018681|Headache|Headache
Drug|Organic Chemical|SIMPLE_SEGMENT|9998,10008|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9998,10008|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Organic Chemical|SIMPLE_SEGMENT|9998,10018|false|false|false|C0724633|metoprolol succinate|Metoprolol Succinate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9998,10018|false|false|false|C0724633|metoprolol succinate|Metoprolol Succinate
Drug|Organic Chemical|SIMPLE_SEGMENT|10009,10018|false|false|false|C0038617;C0220918|Succinates;succinate|Succinate
Event|Event|SIMPLE_SEGMENT|10009,10018|false|false|false|||Succinate
Drug|Organic Chemical|SIMPLE_SEGMENT|10042,10053|false|false|false|C2746078|linagliptin|linaGLIPtin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10042,10053|false|false|false|C2746078|linagliptin|linaGLIPtin
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|10059,10063|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10059,10063|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|10059,10063|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|10059,10063|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Event|Event|SIMPLE_SEGMENT|10064,10069|false|false|false|||DAILY
Drug|Organic Chemical|SIMPLE_SEGMENT|10074,10086|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10074,10086|false|false|false|C0286651|atorvastatin|Atorvastatin
Event|Event|SIMPLE_SEGMENT|10096,10099|false|false|false|||QPM
Drug|Organic Chemical|SIMPLE_SEGMENT|10104,10114|false|false|false|C0016860|furosemide|Furosemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10104,10114|false|false|false|C0016860|furosemide|Furosemide
Drug|Organic Chemical|SIMPLE_SEGMENT|10134,10144|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10134,10144|false|false|false|C0022251|isosorbide|Isosorbide
Event|Event|SIMPLE_SEGMENT|10134,10144|false|false|false|||Isosorbide
Drug|Organic Chemical|SIMPLE_SEGMENT|10134,10156|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10134,10156|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Event|Event|SIMPLE_SEGMENT|10145,10156|false|false|false|||Mononitrate
Drug|Organic Chemical|SIMPLE_SEGMENT|10177,10190|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10177,10190|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Event|Event|SIMPLE_SEGMENT|10177,10190|false|false|false|||Nitroglycerin
Finding|Gene or Genome|SIMPLE_SEGMENT|10210,10213|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10214,10220|false|false|false|C2926611||angina
Event|Event|SIMPLE_SEGMENT|10214,10220|false|false|false|||angina
Finding|Finding|SIMPLE_SEGMENT|10214,10220|false|false|false|C0002962;C2024883|Angina Pectoris|angina
Finding|Sign or Symptom|SIMPLE_SEGMENT|10214,10220|false|false|false|C0002962;C2024883|Angina Pectoris|angina
Drug|Organic Chemical|SIMPLE_SEGMENT|10226,10236|false|false|false|C0244821|ropinirole|rOPINIRole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10226,10236|false|false|false|C0244821|ropinirole|rOPINIRole
Finding|Sign or Symptom|SIMPLE_SEGMENT|10251,10259|false|false|false|C0085631;C3887611|Agitation;Restlessness|restless
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10251,10263|false|false|false|C0035258|Restless Legs Syndrome|restless leg
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10251,10272|false|true|false|C0035258|Restless Legs Syndrome|restless leg syndrome
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10260,10263|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10264,10272|false|false|false|C0039082|Syndrome|syndrome
Event|Event|SIMPLE_SEGMENT|10264,10272|false|false|false|||syndrome
Drug|Organic Chemical|SIMPLE_SEGMENT|10278,10287|false|false|false|C0030049|oxycodone|OxyCODONE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10278,10287|false|false|false|C0030049|oxycodone|OxyCODONE
Event|Event|SIMPLE_SEGMENT|10278,10287|false|false|false|||OxyCODONE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10278,10287|false|false|false|C0524222|Oxycodone measurement|OxyCODONE
Drug|Organic Chemical|SIMPLE_SEGMENT|10289,10302|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10289,10302|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|SIMPLE_SEGMENT|10289,10302|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10289,10302|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10317,10320|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|SIMPLE_SEGMENT|10317,10320|false|false|false|||TAB
Finding|Gene or Genome|SIMPLE_SEGMENT|10328,10331|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10332,10336|false|false|false|C2598155||Pain
Finding|Functional Concept|SIMPLE_SEGMENT|10332,10336|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|10332,10336|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Finding|SIMPLE_SEGMENT|10340,10346|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|Severe
Finding|Intellectual Product|SIMPLE_SEGMENT|10340,10346|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|Severe
Drug|Organic Chemical|SIMPLE_SEGMENT|10352,10363|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10352,10363|false|false|false|C0082607|fluticasone|Fluticasone
Event|Event|SIMPLE_SEGMENT|10352,10363|false|false|false|||Fluticasone
Drug|Organic Chemical|SIMPLE_SEGMENT|10352,10374|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10352,10374|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Organic Chemical|SIMPLE_SEGMENT|10364,10374|false|false|false|C0033474;C0392214|Propionates;propionate|Propionate
Event|Event|SIMPLE_SEGMENT|10384,10388|false|false|false|||PUFF
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|10392,10395|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10392,10395|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|10392,10395|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|10392,10395|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|10392,10395|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|10401,10413|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10401,10413|false|false|false|C0081876|pantoprazole|Pantoprazole
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|10423,10426|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10423,10426|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|10423,10426|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|10423,10426|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|10423,10426|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|10432,10439|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10432,10439|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|SIMPLE_SEGMENT|10461,10470|false|false|false|C0040805|trazodone|TraZODone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10461,10470|false|false|false|C0040805|trazodone|TraZODone
Finding|Gene or Genome|SIMPLE_SEGMENT|10484,10487|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10488,10496|false|false|false|C1950154|Insomnia homeopathic medication|insomnia
Event|Event|SIMPLE_SEGMENT|10488,10496|false|false|false|||insomnia
Finding|Sign or Symptom|SIMPLE_SEGMENT|10488,10496|false|false|false|C0917801|Sleeplessness|insomnia
Drug|Organic Chemical|SIMPLE_SEGMENT|10502,10515|false|false|false|C2974540|canagliflozin|canagliflozin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10502,10515|false|false|false|C2974540|canagliflozin|canagliflozin
Event|Event|SIMPLE_SEGMENT|10502,10515|false|false|false|||canagliflozin
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|10523,10527|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10523,10527|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|10523,10527|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|10523,10527|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Event|Event|SIMPLE_SEGMENT|10528,10533|false|false|false|||DAILY
Drug|Organic Chemical|SIMPLE_SEGMENT|10539,10548|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10539,10548|false|false|false|C0001927|albuterol|albuterol
Event|Event|SIMPLE_SEGMENT|10539,10548|false|false|false|||albuterol
Drug|Organic Chemical|SIMPLE_SEGMENT|10539,10556|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10539,10556|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|10549,10556|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Inorganic Chemical|SIMPLE_SEGMENT|10549,10556|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10549,10556|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Event|Event|SIMPLE_SEGMENT|10549,10556|false|false|false|||sulfate
Finding|Functional Concept|SIMPLE_SEGMENT|10574,10584|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Finding|Organism Function|SIMPLE_SEGMENT|10574,10584|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Event|Event|SIMPLE_SEGMENT|10585,10588|false|false|false|||Q8H
Finding|Gene or Genome|SIMPLE_SEGMENT|10589,10592|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Organic Chemical|SIMPLE_SEGMENT|10598,10607|false|false|false|C0023660|lidocaine|Lidocaine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10598,10607|false|false|false|C0023660|lidocaine|Lidocaine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10598,10607|false|false|false|C0202404|Lidocaine measurement|Lidocaine
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10611,10616|false|false|false|C0445403;C1533128;C1707974|Body tissue patch material;Human patch material;Patch - Extended Release Film|Patch
Event|Event|SIMPLE_SEGMENT|10611,10616|false|false|false|||Patch
Finding|Finding|SIMPLE_SEGMENT|10611,10616|false|false|false|C0332461|Plaque (lesion)|Patch
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10619,10623|false|false|false|C4308013|PTCH1 protein, human|PTCH
Event|Event|SIMPLE_SEGMENT|10619,10623|false|false|false|||PTCH
Finding|Gene or Genome|SIMPLE_SEGMENT|10619,10623|false|false|false|C0694887;C1705339;C1826732;C4308013|PTCH gene;PTCH1 gene;PTCH1 protein, human;PTCH1 wt Allele|PTCH
Finding|Receptor|SIMPLE_SEGMENT|10619,10623|false|false|false|C0694887;C1705339;C1826732;C4308013|PTCH gene;PTCH1 gene;PTCH1 protein, human;PTCH1 wt Allele|PTCH
Event|Event|SIMPLE_SEGMENT|10627,10630|false|false|false|||QPM
Event|Event|SIMPLE_SEGMENT|10635,10644|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|10635,10644|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|10635,10644|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|10635,10644|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|10635,10644|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|10635,10656|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10645,10656|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10645,10656|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|10645,10656|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|10645,10656|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|SIMPLE_SEGMENT|10662,10675|false|false|false|C0008809|ciprofloxacin|Ciprofloxacin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10662,10675|false|false|false|C0008809|ciprofloxacin|Ciprofloxacin
Drug|Antibiotic|SIMPLE_SEGMENT|10662,10679|false|false|false|C0282104|ciprofloxacin hydrochloride|Ciprofloxacin HCl
Drug|Organic Chemical|SIMPLE_SEGMENT|10662,10679|false|false|false|C0282104|ciprofloxacin hydrochloride|Ciprofloxacin HCl
Disorder|Neoplastic Process|SIMPLE_SEGMENT|10676,10679|false|false|false|C0023443|Hairy Cell Leukemia|HCl
Drug|Immunologic Factor|SIMPLE_SEGMENT|10676,10679|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Inorganic Chemical|SIMPLE_SEGMENT|10676,10679|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10676,10679|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Event|Event|SIMPLE_SEGMENT|10676,10679|false|false|false|||HCl
Drug|Organic Chemical|SIMPLE_SEGMENT|10700,10713|false|false|false|C0008809|ciprofloxacin|ciprofloxacin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10700,10713|false|false|false|C0008809|ciprofloxacin|ciprofloxacin
Drug|Antibiotic|SIMPLE_SEGMENT|10700,10717|false|false|false|C0282104|ciprofloxacin hydrochloride|ciprofloxacin HCl
Drug|Organic Chemical|SIMPLE_SEGMENT|10700,10717|false|false|false|C0282104|ciprofloxacin hydrochloride|ciprofloxacin HCl
Disorder|Neoplastic Process|SIMPLE_SEGMENT|10714,10717|false|false|false|C0023443|Hairy Cell Leukemia|HCl
Drug|Immunologic Factor|SIMPLE_SEGMENT|10714,10717|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Inorganic Chemical|SIMPLE_SEGMENT|10714,10717|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10714,10717|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Event|Event|SIMPLE_SEGMENT|10714,10717|false|false|false|||HCl
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10727,10733|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|SIMPLE_SEGMENT|10737,10745|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|10740,10745|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|10740,10745|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Idea or Concept|SIMPLE_SEGMENT|10754,10757|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|10754,10757|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10769,10775|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|10776,10783|false|false|false|||Refills
Finding|Idea or Concept|SIMPLE_SEGMENT|10776,10783|false|false|false|C0807726|refill|Refills
Drug|Antibiotic|SIMPLE_SEGMENT|10792,10803|false|false|false|C0008947|clindamycin|Clindamycin
Drug|Organic Chemical|SIMPLE_SEGMENT|10792,10803|false|false|false|C0008947|clindamycin|Clindamycin
Drug|Antibiotic|SIMPLE_SEGMENT|10823,10834|false|false|false|C0008947|clindamycin|clindamycin
Drug|Organic Chemical|SIMPLE_SEGMENT|10823,10834|false|false|false|C0008947|clindamycin|clindamycin
Drug|Antibiotic|SIMPLE_SEGMENT|10823,10838|false|false|false|C0282105|clindamycin hydrochloride|clindamycin HCl
Drug|Organic Chemical|SIMPLE_SEGMENT|10823,10838|false|false|false|C0282105|clindamycin hydrochloride|clindamycin HCl
Disorder|Neoplastic Process|SIMPLE_SEGMENT|10835,10838|false|false|false|C0023443|Hairy Cell Leukemia|HCl
Drug|Immunologic Factor|SIMPLE_SEGMENT|10835,10838|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Inorganic Chemical|SIMPLE_SEGMENT|10835,10838|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10835,10838|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Event|Event|SIMPLE_SEGMENT|10835,10838|false|false|false|||HCl
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10848,10855|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Anatomy|Cell Component|SIMPLE_SEGMENT|10848,10855|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10848,10855|false|false|false|C0006935|capsule (pharmacologic)|capsule
Finding|Functional Concept|SIMPLE_SEGMENT|10859,10867|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|10862,10867|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|10862,10867|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10873,10878|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|SIMPLE_SEGMENT|10884,10887|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|10884,10887|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10898,10905|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|SIMPLE_SEGMENT|10898,10905|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10898,10905|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Event|Event|SIMPLE_SEGMENT|10906,10913|false|false|false|||Refills
Finding|Idea or Concept|SIMPLE_SEGMENT|10906,10913|false|false|false|C0807726|refill|Refills
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10922,10930|false|false|false|C0907402|insulin glargine|Glargine
Drug|Hormone|SIMPLE_SEGMENT|10922,10930|false|false|false|C0907402|insulin glargine|Glargine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10922,10930|false|false|false|C0907402|insulin glargine|Glargine
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10948,10955|false|false|false|C0528249|Humalog|Humalog
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10948,10955|false|false|false|C0528249|Humalog|Humalog
Event|Event|SIMPLE_SEGMENT|10965,10974|false|false|false|||Breakfast
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|10965,10974|false|false|false|C2698559|Breakfast|Breakfast
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10975,10982|false|false|false|C0528249|Humalog|Humalog
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10975,10982|false|false|false|C0528249|Humalog|Humalog
Event|Event|SIMPLE_SEGMENT|10992,10997|false|false|false|||Lunch
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|10992,10997|false|false|false|C2697949|Lunch|Lunch
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10998,11005|false|false|false|C0528249|Humalog|Humalog
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10998,11005|false|false|false|C0528249|Humalog|Humalog
Event|Event|SIMPLE_SEGMENT|11015,11021|false|false|false|||Dinner
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|11015,11021|false|false|false|C4048877|Dinner|Dinner
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|11022,11029|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Hormone|SIMPLE_SEGMENT|11022,11029|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11022,11029|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Event|Event|SIMPLE_SEGMENT|11022,11029|false|false|false|||Insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|11022,11029|false|false|false|C1337112|INS gene|Insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|11022,11029|false|false|false|C0202098|Insulin measurement|Insulin
Event|Event|SIMPLE_SEGMENT|11033,11040|false|false|false|||Sliding
Finding|Functional Concept|SIMPLE_SEGMENT|11033,11040|false|false|false|C0332246|Sliding|Sliding
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11033,11046|false|false|false|C2937251|sliding scale|Sliding Scale
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11041,11046|false|false|false|C0222045|Integumentary scale|Scale
Event|Activity|SIMPLE_SEGMENT|11041,11046|false|false|false|C1947916|Scaling|Scale
Finding|Conceptual Entity|SIMPLE_SEGMENT|11041,11046|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|Scale
Finding|Intellectual Product|SIMPLE_SEGMENT|11041,11046|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|Scale
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|11057,11064|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Hormone|SIMPLE_SEGMENT|11057,11064|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11057,11064|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Event|Event|SIMPLE_SEGMENT|11057,11064|false|false|false|||Insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|11057,11064|false|false|false|C1337112|INS gene|Insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|11057,11064|false|false|false|C0202098|Insulin measurement|Insulin
Drug|Organic Chemical|SIMPLE_SEGMENT|11070,11080|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11070,11080|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Organic Chemical|SIMPLE_SEGMENT|11070,11090|false|false|false|C0724633|metoprolol succinate|Metoprolol Succinate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11070,11090|false|false|false|C0724633|metoprolol succinate|Metoprolol Succinate
Drug|Organic Chemical|SIMPLE_SEGMENT|11081,11090|false|false|false|C0038617;C0220918|Succinates;succinate|Succinate
Event|Event|SIMPLE_SEGMENT|11081,11090|false|false|false|||Succinate
Drug|Organic Chemical|SIMPLE_SEGMENT|11115,11125|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11115,11125|false|false|false|C0025859|metoprolol|metoprolol
Drug|Organic Chemical|SIMPLE_SEGMENT|11115,11135|false|false|false|C0724633|metoprolol succinate|metoprolol succinate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11115,11135|false|false|false|C0724633|metoprolol succinate|metoprolol succinate
Drug|Organic Chemical|SIMPLE_SEGMENT|11126,11135|false|false|false|C0038617;C0220918|Succinates;succinate|succinate
Event|Event|SIMPLE_SEGMENT|11126,11135|false|false|false|||succinate
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|11145,11151|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|SIMPLE_SEGMENT|11155,11163|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|11158,11163|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|11158,11163|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Event|Activity|SIMPLE_SEGMENT|11170,11174|false|false|false|C1880359|Dispense (activity)|Disp
Finding|Gene or Genome|SIMPLE_SEGMENT|11170,11174|false|false|false|C2828567|PRSS30P gene|Disp
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|11181,11187|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|11188,11195|false|false|false|||Refills
Finding|Idea or Concept|SIMPLE_SEGMENT|11188,11195|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|11204,11213|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11204,11213|false|false|false|C0001927|albuterol|albuterol
Event|Event|SIMPLE_SEGMENT|11204,11213|false|false|false|||albuterol
Drug|Organic Chemical|SIMPLE_SEGMENT|11204,11221|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11204,11221|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|11214,11221|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Inorganic Chemical|SIMPLE_SEGMENT|11214,11221|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11214,11221|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Event|Event|SIMPLE_SEGMENT|11214,11221|false|false|false|||sulfate
Finding|Functional Concept|SIMPLE_SEGMENT|11239,11249|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Finding|Organism Function|SIMPLE_SEGMENT|11239,11249|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Event|Event|SIMPLE_SEGMENT|11250,11253|false|false|false|||Q8H
Finding|Gene or Genome|SIMPLE_SEGMENT|11254,11257|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Organic Chemical|SIMPLE_SEGMENT|11264,11271|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11264,11271|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|SIMPLE_SEGMENT|11294,11306|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11294,11306|false|false|false|C0286651|atorvastatin|Atorvastatin
Event|Event|SIMPLE_SEGMENT|11316,11319|false|false|false|||QPM
Drug|Organic Chemical|SIMPLE_SEGMENT|11326,11337|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11326,11337|false|false|false|C0082607|fluticasone|Fluticasone
Event|Event|SIMPLE_SEGMENT|11326,11337|false|false|false|||Fluticasone
Drug|Organic Chemical|SIMPLE_SEGMENT|11326,11348|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11326,11348|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Organic Chemical|SIMPLE_SEGMENT|11338,11348|false|false|false|C0033474;C0392214|Propionates;propionate|Propionate
Event|Event|SIMPLE_SEGMENT|11358,11362|false|false|false|||PUFF
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|11366,11369|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|11366,11369|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|11366,11369|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|11366,11369|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|11366,11369|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|11376,11386|false|false|false|C0016860|furosemide|Furosemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11376,11386|false|false|false|C0016860|furosemide|Furosemide
Drug|Organic Chemical|SIMPLE_SEGMENT|11409,11419|false|false|false|C0060926|gabapentin|Gabapentin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11409,11419|false|false|false|C0060926|gabapentin|Gabapentin
Finding|Gene or Genome|SIMPLE_SEGMENT|11434,11437|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|SIMPLE_SEGMENT|11438,11446|false|false|false|||Headache
Finding|Sign or Symptom|SIMPLE_SEGMENT|11438,11446|false|false|false|C0018681|Headache|Headache
Drug|Organic Chemical|SIMPLE_SEGMENT|11454,11465|false|false|false|C2746078|linagliptin|linaGLIPtin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11454,11465|false|false|false|C2746078|linagliptin|linaGLIPtin
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|11471,11475|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|11471,11475|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|11471,11475|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|11471,11475|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Event|Event|SIMPLE_SEGMENT|11476,11481|false|false|false|||DAILY
Drug|Organic Chemical|SIMPLE_SEGMENT|11489,11497|false|false|false|C0126174|losartan|Losartan
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11489,11497|false|false|false|C0126174|losartan|Losartan
Event|Event|SIMPLE_SEGMENT|11489,11497|false|false|false|||Losartan
Drug|Organic Chemical|SIMPLE_SEGMENT|11489,11507|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11489,11507|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|11498,11507|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|11498,11507|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Food|SIMPLE_SEGMENT|11498,11507|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|11498,11507|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11498,11507|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Event|Event|SIMPLE_SEGMENT|11498,11507|false|false|false|||Potassium
Finding|Physiologic Function|SIMPLE_SEGMENT|11498,11507|false|false|false|C4553027|Potassium metabolic function|Potassium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|11498,11507|false|false|false|C0202194|Potassium measurement|Potassium
Drug|Organic Chemical|SIMPLE_SEGMENT|11530,11543|false|false|false|C0025872|metronidazole|MetronidAZOLE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11530,11543|false|false|false|C0025872|metronidazole|MetronidAZOLE
Event|Event|SIMPLE_SEGMENT|11530,11543|false|false|false|||MetronidAZOLE
Drug|Clinical Drug|SIMPLE_SEGMENT|11530,11551|false|false|false|C0360349||MetronidAZOLE Topical
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|11544,11551|false|false|false|C1710439|Topical Dosage Form|Topical
Event|Event|SIMPLE_SEGMENT|11544,11551|false|false|false|||Topical
Finding|Functional Concept|SIMPLE_SEGMENT|11544,11551|false|false|false|C1522168|Topical Route of Administration|Topical
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|11556,11559|false|false|false|C0017243;C0972569;C1382104;C1551386|Electrophoresis Gel;Gel;Gel - ContainerSeparator;Gel physical state|Gel
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|11556,11559|false|false|false|C0017243;C0972569;C1382104;C1551386|Electrophoresis Gel;Gel;Gel - ContainerSeparator;Gel physical state|Gel
Drug|Substance|SIMPLE_SEGMENT|11556,11559|false|false|false|C0017243;C0972569;C1382104;C1551386|Electrophoresis Gel;Gel;Gel - ContainerSeparator;Gel physical state|Gel
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|11556,11559|false|false|false|C5977403|Blood group antibody screen.GEL|Gel
Finding|Gene or Genome|SIMPLE_SEGMENT|11562,11566|false|false|false|C1858559|APPL1 gene|Appl
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|11570,11573|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|11570,11573|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|11570,11573|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|11570,11573|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|11570,11573|false|false|false|C1332410|BID gene|BID
Event|Event|SIMPLE_SEGMENT|11574,11577|false|false|false|||PRN
Finding|Gene or Genome|SIMPLE_SEGMENT|11574,11577|false|false|false|C1422467|CIAO3 gene|PRN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11578,11585|false|false|false|C0035854|Rosacea|Rosacea
Event|Event|SIMPLE_SEGMENT|11578,11585|false|false|false|||Rosacea
Drug|Organic Chemical|SIMPLE_SEGMENT|11593,11606|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11593,11606|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Event|Event|SIMPLE_SEGMENT|11593,11606|false|false|false|||Nitroglycerin
Finding|Gene or Genome|SIMPLE_SEGMENT|11626,11629|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11630,11636|false|false|false|C2926611||angina
Event|Event|SIMPLE_SEGMENT|11630,11636|false|false|false|||angina
Finding|Finding|SIMPLE_SEGMENT|11630,11636|false|false|false|C0002962;C2024883|Angina Pectoris|angina
Finding|Sign or Symptom|SIMPLE_SEGMENT|11630,11636|false|false|false|C0002962;C2024883|Angina Pectoris|angina
Drug|Organic Chemical|SIMPLE_SEGMENT|11644,11653|false|false|false|C0030049|oxycodone|OxyCODONE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11644,11653|false|false|false|C0030049|oxycodone|OxyCODONE
Event|Event|SIMPLE_SEGMENT|11644,11653|false|false|false|||OxyCODONE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|11644,11653|false|false|false|C0524222|Oxycodone measurement|OxyCODONE
Drug|Organic Chemical|SIMPLE_SEGMENT|11655,11668|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11655,11668|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|SIMPLE_SEGMENT|11655,11668|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|11655,11668|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|11683,11686|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|SIMPLE_SEGMENT|11683,11686|false|false|false|||TAB
Finding|Gene or Genome|SIMPLE_SEGMENT|11694,11697|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11698,11702|false|false|false|C2598155||Pain
Event|Event|SIMPLE_SEGMENT|11698,11702|false|false|false|||Pain
Finding|Functional Concept|SIMPLE_SEGMENT|11698,11702|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|11698,11702|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Finding|SIMPLE_SEGMENT|11706,11712|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|Severe
Finding|Intellectual Product|SIMPLE_SEGMENT|11706,11712|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|Severe
Drug|Organic Chemical|SIMPLE_SEGMENT|11718,11727|false|false|false|C0030049|oxycodone|oxycodone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11718,11727|false|false|false|C0030049|oxycodone|oxycodone
Event|Event|SIMPLE_SEGMENT|11718,11727|false|false|false|||oxycodone
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|11718,11727|false|false|false|C0524222|Oxycodone measurement|oxycodone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11718,11741|false|false|false|C0717368|acetaminophen / oxycodone|oxycodone-acetaminophen
Drug|Organic Chemical|SIMPLE_SEGMENT|11728,11741|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11728,11741|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Event|Event|SIMPLE_SEGMENT|11728,11741|false|false|false|||acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|11728,11741|false|false|false|C0373527|Acetaminophen measurement|acetaminophen
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|11756,11762|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|SIMPLE_SEGMENT|11766,11774|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|11769,11774|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|11769,11774|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11782,11787|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Event|Event|SIMPLE_SEGMENT|11782,11787|false|false|false|||times
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|11804,11810|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|11811,11818|false|false|false|||Refills
Finding|Idea or Concept|SIMPLE_SEGMENT|11811,11818|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|11828,11840|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11828,11840|false|false|false|C0081876|pantoprazole|Pantoprazole
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|11850,11853|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|11850,11853|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|11850,11853|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|11850,11853|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|11850,11853|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|11861,11871|false|false|false|C0244821|ropinirole|rOPINIRole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11861,11871|false|false|false|C0244821|ropinirole|rOPINIRole
Finding|Sign or Symptom|SIMPLE_SEGMENT|11886,11894|false|false|false|C0085631;C3887611|Agitation;Restlessness|restless
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11886,11898|false|false|false|C0035258|Restless Legs Syndrome|restless leg
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11886,11907|false|true|false|C0035258|Restless Legs Syndrome|restless leg syndrome
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11895,11898|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11899,11907|false|false|false|C0039082|Syndrome|syndrome
Event|Event|SIMPLE_SEGMENT|11899,11907|false|false|false|||syndrome
Drug|Organic Chemical|SIMPLE_SEGMENT|11915,11924|false|false|false|C0040805|trazodone|TraZODone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11915,11924|false|false|false|C0040805|trazodone|TraZODone
Finding|Gene or Genome|SIMPLE_SEGMENT|11938,11941|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11942,11950|false|false|false|C1950154|Insomnia homeopathic medication|insomnia
Event|Event|SIMPLE_SEGMENT|11942,11950|false|false|false|||insomnia
Finding|Sign or Symptom|SIMPLE_SEGMENT|11942,11950|false|false|false|C0917801|Sleeplessness|insomnia
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|11957,11961|false|false|false|C0675390|ARID1A protein, human|HELD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|11957,11961|false|false|false|C0675390|ARID1A protein, human|HELD
Event|Event|SIMPLE_SEGMENT|11957,11961|false|false|false|||HELD
Finding|Gene or Genome|SIMPLE_SEGMENT|11957,11961|false|false|false|C1948036;C2985160|ARID1A wt Allele;Held - activity status|HELD
Finding|Idea or Concept|SIMPLE_SEGMENT|11957,11961|false|false|false|C1948036;C2985160|ARID1A wt Allele;Held - activity status|HELD
Drug|Organic Chemical|SIMPLE_SEGMENT|11963,11976|false|false|false|C2974540|canagliflozin|canagliflozin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11963,11976|false|false|false|C2974540|canagliflozin|canagliflozin
Event|Event|SIMPLE_SEGMENT|11963,11976|false|false|false|||canagliflozin
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|11984,11988|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|11984,11988|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|11984,11988|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|11984,11988|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12001,12011|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|12001,12011|false|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|12001,12011|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|SIMPLE_SEGMENT|12017,12021|false|false|false|||held
Event|Event|SIMPLE_SEGMENT|12030,12037|true|false|false|||restart
Drug|Organic Chemical|SIMPLE_SEGMENT|12038,12051|true|false|false|C2974540|canagliflozin|canagliflozin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12038,12051|true|false|false|C2974540|canagliflozin|canagliflozin
Event|Event|SIMPLE_SEGMENT|12038,12051|true|false|false|||canagliflozin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|12099,12103|false|false|false|C0675390|ARID1A protein, human|HELD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|12099,12103|false|false|false|C0675390|ARID1A protein, human|HELD
Event|Event|SIMPLE_SEGMENT|12099,12103|false|false|false|||HELD
Finding|Gene or Genome|SIMPLE_SEGMENT|12099,12103|false|false|false|C1948036;C2985160|ARID1A wt Allele;Held - activity status|HELD
Finding|Idea or Concept|SIMPLE_SEGMENT|12099,12103|false|false|false|C1948036;C2985160|ARID1A wt Allele;Held - activity status|HELD
Drug|Organic Chemical|SIMPLE_SEGMENT|12105,12114|false|false|false|C0023660|lidocaine|Lidocaine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12105,12114|false|false|false|C0023660|lidocaine|Lidocaine
Event|Event|SIMPLE_SEGMENT|12105,12114|false|false|false|||Lidocaine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|12105,12114|false|false|false|C0202404|Lidocaine measurement|Lidocaine
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|12118,12123|false|false|false|C0445403;C1533128;C1707974|Body tissue patch material;Human patch material;Patch - Extended Release Film|Patch
Event|Event|SIMPLE_SEGMENT|12118,12123|false|false|false|||Patch
Finding|Finding|SIMPLE_SEGMENT|12118,12123|false|false|false|C0332461|Plaque (lesion)|Patch
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|12126,12130|false|false|false|C4308013|PTCH1 protein, human|PTCH
Event|Event|SIMPLE_SEGMENT|12126,12130|false|false|false|||PTCH
Finding|Gene or Genome|SIMPLE_SEGMENT|12126,12130|false|false|false|C0694887;C1705339;C1826732;C4308013|PTCH gene;PTCH1 gene;PTCH1 protein, human;PTCH1 wt Allele|PTCH
Finding|Receptor|SIMPLE_SEGMENT|12126,12130|false|false|false|C0694887;C1705339;C1826732;C4308013|PTCH gene;PTCH1 gene;PTCH1 protein, human;PTCH1 wt Allele|PTCH
Event|Event|SIMPLE_SEGMENT|12134,12137|false|false|false|||QPM
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12144,12154|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|12144,12154|false|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|12144,12154|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|SIMPLE_SEGMENT|12160,12164|false|false|false|||held
Event|Event|SIMPLE_SEGMENT|12173,12180|true|false|false|||restart
Drug|Organic Chemical|SIMPLE_SEGMENT|12181,12190|true|false|false|C0023660|lidocaine|Lidocaine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12181,12190|true|false|false|C0023660|lidocaine|Lidocaine
Event|Event|SIMPLE_SEGMENT|12181,12190|true|false|false|||Lidocaine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|12181,12190|true|false|false|C0202404|Lidocaine measurement|Lidocaine
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|12194,12199|true|false|false|C0445403;C1533128;C1707974|Body tissue patch material;Human patch material;Patch - Extended Release Film|Patch
Event|Event|SIMPLE_SEGMENT|12194,12199|true|false|false|||Patch
Finding|Finding|SIMPLE_SEGMENT|12194,12199|true|false|false|C0332461|Plaque (lesion)|Patch
Event|Event|SIMPLE_SEGMENT|12210,12215|false|false|false|||speak
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12227,12230|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|12227,12230|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|12227,12230|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|12227,12230|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|SIMPLE_SEGMENT|12227,12230|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|12227,12230|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|SIMPLE_SEGMENT|12227,12230|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12227,12230|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|SIMPLE_SEGMENT|12227,12230|false|false|false|||PCP
Finding|Gene or Genome|SIMPLE_SEGMENT|12227,12230|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|SIMPLE_SEGMENT|12227,12230|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Event|SIMPLE_SEGMENT|12239,12243|false|false|false|||Home
Finding|Idea or Concept|SIMPLE_SEGMENT|12239,12243|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|SIMPLE_SEGMENT|12239,12243|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|SIMPLE_SEGMENT|12239,12243|false|false|false|C1553498|home health encounter|Home
Event|Occupational Activity|SIMPLE_SEGMENT|12249,12256|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|12249,12256|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Event|Event|SIMPLE_SEGMENT|12259,12267|false|false|false|||Facility
Finding|Intellectual Product|SIMPLE_SEGMENT|12259,12267|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|SIMPLE_SEGMENT|12275,12284|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|12275,12284|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|12275,12284|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|12275,12284|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|12275,12284|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|12275,12294|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12285,12294|false|false|false|C0945731||Diagnosis
Event|Event|SIMPLE_SEGMENT|12285,12294|false|false|false|||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|12285,12294|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|12285,12294|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|12285,12294|false|false|false|C0011900|Diagnosis|Diagnosis
Finding|Finding|SIMPLE_SEGMENT|12312,12320|false|false|false|C0241863|Diabetic|Diabetic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12312,12325|false|false|false|C0206172|Diabetic Foot|Diabetic foot
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12312,12331|false|false|false|C1456868|Diabetic foot ulcer|Diabetic foot ulcer
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|12321,12325|false|false|false|C0016504;C4299097|Foot;Lower extremity>Foot|foot
Finding|Finding|SIMPLE_SEGMENT|12321,12325|false|false|false|C0555980|Foot problem|foot
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12321,12331|false|false|false|C0085119|Foot Ulcer|foot ulcer
Event|Event|SIMPLE_SEGMENT|12326,12331|false|false|false|||ulcer
Finding|Body Substance|SIMPLE_SEGMENT|12326,12331|false|false|false|C0041582;C1547940;C1550672|Specimen Type - Ulcer;Ulcer|ulcer
Finding|Intellectual Product|SIMPLE_SEGMENT|12326,12331|false|false|false|C0041582;C1547940;C1550672|Specimen Type - Ulcer;Ulcer|ulcer
Finding|Pathologic Function|SIMPLE_SEGMENT|12326,12331|false|false|false|C0041582;C1547940;C1550672|Specimen Type - Ulcer;Ulcer|ulcer
Finding|Finding|SIMPLE_SEGMENT|12332,12340|false|false|false|C0241863|Diabetic|Diabetic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12332,12353|false|false|false|C0011880|Diabetic Ketoacidosis|Diabetic ketoacidosis
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12332,12353|false|false|false|C1504665|Products Used to Treat Diabetic Ketoacidosis|Diabetic ketoacidosis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12341,12353|false|false|false|C0220982|Ketoacidosis|ketoacidosis
Event|Event|SIMPLE_SEGMENT|12341,12353|false|false|false|||ketoacidosis
Anatomy|Body Location or Region|SIMPLE_SEGMENT|12355,12360|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|SIMPLE_SEGMENT|12355,12360|false|false|false|C0741025|Chest problem|Chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12355,12365|false|false|false|C2926613||Chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|12355,12365|false|false|false|C0008031|Chest Pain|Chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12361,12365|false|true|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|12361,12365|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|12361,12365|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|12361,12365|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Disorder|Neoplastic Process|SIMPLE_SEGMENT|12368,12377|false|false|false|C0027627|Neoplasm Metastasis|SECONDARY
Event|Event|SIMPLE_SEGMENT|12368,12377|false|false|false|||SECONDARY
Finding|Functional Concept|SIMPLE_SEGMENT|12368,12377|false|false|false|C1522484|metastatic qualifier|SECONDARY
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12388,12396|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|DIABETES
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12388,12405|false|false|false|C0011849|Diabetes Mellitus|DIABETES MELLITUS
Event|Event|SIMPLE_SEGMENT|12397,12405|false|false|false|||MELLITUS
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|12407,12414|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|INSULIN
Drug|Hormone|SIMPLE_SEGMENT|12407,12414|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|INSULIN
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12407,12414|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|INSULIN
Event|Event|SIMPLE_SEGMENT|12407,12414|false|false|false|||INSULIN
Finding|Gene or Genome|SIMPLE_SEGMENT|12407,12414|false|false|false|C1337112|INS gene|INSULIN
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|12407,12414|false|false|false|C0202098|Insulin measurement|INSULIN
Finding|Functional Concept|SIMPLE_SEGMENT|12415,12424|false|false|false|C3244310|dependent|DEPENDENT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12426,12430|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12426,12430|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|SIMPLE_SEGMENT|12426,12430|false|false|false|||COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|12426,12430|false|false|false|C1412502|ARCN1 gene|COPD
Event|Event|SIMPLE_SEGMENT|12434,12443|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|12434,12443|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|12434,12443|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|12434,12443|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|12434,12443|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12444,12453|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12444,12453|false|false|false|C0012634|Disease|Condition
Event|Event|SIMPLE_SEGMENT|12444,12453|false|false|false|||Condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|12444,12453|false|false|false|C1705253|Logical Condition|Condition
Finding|Mental Process|SIMPLE_SEGMENT|12455,12461|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12455,12468|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|SIMPLE_SEGMENT|12455,12468|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12462,12468|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|12462,12468|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|12470,12475|false|false|false|||Clear
Finding|Idea or Concept|SIMPLE_SEGMENT|12470,12475|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|SIMPLE_SEGMENT|12480,12488|false|false|false|||coherent
Finding|Finding|SIMPLE_SEGMENT|12480,12488|false|false|false|C4068804|Coherent|coherent
Event|Event|SIMPLE_SEGMENT|12490,12495|false|false|false|||Level
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12490,12512|false|false|false|C4050479||Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|12490,12512|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|SIMPLE_SEGMENT|12499,12512|false|false|false|||Consciousness
Finding|Finding|SIMPLE_SEGMENT|12499,12512|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|SIMPLE_SEGMENT|12499,12512|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12514,12519|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|12514,12519|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12514,12519|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|SIMPLE_SEGMENT|12514,12519|false|false|false|||Alert
Finding|Finding|SIMPLE_SEGMENT|12514,12519|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|12514,12519|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|12514,12519|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|SIMPLE_SEGMENT|12524,12535|false|false|false|||interactive
Finding|Functional Concept|SIMPLE_SEGMENT|12524,12535|false|false|false|C1704675|Interaction|interactive
Event|Activity|SIMPLE_SEGMENT|12537,12545|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|12537,12545|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|SIMPLE_SEGMENT|12537,12545|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12546,12552|false|false|false|C5889824||Status
Event|Event|SIMPLE_SEGMENT|12546,12552|false|false|false|||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|12546,12552|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|12554,12564|false|false|false|||Ambulatory
Finding|Functional Concept|SIMPLE_SEGMENT|12554,12564|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|SIMPLE_SEGMENT|12554,12564|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|SIMPLE_SEGMENT|12554,12564|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|SIMPLE_SEGMENT|12554,12564|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|SIMPLE_SEGMENT|12567,12578|false|false|false|||Independent
Finding|Finding|SIMPLE_SEGMENT|12567,12578|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|SIMPLE_SEGMENT|12567,12578|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Event|Event|SIMPLE_SEGMENT|12583,12592|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|12583,12592|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|12583,12592|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|12583,12592|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|12583,12592|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12583,12605|false|false|false|C3669312||Discharge Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|12583,12605|false|false|false|C4282220|Discharge instructions|Discharge Instructions
Procedure|Health Care Activity|SIMPLE_SEGMENT|12583,12605|false|false|false|C2266673|hospital discharge instructions (treatment)|Discharge Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12593,12605|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|12593,12605|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|12593,12605|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Finding|Gene or Genome|SIMPLE_SEGMENT|12607,12611|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Event|Event|SIMPLE_SEGMENT|12632,12640|false|false|false|||pleasure
Finding|Intellectual Product|SIMPLE_SEGMENT|12632,12640|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|SIMPLE_SEGMENT|12632,12640|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|SIMPLE_SEGMENT|12648,12652|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|12648,12652|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|12648,12652|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|12648,12652|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|12648,12655|false|false|false|C1555558|care of - AddressPartType|care of
Event|Event|SIMPLE_SEGMENT|12684,12687|false|false|false|||WAS
Event|Event|SIMPLE_SEGMENT|12697,12705|false|false|false|||HOSPITAL
Finding|Idea or Concept|SIMPLE_SEGMENT|12697,12705|false|false|false|C1547192|Organization unit type - Hospital|HOSPITAL
Event|Event|SIMPLE_SEGMENT|12750,12758|false|false|false|||admitted
Anatomy|Body Location or Region|SIMPLE_SEGMENT|12775,12780|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|12775,12780|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12775,12785|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|12775,12785|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12781,12785|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|12781,12785|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|12781,12785|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|12781,12785|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|12806,12813|true|false|false|C1184743|bony process|process
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12806,12813|true|false|false|C1951340|Process Pharmacologic Substance|process
Event|Event|SIMPLE_SEGMENT|12806,12813|true|false|false|||process
Finding|Functional Concept|SIMPLE_SEGMENT|12806,12813|true|false|false|C4521054|Process (qualifier value)|process
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|12806,12813|true|false|false|C1522240|Process|process
Event|Event|SIMPLE_SEGMENT|12814,12820|true|false|false|||called
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12821,12824|true|false|false|C0011880|Diabetic Ketoacidosis|DKA
Event|Event|SIMPLE_SEGMENT|12821,12824|true|false|false|||DKA
Event|Event|SIMPLE_SEGMENT|12834,12840|true|false|false|||taking
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|12849,12856|true|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|SIMPLE_SEGMENT|12849,12856|true|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12849,12856|true|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|SIMPLE_SEGMENT|12849,12856|true|false|false|||insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|12849,12856|true|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|12849,12856|true|false|false|C0202098|Insulin measurement|insulin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12876,12879|false|false|false|C4522181|Brachial Amyotrophic Diplegia|bad
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|12876,12879|false|false|false|C1530798|BAD protein, human|bad
Drug|Biologically Active Substance|SIMPLE_SEGMENT|12876,12879|false|false|false|C1530798|BAD protein, human|bad
Event|Event|SIMPLE_SEGMENT|12876,12879|false|false|false|||bad
Finding|Gene or Genome|SIMPLE_SEGMENT|12876,12879|false|false|false|C1366450|BAD gene|bad
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12880,12889|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|SIMPLE_SEGMENT|12880,12889|false|false|false|||infection
Finding|Pathologic Function|SIMPLE_SEGMENT|12880,12889|false|false|false|C3714514|Infection|infection
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|12898,12902|false|false|false|C0016504;C4299097|Foot;Lower extremity>Foot|foot
Finding|Finding|SIMPLE_SEGMENT|12898,12902|false|false|false|C0555980|Foot problem|foot
Event|Activity|SIMPLE_SEGMENT|12911,12919|false|false|false|C1709305|Occur (action)|HAPPENED
Event|Event|SIMPLE_SEGMENT|12911,12919|false|false|false|||HAPPENED
Finding|Idea or Concept|SIMPLE_SEGMENT|12927,12935|false|false|false|C1547192|Organization unit type - Hospital|HOSPITAL
Event|Event|SIMPLE_SEGMENT|12991,12996|false|false|false|||tests
Finding|Intellectual Product|SIMPLE_SEGMENT|12991,12996|false|false|false|C0392366|Tests (qualifier value)|tests
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|12991,12996|false|false|false|C0022885|Laboratory Procedures|tests
Event|Event|SIMPLE_SEGMENT|13000,13006|false|false|false|||figure
Anatomy|Body Location or Region|SIMPLE_SEGMENT|13019,13024|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|13019,13024|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13019,13029|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|13019,13029|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13025,13029|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|13025,13029|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|13025,13029|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|13025,13029|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|13035,13041|false|false|false|||caused
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|13047,13052|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|13047,13052|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|13047,13052|false|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13047,13059|false|false|false|C0027051|Myocardial Infarction|heart attack
Event|Event|SIMPLE_SEGMENT|13053,13059|false|false|false|||attack
Finding|Finding|SIMPLE_SEGMENT|13053,13059|false|false|false|C1261512;C1304680|Attack (finding);Attack behavior|attack
Finding|Social Behavior|SIMPLE_SEGMENT|13053,13059|false|false|false|C1261512;C1304680|Attack (finding);Attack behavior|attack
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13077,13083|false|false|false|C1718621|W stress|stress
Drug|Organic Chemical|SIMPLE_SEGMENT|13077,13083|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13077,13083|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Finding|Finding|SIMPLE_SEGMENT|13077,13083|false|false|false|C0038435|Stress|stress
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|13077,13088|false|false|false|C0015260;C3494508|Exercise stress test;Stress Test|stress test
Anatomy|Body Location or Region|SIMPLE_SEGMENT|13084,13088|false|false|false|C4318744|Test - temporal region|test
Event|Event|SIMPLE_SEGMENT|13084,13088|false|false|false|||test
Finding|Functional Concept|SIMPLE_SEGMENT|13084,13088|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Finding|Intellectual Product|SIMPLE_SEGMENT|13084,13088|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|13084,13088|false|false|false|C0456984|Test Result|test
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|13084,13088|false|false|false|C0022885|Laboratory Procedures|test
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|13103,13111|false|false|false|C4727483|BRAF Gene Rearrangement|positive
Event|Event|SIMPLE_SEGMENT|13103,13111|false|false|false|||positive
Finding|Classification|SIMPLE_SEGMENT|13103,13111|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|SIMPLE_SEGMENT|13103,13111|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Event|Event|SIMPLE_SEGMENT|13112,13119|false|false|false|||results
Finding|Intellectual Product|SIMPLE_SEGMENT|13124,13128|false|false|false|C1720594|Then - dosing instruction fragment|then
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13135,13144|false|false|false|C0945766||procedure
Event|Event|SIMPLE_SEGMENT|13135,13144|false|false|false|||procedure
Event|Occupational Activity|SIMPLE_SEGMENT|13135,13144|false|false|false|C1546467|Act Class - procedure|procedure
Finding|Functional Concept|SIMPLE_SEGMENT|13135,13144|false|false|false|C2700391|Procedure (set of actions)|procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|13135,13144|false|false|false|C0184661|Interventional procedure|procedure
Event|Event|SIMPLE_SEGMENT|13145,13151|false|false|false|||called
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|13154,13161|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|13154,13161|false|false|false|C1314974|Cardiac attachment|cardiac
Event|Event|SIMPLE_SEGMENT|13163,13167|false|false|false|||cath
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|13163,13167|false|false|false|C0007430|Catheterization|cath
Event|Event|SIMPLE_SEGMENT|13175,13181|true|false|false|||showed
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|13206,13211|true|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|13206,13211|true|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|13206,13211|true|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13206,13218|true|true|false|C0027051|Myocardial Infarction|heart attack
Event|Event|SIMPLE_SEGMENT|13212,13218|true|false|false|||attack
Finding|Finding|SIMPLE_SEGMENT|13212,13218|true|false|false|C1261512;C1304680|Attack (finding);Attack behavior|attack
Finding|Social Behavior|SIMPLE_SEGMENT|13212,13218|true|false|false|C1261512;C1304680|Attack (finding);Attack behavior|attack
Event|Event|SIMPLE_SEGMENT|13228,13239|false|false|false|||podiatrists
Event|Event|SIMPLE_SEGMENT|13246,13257|false|false|false|||debridement
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|13246,13257|false|false|false|C0011079;C3245462|Debridement;Sterile maggot wound debridement|debridement
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|13266,13270|false|false|false|C0016504;C4299097|Foot;Lower extremity>Foot|foot
Finding|Finding|SIMPLE_SEGMENT|13266,13270|false|false|false|C0555980|Foot problem|foot
Event|Event|SIMPLE_SEGMENT|13279,13283|false|false|false|||gave
Drug|Antibiotic|SIMPLE_SEGMENT|13288,13299|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|SIMPLE_SEGMENT|13288,13299|false|false|false|||antibiotics
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|13309,13313|false|false|false|C0016504;C4299097|Foot;Lower extremity>Foot|foot
Finding|Finding|SIMPLE_SEGMENT|13309,13313|false|false|false|C0555980|Foot problem|foot
Event|Event|SIMPLE_SEGMENT|13322,13330|false|false|false|||adjusted
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|13336,13343|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|SIMPLE_SEGMENT|13336,13343|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13336,13343|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|SIMPLE_SEGMENT|13336,13343|false|false|false|||insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|13336,13343|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|13336,13343|false|false|false|C0202098|Insulin measurement|insulin
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|13336,13350|false|false|false|C0428405|Insulin level|insulin levels
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|13336,13350|false|false|false|C0202098|Insulin measurement|insulin levels
Event|Event|SIMPLE_SEGMENT|13344,13350|false|false|false|||levels
Event|Event|SIMPLE_SEGMENT|13371,13375|false|false|false|||WHEN
Event|Event|SIMPLE_SEGMENT|13381,13385|false|false|false|||HOME
Finding|Idea or Concept|SIMPLE_SEGMENT|13381,13385|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|HOME
Finding|Intellectual Product|SIMPLE_SEGMENT|13381,13385|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|HOME
Procedure|Health Care Activity|SIMPLE_SEGMENT|13381,13385|false|false|false|C1553498|home health encounter|HOME
Event|Event|SIMPLE_SEGMENT|13426,13430|false|false|false|||Take
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13443,13454|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13443,13454|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|13443,13454|false|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|13443,13454|false|false|false|C4284232|Medications|medications
Drug|Antibiotic|SIMPLE_SEGMENT|13479,13490|false|false|false|C0008947|clindamycin|Clindamycin
Drug|Organic Chemical|SIMPLE_SEGMENT|13479,13490|false|false|false|C0008947|clindamycin|Clindamycin
Event|Event|SIMPLE_SEGMENT|13479,13490|false|false|false|||Clindamycin
Drug|Antibiotic|SIMPLE_SEGMENT|13495,13506|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|SIMPLE_SEGMENT|13495,13506|false|false|false|||antibiotics
Event|Event|SIMPLE_SEGMENT|13511,13515|false|false|false|||need
Event|Event|SIMPLE_SEGMENT|13520,13524|false|false|false|||take
Event|Event|SIMPLE_SEGMENT|13535,13546|false|false|false|||podiatrists
Event|Event|SIMPLE_SEGMENT|13574,13583|false|false|false|||scheduled
Event|Event|SIMPLE_SEGMENT|13588,13591|false|false|false|||see
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|13610,13617|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|SIMPLE_SEGMENT|13610,13617|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13610,13617|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|SIMPLE_SEGMENT|13610,13617|false|false|false|||insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|13610,13617|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|13610,13617|false|false|false|C0202098|Insulin measurement|insulin
Event|Event|SIMPLE_SEGMENT|13618,13625|false|false|false|||regimen
Finding|Intellectual Product|SIMPLE_SEGMENT|13618,13625|false|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|13618,13625|false|false|false|C0040808|Treatment Protocols|regimen
Event|Event|SIMPLE_SEGMENT|13643,13652|false|false|false|||different
Event|Event|SIMPLE_SEGMENT|13664,13667|false|false|false|||old
Event|Event|SIMPLE_SEGMENT|13668,13675|false|false|false|||regimen
Finding|Intellectual Product|SIMPLE_SEGMENT|13668,13675|false|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|13668,13675|false|false|false|C0040808|Treatment Protocols|regimen
Event|Event|SIMPLE_SEGMENT|13686,13690|false|false|false|||need
Event|Event|SIMPLE_SEGMENT|13694,13698|false|false|false|||take
Drug|Organic Chemical|SIMPLE_SEGMENT|13699,13706|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13699,13706|false|false|false|C0004057|aspirin|aspirin
Event|Event|SIMPLE_SEGMENT|13699,13706|false|false|false|||aspirin
Drug|Organic Chemical|SIMPLE_SEGMENT|13711,13723|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13711,13723|false|false|false|C0286651|atorvastatin|Atorvastatin
Finding|Idea or Concept|SIMPLE_SEGMENT|13730,13733|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|13730,13733|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|13746,13755|false|false|false|||blockages
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|13764,13769|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|13764,13769|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Event|Event|SIMPLE_SEGMENT|13764,13769|false|false|false|||heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|13764,13769|false|false|false|C0795691|HEART PROBLEM|heart
Event|Event|SIMPLE_SEGMENT|13775,13782|false|false|false|||forming
Event|Activity|SIMPLE_SEGMENT|13807,13819|false|false|false|C0003629|Appointments|appointments
Event|Event|SIMPLE_SEGMENT|13807,13819|false|false|false|||appointments
Finding|Idea or Concept|SIMPLE_SEGMENT|13827,13831|false|false|false|C1552851|next - HtmlLinkType|next
Finding|Intellectual Product|SIMPLE_SEGMENT|13832,13836|false|false|false|C1561540|Transaction counts and value totals - week|week
Event|Event|SIMPLE_SEGMENT|13850,13859|false|false|false|||important
Event|Event|SIMPLE_SEGMENT|13869,13871|false|false|false|||go
Event|Event|SIMPLE_SEGMENT|13897,13900|false|false|false|||get
Event|Event|SIMPLE_SEGMENT|13906,13912|false|false|false|||health
Finding|Idea or Concept|SIMPLE_SEGMENT|13906,13912|false|false|false|C0018684|Health|health
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13933,13939|false|false|false|C0944911||weight
Event|Event|SIMPLE_SEGMENT|13933,13939|false|false|false|||weight
Finding|Finding|SIMPLE_SEGMENT|13933,13939|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|SIMPLE_SEGMENT|13933,13939|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|SIMPLE_SEGMENT|13933,13939|false|false|false|C1305866|Weighing patient|weight
Event|Event|SIMPLE_SEGMENT|13943,13952|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|13943,13952|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|13943,13952|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|13943,13952|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|13943,13952|false|false|false|C0030685|Patient Discharge|discharge
Finding|Finding|SIMPLE_SEGMENT|14009,14016|false|false|false|C4534363|At home|at home
Event|Event|SIMPLE_SEGMENT|14012,14016|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|14012,14016|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|14012,14016|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|14012,14016|false|false|false|C1553498|home health encounter|home
Event|Event|SIMPLE_SEGMENT|14021,14024|false|false|false|||use
Finding|Finding|SIMPLE_SEGMENT|14038,14041|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|14038,14041|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|14042,14050|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|SIMPLE_SEGMENT|14042,14050|false|false|false|||baseline
Finding|Idea or Concept|SIMPLE_SEGMENT|14042,14050|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Event|Event|SIMPLE_SEGMENT|14062,14067|false|false|false|||weigh
Finding|Idea or Concept|SIMPLE_SEGMENT|14083,14086|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|14083,14086|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|14103,14107|false|false|false|||Call
Event|Event|SIMPLE_SEGMENT|14114,14120|false|false|false|||doctor
Finding|Intellectual Product|SIMPLE_SEGMENT|14114,14120|false|false|false|C2348314|Doctor - Title|doctor
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14129,14135|false|false|false|C0944911||weight
Event|Event|SIMPLE_SEGMENT|14129,14135|false|false|false|||weight
Finding|Finding|SIMPLE_SEGMENT|14129,14135|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|SIMPLE_SEGMENT|14129,14135|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|SIMPLE_SEGMENT|14129,14135|false|false|false|C1305866|Weighing patient|weight
Event|Event|SIMPLE_SEGMENT|14136,14140|false|false|false|||goes
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|14159,14162|false|false|false|C3161851|liquid-based cytology (procedure)|lbs
Finding|Intellectual Product|SIMPLE_SEGMENT|14169,14173|false|false|false|C5239649|PANEL.SURVEY.SEEK|Seek
Finding|Functional Concept|SIMPLE_SEGMENT|14174,14181|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Idea or Concept|SIMPLE_SEGMENT|14174,14181|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Intellectual Product|SIMPLE_SEGMENT|14174,14181|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|14174,14181|false|false|false|C0199168|Medical service|medical
Event|Event|SIMPLE_SEGMENT|14182,14191|false|false|false|||attention
Finding|Intellectual Product|SIMPLE_SEGMENT|14182,14191|false|false|false|C0004268;C4281780|Attention;Attention - G-code|attention
Finding|Mental Process|SIMPLE_SEGMENT|14182,14191|false|false|false|C0004268;C4281780|Attention;Attention - G-code|attention
Finding|Finding|SIMPLE_SEGMENT|14204,14207|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|14204,14207|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Event|Event|SIMPLE_SEGMENT|14222,14230|false|false|false|||symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|14222,14230|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|14222,14230|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|SIMPLE_SEGMENT|14247,14255|false|false|false|||swelling
Finding|Finding|SIMPLE_SEGMENT|14247,14255|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|SIMPLE_SEGMENT|14247,14255|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|14264,14268|false|false|false|C1140621|Leg|legs
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14264,14268|false|false|false|C5781420||legs
Anatomy|Body Location or Region|SIMPLE_SEGMENT|14270,14279|false|false|false|C0000726|Abdomen|abdominal
Finding|Finding|SIMPLE_SEGMENT|14270,14290|false|false|false|C0000731|Abdomen distended|abdominal distention
Event|Event|SIMPLE_SEGMENT|14280,14290|false|false|false|||distention
Finding|Finding|SIMPLE_SEGMENT|14280,14290|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distention
Finding|Pathologic Function|SIMPLE_SEGMENT|14280,14290|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distention
Event|Event|SIMPLE_SEGMENT|14296,14305|false|false|false|||shortness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14296,14315|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|SIMPLE_SEGMENT|14296,14315|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|SIMPLE_SEGMENT|14309,14315|false|false|false|C0225386|Breath|breath
Event|Event|SIMPLE_SEGMENT|14329,14338|false|false|false|||worsening
Finding|Idea or Concept|SIMPLE_SEGMENT|14329,14338|false|false|false|C1546960|Patient Outcome - Worsening|worsening
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14339,14343|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|14339,14343|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|14339,14343|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|14339,14343|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14347,14354|false|false|false|C0041834|Erythema|redness
Event|Event|SIMPLE_SEGMENT|14347,14354|false|false|false|||redness
Finding|Finding|SIMPLE_SEGMENT|14347,14354|false|false|false|C0332575|Redness|redness
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|14364,14368|false|false|false|C0016504;C4299097|Foot;Lower extremity>Foot|foot
Finding|Finding|SIMPLE_SEGMENT|14364,14368|false|false|false|C0555980|Foot problem|foot
Event|Event|SIMPLE_SEGMENT|14370,14379|false|false|false|||urinating
Event|Event|SIMPLE_SEGMENT|14399,14406|false|false|false|||thirsty
Finding|Finding|SIMPLE_SEGMENT|14399,14406|false|false|false|C0232471|Thirsty|thirsty
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14420,14425|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|14420,14425|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|14420,14425|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Drug|Organic Chemical|SIMPLE_SEGMENT|14420,14431|false|false|false|C0005802|Blood Glucose|blood sugar
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|14420,14431|false|false|false|C0392201|Blood glucose measurement|blood sugar
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|14426,14431|false|false|false|C0007004;C0242209;C3665462|Carbohydrates;Sugars;raw sugar|sugar
Drug|Organic Chemical|SIMPLE_SEGMENT|14426,14431|false|false|false|C0007004;C0242209;C3665462|Carbohydrates;Sugars;raw sugar|sugar
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14426,14431|false|false|false|C0007004;C0242209;C3665462|Carbohydrates;Sugars;raw sugar|sugar
Event|Event|SIMPLE_SEGMENT|14426,14431|false|false|false|||sugar
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|14477,14480|false|false|false|C0228225|Structure of calcar avis|cal
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|14477,14480|false|false|false|C1135160|monoclonal antibody CAL|cal
Drug|Immunologic Factor|SIMPLE_SEGMENT|14477,14480|false|false|false|C1135160|monoclonal antibody CAL|cal
Finding|Gene or Genome|SIMPLE_SEGMENT|14477,14480|false|false|false|C1425021;C1825283;C3273482;C5890925|FBLIM1 wt Allele;FBLP1 gene;GOPC gene;GOPC wt Allele|cal
Event|Event|SIMPLE_SEGMENT|14487,14493|false|false|false|||doctor
Finding|Intellectual Product|SIMPLE_SEGMENT|14487,14493|false|false|false|C2348314|Doctor - Title|doctor
Event|Event|SIMPLE_SEGMENT|14507,14515|false|false|false|||pleasure
Finding|Intellectual Product|SIMPLE_SEGMENT|14507,14515|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|SIMPLE_SEGMENT|14507,14515|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Event|SIMPLE_SEGMENT|14516,14529|false|false|false|||participating
Event|Activity|SIMPLE_SEGMENT|14538,14542|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|14538,14542|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|14538,14542|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|14538,14542|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Event|Activity|SIMPLE_SEGMENT|14579,14583|false|false|false|C1947933|care activity|Care
Finding|Finding|SIMPLE_SEGMENT|14579,14583|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|SIMPLE_SEGMENT|14579,14583|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14579,14588|false|false|false|C4321316||Care Team
Finding|Finding|SIMPLE_SEGMENT|14579,14588|false|false|false|C4321315|Care team|Care Team
Procedure|Health Care Activity|SIMPLE_SEGMENT|14595,14603|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14604,14616|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|14604,14616|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|14604,14616|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

