CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Neurosurgical Procedures|Procedure|false|false||NEUROSURGERYnull|Science of neurosurgery|Title|false|false||NEUROSURGERYnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|Known|Modifier|false|false||Knownnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|Adverse reaction to drug|Finding|true|false||Adverse Drug Reactionsnull|Adverse reaction to drug|Finding|true|false||Drug Reactionsnull|Pharmaceutical Preparations|Drug|false|false||Drug
null|Pharmacologic Substance|Drug|false|false||Drugnull|Drug problem|Finding|false|false||Drugnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Chief complaint (finding)|Finding|false|false||Chief Complaintnull|Complaint (finding)|Finding|false|false||Complaintnull|null|Attribute|false|false||Complaintnull|Headache|Finding|false|false||Headachesnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|suboccipital craniotomy|Procedure|false|false||Suboccipital craniotomynull|Suboccipital approach|Modifier|false|false||Suboccipitalnull|Craniotomy|Procedure|false|false||craniotomynull|removal technique|Procedure|false|false||resection
null|Excision|Procedure|false|false||resectionnull|Cerebellum|Anatomy|false|false||cerebellarnull|Lesion|Finding|false|false||lesion
null|null|Finding|false|false||lesionnull|History of present illness (finding)|Finding|false|false||History of Present Illnessnull|null|Attribute|false|false||History of Present Illnessnull|Medical History|Finding|false|false||History ofnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Present illness|Finding|false|false||Present Illnessnull|Present|Finding|false|false||Present
null|Presentation|Finding|false|false||Presentnull|Illness (finding)|Finding|false|false||Illnessnull|Females|Subject|false|false||female
null|Woman|Subject|false|false||femalenull|Female, Self-Report|Modifier|false|false||female
null|Female Phenotype|Modifier|false|false||femalenull|Cerebral Aneurysm|Disorder|false|false|C0228174;C0006104|cerebral aneurysmnull|Cerebral hemisphere structure (body structure)|Anatomy|false|false|C0917996;C0002940|cerebral
null|Brain|Anatomy|false|false|C0917996;C0002940|cerebralnull|Aneurysm|Finding|false|false|C0228174;C0006104|aneurysmnull|Closure by clip (procedure)|Procedure|false|false||clippingnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Cerebellum|Anatomy|false|false||cerebellarnull|Lesion|Finding|false|false||lesion
null|null|Finding|false|false||lesionnull|Patient-Reported|Finding|false|false||Patient reportsnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Report (document)|Finding|false|false||reportsnull|Reporting|Procedure|false|false||reportsnull|Three weeks|Time|false|false||three weeksnull|week|Time|false|false||weeksnull|FBXW7 wt Allele|Finding|false|false||ago
null|FBXW7 gene|Finding|false|false||agonull|Headache|Finding|false|false||headachesnull|Observation Interpretation - Abnormal|Finding|false|false||abnormal
null|Abnormal|Finding|false|false||abnormalnull|Headache|Finding|false|false||headachesnull|Global|Modifier|false|false||global
null|Generalized|Modifier|false|false||globalnull|Tylenol|Drug|false|false||Tylenol
null|Tylenol|Drug|false|false||Tylenolnull|Worst|Modifier|false|false||worstnull|Difficulty walking|Finding|false|false||difficulty walkingnull|Has difficulty doing (qualifier value)|Finding|false|false||difficultynull|history of recreational walking|Finding|false|false||walking
null|walking - neurological symptom|Finding|false|false||walking
null|Walking (function)|Finding|false|false||walkingnull|Three weeks|Time|false|false||three weeksnull|week|Time|false|false||weeksnull|FBXW7 wt Allele|Finding|false|false||ago
null|FBXW7 gene|Finding|false|false||agonull|history of recreational walking|Finding|false|false||walking
null|walking - neurological symptom|Finding|false|false||walking
null|Walking (function)|Finding|false|false||walkingnull|Cerebellar decompression injury|Disorder|false|false||staggeringnull|Staggering gait|Finding|false|false||staggeringnull|Side|Modifier|false|false||sidenull|side to side|Finding|false|false||to sidenull|Side|Modifier|false|false||sidenull|Vision|Finding|false|false||visionnull|null|Attribute|false|false||visionnull|Specialized Stand Alone Plan - Vision|Entity|false|false||visionnull|Changing|Finding|true|false||changesnull|Changed status|LabModifier|false|false||changesnull|Nausea|Finding|true|false||nauseanull|null|Attribute|true|false||nauseanull|Vomiting|Finding|true|false||vomitingnull|Confusion|Disorder|false|false||confusionnull|Clouded consciousness|Finding|false|false||confusionnull|Word finding difficulty (disorder)|Disorder|false|false||word finding difficultynull|Term (lexical)|Finding|false|false||wordnull|Experimental Finding|Finding|false|false||finding
null|Signs and Symptoms|Finding|false|false||finding
null|Finding|Finding|false|false||findingnull|Has difficulty doing (qualifier value)|Finding|false|false||difficultynull|Carcinoma in situ of eye|Disorder|false|false|C4266572;C0015392;C0700042|eye
null|Disorder of eye|Disorder|false|false|C4266572;C0015392;C0700042|eyenull|Eye - Specimen Source Code|Finding|false|false|C4266572;C0015392;C0700042|eye
null|Eye problem|Finding|false|false|C4266572;C0015392;C0700042|eye
null|Eye Specimen|Finding|false|false|C4266572;C0015392;C0700042|eyenull|Head>Eye|Anatomy|false|false|C2348314;C1550636;C1546630;C0262477;C0154094;C0015397|eye
null|Eye|Anatomy|false|false|C2348314;C1550636;C1546630;C0262477;C0154094;C0015397|eye
null|Orbital region|Anatomy|false|false|C2348314;C1550636;C1546630;C0262477;C0154094;C0015397|eyenull|Doctor - Title|Finding|false|false|C4266572;C0015392;C0700042|doctornull|Physicians|Subject|false|false||doctornull|Morning|Time|false|false||morningnull|Extended Priority Codes - Routine|Finding|false|false||routine
null|Report priority - Routine|Finding|false|false||routine
null|Admission Type - Routine|Finding|false|false||routine
null|Level of Care - Routine|Finding|false|false||routine
null|Processing priority - Routine|Finding|false|false||routine
null|Referral priority - Routine|Finding|false|false||routinenull|Routine coag|Procedure|false|false||routinenull|Priority - Routine|Time|false|false||routinenull|Routine|Modifier|false|false||routinenull|Visit|Finding|false|false||visitnull|Processing type - Evaluation|Finding|false|false||evaluationnull|Evaluation procedure|Procedure|false|false||evaluation
null|Evaluation|Procedure|false|false||evaluationnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Academic Research Enhancement Awards|Event|false|false||areanull|Geographic Locations|Entity|false|false||areanull|Area|Modifier|false|false||areanull|Table Cell Horizontal Align - left|Finding|false|false|C0007765|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Malignant neoplasm of cerebellum|Disorder|false|false|C0007765|cerebellumnull|Cerebellum|Anatomy|false|false|C0153640;C1552822|cerebellumnull|Underlying|Finding|false|false||underlyingnull|Lesion|Finding|false|false||lesion
null|null|Finding|false|false||lesionnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Aneurysm clip|Device|true|false||aneurysm clipnull|Aneurysm|Finding|false|false||aneurysmnull|CLIP - Codes for radiology reports|Finding|false|false||clip
null|CD74 gene|Finding|false|false||clip
null|CLIP2 gene|Finding|false|false||clip
null|CLIP1 gene|Finding|false|false||clip
null|POMC gene|Finding|false|false||clip
null|POMC wt Allele|Finding|false|false||clip
null|CLIP1 wt Allele|Finding|false|false||clipnull|Comprehensive Lifestyle Intervention Program|Procedure|false|false||clipnull|Clip|Device|false|false||clipnull|CYREN gene|Finding|true|false||MRInull|Magnetic resonance imaging service|Procedure|true|false||MRI
null|Magnetic Resonance Imaging|Procedure|true|false||MRInull|Maori Language|Entity|true|false||MRInull|Consistent with|Finding|false|false||compatiblenull|Compatible|Modifier|false|false||compatiblenull|PMH - past medical history|Finding|false|false||Past Medical History
null|Medical History|Finding|false|false||Past Medical Historynull|Medical History|Finding|false|false||Medical Historynull|Medical referral type|Finding|false|false||Medical
null|Medical|Finding|false|false||Medical
null|Medical school type|Finding|false|false||Medicalnull|Medical service|Procedure|false|false||Medicalnull|Medical History|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|History of present illness (finding)|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Hypertensive disease|Disorder|false|false||Hypertensionnull|Clipping arterial aneurysm|Procedure|false|false||aneurysm clippingnull|Aneurysm|Finding|false|false||aneurysmnull|Closure by clip (procedure)|Procedure|false|false||clippingnull|Social and personal history|Finding|false|false||Social History
null|Social History|Finding|false|false||Social Historynull|Social|Finding|false|false||Socialnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Family Medical History|Finding|false|false||Family Historynull|Entity Name Part Type - family|Finding|false|false||Family
null|Last Name|Finding|false|false||Family
null|Living Arrangement - Family|Finding|false|false||Family
null|Family (taxonomic)|Finding|false|false||Family
null|Family Collection|Finding|false|false||Familynull|Family|Subject|false|false||Familynull|History of present illness (finding)|Finding|false|true||History
null|History of previous events|Finding|false|true||History
null|Historical aspects qualifier|Finding|false|true||History
null|Medical History|Finding|false|true||History
null|Concept History|Finding|false|true||Historynull|History|Subject|false|false||Historynull|Known|Modifier|false|false||knownnull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Cerebrovascular accident|Disorder|false|false||strokenull|Stroke (heart beat)|Finding|false|false||strokenull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Aneurysm|Finding|true|false||aneurysmnull|physical examination (physical finding)|Finding|false|false||Physical Examnull|Physical Examination|Procedure|false|false||Physical Examnull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|On admission|Time|false|false||ON ADMISSIONnull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||Gen
null|GEN1 wt Allele|Finding|false|false||Gen
null|GEN1 gene|Finding|false|false||Gennull|Feeling comfortable|Finding|false|false||comfortablenull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|HEENT|Anatomy|false|false||HEENTnull|Pupil|Anatomy|false|false||Pupilsnull|Extraocular|Finding|false|false||EOMsnull|Full|Modifier|false|false||fullnull|Passive joint movement of neck (finding)|Finding|false|false|C0027530;C3159206|Neck
null|Neck problem|Finding|false|false|C0027530;C3159206|Necknull|dendritic spine neck|Anatomy|false|false|C0812434;C0684335|Neck
null|Neck|Anatomy|false|false|C0812434;C0684335|Necknull|Supple|Finding|false|false||Supplenull|Feels warm|Finding|false|false||Warmnull|warming process|Phenomenon|false|false||Warmnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Neurology speciality|Title|false|false||Neuronull|Neurologic (qualifier value)|Modifier|false|false||Neuronull|Mental state|Finding|false|false||Mental statusnull|null|Attribute|false|false||Mental status
null|null|Attribute|false|false||Mental statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||statusnull|null|Attribute|false|false||statusnull|Social status|Modifier|false|false||status
null|Status|Modifier|false|false||statusnull|Alert brand of caffeine|Drug|false|false||alert
null|Alert brand of caffeine|Drug|false|false||alertnull|Mentally alert|Finding|false|false||alert
null|Consciousness clear|Finding|false|false||alert
null|Alert note|Finding|false|false||alert
null|Alert|Finding|false|false||alertnull|null|Attribute|false|false||alertnull|cooperative|Entity|false|false||cooperativenull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Affect (mental function)|Finding|false|false||affectnull|assessment of affect|Procedure|false|false||affectnull|Mental Orientation|Finding|false|false||Orientationnull|Orientation, Spatial|Modifier|false|false||Orientation
null|Genomic Orientation|Modifier|false|false||Orientation
null|Orientation|Modifier|false|false||Orientationnull|Oriented to person|Finding|false|false||Oriented to personnull|Oriented to place|Finding|false|false||Orientednull|Orientation, Spatial|Modifier|false|false||Orientednull|Person Info|Finding|false|false||personnull|null|Attribute|false|false||personnull|Persons|Subject|false|false||personnull|Place - dosing instruction imperative|Finding|false|false||placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|Programming Languages|Finding|false|false||Languagenull|null|Attribute|false|false||Languagenull|Languages|Entity|false|false||Languagenull|Speech|Finding|false|false||Speechnull|Speech assessment|Procedure|false|false||Speechnull|Language Ability Proficiency - Good|Finding|false|false||good
null|Language Proficiency - Good|Finding|false|false||goodnull|Specimen Quality - Good|Modifier|false|false||good
null|Good|Modifier|false|false||goodnull|Comprehension|Finding|false|false||comprehensionnull|speech fluency repetition (physical finding)|Finding|false|false||repetition
null|Repeat|Finding|false|false||repetitionnull|Naming (function)|Finding|false|false||Namingnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Dysarthria|Disorder|true|false||dysarthrianull|error|Modifier|false|false||errorsnull|Neoplasm of uncertain or unknown behavior of cranial nerves|Disorder|false|false|C0027740;C0010268;C0037303|Cranial Nerves
null|Benign neoplasm of cranial nerves|Disorder|false|false|C0027740;C0010268;C0037303|Cranial Nervesnull|Cranial Nerves|Anatomy|false|false|C0004992;C0496937|Cranial Nervesnull|Bone structure of cranium|Anatomy|false|false|C0004992;C0496937|Cranialnull|Cranial|Modifier|false|false||Cranialnull|Nerve|Anatomy|false|false|C0004992;C0496937|Nervesnull|Structure of pupil of left eye|Anatomy|false|false|C1552822;C1552823|Left pupilnull|Table Cell Horizontal Align - left|Finding|false|false|C0034121;C1305618;C0229187|Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|null|Anatomy|false|false|C1552822|pupil
null|Pupil|Anatomy|false|false|C1552822|pupilnull|Table Cell Horizontal Align - right|Finding|false|false|C0229187|rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Reactive Therapy|Procedure|false|false||reactivenull|Reactive|Modifier|false|false||reactivenull|TNFSF14 protein, human|Drug|false|false||light
null|TNFSF14 protein, human|Drug|false|false||lightnull|Light - subjective measurement|Finding|false|false||light
null|TNFSF14 wt Allele|Finding|false|false||light
null|TNFSF14 gene|Finding|false|false||light
null|Light color|Finding|false|false||lightnull|Phototherapy|Procedure|false|false||lightnull|Light|Phenomenon|false|false||lightnull|Light (qualifier)|Modifier|false|false||lightnull|examination of extraocular movements|Procedure|false|false||Extraocular movementsnull|Extraocular|Finding|false|false||Extraocularnull|Movement|Finding|false|false||movementsnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Nystagmus|Disorder|false|false||nystagmusnull|Roman numeral VII|Finding|false|false|C2338708;C3496273;C3496274|VIInull|Lamina VII of gray matter of spinal cord|Anatomy|false|false|C0445385|VII
null|lobule VII|Anatomy|false|false|C0445385|VII
null|layer VII (Cajal)|Anatomy|false|false|C0445385|VIInull|Face|Anatomy|false|false|C0808080|Facialnull|Facial|Modifier|false|false||Facialnull|Strength (attribute)|Finding|false|false|C0015450|strengthnull|Pharmaceutical Strength|LabModifier|false|false||strength
null|Physical Strength|LabModifier|false|false||strengthnull|Observation of Sensation|Finding|false|false||sensation
null|Sensory perception|Finding|false|false||sensationnull|sensory exam|Procedure|false|false||sensationnull|Sensation quality|Modifier|false|false||sensationnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Symmetric Relationship|Finding|false|false||symmetric
null|Symmetrical|Finding|false|false||symmetricnull|Structure of sternocleidomastoid muscle|Anatomy|false|false||Sternocleidomastoidnull|Structure of trapezius muscle|Anatomy|false|false||trapeziusnull|tongue midline|Finding|false|false|C1660780;C0040408|Tongue midlinenull|Benign neoplasm of tongue|Disorder|false|false|C1660780;C0040408|Tonguenull|Procedure on tongue|Procedure|false|false|C0040408;C1660780|Tonguenull|Tongue|Anatomy|false|false|C0015644;C3693372;C0153933;C0872394|Tonguenull|midline cell component|Anatomy|false|false|C0153933;C3693372;C0015644;C0872394|midlinenull|Midline (qualifier value)|Modifier|false|false||midlinenull|Muscular fasciculation|Finding|true|false|C0040408;C1660780|fasciculationsnull|motor movement|Finding|false|false||Motornull|Motor Device|Device|false|false||Motornull|Bulk (conceptual)|Drug|false|false||bulk
null|Dietary Fiber|Drug|false|false||bulknull|Dyskinetic syndrome|Disorder|true|false||abnormal movementsnull|Abnormal movement|Finding|true|false||abnormal movementsnull|Observation Interpretation - Abnormal|Finding|false|false||abnormal
null|Abnormal|Finding|false|false||abnormalnull|Movement|Finding|true|false||movementsnull|Tremor|Finding|false|false||tremorsnull|Strength (attribute)|Finding|false|false||Strengthnull|Pharmaceutical Strength|LabModifier|false|false||Strength
null|Physical Strength|LabModifier|false|false||Strengthnull|Full|Modifier|false|false||fullnull|Power (Psychology)|Finding|false|false||powernull|Power|LabModifier|false|false||powernull|Intensity and Distress 1|Finding|false|false||Slightnull|Slight (qualifier value)|Modifier|false|false||Slight
null|Mild (qualifier value)|Modifier|false|false||Slightnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Upward|Modifier|false|false||upwardnull|Observation of Sensation|Finding|false|false||Sensation
null|Sensory perception|Finding|false|false||Sensationnull|sensory exam|Procedure|false|false||Sensationnull|Sensation quality|Modifier|false|false||Sensationnull|Gender Status - Intact|Finding|false|false||Intactnull|Intact|Modifier|false|false||Intactnull|Light touch|Finding|false|false||light touchnull|TNFSF14 protein, human|Drug|false|false||light
null|TNFSF14 protein, human|Drug|false|false||lightnull|Light - subjective measurement|Finding|false|false||light
null|TNFSF14 wt Allele|Finding|false|false||light
null|TNFSF14 gene|Finding|false|false||light
null|Light color|Finding|false|false||lightnull|Phototherapy|Procedure|false|false||lightnull|Light|Phenomenon|false|false||lightnull|Light (qualifier)|Modifier|false|false||lightnull|Touch Perception|Finding|false|false||touch
null|Touch sensation|Finding|false|false||touchnull|Therapeutic Touch|Procedure|false|false||touchnull|Tactile|Modifier|false|false||touchnull|Coordination of Benefits - Coordination|Finding|false|false||Coordination
null|Coordinated|Finding|false|false||Coordination
null|Physiologic Coordination|Finding|false|false||Coordinationnull|Upper extremity>Finger|Anatomy|false|false||finger
null|Fingers|Anatomy|false|false||finger
null|Fingers not including thumb|Anatomy|false|false||fingernull|Upper extremity>Finger|Anatomy|false|false||finger
null|Fingers|Anatomy|false|false||finger
null|Fingers not including thumb|Anatomy|false|false||fingernull|Heel|Anatomy|false|false||heelnull|Shin|Anatomy|false|false||shinnull|On discharge|Time|false|false||ON DISCHARGEnull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|Eye|Anatomy|false|false|C5848506|eyesnull|null|Attribute|false|false|C0015392|eyesnull|Mental Orientation|Finding|false|false||Orientationnull|Orientation, Spatial|Modifier|false|false||Orientation
null|Genomic Orientation|Modifier|false|false||Orientation
null|Orientation|Modifier|false|false||Orientationnull|Person Info|Finding|false|false||Personnull|null|Attribute|false|false||Personnull|Persons|Subject|false|false||Personnull|Place - dosing instruction imperative|Finding|false|false||Placenull|null|Procedure|false|false||Placenull|put - instruction imperative|Event|false|false||Placenull|Place|Modifier|false|false||Placenull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||Time
null|Time (foundation metadata concept)|Finding|false|false||Time
null|Value type - Time|Finding|false|false||Time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||Time
null|Data types - Time|Finding|false|false||Time
null|null|Finding|false|false||Timenull|Time|Time|false|false||Timenull|LITAF gene|Finding|false|false||Simplenull|Simple|Modifier|false|false||Simplenull|complex (molecular entity)|Drug|false|false||Complexnull|Complex|Modifier|false|false||Complexnull|Pupil|Anatomy|false|false||Pupilsnull|Table Cell Horizontal Align - right|Finding|false|false||Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|Table Cell Horizontal Align - left|Finding|false|false||Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Extraocular|Finding|false|false|C0028863|EOMnull|Muscle of orbit|Anatomy|false|false|C0241886|EOMnull|Full|Modifier|false|false||Fullnull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Prominent|Modifier|false|false||prominentnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Lateral|Modifier|false|false||lateralnull|FANCONI ANEMIA, COMPLEMENTATION GROUP E|Disorder|false|false|C0015450;C4266571|Facenull|FANCE wt Allele|Finding|false|false|C0015450;C4266571|Face
null|FANCE gene|Finding|false|false|C0015450;C4266571|Face
null|ELOVL6 gene|Finding|false|false|C0015450;C4266571|Facenull|Head>Face|Anatomy|false|false|C3160739;C1423759;C2828055;C1414531;C0332516;C2699744|Face
null|Face|Anatomy|false|false|C3160739;C1423759;C2828055;C1414531;C0332516;C2699744|Facenull|Face (spatial concept)|Modifier|false|false||Facenull|Symmetric Relationship|Finding|false|false|C0015450;C4266571|Symmetric
null|Symmetrical|Finding|false|false|C0015450;C4266571|Symmetricnull|Yes - Expanded yes/no indicator|Finding|false|false||Yes
null|Yes (qualifier value)|Finding|false|false||Yes
null|Yes - Identity May Be Divulged|Finding|false|false||Yes
null|Yes (indicator)|Finding|false|false||Yes
null|Yes|Finding|false|false||Yes
null|Yes - Yes/no indicator|Finding|false|false||Yes
null|Yes - Event Expected|Finding|false|false||Yes
null|Yes - Assignment of Benefits|Finding|false|false||Yes
null|YES1 wt Allele|Finding|false|false||Yes
null|YES1 gene|Finding|false|false||Yes
null|Yes - Release Information|Finding|false|false||Yes
null|YES Portal|Finding|false|false||Yes
null|Yes - Notify Clergy Code|Finding|false|false||Yesnull|Yes - Event Seriousness|Modifier|false|false||Yesnull|midline cell component|Anatomy|false|false||Midlinenull|Midline (qualifier value)|Modifier|false|false||Midlinenull|Yes - Expanded yes/no indicator|Finding|false|false||Yes
null|Yes (qualifier value)|Finding|false|false||Yes
null|Yes - Identity May Be Divulged|Finding|false|false||Yes
null|Yes (indicator)|Finding|false|false||Yes
null|Yes|Finding|false|false||Yes
null|Yes - Yes/no indicator|Finding|false|false||Yes
null|Yes - Event Expected|Finding|false|false||Yes
null|Yes - Assignment of Benefits|Finding|false|false||Yes
null|YES1 wt Allele|Finding|false|false||Yes
null|YES1 gene|Finding|false|false||Yes
null|Yes - Release Information|Finding|false|false||Yes
null|YES Portal|Finding|false|false||Yes
null|Yes - Notify Clergy Code|Finding|false|false||Yesnull|Yes - Event Seriousness|Modifier|false|false||Yesnull|Pronator drift|Finding|false|false||Pronator Driftnull|Yes - Expanded yes/no indicator|Finding|false|false||Yes
null|Yes (qualifier value)|Finding|false|false||Yes
null|Yes - Identity May Be Divulged|Finding|false|false||Yes
null|Yes (indicator)|Finding|false|false||Yes
null|Yes|Finding|false|false||Yes
null|Yes - Yes/no indicator|Finding|false|false||Yes
null|Yes - Event Expected|Finding|false|false||Yes
null|Yes - Assignment of Benefits|Finding|false|false||Yes
null|YES1 wt Allele|Finding|false|false||Yes
null|YES1 gene|Finding|false|false||Yes
null|Yes - Release Information|Finding|false|false||Yes
null|YES Portal|Finding|false|false||Yes
null|Yes - Notify Clergy Code|Finding|false|false||Yesnull|Yes - Event Seriousness|Modifier|false|false||Yesnull|Speech|Finding|true|false||Speechnull|Speech assessment|Procedure|true|false||Speechnull|Yes - Expanded yes/no indicator|Finding|false|false||Yes
null|Yes (qualifier value)|Finding|false|false||Yes
null|Yes - Identity May Be Divulged|Finding|false|false||Yes
null|Yes (indicator)|Finding|false|false||Yes
null|Yes|Finding|false|false||Yes
null|Yes - Yes/no indicator|Finding|false|false||Yes
null|Yes - Event Expected|Finding|false|false||Yes
null|Yes - Assignment of Benefits|Finding|false|false||Yes
null|YES1 wt Allele|Finding|false|false||Yes
null|YES1 gene|Finding|false|false||Yes
null|Yes - Release Information|Finding|false|false||Yes
null|YES Portal|Finding|false|false||Yes
null|Yes - Notify Clergy Code|Finding|false|false||Yesnull|Yes - Event Seriousness|Modifier|false|false||Yesnull|Comprehension|Finding|false|false||Comprehensionnull|Gender Status - Intact|Finding|false|false||Intactnull|Intact|Modifier|false|false||Intactnull|Yes - Expanded yes/no indicator|Finding|false|false||Yes
null|Yes (qualifier value)|Finding|false|false||Yes
null|Yes - Identity May Be Divulged|Finding|false|false||Yes
null|Yes (indicator)|Finding|false|false||Yes
null|Yes|Finding|false|false||Yes
null|Yes - Yes/no indicator|Finding|false|false||Yes
null|Yes - Event Expected|Finding|false|false||Yes
null|Yes - Assignment of Benefits|Finding|false|false||Yes
null|YES1 wt Allele|Finding|false|false||Yes
null|YES1 gene|Finding|false|false||Yes
null|Yes - Release Information|Finding|false|false||Yes
null|YES Portal|Finding|false|false||Yes
null|Yes - Notify Clergy Code|Finding|false|false||Yesnull|Yes - Event Seriousness|Modifier|false|false||Yesnull|motor movement|Finding|false|false||Motornull|Motor Device|Device|false|false||Motornull|Table Cell Horizontal Align - right|Finding|false|false||Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|Table Cell Horizontal Align - left|Finding|false|false||Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|Observation of Sensation|Finding|false|false||Sensation
null|Sensory perception|Finding|false|false||Sensationnull|sensory exam|Procedure|false|false||Sensationnull|Sensation quality|Modifier|false|false||Sensationnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Light touch|Finding|false|false||light touchnull|TNFSF14 protein, human|Drug|false|false||light
null|TNFSF14 protein, human|Drug|false|false||lightnull|Light - subjective measurement|Finding|false|false||light
null|TNFSF14 wt Allele|Finding|false|false||light
null|TNFSF14 gene|Finding|false|false||light
null|Light color|Finding|false|false||lightnull|Phototherapy|Procedure|false|false||lightnull|Light|Phenomenon|false|false||lightnull|Light (qualifier)|Modifier|false|false||lightnull|Touch sensation|Finding|false|false||touch
null|Touch Perception|Finding|false|false||touchnull|Therapeutic Touch|Procedure|false|false||touchnull|Tactile|Modifier|false|false||touchnull|ATP5F1A gene|Finding|false|false||OMRnull|AML Lab Table|Finding|false|false||lab
null|LAT2 gene|Finding|false|false||lab
null|EWS Lab Table|Finding|false|false||labnull|Laboratory|Device|false|false||labnull|Labrador retriever|Entity|false|false||lab
null|Laboratory|Entity|false|false||labnull|Imaging problem|Finding|false|false||imagingnull|Diagnostic Imaging|Procedure|false|false||imaging
null|Imaging Techniques|Procedure|false|false||imagingnull|Imaging Technology|Title|false|false||imagingnull|BRIEF Health Literacy Screening Tool|Finding|false|false||Brief
null|Behavior Rating Inventory of Executive Function|Finding|false|false||Briefnull|Brief|Time|false|false||Briefnull|Shortened|Modifier|false|false||Briefnull|Hospital course|Finding|false|false||Hospital Coursenull|null|Attribute|false|false||Hospital Coursenull|Organization unit type - Hospital|Finding|false|false||Hospitalnull|Hospitals|Device|false|false||Hospitalnull|Hospitals|Entity|false|false||Hospitalnull|Hospital environment|Modifier|false|false||Hospitalnull|Course|Time|false|false||Coursenull|Lesion of brain|Finding|false|false|C4266577;C0006104|Brain lesionnull|Brain Diseases|Disorder|false|false|C4266577;C0006104|Brainnull|Head>Brain|Anatomy|false|false|C0221505;C1546698;C0221198;C0006111|Brain
null|Brain|Anatomy|false|false|C0221505;C1546698;C0221198;C0006111|Brainnull|Lesion|Finding|false|false|C4266577;C0006104|lesion
null|null|Finding|false|false|C4266577;C0006104|lesionnull|Relationship modifier - Patient|Finding|false|false|C0007765|Patient
null|Specimen Type - Patient|Finding|false|false|C0007765|Patient
null|Mail Claim Party - Patient|Finding|false|false|C0007765|Patient
null|Report source - Patient|Finding|false|false|C0007765|Patient
null|null|Finding|false|false|C0007765|Patient
null|Disabled Person Code - Patient|Finding|false|false|C0007765|Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Cerebellum|Anatomy|false|false|C1578483;C1550655;C1578481;C1578486;C1578484;C1578485|cerebellarnull|National Center for Health Care Technology, U.S.|Entity|false|false||NCHCTnull|Contrast Media|Drug|false|false||contrastnull|Contrast|Modifier|false|false||contrastnull|mass lesion|Disorder|false|false||mass lesionnull|Morphology, Attenuation, Size, and Structure Criteria|Finding|false|false||mass
null|null|Finding|false|false||mass
null|FBN1 wt Allele|Finding|false|false||mass
null|FBN1 gene|Finding|false|false||mass
null|Mass of body region|Finding|false|false||mass
null|Mass of body structure|Finding|false|false||massnull|Mass, a measure of quantity of matter|LabModifier|false|false||mass
null|Molecular Mass|LabModifier|false|false||massnull|Lesion|Finding|false|false||lesion
null|null|Finding|false|false||lesionnull|Hydrocephalus|Disorder|false|false||hydrocephalusnull|Unable|Finding|false|false||unablenull|CYREN gene|Finding|false|false||MRInull|Magnetic resonance imaging service|Procedure|false|false||MRI
null|Magnetic Resonance Imaging|Procedure|false|false||MRInull|Maori Language|Entity|false|false||MRInull|Aneurysm clip|Device|false|false||aneurysm clipnull|Aneurysm|Finding|false|false||aneurysmnull|CLIP - Codes for radiology reports|Finding|false|false||clip
null|CD74 gene|Finding|false|false||clip
null|CLIP2 gene|Finding|false|false||clip
null|CLIP1 gene|Finding|false|false||clip
null|POMC gene|Finding|false|false||clip
null|POMC wt Allele|Finding|false|false||clip
null|CLIP1 wt Allele|Finding|false|false||clipnull|Comprehensive Lifestyle Intervention Program|Procedure|false|false||clipnull|Clip|Device|false|false||clipnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Close|Finding|false|false||close
null|Closed|Finding|false|false||closenull|Preventive monitoring|Procedure|false|false||monitoringnull|null|Event|false|false||monitoringnull|Operative Surgical Procedures|Procedure|false|false||surgical
null|Surgical service|Procedure|false|false||surgicalnull|null|Finding|false|false||planning
null|Planned|Finding|false|false||planningnull|dexamethasone|Drug|false|false||dexamethasone
null|dexamethasone|Drug|false|false||dexamethasonenull|Mass Effect|Finding|false|false||mass effectnull|Mass of body structure|Finding|false|false||mass
null|Morphology, Attenuation, Size, and Structure Criteria|Finding|false|false||mass
null|null|Finding|false|false||mass
null|FBN1 wt Allele|Finding|false|false||mass
null|FBN1 gene|Finding|false|false||mass
null|Mass of body region|Finding|false|false||massnull|Mass, a measure of quantity of matter|LabModifier|false|false||mass
null|Molecular Mass|LabModifier|false|false||massnull|Effect, Appearance|Modifier|false|false||effect
null|Effect|Modifier|false|false||effectnull|Trunk structure|Anatomy|false|false||torsonull|null|Finding|false|false|C4037972;C0024109|lung nodulesnull|Lung diseases|Disorder|false|false|C4037972;C0024109|lungnull|Lung Problem|Finding|false|false|C4037972;C0024109|lungnull|Chest>Lung|Anatomy|false|false|C0024115;C0740941;C0034079|lung
null|Lung|Anatomy|false|false|C0024115;C0740941;C0034079|lungnull|More|LabModifier|false|false||morenull|Acknowledgement Detail Type - Information|Finding|false|false||information
null|Error severity - Information|Finding|false|false||information
null|Information|Finding|false|false||information
null|control act - information|Finding|false|false||informationnull|Neurology speciality|Title|false|false||Neuronull|Neurologic (qualifier value)|Modifier|false|false||Neuronull|diagnostic service sources radiology labs radiation oncology|Procedure|false|false||radiation oncologynull|Radiation Oncology specialty|Title|false|false||radiation oncologynull|Radiation Ionizing Radiotherapy|Procedure|false|false||radiation
null|Radiotherapy Research|Procedure|false|false||radiation
null|Radiation therapy (procedure)|Procedure|false|false||radiationnull|Electromagnetic Radiation|Phenomenon|false|false||radiation
null|Radiation|Phenomenon|false|false||radiationnull|Unit of radiation dose|LabModifier|false|false||radiationnull|Neoplasms|Disorder|false|false||oncologynull|oncology services|Procedure|false|false||oncologynull|oncology (field)|Title|false|false||oncologynull|Infantile Neuroaxonal Dystrophy|Disorder|false|false||Plannull|Treatment Plan|Finding|false|false||Plan
null|Planned|Finding|false|false||Plan
null|null|Finding|false|false||Plannull|removal technique|Procedure|false|false||surgical resection
null|Excision|Procedure|false|false||surgical resectionnull|Operative Surgical Procedures|Procedure|false|false||surgical
null|Surgical service|Procedure|false|false||surgicalnull|removal technique|Procedure|false|false||resection
null|Excision|Procedure|false|false||resectionnull|Lesion|Finding|false|false||lesion
null|null|Finding|false|false||lesionnull|Aneurysm clip|Device|false|false||aneurysm clipnull|Aneurysm|Finding|false|false||aneurysmnull|CLIP - Codes for radiology reports|Finding|false|false||clip
null|CD74 gene|Finding|false|false||clip
null|CLIP2 gene|Finding|false|false||clip
null|CLIP1 gene|Finding|false|false||clip
null|POMC gene|Finding|false|false||clip
null|POMC wt Allele|Finding|false|false||clip
null|CLIP1 wt Allele|Finding|false|false||clipnull|Comprehensive Lifestyle Intervention Program|Procedure|false|false||clipnull|Clip|Device|false|false||clipnull|CYREN gene|Finding|false|false||MRInull|Magnetic resonance imaging service|Procedure|false|false||MRI
null|Magnetic Resonance Imaging|Procedure|false|false||MRInull|Maori Language|Entity|false|false||MRInull|Consistent with|Finding|false|false||compatiblenull|Compatible|Modifier|false|false||compatiblenull|Able (qualifier value)|Finding|false|false||ablenull|Ability|Subject|false|false||ablenull|Nuclear magnetic resonance imaging brain|Procedure|false|false|C4266577;C0006104|MRI Brainnull|CYREN gene|Finding|false|false|C4266577;C0006104|MRInull|Magnetic resonance imaging service|Procedure|false|false|C4266577;C0006104|MRI
null|Magnetic Resonance Imaging|Procedure|false|false|C4266577;C0006104|MRInull|Maori Language|Entity|false|false||MRInull|Brain Diseases|Disorder|false|false|C4266577;C0006104|Brainnull|Head>Brain|Anatomy|false|false|C4028269;C0006111;C1824234;C1301732;C0032074;C0024485;C0587658;C0543467;C0587668|Brain
null|Brain|Anatomy|false|false|C4028269;C0006111;C1824234;C1301732;C0032074;C0024485;C0587658;C0543467;C0587668|Brainnull|Operative Surgical Procedures|Procedure|false|false|C4266577;C0006104|surgical
null|Surgical service|Procedure|false|false|C4266577;C0006104|surgicalnull|null|Finding|false|false|C4266577;C0006104|planning
null|Planned|Finding|false|false|C4266577;C0006104|planningnull|Evening|Time|false|false||eveningnull|suboccipital craniotomy|Procedure|false|false||suboccipital craniotomynull|Suboccipital approach|Modifier|false|false||suboccipitalnull|Craniotomy|Procedure|false|false||craniotomynull|removal technique|Procedure|false|false||resection
null|Excision|Procedure|false|false||resectionnull|null|Disorder|false|false|C0007765|cerebellar lesionnull|Cerebellum|Anatomy|false|false|C0742035;C1546698;C0221198|cerebellarnull|Lesion|Finding|false|false|C0007765|lesion
null|null|Finding|false|false|C0007765|lesionnull|Neurology speciality|Title|false|false||Neuronull|Neurologic (qualifier value)|Modifier|false|false||Neuronull|Inventory of Callous-Unemotional Traits|Finding|false|false|C0228479|ICUnull|Structure of intraculminate fissure|Anatomy|false|false|C4554035|ICUnull|intensive care unit|Device|false|false||ICUnull|intensive care unit|Entity|false|false||ICUnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Floor (anatomic)|Anatomy|false|false||floornull|floor (object)|Device|false|false||floornull|Floor - story of building|Entity|false|false||floornull|What subject filter - Status|Finding|false|false||statusnull|null|Attribute|false|false||statusnull|Social status|Modifier|false|false||status
null|Status|Modifier|false|false||statusnull|dexamethasone|Drug|false|false||Dexamethasone
null|dexamethasone|Drug|false|false||Dexamethasonenull|Maintenance dose|LabModifier|false|false||maintenance dosenull|Maintenance|Event|false|false||maintenancenull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Course|Time|false|false||coursenull|1 Week|Time|false|false||one weeknull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|Pathology processes|Finding|false|false||pathology
null|Pathological aspects|Finding|false|false||pathologynull|Pathology procedure|Procedure|false|false||pathologynull|Pathology|Title|false|false||pathologynull|Small cell carcinoma of lung|Disorder|false|false|C0007634;C4037972;C0024109|small cell lung carcinomanull|Small|LabModifier|false|false||smallnull|CELP gene|Finding|false|false|C0007634|cell
null|CEL gene|Finding|false|false|C0007634|cellnull|Cells|Anatomy|false|false|C0007097;C0684249;C1413336;C1413337;C0149925;C0740941;C0024115|cellnull|Cell Device|Device|false|false||cell
null|Cellular Phone|Device|false|false||cellnull|Cell (compartment)|Modifier|false|false||cellnull|Carcinoma of lung|Disorder|false|false|C0007634;C4037972;C0024109|lung carcinomanull|Lung diseases|Disorder|false|false|C4037972;C0024109;C0007634|lungnull|Lung Problem|Finding|false|false|C4037972;C0024109;C0007634|lungnull|Chest>Lung|Anatomy|false|false|C0740941;C0684249;C0024115;C0149925|lung
null|Lung|Anatomy|false|false|C0740941;C0684249;C0024115;C0149925|lungnull|Carcinoma|Disorder|false|false|C0007634|carcinomanull|Lung diseases|Disorder|false|false|C4037972;C0024109|Lungnull|Lung Problem|Finding|false|false|C4037972;C0024109|Lungnull|Chest>Lung|Anatomy|false|false|C0221198;C0740941;C0024115|Lung
null|Lung|Anatomy|false|false|C0221198;C0740941;C0024115|Lungnull|Lesion|Finding|false|false|C4037972;C0024109|lesionsnull|Trunk structure|Anatomy|false|false|C0740941;C0034079;C0024115|torsonull|null|Finding|false|false|C4037972;C0024109;C0460005|lung nodulesnull|Lung diseases|Disorder|false|false|C0460005;C4037972;C0024109|lungnull|Lung Problem|Finding|false|false|C0460005;C4037972;C0024109|lungnull|Chest>Lung|Anatomy|false|false|C0034079;C0740941;C0024115|lung
null|Lung|Anatomy|false|false|C0034079;C0740941;C0024115|lungnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Paramedian approach|Modifier|false|false||paramediannull|Aortic arch malformation|Disorder|false|false|C0003483;C0003741;C0230467;C0741204;C0003489;C4037976|aortic archnull|Aortic arch structure|Anatomy|false|false|C4722404;C1538146;C4759703|aortic arch
null|Chest>Aortic arch|Anatomy|false|false|C4722404;C1538146;C4759703|aortic archnull|Aorta|Anatomy|false|false|C4759703|aorticnull|Age-Related Clonal Hematopoiesis|Finding|false|false|C0003741;C0230467;C0741204;C0003489;C4037976|arch
null|ZBTB8OS gene|Finding|false|false|C0003741;C0230467;C0741204;C0003489;C4037976|archnull|Arch of foot|Anatomy|false|false|C4722404;C1538146;C4759703|arch
null|Structure of nucleus infundibularis hypothalami|Anatomy|false|false|C4722404;C1538146;C4759703|arch
null|ARCH|Anatomy|false|false|C4722404;C1538146;C4759703|archnull|Structure of right upper lobe of lung|Anatomy|false|false|C3539671;C1428707;C1552823|right upper lobenull|Table Cell Horizontal Align - right|Finding|false|false|C0225756;C0796494;C1261074|rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Structure of upper lobe of lung|Anatomy|false|false|C1552823;C3539671;C1428707|upper lobenull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|AKT1S1 wt Allele|Finding|false|false|C0796494;C0225756;C1261074|lobe
null|AKT1S1 gene|Finding|false|false|C0796494;C0225756;C1261074|lobenull|lobe|Anatomy|false|false|C3539671;C1428707;C1552823|lobenull|Pulmonary (intended site)|Finding|false|false|C0024109|Pulmonarynull|Lung|Anatomy|false|false|C2707265;C4522268|Pulmonarynull|null|Attribute|false|false|C0024109|Pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||Pulmonarynull|Further|Modifier|false|false||furthernull|Intervention regimes|Procedure|false|false||intervention
null|Nursing interventions|Procedure|false|false||intervention
null|Interventional procedure|Procedure|false|false||interventionnull|Diagnosis Type - Final|Finding|false|false||finalnull|Final|Time|false|false||finalnull|End-stage|Modifier|false|false||finalnull|Pathology processes|Finding|false|false||pathology
null|Pathological aspects|Finding|false|false||pathologynull|Pathology procedure|Procedure|false|false||pathologynull|Pathology|Title|false|false||pathologynull|Heme|Drug|false|false||Heme
null|Heme|Drug|false|false||Hemenull|Assistant Secretary for Technology Policy/Office of the National Coordinator for Health Information Technology|Entity|false|false||Oncnull|Recommendation|Finding|false|false||recommendationsnull|Further|Modifier|false|false||furthernull|Radioisotope scan of lung|Procedure|true|false|C4037972;C0024109|lung imagingnull|Lung diseases|Disorder|false|false|C4037972;C0024109|lungnull|Lung Problem|Finding|false|false|C4037972;C0024109|lungnull|Chest>Lung|Anatomy|false|false|C0203683;C0079595;C0011923;C0740941;C0024115|lung
null|Lung|Anatomy|false|false|C0203683;C0079595;C0011923;C0740941;C0024115|lungnull|Imaging problem|Finding|true|false||imagingnull|Diagnostic Imaging|Procedure|true|false|C4037972;C0024109|imaging
null|Imaging Techniques|Procedure|true|false|C4037972;C0024109|imagingnull|Imaging Technology|Title|false|false||imagingnull|Separate|Modifier|false|false||separatenull|Biopsy of lung|Procedure|false|false|C4037972;C0024109|lung biopsynull|Lung diseases|Disorder|false|false|C4037972;C0024109|lungnull|Lung Problem|Finding|false|false|C4037972;C0024109|lungnull|Chest>Lung|Anatomy|false|false|C0740941;C0189485;C0024115|lung
null|Lung|Anatomy|false|false|C0740941;C0189485;C0024115|lungnull|biopsy characteristics|Finding|false|false||biopsy
null|null|Finding|false|false||biopsynull|Biopsy Procedures on the Pharynx, Adenoids, and Tonsils|Procedure|false|false||biopsy
null|Biopsy|Procedure|false|false||biopsy
null|Consent Type - biopsy|Procedure|false|false||biopsynull|Pulmonary (intended site)|Finding|false|false|C0024109|Pulmonarynull|Lung|Anatomy|false|false|C1533734;C3887704;C0087111;C2707265;C4522268;C0332305|Pulmonarynull|null|Attribute|false|false|C0024109|Pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||Pulmonarynull|Heme|Drug|false|false||Heme
null|Heme|Drug|false|false||Hemenull|Assistant Secretary for Technology Policy/Office of the National Coordinator for Health Information Technology|Entity|false|false||Oncnull|With staging|Finding|false|false|C0024109|stagingnull|Biomaterial Treatment|Finding|false|false||treatment
null|Treating|Finding|false|false||treatment
null|therapeutic aspects|Finding|false|false||treatmentnull|treatment - ActInformationManagementReason|Procedure|false|false|C0024109|treatment
null|Administration (procedure)|Procedure|false|false|C0024109|treatment
null|Therapeutic procedure|Procedure|false|false|C0024109|treatmentnull|Tissue Specimen Code|Finding|false|false|C0040300|tissuenull|Body tissue|Anatomy|false|false|C1547928;C0205469;C0677042|tissuenull|Pathology processes|Finding|false|false|C0040300|pathology
null|Pathological aspects|Finding|false|false|C0040300|pathologynull|Pathology procedure|Procedure|false|false||pathologynull|Pathology|Title|false|false||pathologynull|removal technique|Procedure|false|false||resection
null|Excision|Procedure|false|false||resectionnull|Lesion of brain|Finding|false|false|C4266577;C0006104|brain lesionnull|Brain Diseases|Disorder|false|false|C4266577;C0006104|brainnull|Head>Brain|Anatomy|false|false|C0221505;C0006111;C1546698;C0221198|brain
null|Brain|Anatomy|false|false|C0221505;C0006111;C1546698;C0221198|brainnull|Lesion|Finding|false|false|C4266577;C0006104|lesion
null|null|Finding|false|false|C4266577;C0006104|lesionnull|Diagnosis Type - Final|Finding|false|false||finalnull|Final|Time|false|false||finalnull|End-stage|Modifier|false|false||finalnull|Pathology processes|Finding|false|false||pathology
null|Pathological aspects|Finding|false|false||pathologynull|Pathology procedure|Procedure|false|false||pathologynull|Pathology|Title|false|false||pathologynull|Small|LabModifier|false|false||smallnull|CELP gene|Finding|false|false|C0007634|cell
null|CEL gene|Finding|false|false|C0007634|cellnull|Cells|Anatomy|false|false|C1413336;C1413337|cellnull|Cell Device|Device|false|false||cell
null|Cellular Phone|Device|false|false||cellnull|Cell (compartment)|Modifier|false|false||cellnull|Carcinoma of lung|Disorder|false|false|C4037972;C0024109|lung carcinomanull|Lung diseases|Disorder|false|false|C4037972;C0024109|lungnull|Lung Problem|Finding|false|false|C4037972;C0024109|lungnull|Chest>Lung|Anatomy|false|false|C0740941;C0684249;C0007097;C0024115|lung
null|Lung|Anatomy|false|false|C0740941;C0684249;C0007097;C0024115|lungnull|Carcinoma|Disorder|false|false|C4037972;C0024109|carcinomanull|Dissecting Thoracic Aortic Aneurysm|Disorder|false|false|C0817096|thoracicnull|Chest|Anatomy|false|false|C5779551|thoracicnull|Oncologists|Subject|false|false||oncologistnull|Hyperglycemia steroid-induced|Disorder|false|false||Steroid-induced hyperglycemianull|Steroid [EPC]|Drug|false|false||Steroid
null|Steroids|Drug|false|false||Steroid
null|Steroids|Drug|false|false||Steroidnull|Hyperglycemia|Disorder|false|false||hyperglycemianull|Glucose in blood specimen above reference range|Finding|false|false||hyperglycemianull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Scale, LOINC Axis 5|Finding|false|false|C0222045|scale
null|Base Number|Finding|false|false|C0222045|scale
null|Scale - rank|Finding|false|false|C0222045|scalenull|Integumentary scale|Anatomy|false|false|C1947916;C0005768;C0229664;C0005767;C0851353;C0349674;C2981742;C1522412;C0202098;C1337112;C1533581;C0795635;C4721402;C1579433;C0021641;C3714501;C2239291|scalenull|Weight measurement scales|Device|false|false||scalenull|Scaling|Event|false|false|C0222045|scalenull|insulin, regular, human|Drug|false|false|C0222045|Insulin
null|Insulin [EPC]|Drug|false|false|C0222045|Insulin
null|INS protein, human|Drug|false|false|C0222045|Insulin
null|INS protein, human|Drug|false|false|C0222045|Insulin
null|Insulin|Drug|false|false|C0222045|Insulin
null|Insulin|Drug|false|false|C0222045|Insulin
null|Insulin|Drug|false|false|C0222045|Insulin
null|Therapeutic Insulin|Drug|false|false|C0222045|Insulin
null|Therapeutic Insulin|Drug|false|false|C0222045|Insulin
null|Therapeutic Insulin|Drug|false|false|C0222045|Insulin
null|Insulin Drug Class|Drug|false|false|C0222045|Insulin
null|Insulin Drug Class|Drug|false|false|C0222045|Insulin
null|insulin, regular, human|Drug|false|false|C0222045|Insulin
null|insulin, regular, human|Drug|false|false|C0222045|Insulinnull|INS gene|Finding|false|false|C0222045|Insulinnull|Insulin measurement|Procedure|false|false|C0222045|Insulinnull|Elevated|Modifier|false|false||elevated
null|High|Modifier|false|false||elevatednull|Blood Glucose|Drug|false|false||blood sugarsnull|Blood and lymphatic system disorders|Disorder|false|false|C0222045|bloodnull|peripheral blood|Finding|false|false|C0222045|blood
null|Blood|Finding|false|false|C0222045|blood
null|In Blood|Finding|false|false|C0222045|bloodnull|Sugars|Drug|false|false||sugars
null|Sugars|Drug|false|false||sugarsnull|sugars (lab test)|Procedure|false|false|C0222045|sugarsnull|dexamethasone|Drug|false|false||Dexamethasone
null|dexamethasone|Drug|false|false||Dexamethasonenull|Referral category - Inpatient|Finding|false|false||inpatient
null|Patient Class - Inpatient|Finding|false|false||inpatientnull|inpatient encounter|Procedure|false|false||inpatientnull|inpatient|Subject|false|false||inpatientnull|Team|Subject|false|false||teamnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|insulin, regular, human|Drug|false|false||Insulin
null|Insulin [EPC]|Drug|false|false||Insulin
null|INS protein, human|Drug|false|false||Insulin
null|INS protein, human|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Insulin Drug Class|Drug|false|false||Insulin
null|Insulin Drug Class|Drug|false|false||Insulin
null|insulin, regular, human|Drug|false|false||Insulin
null|insulin, regular, human|Drug|false|false||Insulinnull|INS gene|Finding|false|false||Insulinnull|Insulin measurement|Procedure|false|false||Insulinnull|Blood glucose meters (device)|Device|false|false||glucometernull|Blood Glucose|Drug|false|false||blood sugarsnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Sugars|Drug|false|false||sugars
null|Sugars|Drug|false|false||sugarsnull|sugars (lab test)|Procedure|false|false||sugarsnull|Daily|Time|false|false||dailynull|objective (goal)|Finding|false|false||goal
null|Act Mood - Goal|Finding|false|false||goalnull|Blood Glucose|Drug|false|false||blood sugarnull|Blood glucose measurement|Procedure|false|false||blood sugarnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|raw sugar|Drug|false|false||sugar
null|raw sugar|Drug|false|false||sugar
null|Sugars|Drug|false|false||sugar
null|Sugars|Drug|false|false||sugar
null|Carbohydrates|Drug|false|false||sugarnull|Smaller|Modifier|false|false||lessnull|Less Than|LabModifier|false|false||lessnull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|Bradycardia by ECG Finding|Finding|false|false||Bradycardia
null|Bradycardia|Finding|false|false||Bradycardianull|Transfer - product ownership|Finding|false|false||transfer
null|Transfer Technique|Finding|false|false||transfer
null|ActClass - transfer|Finding|false|false||transfer
null|null|Finding|false|false||transfernull|Transfer (immobility management)|Procedure|false|false||transfernull|TCF21 wt Allele|Finding|false|false||POD1
null|CORO7 gene|Finding|false|false||POD1
null|TCF21 gene|Finding|false|false||POD1null|Inventory of Callous-Unemotional Traits|Finding|false|false|C0228479|ICUnull|Structure of intraculminate fissure|Anatomy|false|false|C4554035;C0741624|ICUnull|intensive care unit|Device|false|false||ICUnull|intensive care unit|Entity|false|false||ICUnull|Asymptomatic bradycardia|Disorder|false|false|C0228479|asymptomatic bradycardianull|Asymptomatic diagnosis of|Finding|false|false||asymptomatic
null|Asymptomatic (finding)|Finding|false|false||asymptomaticnull|Bradycardia by ECG Finding|Finding|false|false||bradycardia
null|Bradycardia|Finding|false|false||bradycardianull|Asymptomatic diagnosis of|Finding|false|false||asymptomatic
null|Asymptomatic (finding)|Finding|false|false||asymptomaticnull|Liquid substance|Drug|false|false||fluidsnull|Mouse Body Fluid or Substance|Finding|false|false||fluidsnull|Fluid Therapy|Procedure|false|false||fluidsnull|Administration (procedure)|Procedure|false|false||administrationnull|Administration occupational activities|Event|false|false||administrationnull|Synthetic Levothyroxine|Drug|false|false||levothyroxine
null|Synthetic Levothyroxine|Drug|false|false||levothyroxine
null|levothyroxine|Drug|false|false||levothyroxine
null|levothyroxine|Drug|false|false||levothyroxine
null|levothyroxine|Drug|false|false||levothyroxinenull|Asymptomatic diagnosis of|Finding|false|false||asymptomatic
null|Asymptomatic (finding)|Finding|false|false||asymptomaticnull|Bell Palsy|Disorder|false|false||Bell's palsy
null|Facial paralysis|Disorder|false|false||Bell's palsynull|Bell Device|Device|false|false||Bellnull|Palsy|Finding|false|false||palsy
null|Paralysed|Finding|false|false||palsynull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|valacyclovir|Drug|false|false||Valacyclovir
null|valacyclovir|Drug|false|false||Valacyclovirnull|Glucose tolerance test|Procedure|false|false||gttsnull|Drop Dosing Unit|LabModifier|false|false||gttsnull|Urgency of micturition|Finding|false|false|C0042027|Urinary urgencynull|Urinary tract|Anatomy|false|false|C0085606|Urinarynull|urinary|Modifier|false|false||Urinarynull|Urgent|Modifier|false|false||urgencynull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Urgency of micturition|Finding|false|false|C0042027|urinary urgencynull|Urinary tract|Anatomy|false|false|C0085606|urinarynull|urinary|Modifier|false|false||urinarynull|Urgent|Modifier|false|false||urgencynull|Frequency|Finding|false|false||frequency
null|How Often|Finding|false|false||frequencynull|With frequency|Time|false|false||frequency
null|Frequencies (time pattern)|Time|false|false||frequencynull|Kind of quantity - Frequency|LabModifier|false|false||frequency
null|Statistical Frequency|LabModifier|false|false||frequency
null|Spatial Frequency|LabModifier|false|false||frequencynull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Culture Dose Form|Drug|false|false||culturenull|Culture (Anthropological)|Finding|false|false||culture
null|Cultural aspects|Finding|false|false||culturenull|Microbial culture (procedure)|Procedure|false|false||culture
null|Laboratory culture|Procedure|false|false||culturenull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Clinical Service|Procedure|false|false||servicesnull|Services|Event|false|false||servicesnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Disease|Disorder|false|false||conditionnull|Logical Condition|Finding|false|false||conditionnull|null|Attribute|false|false||conditionnull|Condition|Modifier|false|false||conditionnull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|Arylsulfatase A, human|Drug|false|false||ASA
null|Arylsulfatase A, human|Drug|false|false||ASA
null|aspirin|Drug|false|false||ASA
null|aspirin|Drug|false|false||ASAnull|ARSA gene|Finding|false|false||ASAnull|alendronate|Drug|false|false||Alendronate
null|alendronate|Drug|false|false||Alendronatenull|Weekly|Time|false|false||weeklynull|vitamin D3|Drug|false|false||Vitamin D3
null|vitamin D3|Drug|false|false||Vitamin D3
null|cholecalciferol|Drug|false|false||Vitamin D3
null|cholecalciferol|Drug|false|false||Vitamin D3
null|cholecalciferol|Drug|false|false||Vitamin D3null|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitaminnull|Unit - NCI Thesaurus Property|LabModifier|false|false||units
null|Unit of Measure|LabModifier|false|false||units
null|Unit|LabModifier|false|false||unitsnull|Daily|Time|false|false||dailynull|Synthetic Levothyroxine|Drug|false|false||Levothyroxine
null|Synthetic Levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxinenull|Daily|Time|false|false||dailynull|lisinopril|Drug|false|false||Lisinopril
null|lisinopril|Drug|false|false||Lisinoprilnull|Daily|Time|false|false||dailynull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Mild Severity of Illness Code|Finding|false|false||Mildnull|Mild (qualifier value)|Modifier|false|false||Mild
null|Mild Allergy Severity|Modifier|false|false||Mildnull|Fever symptoms (finding)|Finding|false|false||Fever
null|Fever|Finding|false|false||Fevernull|bisacodyl|Drug|false|false||Bisacodyl
null|bisacodyl|Drug|false|false||Bisacodylnull|Daily|Time|false|false||DAILYnull|dexamethasone|Drug|false|false||Dexamethasone
null|dexamethasone|Drug|false|false||Dexamethasonenull|Every eight hours|Time|false|false||Q8Hnull|Duration brand of oxymetazoline|Drug|false|false||Durationnull|Duration (temporal concept)|Time|false|false||Durationnull|Dosage|LabModifier|false|false||Dosesnull|Maintenance dose|LabModifier|false|false||maintenance dosenull|Maintenance|Event|false|false||maintenancenull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|null|Attribute|false|false||dose #null|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Dosage|LabModifier|false|false||dosesnull|dexamethasone|Drug|false|false||dexamethasone
null|dexamethasone|Drug|false|false||dexamethasonenull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false|C0230028;C0226896|by mouthnull|Oral cavity|Anatomy|false|false|C1527415|mouth
null|Oral region|Anatomy|false|false|C1527415|mouthnull|Hour|Time|false|false||hoursnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|docusate sodium|Drug|false|false||Docusate Sodium
null|docusate sodium|Drug|false|false||Docusate Sodiumnull|docusate|Drug|false|false||Docusate
null|docusate|Drug|false|false||Docusatenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|famotidine|Drug|false|false||Famotidine
null|famotidine|Drug|false|false||Famotidinenull|Every twenty four hours|Time|false|false||Q24Hnull|famotidine|Drug|false|false||famotidine
null|famotidine|Drug|false|false||famotidinenull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false|C0230028;C0226896|by mouthnull|Oral cavity|Anatomy|false|false|C1527415;C1561538;C1561539|mouth
null|Oral region|Anatomy|false|false|C1527415;C1561538;C1561539|mouthnull|Twice a day|Time|false|false||twice a daynull|Transaction counts and value totals - day|Finding|false|false|C0230028;C0226896|day
null|Precision - day|Finding|false|false|C0230028;C0226896|daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|polyethylene glycols|Drug|false|false||Polyethylene Glycol
null|polyethylene glycols|Drug|false|false||Polyethylene Glycolnull|high-density polyethylene|Drug|false|false||Polyethylene
null|high-density polyethylene|Drug|false|false||Polyethylene
null|polyethylenes|Drug|false|false||Polyethylene
null|polyethylenes|Drug|false|false||Polyethylene
null|Polyethylene|Drug|false|false||Polyethylene
null|Polyethylene|Drug|false|false||Polyethylenenull|ethylene glycol|Drug|false|false||Glycol
null|Glycol|Drug|false|false||Glycol
null|ethylene glycol|Drug|false|false||Glycol
null|Glycols|Drug|false|false||Glycolnull|Daily|Time|false|false||DAILYnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Constipation|Finding|false|false||Constipationnull|Firstly|Modifier|false|false||Firstnull|First (number)|LabModifier|false|false||Firstnull|Line Specimen|Drug|false|false||Line
null|Long Interspersed Elements|Drug|false|false||Line
null|Long Interspersed Elements|Drug|false|false||Linenull|line source specimen code|Finding|false|false||Linenull|Intravascular line|Device|false|false||Linenull|Linear|Modifier|false|false||Linenull|Line Unit of Length|LabModifier|false|false||Linenull|sennosides, USP|Drug|false|false||Senna
null|sennosides, USP|Drug|false|false||Sennanull|Senna alexandrina|Entity|false|false||Senna
null|Senna Plant|Entity|false|false||Sennanull|levothyroxine sodium|Drug|false|false||Levothyroxine Sodium
null|levothyroxine sodium|Drug|false|false||Levothyroxine Sodium
null|levothyroxine sodium|Drug|false|false||Levothyroxine Sodiumnull|Synthetic Levothyroxine|Drug|false|false||Levothyroxine
null|Synthetic Levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxinenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|microgram|LabModifier|false|false||mcgnull|Daily|Time|false|false||DAILYnull|lisinopril|Drug|false|false||Lisinopril
null|lisinopril|Drug|false|false||Lisinoprilnull|Daily|Time|false|false||DAILYnull|prednisolone acetate|Drug|false|false||PrednisoLONE Acetate
null|prednisolone acetate|Drug|false|false||PrednisoLONE Acetatenull|prednisolone|Drug|false|false||PrednisoLONE
null|prednisolone|Drug|false|false||PrednisoLONEnull|acetate|Drug|false|false||Acetate
null|acetate|Drug|false|false||Acetatenull|Ophthalmic Route of Administration|Finding|false|false||Ophthnull|Drops - Drug Form|Drug|false|false|C0229090|DROPnull|Dropping|Event|false|false|C0229090|DROPnull|Drop (unit of presentation)|LabModifier|false|false||DROP
null|Drop British|LabModifier|false|false||DROP
null|Drop Dosing Unit|LabModifier|false|false||DROP
null|Medical Drop|LabModifier|false|false||DROP
null|Drop Unit of Volume|LabModifier|false|false||DROPnull|examination of left eye|Procedure|false|false|C4266572;C0015392;C0700042;C0229090|LEFT EYEnull|Left eye structure|Anatomy|false|false|C0154094;C0015397;C0991568;C1705648;C1552822;C2141124;C1550636;C1546630;C0262477|LEFT EYEnull|Table Cell Horizontal Align - left|Finding|false|false|C0229090;C4266572;C0015392;C0700042|LEFTnull|Left sided|Modifier|false|false||LEFT
null|Left|Modifier|false|false||LEFTnull|Carcinoma in situ of eye|Disorder|false|false|C0229090;C4266572;C0015392;C0700042|EYE
null|Disorder of eye|Disorder|false|false|C0229090;C4266572;C0015392;C0700042|EYEnull|Eye - Specimen Source Code|Finding|false|false|C4266572;C0015392;C0700042;C0229090|EYE
null|Eye problem|Finding|false|false|C4266572;C0015392;C0700042;C0229090|EYE
null|Eye Specimen|Finding|false|false|C4266572;C0015392;C0700042;C0229090|EYEnull|Head>Eye|Anatomy|false|false|C2141124;C1550636;C1546630;C0262477;C0154094;C0015397;C1552822|EYE
null|Eye|Anatomy|false|false|C2141124;C1550636;C1546630;C0262477;C0154094;C0015397;C1552822|EYE
null|Orbital region|Anatomy|false|false|C2141124;C1550636;C1546630;C0262477;C0154094;C0015397;C1552822|EYEnull|Four times daily|Time|false|false||QIDnull|valacyclovir|Drug|false|false||ValACYclovir
null|valacyclovir|Drug|false|false||ValACYclovirnull|Every eight hours|Time|false|false||Q8Hnull|Vitamin D Drug Class|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|D Vitamin|Drug|false|false||Vitamin D
null|Vitamin D [EPC]|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|Vitamin D Drug Class|Drug|false|false||Vitamin Dnull|Vitamin D measurement|Procedure|false|false||Vitamin Dnull|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitaminnull|Storage Unit|Device|false|false||UNIT
null|Unit device|Device|false|false||UNITnull|Unit - NCI Thesaurus Property|LabModifier|false|false||UNIT
null|Unit of Measure|LabModifier|false|false||UNIT
null|Unit|LabModifier|false|false||UNIT
null|Enzyme Unit|LabModifier|false|false||UNITnull|Daily|Time|false|false||DAILYnull|ARID1A protein, human|Drug|false|false||HELD
null|ARID1A protein, human|Drug|false|false||HELDnull|Held - activity status|Finding|false|false||HELD
null|ARID1A wt Allele|Finding|false|false||HELDnull|alendronate sodium|Drug|false|false||Alendronate Sodium
null|alendronate sodium|Drug|false|false||Alendronate Sodiumnull|alendronate|Drug|false|false||Alendronate
null|alendronate|Drug|false|false||Alendronatenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|Weekly|Time|false|false||/WEEKnull|Transaction counts and value totals - week|Finding|false|false||WEEKnull|week|Time|false|false||WEEKnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|alendronate sodium|Drug|false|false||Alendronate Sodium
null|alendronate sodium|Drug|false|false||Alendronate Sodiumnull|alendronate|Drug|false|false||Alendronate
null|alendronate|Drug|false|false||Alendronatenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|ARID1A protein, human|Drug|false|false||HELD
null|ARID1A protein, human|Drug|false|false||HELDnull|Held - activity status|Finding|false|false||HELD
null|ARID1A wt Allele|Finding|false|false||HELDnull|aspirin|Drug|false|false||Aspirin
null|aspirin|Drug|false|false||Aspirinnull|Daily|Time|false|false||DAILYnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|aspirin|Drug|false|false||Aspirin
null|aspirin|Drug|false|false||Aspirinnull|Blood glucose meters (device)|Device|false|false||glucometernull|Blood glucose meters (device)|Device|false|false||glucometernull|Blood Glucose|Drug|false|false||blood sugarsnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Sugars|Drug|false|false||sugars
null|Sugars|Drug|false|false||sugarsnull|sugars (lab test)|Procedure|false|false||sugarsnull|Hour|Time|false|false||hoursnull|Meal (occasion for eating)|Finding|false|false||mealnull|Records|Finding|false|false||Recordnull|Record - QueryRequestLimit|LabModifier|false|false||Recordnull|Numbers|LabModifier|false|false||numbers
null|Count of entities|LabModifier|false|false||numbersnull|Oncologists|Subject|false|false||Oncologistnull|Test Strip Device|Device|false|false||test stripsnull|Tests (qualifier value)|Finding|false|false|C4318744|test
null|Testing|Finding|false|false|C4318744|testnull|Laboratory Procedures|Procedure|false|false|C4318744|testnull|Test - temporal region|Anatomy|false|false|C0456984;C0039593;C0392366;C0022885|testnull|Test Result|Lab|false|false|C4318744|testnull|Test Dosing Unit|LabModifier|false|false||testnull|strip medical device|Device|false|false||stripsnull|Blood Glucose|Drug|false|false||blood sugarsnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Sugars|Drug|false|false||sugars
null|Sugars|Drug|false|false||sugarsnull|sugars (lab test)|Procedure|false|false||sugarsnull|refill|Finding|false|false||refillsnull|Lancet|Device|false|false||Lancetsnull|Blood Glucose|Drug|false|false||blood sugarsnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Sugars|Drug|false|false||sugars
null|Sugars|Drug|false|false||sugarsnull|sugars (lab test)|Procedure|false|false||sugarsnull|refill|Finding|false|false||refillsnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|ADMIN.FACILITY|Finding|false|false||Facilitynull|Facility (object)|Device|false|false||Facilitynull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Brain Neoplasms|Disorder|false|false|C4266577;C0006104|Brain tumornull|Brain Diseases|Disorder|false|false|C4266577;C0006104|Brainnull|Head>Brain|Anatomy|false|false|C0006118;C0006111;C3273930;C1578706;C0027651|Brain
null|Brain|Anatomy|false|false|C0006118;C0006111;C3273930;C1578706;C0027651|Brainnull|Neoplasms|Disorder|false|false|C4266577;C0006104|tumornull|Tumor Mass|Finding|false|false|C4266577;C0006104|tumor
null|null|Finding|false|false|C4266577;C0006104|tumornull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Disease|Disorder|false|false||Conditionnull|Logical Condition|Finding|false|false||Conditionnull|null|Attribute|false|false||Conditionnull|Condition|Modifier|false|false||Conditionnull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Helping Behavior|Finding|false|false||assistancenull|Assisted (qualifier value)|Modifier|false|false||assistancenull|AICDA protein, human|Drug|false|false||aid
null|AICDA protein, human|Drug|false|false||aidnull|AICDA wt Allele|Finding|false|false||aid
null|AICDA gene|Finding|false|false||aidnull|AID - Artificial insemination by donor|Procedure|false|false||aid
null|dacarbazine/doxorubicin/ifosfamide protocol|Procedure|false|false||aidnull|Aid (attribute)|Modifier|false|false||aid
null|Assisted (qualifier value)|Modifier|false|false||aidnull|Discharge instructions|Finding|false|false||Discharge Instructionsnull|hospital discharge instructions (treatment)|Procedure|false|false||Discharge Instructionsnull|null|Attribute|false|false||Discharge Instructionsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructionsnull|Level of Care - Surgery|Finding|false|false||Surgery
null|Surgical procedure finding|Finding|false|false||Surgery
null|Surgical aspects|Finding|false|false||Surgerynull|Operative Surgical Procedures|Procedure|false|false||Surgerynull|General surgery specialty|Title|false|false||Surgery
null|Surgery specialty|Title|false|false||Surgerynull|Level of Care - Surgery|Finding|false|false|C4266577;C0006104|surgery
null|Surgical procedure finding|Finding|false|false|C4266577;C0006104|surgery
null|Surgical aspects|Finding|false|false|C4266577;C0006104|surgerynull|Operative Surgical Procedures|Procedure|false|false|C4266577;C0006104|surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Lesion of brain|Finding|false|false|C4266577;C0006104|brain lesionnull|Brain Diseases|Disorder|false|false|C4266577;C0006104|brainnull|Head>Brain|Anatomy|false|false|C1546698;C0221198;C0038895;C1457907;C1547138;C0543467;C0006111;C0221505|brain
null|Brain|Anatomy|false|false|C1546698;C0221198;C0038895;C1457907;C1547138;C0543467;C0006111;C0221505|brainnull|Lesion|Finding|false|false|C4266577;C0006104|lesion
null|null|Finding|false|false|C4266577;C0006104|lesionnull|Brain Diseases|Disorder|false|false|C4266577;C0006104|brainnull|Head>Brain|Anatomy|false|false|C0006111|brain
null|Brain|Anatomy|false|false|C0006111|brainnull|Specimen|Drug|false|false||samplenull|Nucleotide Sequence Sample Name|Finding|false|false|C4266577;C0006104;C0040300|sample
null|Biospecimen|Finding|false|false|C4266577;C0006104;C0040300|samplenull|Tissue Specimen Code|Finding|false|false|C4266577;C0006104;C0040300|tissuenull|Body tissue|Anatomy|false|false|C0006111;C1547928;C1546698;C0221198;C5551027;C2347026|tissuenull|Lesion|Finding|false|false|C4266577;C0006104;C0040300|lesion
null|null|Finding|false|false|C4266577;C0006104;C0040300|lesionnull|Brain Diseases|Disorder|false|false|C0040300;C4266577;C0006104|brainnull|Head>Brain|Anatomy|false|false|C5551027;C2347026;C1546698;C0221198;C1547928;C0006111|brain
null|Brain|Anatomy|false|false|C5551027;C2347026;C1546698;C0221198;C1547928;C0006111|brainnull|Pathology processes|Finding|false|false||pathology
null|Pathological aspects|Finding|false|false||pathologynull|Pathology procedure|Procedure|false|false||pathologynull|Pathology|Title|false|false||pathologynull|Testing|Finding|false|false||testing
null|Tests (qualifier value)|Finding|false|false||testingnull|Surgical wound|Disorder|false|false|C2338258|incisionnull|Surgical incisions|Procedure|false|false|C2338258|incisionnull|Cranial incision point|Anatomy|false|false|C0184898;C0332803|incisionnull|Suture Joint|Anatomy|false|false||suturesnull|Surgical sutures|Device|false|false||suturesnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Surgical wound|Disorder|false|false|C2338258|incisionnull|Surgical incisions|Procedure|false|false|C2338258|incisionnull|Cranial incision point|Anatomy|false|false|C0184898;C0332803|incisionnull|Vitelliform Macular Dystrophy|Disorder|false|false|C2338258|bestnull|BEST1 wt Allele|Finding|false|false||best
null|BEST1 gene|Finding|false|false||bestnull|best (quality)|Modifier|false|false||bestnull|Surgical wound|Disorder|false|false|C2338258|incisionnull|Surgical incisions|Procedure|false|false|C2338258|incisionnull|Cranial incision point|Anatomy|false|false|C0339510;C0332803;C0184898|incisionnull|Open|Modifier|false|false||opennull|Air (substance)|Drug|false|false||air
null|air|Drug|false|false||air
null|air|Drug|false|false||airnull|ACUTE INSULIN RESPONSE|Finding|false|false||air
null|AIRN gene|Finding|false|false||air
null|AI/RHEUM|Finding|false|false||airnull|Call - dosing instruction fragment|Finding|false|false||Call
null|Call (Instruction)|Finding|false|false||Call
null|Decision|Finding|false|false||Call
null|CHL1 gene|Finding|false|false||Callnull|null|Attribute|false|false||surgeonnull|Surgeon|Subject|false|false||surgeonnull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|Erythema|Disorder|false|false||rednessnull|Redness|Finding|false|false||rednessnull|Red color|Modifier|false|false||rednessnull|Fever symptoms (finding)|Finding|false|false||fever
null|Fever|Finding|false|false||fevernull|Body Substance Discharge|Finding|false|false||drainage
null|Body Fluid Discharge|Finding|false|false||drainagenull|Drainage procedure|Procedure|false|false||drainagenull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|Heavy (weight) (qualifier value)|Modifier|false|false||heavy
null|Heavy (amount)|Modifier|false|false||heavynull|Lifting|Event|false|false||liftingnull|Go Jogging or Running Question|Finding|false|false||running
null|Running (physical activity)|Finding|false|false||running
null|running (history)|Finding|false|false||runningnull|climbing (history)|Finding|false|false||climbing
null|Climbing|Finding|false|false||climbing
null|Does climb|Finding|false|false||climbingnull|Strenuous Exercise|Finding|false|false||strenuous exercisenull|Strenuous|Modifier|false|false||strenuousnull|Exercise|Finding|false|false||exercisenull|Exercise Pain Management|Procedure|false|false||exercisenull|Follow-up status|Finding|false|false||follow-upnull|follow-up|Procedure|false|false||follow-upnull|Follow - dosing instruction imperative|Finding|false|false||follow
null|Follow|Finding|false|false||follownull|Followed by|Time|false|false||follownull|Appointments|Event|false|false||appointmentnull|Does walk|Finding|false|false||walksnull|Slow|Modifier|false|false||slowlynull|Activity (animal life circumstance)|Finding|false|false||activity
null|Physical activity|Finding|false|false||activitynull|Activities|Event|false|false||activitynull|null|Modifier|false|false||activitynull|Own|Finding|false|false||ownnull|cyclophosphamide/doxorubicin/etoposide/prednisone|Drug|false|false||pace
null|cisplatin/cyclophosphamide/doxorubicin/etoposide|Drug|false|false||pace
null|FURIN protein, human|Drug|false|false||pace
null|FURIN protein, human|Drug|false|false||pacenull|furin activity|Finding|false|false||pace
null|FURIN gene|Finding|false|false||pace
null|Patient Assessment of Cancer Communication Experiences|Finding|false|false||pacenull|cisplatin/cyclophosphamide/doxorubicin/vindesine protocol|Procedure|false|false||pacenull|Program of All-Inclusive Care for the Elderly (PACE)|Subject|false|false||pacenull|Pace Unit of Measure|LabModifier|false|false||pacenull|Symptoms|Finding|false|false||symptomnull|null|Attribute|false|false||symptomnull|Free of (attribute)|Finding|false|false||freenull|Empty (qualifier)|Modifier|false|false||freenull|At rest (qualifier value)|Finding|false|false||at restnull|REST protein, human|Drug|false|false||rest
null|REST protein, human|Drug|false|false||restnull|site-specific telomere resolvase activity|Finding|false|false||rest
null|Rest|Finding|false|false||rest
null|REST gene|Finding|false|false||restnull|Too much|Finding|false|false||too muchnull|Much|Finding|false|false||muchnull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Automobile Driving|Finding|false|false||drivingnull|Narcotics|Drug|true|false||narcotic
null|Narcotics|Drug|true|false||narcoticnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Seizures|Finding|false|false||seizurenull|Law (document)|Finding|false|false||lawnull|Law Profession|Subject|false|false||lawnull|Rules of conduct|Entity|false|false||law
null|aspects of laws|Entity|false|false||law
null|Legal system|Entity|false|false||lawnull|Law (view)|Modifier|false|false||lawnull|Contact - HL7 Attribution|Finding|false|false||contact
null|Contact with|Finding|false|false||contact
null|Communication Contact|Finding|false|false||contactnull|contact person|Subject|false|false||contactnull|Physical contact|Phenomenon|false|false||contactnull|Personal Contact|Event|false|false||contactnull|Sports|Finding|false|false||sportsnull|Neurosurgeon|Subject|false|false||neurosurgeonnull|Contact - HL7 Attribution|Finding|false|false||contact
null|Contact with|Finding|false|false||contact
null|Communication Contact|Finding|false|false||contactnull|contact person|Subject|false|false||contactnull|Physical contact|Phenomenon|false|false||contactnull|Personal Contact|Event|false|false||contactnull|Sports|Finding|false|false||sportsnull|6 months|Time|false|false||6 monthsnull|month|Time|false|false||monthsnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Thinning Weight Loss|Finding|false|false||thinningnull|Decreased thickness|Modifier|false|false||thinningnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|aspirin|Drug|false|false||Aspirin
null|aspirin|Drug|false|false||Aspirinnull|ibuprofen|Drug|false|false||Ibuprofen
null|ibuprofen|Drug|false|false||Ibuprofennull|Plavix|Drug|false|false||Plavix
null|Plavix|Drug|false|false||Plavixnull|Coumadin|Drug|false|false||Coumadin
null|Coumadin|Drug|false|false||Coumadinnull|Neurosurgeon|Subject|false|false||neurosurgeonnull|aspirin|Drug|false|false||Aspirin
null|aspirin|Drug|false|false||Aspirinnull|Daily|Time|false|false||dailynull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|alendronate|Drug|false|false||Alendronate
null|alendronate|Drug|false|false||Alendronatenull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Tylenol|Drug|false|false||Tylenol
null|Tylenol|Drug|false|false||Tylenolnull|minor (disease)|Disorder|false|false||minornull|NR4A3 wt Allele|Finding|false|false||minor
null|NR4A3 gene|Finding|false|false||minornull|Minor (person)|Subject|false|false||minornull|Minor (value)|Modifier|false|false||minornull|Discomfort|Finding|false|false||discomfortnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|dexamethasone|Drug|false|false||Dexamethasone
null|dexamethasone|Drug|false|false||Dexamethasonenull|Steroid [EPC]|Drug|false|false||steroid
null|Steroids|Drug|false|false||steroid
null|Steroids|Drug|false|false||steroidnull|Treats (attribute)|Finding|false|false||treats
null|Intent To Treat|Finding|false|false||treatsnull|Brain Edema|Finding|false|false|C0524466|intracranial swellingnull|Intracranial Route of Administration|Finding|false|false|C0524466|intracranialnull|Intracranial|Anatomy|false|false|C0013604;C0038999;C1527311;C1522213|intracranialnull|Swelling|Finding|false|false|C0524466|swelling
null|Edema|Finding|false|false|C0524466|swellingnull|dexamethasone|Drug|false|false||Dexamethasone
null|dexamethasone|Drug|false|false||Dexamethasonenull|Maintenance dose|LabModifier|false|false||maintenance dosenull|Maintenance|Event|false|false||maintenancenull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Hyperglycemia|Disorder|false|false||elevated blood glucosenull|elevated random blood glucose level|Finding|false|false||elevated blood glucose
null|Blood glucose increased|Finding|false|false||elevated blood glucosenull|Elevated|Modifier|false|false||elevated
null|High|Modifier|false|false||elevatednull|Finding of blood glucose level|Lab|false|false||blood glucose levelsnull|Blood Glucose|Drug|false|false||blood glucosenull|Blood glucose measurement|Procedure|false|false||blood glucosenull|Finding of blood glucose level|Lab|false|false||blood glucosenull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|null|Lab|false|false||glucose levelsnull|glucose|Drug|false|false||glucose
null|glucose|Drug|false|false||glucose
null|glucose|Drug|false|false||glucosenull|Glucose measurement|Procedure|false|false||glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||glucosenull|Levels (qualifier value)|Modifier|false|false||levelsnull|insulin, regular, human|Drug|false|false||Insulin
null|Insulin [EPC]|Drug|false|false||Insulin
null|INS protein, human|Drug|false|false||Insulin
null|INS protein, human|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Insulin Drug Class|Drug|false|false||Insulin
null|Insulin Drug Class|Drug|false|false||Insulin
null|insulin, regular, human|Drug|false|false||Insulin
null|insulin, regular, human|Drug|false|false||Insulinnull|INS gene|Finding|false|false||Insulinnull|Insulin measurement|Procedure|false|false||Insulinnull|Check|Finding|false|false||checknull|null|Event|false|false||checknull|Blood Glucose|Drug|false|false||blood sugarsnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Sugars|Drug|false|false||sugars
null|Sugars|Drug|false|false||sugarsnull|sugars (lab test)|Procedure|false|false||sugarsnull|Daily|Time|false|false||dailynull|At home|Finding|false|false||at homenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Blood glucose meters (device)|Device|false|false||glucometernull|Nurses|Subject|false|false||nursenull|Participation Type - device|Finding|false|false||devicenull|Medical Devices|Device|false|false||device
null|Devices|Device|false|false||devicenull|Kind of quantity - Device|LabModifier|false|false||devicenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Blood Glucose|Drug|false|false||blood sugarsnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Sugars|Drug|false|false||sugars
null|Sugars|Drug|false|false||sugarsnull|sugars (lab test)|Procedure|false|false||sugarsnull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|objective (goal)|Finding|false|false||goal
null|Act Mood - Goal|Finding|false|false||goalnull|Blood Glucose|Drug|false|false||blood sugarnull|Blood glucose measurement|Procedure|false|false||blood sugarnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|raw sugar|Drug|false|false||sugar
null|raw sugar|Drug|false|false||sugar
null|Sugars|Drug|false|false||sugar
null|Sugars|Drug|false|false||sugar
null|Carbohydrates|Drug|false|false||sugarnull|Less Than|LabModifier|false|false||less thannull|Smaller|Modifier|false|false||lessnull|Less Than|LabModifier|false|false||lessnull|Experience (Practice)|Finding|false|false||Experience
null|Experience|Finding|false|false||Experiencenull|Headache|Finding|false|false||headachesnull|Incisional pain|Finding|false|false||incisional painnull|Surgical incisions|Procedure|false|false||incisionalnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Postoperative Period|Time|false|false||post-operativenull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|FANCONI ANEMIA, COMPLEMENTATION GROUP E|Disorder|false|false|C0015450;C4266571;C0015392|facenull|FANCE wt Allele|Finding|false|false|C0015450;C4266571;C0015392|face
null|FANCE gene|Finding|false|false|C0015450;C4266571;C0015392|face
null|ELOVL6 gene|Finding|false|false|C0015450;C4266571;C0015392|facenull|Head>Face|Anatomy|false|false|C1423759;C2828055;C1414531;C5848506;C3160739|face
null|Face|Anatomy|false|false|C1423759;C2828055;C1414531;C5848506;C3160739|facenull|Face (spatial concept)|Modifier|false|false||facenull|Eye|Anatomy|false|false|C1423759;C2828055;C1414531;C5848506;C3160739|eyesnull|null|Attribute|false|false|C0015450;C4266571;C0015392|eyesnull|post operative (finding)|Finding|false|false||after surgerynull|Postoperative Period|Time|false|false||after surgerynull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Precision - second|Finding|false|false||second
null|metastatic qualifier|Finding|false|false||second
null|Second Suffix|Finding|false|false||secondnull|seconds|Time|false|false||secondnull|Second Unit of Plane Angle|LabModifier|false|false||second
null|second (number)|LabModifier|false|false||secondnull|III (suffix)|Modifier|false|false||thirdnull|Third|LabModifier|false|false||thirdnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Apply (administration method)|Finding|false|false||apply
null|Apply (instruction)|Finding|false|false||apply
null|null|Finding|false|false||apply
null|Apply|Finding|false|false||applynull|Ice Pharmaceutical|Drug|false|false|C3496566;C0228434|ice
null|Ice Pharmaceutical|Drug|false|false|C3496566;C0228434|ice
null|Ice|Drug|false|false|C3496566;C0228434|ice
null|methamphetamine|Drug|false|false|C3496566;C0228434|ice
null|methamphetamine|Drug|false|false|C3496566;C0228434|ice
null|methamphetamine|Drug|false|false|C3496566;C0228434|ice
null|Caspase-1, human|Drug|false|false|C3496566;C0228434|ice
null|Caspase-1, human|Drug|false|false|C3496566;C0228434|icenull|caspase-1 activity|Finding|false|false|C3496566;C0228434|ice
null|CASP1 wt Allele|Finding|false|false|C3496566;C0228434|ice
null|CES2 gene|Finding|false|false|C3496566;C0228434|ice
null|CES2 wt Allele|Finding|false|false|C3496566;C0228434|ice
null|CASP1 gene|Finding|false|false|C3496566;C0228434|icenull|cryotherapy using ice|Procedure|false|false|C3496566;C0228434|ice
null|cytarabine/etoposide/idarubicin|Procedure|false|false|C3496566;C0228434|ice
null|AIE Regimen|Procedure|false|false|C3496566;C0228434|ice
null|carboplatin/etoposide/ifosfamide|Procedure|false|false|C3496566;C0228434|icenull|Structure of inferior central nucleus of pons|Anatomy|false|false|C0020746;C1873773;C4721557;C0025611;C0582051;C1705786;C3889432;C1366479;C1150137;C1413348;C0678568;C0249492;C1879508;C0280697;C0556917|ice
null|intracentral fissure|Anatomy|false|false|C0020746;C1873773;C4721557;C0025611;C0582051;C1705786;C3889432;C1366479;C1150137;C1413348;C0678568;C0249492;C1879508;C0280697;C0556917|icenull|null|Phenomenon|false|false|C3496566;C0228434|coolnull|Specimen Condition - Cool|Modifier|false|false||coolnull|Feels warm|Finding|false|false|C3496566;C0228434|warmnull|warming process|Phenomenon|false|false||warmnull|Eye|Anatomy|false|false|C5848506|eyesnull|null|Attribute|false|false|C0015392|eyesnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|Observation Interpretation - worse|Finding|false|false||worse
null|Worse|Finding|false|false||worsenull|Worsening (qualifier value)|Modifier|false|false||worsenull|Morning|Time|false|false||in the morningnull|Morning After|Drug|false|false||morning after
null|Morning After|Drug|false|false||morning afternull|Morning After Time Pattern|Time|false|false||morning afternull|Morning|Time|false|false||morningnull|Residential flat|Device|false|false||flatnull|Flat shape|Modifier|false|false||flatnull|Sore to touch|Finding|false|false||sorenessnull|outcomes otolaryngology chewing|Finding|false|false||chewing
null|Chewing|Finding|false|false||chewingnull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|With time|Time|false|false||with timenull|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Food|Drug|false|false||foodsnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|More|LabModifier|false|false||morenull|Feeling tired|Finding|false|false||tired
null|Feel Tired question|Finding|false|false||tired
null|Fatigue|Finding|false|false||tirednull|Restlessness|Finding|false|false||restlessness
null|Psychomotor Agitation|Finding|false|false||restlessness
null|Agitation|Finding|false|false||restlessnessnull|Common Specifications in HL7 V3 Publishing|Finding|false|false||common
null|shared attribute|Finding|false|false||commonnull|Common (qualifier value)|LabModifier|false|false||commonnull|Constipation|Finding|false|false||Constipationnull|Common Specifications in HL7 V3 Publishing|Finding|false|false||common
null|shared attribute|Finding|false|false||commonnull|Common (qualifier value)|LabModifier|false|false||commonnull|SURE Test|Finding|false|false||surenull|Certain (qualifier value)|Modifier|false|false||surenull|Drink (dietary substance)|Drug|false|false||drinknull|Liquid substance|Drug|false|false||fluidsnull|Mouse Body Fluid or Substance|Finding|false|false||fluidsnull|Fluid Therapy|Procedure|false|false||fluidsnull|High residue diet|Procedure|false|false|C1304649|high-fiber dietnull|Message Waiting Priority - High|Finding|false|false||high
null|high - ActExposureLevelCode|Finding|false|false||high
null|IPSS Risk Category High|Finding|false|false||high
null|IPSS-R Risk Category High|Finding|false|false||high
null|High (finding)|Finding|false|false||highnull|Observation Value - High|Modifier|false|false||high
null|High|Modifier|false|false||high
null|Abnormally high|Modifier|false|false||highnull|Fiber brand of calcium polycarbophil|Drug|false|false|C1304649|fiber
null|fiber|Drug|false|false|C1304649|fiber
null|fiber|Drug|false|false|C1304649|fiber
null|Fiber brand of calcium polycarbophil|Drug|false|false|C1304649|fibernull|Tissue fiber|Anatomy|false|false|C0012159;C0301568;C1549512;C0225326;C1321801|fibernull|Fiber Device|Device|false|false||fibernull|Animal in fiber production|Entity|false|false||fiber
null|Plant fiber|Entity|false|false||fibernull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false|C1304649|dietnull|Diet therapy|Procedure|false|false|C1304649|dietnull|Narcotics|Drug|false|false||narcotics
null|Narcotics|Drug|false|false||narcoticsnull|prescription document|Finding|false|false||prescriptionnull|Prescription (procedure)|Procedure|false|false||prescriptionnull|Prescription (attribute)|Attribute|false|false||prescriptionnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Drugs, Non-Prescription|Drug|false|false||over-the-counternull|Counter brand of Terbufos|Drug|false|false||counter
null|Counter brand of Terbufos|Drug|false|false||counternull|Counter device|Device|false|false||counternull|Stool Softener brand of docusate sodium|Drug|false|false||stool softener
null|Stool Softener brand of docusate sodium|Drug|false|false||stool softener
null|Stool Softener|Drug|false|false||stool softenernull|Feces|Finding|false|false||stoolnull|Stool seat|Device|false|false||stoolnull|Doctor - Title|Finding|false|false||Doctornull|Physicians|Subject|false|false||Doctornull|Severe Extremity Pain|Finding|false|false||Severe pain
null|Severe pain|Finding|false|false||Severe pain
null|Neck Pain Score 6|Finding|false|false||Severe painnull|Severe - Severity of Illness Code|Finding|false|false||Severe
null|Intensity and Distress 5|Finding|false|false||Severe
null|Severe - Triage Code|Finding|false|false||Severe
null|Severe (severity modifier)|Finding|false|false||Severe
null|Allergy Severity - Severe|Finding|false|false||Severenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|Erythema|Disorder|false|false|C2338258|rednessnull|Redness|Finding|false|false||rednessnull|Red color|Modifier|false|false||rednessnull|Body Substance Discharge|Finding|false|false||drainage
null|Body Fluid Discharge|Finding|false|false||drainagenull|Drainage procedure|Procedure|false|false||drainagenull|Surgical wound|Disorder|false|false|C2338258|incisionnull|Surgical incisions|Procedure|false|false|C2338258|incisionnull|Cranial incision point|Anatomy|false|false|C0332803;C0041834;C0184898|incisionnull|null|Finding|false|false|C1515974|sitenull|Anatomic Site|Anatomy|false|false|C1546778|sitenull|Study Site|Modifier|false|false||site
null|Site|Modifier|false|false||sitenull|Fever symptoms (finding)|Finding|false|false||Fever
null|Fever|Finding|false|false||Fevernull|Greater Than|LabModifier|false|false||greater thannull|Greater|LabModifier|false|false||greaternull|Degrees fahrenheit|LabModifier|false|false||degrees Fahrenheitnull|Academic degree|Finding|false|false||degreesnull|Degree or extent|LabModifier|false|false||degreesnull|Degrees fahrenheit|LabModifier|false|false||Fahrenheitnull|Nausea|Finding|false|false||Nauseanull|null|Attribute|false|false||Nauseanull|Vomiting|Finding|false|false||vomitingnull|Extreme Response|Finding|false|false||Extremenull|Extreme|Modifier|false|false||Extremenull|Somnolence|Disorder|false|false||sleepinessnull|Drowsiness|Finding|false|false||sleepinessnull|Able (qualifier value)|Finding|false|false||ablenull|Ability|Subject|false|false||ablenull|Stay Awake|Drug|false|false||stay awake
null|Stay Awake|Drug|false|false||stay awakenull|Awake (finding)|Finding|false|false||awakenull|Awakening (time frame)|Time|false|false||awakenull|Severe - Severity of Illness Code|Finding|false|false||Severe
null|Intensity and Distress 5|Finding|false|false||Severe
null|Severe - Triage Code|Finding|false|false||Severe
null|Severe (severity modifier)|Finding|false|false||Severe
null|Allergy Severity - Severe|Finding|false|false||Severenull|Headache|Finding|false|false||headachesnull|Pain Relieve brand of acetaminophen|Drug|false|false||pain relievers
null|Pain Relieve brand of acetaminophen|Drug|false|false||pain relievers
null|Analgesics|Drug|false|false||pain relievers
null|Analgesics|Drug|false|false||pain relievers
null|Analgesics|Drug|false|false||pain relieversnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Seizures|Finding|false|false||Seizuresnull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|Problems - What subject filter|Finding|false|false||problemsnull|Vision|Finding|false|false||visionnull|null|Attribute|false|false||visionnull|Specialized Stand Alone Plan - Vision|Entity|false|false||visionnull|Ability to speak|Finding|false|false||ability to speaknull|Ability Question|Finding|false|false||ability tonull|Oral Intake Ability|Finding|false|false||abilitynull|Ability|Subject|false|false||abilitynull|Speak - language ability|Finding|false|false||speak
null|Speaking (function)|Finding|false|false||speak
null|Does speak|Finding|false|false||speaknull|Weakness|Finding|false|false|C0015450;C4266571|Weakness
null|Asthenia|Finding|false|false|C0015450;C4266571|Weaknessnull|Changing|Finding|false|false|C0015450;C4266571|changesnull|Changed status|LabModifier|false|false||changesnull|Observation of Sensation|Finding|false|false|C0015450;C4266571|sensation
null|Sensory perception|Finding|false|false|C0015450;C4266571|sensationnull|sensory exam|Procedure|false|false|C0015450;C4266571|sensationnull|Sensation quality|Modifier|false|false||sensationnull|FANCONI ANEMIA, COMPLEMENTATION GROUP E|Disorder|false|false|C0015450;C4266571|facenull|FANCE wt Allele|Finding|false|false|C0015450;C4266571|face
null|FANCE gene|Finding|false|false|C0015450;C4266571|face
null|ELOVL6 gene|Finding|false|false|C0015450;C4266571|facenull|Head>Face|Anatomy|false|false|C3160739;C1423759;C2828055;C1414531;C3714552;C0004093;C0392747;C0036658;C0542538;C2229507;C0206655;C5575339;C2681631|face
null|Face|Anatomy|false|false|C3160739;C1423759;C2828055;C1414531;C3714552;C0004093;C0392747;C0036658;C0542538;C2229507;C0206655;C5575339;C2681631|facenull|Face (spatial concept)|Modifier|false|false||facenull|Alveolar rhabdomyosarcoma|Disorder|false|false|C0446516;C0015450;C4266571|armsnull|Adherence to Refills and Medications Scale|Finding|false|false|C0446516;C0015450;C4266571|arms
null|KIDINS220 gene|Finding|false|false|C0446516;C0015450;C4266571|armsnull|Upper arm|Anatomy|false|false|C5782111;C5575339;C2681631;C0206655|armsnull|null|Attribute|false|false|C0446516|armsnull|Leg|Anatomy|false|false||leg
null|Lower Extremity|Anatomy|false|false||legnull|Call - dosing instruction fragment|Finding|false|false||Call
null|Call (Instruction)|Finding|false|false||Call
null|Decision|Finding|false|false||Call
null|CHL1 gene|Finding|false|false||Callnull|Proximal|Modifier|false|false||nearestnull|Encounter Referral Source - emergency room|Finding|false|false||Emergency Roomnull|Accident and Emergency department|Device|false|false||Emergency Roomnull|Accident and Emergency department|Entity|false|false||Emergency Roomnull|Consent Non-Disclosure Reason - Emergency|Finding|false|false||Emergency
null|Admission Type - Emergency|Finding|false|false||Emergency
null|Referral category - Emergency|Finding|false|false||Emergency
null|Emergencies [Disease/Finding]|Finding|false|false||Emergency
null|Consent Bypass Reason - Emergency|Finding|false|false||Emergency
null|Level of Care - Emergency|Finding|false|false||Emergency
null|Certification patient type - Emergency|Finding|false|false||Emergency
null|Encounter Admission Source - emergency|Finding|false|false||Emergency
null|Patient Class - Emergency|Finding|false|false||Emergency
null|Visit Priority Code - Emergency|Finding|false|false||Emergencynull|emergency encounter|Procedure|false|false||Emergencynull|Emergency Situation|Phenomenon|false|false||Emergencynull|Specialty Type - Emergency|Title|false|false||Emergencynull|Bale out|Time|false|false||Emergencynull|Room - Patient location type|Modifier|false|false||Room
null|Room|Modifier|false|false||Roomnull|Experience (Practice)|Finding|false|false||experience
null|Experience|Finding|false|false||experiencenull|Following|Time|false|false||following
null|Status post|Time|false|false||followingnull|Sudden (qualifier value)|Modifier|false|false||Suddennull|Numbness|Finding|false|false|C0015450;C4266571|numbness
null|Hypesthesia|Finding|false|false|C0015450;C4266571|numbnessnull|Weakness|Finding|false|false|C0015450;C4266571|weakness
null|Asthenia|Finding|false|false|C0015450;C4266571|weaknessnull|FANCONI ANEMIA, COMPLEMENTATION GROUP E|Disorder|false|false|C0015450;C4266571|facenull|FANCE wt Allele|Finding|false|false|C0015450;C4266571|face
null|FANCE gene|Finding|false|false|C0015450;C4266571|face
null|ELOVL6 gene|Finding|false|false|C0015450;C4266571|facenull|Head>Face|Anatomy|false|false|C1824218;C3715044;C3160739;C1423759;C2828055;C1414531;C3714552;C0004093;C0028643;C0020580;C1522541;C5400986;C4761640;C3495676|face
null|Face|Anatomy|false|false|C1824218;C3715044;C3160739;C1423759;C2828055;C1414531;C3714552;C0004093;C0028643;C0020580;C1522541;C5400986;C4761640;C3495676|facenull|Face (spatial concept)|Modifier|false|false||facenull|Anorectal Malformations|Disorder|false|false|C0446516;C1140618;C1269078;C0015450;C4266571|armnull|AKR1A1 wt Allele|Finding|false|false|C0015450;C4266571;C0446516;C1140618;C1269078|arm
null|ARMC9 gene|Finding|false|false|C0015450;C4266571;C0446516;C1140618;C1269078|armnull|Protocol Treatment Arm|Procedure|false|false|C0446516;C1140618;C1269078;C0015450;C4266571|arm
null|Axillary Reverse Mapping|Procedure|false|false|C0446516;C1140618;C1269078;C0015450;C4266571|arm
null|Study Arm|Procedure|false|false|C0446516;C1140618;C1269078;C0015450;C4266571|armnull|Upper arm|Anatomy|false|false|C1522541;C5400986;C4761640;C1824218;C3715044;C3495676|arm
null|null|Anatomy|false|false|C1522541;C5400986;C4761640;C1824218;C3715044;C3495676|arm
null|Upper Extremity|Anatomy|false|false|C1522541;C5400986;C4761640;C1824218;C3715044;C3495676|armnull|Leg|Anatomy|false|false||leg
null|Lower Extremity|Anatomy|false|false||legnull|Sudden (qualifier value)|Modifier|false|false||Suddennull|Confusion|Disorder|false|false||confusionnull|Clouded consciousness|Finding|false|false||confusionnull|Comprehension|Finding|false|false||understandingnull|Sudden (qualifier value)|Modifier|false|false||Suddennull|Dizziness|Finding|false|false||dizziness
null|Vertigo|Finding|false|false||dizzinessnull|Impairment of balance|Finding|false|false||loss of balancenull|Loss (adaptation)|Finding|false|false||lossnull|Loss (quantitative)|LabModifier|false|false||lossnull|Balance (substance)|Drug|false|false||balance
null|Balance (substance)|Drug|false|false||balancenull|Ability to balance|Finding|false|false||balance
null|Equilibrium|Finding|false|false||balancenull|examination of balance|Procedure|false|false||balancenull|balance device|Device|false|false||balancenull|Balanced (qualifier value)|Modifier|false|false||balancenull|Coordination of Benefits - Coordination|Finding|false|false||coordination
null|Coordinated|Finding|false|false||coordination
null|Physiologic Coordination|Finding|false|false||coordinationnull|Sudden (qualifier value)|Modifier|false|false||Suddennull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Headache|Finding|false|false||headachesnull|Known|Modifier|false|false||knownnull|Indication of (contextual qualifier)|Finding|true|false||reasonnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions