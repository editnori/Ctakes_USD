 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|43,52|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|43,52|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|43,57|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|77,86|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|77,86|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|77,91|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|133,136|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|144,151|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|144,151|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|153,161|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|SIMPLE_SEGMENT|164,173|false|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|164,173|false|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|164,173|false|false|false|C0020517|Hypersensitivity|Allergies
Attribute|Clinical Attribute|SIMPLE_SEGMENT|185,194|true|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|185,194|true|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|185,194|true|false|false|C0020517|Hypersensitivity|Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|197,219|true|false|false|C0041755|Adverse reaction to drug|Adverse Drug Reactions
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|205,209|true|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|Drug
Finding|Finding|SIMPLE_SEGMENT|205,209|true|false|false|C0740721|Drug problem|Drug
Finding|Pathologic Function|SIMPLE_SEGMENT|205,219|true|false|false|C0041755|Adverse reaction to drug|Drug Reactions
Event|Event|SIMPLE_SEGMENT|210,219|true|false|false|||Reactions
Event|Event|SIMPLE_SEGMENT|222,231|false|false|false|||Attending
Finding|Functional Concept|SIMPLE_SEGMENT|222,231|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|SIMPLE_SEGMENT|240,255|false|false|false|C0277786|Chief complaint (finding)|Chief Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|246,255|false|false|false|C3864418||Complaint
Event|Event|SIMPLE_SEGMENT|246,255|false|false|false|||Complaint
Finding|Finding|SIMPLE_SEGMENT|246,255|false|false|false|C5441521|Complaint (finding)|Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|257,267|false|false|false|C2979880||subjective
Finding|Finding|SIMPLE_SEGMENT|257,267|false|false|false|C2266644|subjective (symptom)|subjective
Event|Event|SIMPLE_SEGMENT|268,274|false|false|false|||fevers
Finding|Sign or Symptom|SIMPLE_SEGMENT|268,274|false|false|false|C0015967|Fever|fevers
Event|Event|SIMPLE_SEGMENT|276,284|false|false|false|||lethargy
Finding|Sign or Symptom|SIMPLE_SEGMENT|276,284|false|false|false|C0023380|Lethargy|lethargy
Finding|Finding|SIMPLE_SEGMENT|290,296|false|false|false|C4554530|Bloody|bloody
Drug|Substance|SIMPLE_SEGMENT|297,302|false|false|false|C1550628|Drain - SpecimenType|drain
Finding|Intellectual Product|SIMPLE_SEGMENT|297,302|false|false|false|C1546604|Drain Specimen Code|drain
Event|Event|SIMPLE_SEGMENT|303,309|false|false|false|||output
Finding|Conceptual Entity|SIMPLE_SEGMENT|303,309|false|false|false|C1709366|system output|output
Procedure|Health Care Activity|SIMPLE_SEGMENT|303,309|false|false|false|C3251815|Measurement of fluid output|output
Finding|Classification|SIMPLE_SEGMENT|313,318|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|SIMPLE_SEGMENT|319,327|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|319,327|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|331,349|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|340,349|false|false|false|C0945766||Procedure
Event|Event|SIMPLE_SEGMENT|340,349|false|false|false|||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|340,349|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|340,349|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|340,349|false|false|false|C0184661|Interventional procedure|Procedure
Finding|Gene or Genome|SIMPLE_SEGMENT|364,369|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|370,376|false|false|false|C0030797|Pelvis|pelvic
Drug|Substance|SIMPLE_SEGMENT|377,382|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|377,382|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|383,394|false|false|false|||collections
Event|Event|SIMPLE_SEGMENT|399,405|false|false|false|||guided
Event|Event|SIMPLE_SEGMENT|407,420|false|false|false|||repositioning
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|407,420|false|false|false|C0556030|Repositioning (procedure)|repositioning
Drug|Substance|SIMPLE_SEGMENT|433,438|false|false|false|C1550628|Drain - SpecimenType|drain
Event|Event|SIMPLE_SEGMENT|433,438|false|false|false|||drain
Finding|Intellectual Product|SIMPLE_SEGMENT|433,438|false|false|false|C1546604|Drain Specimen Code|drain
Event|Event|SIMPLE_SEGMENT|443,452|false|false|false|||placement
Procedure|Health Care Activity|SIMPLE_SEGMENT|443,452|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|443,452|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Finding|Functional Concept|SIMPLE_SEGMENT|459,469|false|false|false|C1524062|Additional|additional
Drug|Substance|SIMPLE_SEGMENT|471,476|false|false|false|C1550628|Drain - SpecimenType|drain
Event|Event|SIMPLE_SEGMENT|471,476|false|false|false|||drain
Finding|Intellectual Product|SIMPLE_SEGMENT|471,476|false|false|false|C1546604|Drain Specimen Code|drain
Event|Activity|SIMPLE_SEGMENT|484,491|false|false|false|C1883720|Removing (action)|Removal
Event|Event|SIMPLE_SEGMENT|484,491|false|false|false|||Removal
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|484,491|false|false|false|C0015252;C0185115;C0728940|Excision;Extraction;removal technique|Removal
Drug|Substance|SIMPLE_SEGMENT|516,521|false|false|false|C1550628|Drain - SpecimenType|drain
Event|Event|SIMPLE_SEGMENT|516,521|false|false|false|||drain
Finding|Intellectual Product|SIMPLE_SEGMENT|516,521|false|false|false|C1546604|Drain Specimen Code|drain
Event|Event|SIMPLE_SEGMENT|527,534|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|527,534|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|527,534|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|527,534|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|527,537|false|false|false|C0262926|Medical History|History of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|527,553|false|false|false|C0488508||History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|527,553|false|false|false|C0262512|History of present illness (finding)|History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|538,545|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Idea or Concept|SIMPLE_SEGMENT|538,545|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Finding|SIMPLE_SEGMENT|538,553|false|false|false|C4264312|Present illness|Present Illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|546,553|false|false|false|C0221423|Illness (finding)|Illness
Event|Event|SIMPLE_SEGMENT|578,581|false|false|false|||PMH
Finding|Finding|SIMPLE_SEGMENT|578,581|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|PMH
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|585,597|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|SIMPLE_SEGMENT|585,597|false|false|false|||hypertension
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|602,609|false|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|SIMPLE_SEGMENT|602,609|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Event|Event|SIMPLE_SEGMENT|602,609|false|false|false|||bladder
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|602,609|false|false|false|C0872388|Procedures on bladder|bladder
Disorder|Neoplastic Process|SIMPLE_SEGMENT|611,617|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|SIMPLE_SEGMENT|611,617|false|false|false|||cancer
Finding|Finding|SIMPLE_SEGMENT|619,623|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|SIMPLE_SEGMENT|619,623|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|SIMPLE_SEGMENT|619,623|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Finding|SIMPLE_SEGMENT|619,629|false|false|false|C0205082;C4554016|Enneking High Surgical Grade;Severe (severity modifier)|high grade
Finding|Intellectual Product|SIMPLE_SEGMENT|619,629|false|false|false|C0205082;C4554016|Enneking High Surgical Grade;Severe (severity modifier)|high grade
Finding|Classification|SIMPLE_SEGMENT|624,629|false|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|grade
Finding|Finding|SIMPLE_SEGMENT|624,629|false|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|grade
Disorder|Neoplastic Process|SIMPLE_SEGMENT|630,659|false|false|false|C1512751|Invasive Urothelial Carcinoma|invasive urothelial carcinoma
Disorder|Neoplastic Process|SIMPLE_SEGMENT|639,659|false|false|false|C0007138;C2145472|Carcinoma, Transitional Cell;Urothelial Carcinoma|urothelial carcinoma
Disorder|Neoplastic Process|SIMPLE_SEGMENT|650,659|false|false|false|C0007097|Carcinoma|carcinoma
Finding|Finding|SIMPLE_SEGMENT|660,664|false|false|false|C1711132|pT2b TNM Finding|pT2b
Event|Event|SIMPLE_SEGMENT|671,674|false|false|false|||TAH
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|671,674|false|false|false|C0404079|Total abdominal hysterectomy|TAH
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|671,678|false|false|false|C0542407|Total abdominal hysterectomy with bilateral salpingo-oophorectomy|TAH/BSO
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|675,678|false|false|false|C0054252|Buthionine Sulfoximine|BSO
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|675,678|false|false|false|C0054252|Buthionine Sulfoximine|BSO
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|675,678|false|false|false|C0054252|Buthionine Sulfoximine|BSO
Event|Event|SIMPLE_SEGMENT|675,678|false|false|false|||BSO
Drug|Chemical Viewed Structurally|SIMPLE_SEGMENT|680,687|false|false|false|C0302912|Radicals (chemistry)|radical
Event|Event|SIMPLE_SEGMENT|680,687|false|false|false|||radical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|680,698|false|false|false|C0194401|Complete cystectomy|radical cystectomy
Event|Event|SIMPLE_SEGMENT|688,698|false|false|false|||cystectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|688,698|false|false|false|C0010651|Cystectomy|cystectomy
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|701,706|false|false|false|C0020885|ileum|ileal
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|701,714|false|false|false|C0441253|Structure of ileal conduit|ileal conduit
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|701,714|false|false|false|C0348002|Ileal conduit procedure|ileal conduit
Event|Event|SIMPLE_SEGMENT|707,714|false|false|false|||conduit
Event|Event|SIMPLE_SEGMENT|719,734|false|false|false|||intra-abdominal
Finding|Functional Concept|SIMPLE_SEGMENT|719,734|false|false|false|C1512911|Intraabdominal Route of Administration|intra-abdominal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|736,745|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|SIMPLE_SEGMENT|736,745|false|false|false|||infection
Finding|Pathologic Function|SIMPLE_SEGMENT|736,745|false|false|false|C3714514|Infection|infection
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|750,756|false|false|false|C0030797|Pelvis|pelvic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|750,773|false|false|false|C1697454|Pelvic fluid collection|pelvic fluid collection
Drug|Substance|SIMPLE_SEGMENT|757,762|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|757,762|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|763,773|false|false|false|||collection
Finding|Conceptual Entity|SIMPLE_SEGMENT|763,773|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|SIMPLE_SEGMENT|763,773|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|SIMPLE_SEGMENT|763,773|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|SIMPLE_SEGMENT|763,773|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Drug|Substance|SIMPLE_SEGMENT|789,794|false|false|false|C1550628|Drain - SpecimenType|drain
Event|Event|SIMPLE_SEGMENT|789,794|false|false|false|||drain
Finding|Intellectual Product|SIMPLE_SEGMENT|789,794|false|false|false|C1546604|Drain Specimen Code|drain
Event|Event|SIMPLE_SEGMENT|796,805|false|false|false|||placement
Procedure|Health Care Activity|SIMPLE_SEGMENT|796,805|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|796,805|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Event|Event|SIMPLE_SEGMENT|814,822|false|false|false|||presents
Event|Event|SIMPLE_SEGMENT|851,858|false|false|false|||malaise
Finding|Sign or Symptom|SIMPLE_SEGMENT|851,858|false|false|false|C0231218|Malaise|malaise
Finding|Idea or Concept|SIMPLE_SEGMENT|865,868|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|865,868|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|872,878|false|false|false|||fevers
Finding|Sign or Symptom|SIMPLE_SEGMENT|872,878|false|false|false|C0015967|Fever|fevers
Finding|Body Substance|SIMPLE_SEGMENT|883,890|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|883,890|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|883,890|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Substance|SIMPLE_SEGMENT|915,920|false|false|false|C1550628|Drain - SpecimenType|drain
Event|Event|SIMPLE_SEGMENT|915,920|false|false|false|||drain
Finding|Intellectual Product|SIMPLE_SEGMENT|915,920|false|false|false|C1546604|Drain Specimen Code|drain
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|915,930|false|false|false|C3495845|Drain placement|drain placement
Event|Event|SIMPLE_SEGMENT|921,930|false|false|false|||placement
Procedure|Health Care Activity|SIMPLE_SEGMENT|921,930|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|921,930|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Finding|Functional Concept|SIMPLE_SEGMENT|936,951|false|false|false|C1512911|Intraabdominal Route of Administration|intra-abdominal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|936,968|false|false|false|C4285843|Intra-abdominal fluid collection|intra-abdominal fluid collection
Drug|Substance|SIMPLE_SEGMENT|952,957|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|952,957|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|952,957|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|958,968|false|false|false|||collection
Finding|Conceptual Entity|SIMPLE_SEGMENT|958,968|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|SIMPLE_SEGMENT|958,968|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|SIMPLE_SEGMENT|958,968|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|SIMPLE_SEGMENT|958,968|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|973,982|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|SIMPLE_SEGMENT|973,982|false|false|false|||infection
Finding|Pathologic Function|SIMPLE_SEGMENT|973,982|false|false|false|C3714514|Infection|infection
Event|Event|SIMPLE_SEGMENT|984,991|false|false|false|||thought
Finding|Idea or Concept|SIMPLE_SEGMENT|984,991|false|false|true|C0039869;C4319827|Thought|thought
Finding|Mental Process|SIMPLE_SEGMENT|984,991|false|false|true|C0039869;C4319827|Thought|thought
Event|Event|SIMPLE_SEGMENT|999,1010|false|false|false|||complicated
Event|Event|SIMPLE_SEGMENT|1021,1024|false|false|false|||TAH
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1021,1024|false|false|false|C0404079|Total abdominal hysterectomy|TAH
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1021,1028|false|false|false|C0542407|Total abdominal hysterectomy with bilateral salpingo-oophorectomy|TAH/BSO
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1025,1028|false|false|false|C0054252|Buthionine Sulfoximine|BSO
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|1025,1028|false|false|false|C0054252|Buthionine Sulfoximine|BSO
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1025,1028|false|false|false|C0054252|Buthionine Sulfoximine|BSO
Event|Event|SIMPLE_SEGMENT|1025,1028|false|false|false|||BSO
Drug|Chemical Viewed Structurally|SIMPLE_SEGMENT|1030,1037|false|false|false|C0302912|Radicals (chemistry)|radical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1030,1048|false|false|false|C0194401|Complete cystectomy|radical cystectomy
Event|Event|SIMPLE_SEGMENT|1038,1048|false|false|false|||cystectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1038,1048|false|false|false|C0010651|Cystectomy|cystectomy
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1053,1059|false|false|false|C0030797|Pelvis|pelvic
Finding|Body Substance|SIMPLE_SEGMENT|1061,1066|false|false|false|C0024202|Lymph|lymph
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1061,1071|false|false|false|C0024204|lymph nodes|lymph node
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1061,1078|false|false|false|C0193842|Biopsy of lymph node|lymph node biopsy
Event|Event|SIMPLE_SEGMENT|1072,1078|false|false|false|||biopsy
Finding|Finding|SIMPLE_SEGMENT|1072,1078|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Finding|Intellectual Product|SIMPLE_SEGMENT|1072,1078|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1072,1078|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Procedure|Health Care Activity|SIMPLE_SEGMENT|1072,1078|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1085,1094|false|false|false|C0945766||procedure
Event|Event|SIMPLE_SEGMENT|1085,1094|false|false|false|||procedure
Event|Occupational Activity|SIMPLE_SEGMENT|1085,1094|false|false|false|C1546467|Act Class - procedure|procedure
Finding|Functional Concept|SIMPLE_SEGMENT|1085,1094|false|false|false|C2700391|Procedure (set of actions)|procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1085,1094|false|false|false|C0184661|Interventional procedure|procedure
Event|Event|SIMPLE_SEGMENT|1142,1149|false|false|false|||noticed
Event|Event|SIMPLE_SEGMENT|1162,1169|false|false|false|||malaise
Finding|Sign or Symptom|SIMPLE_SEGMENT|1162,1169|false|false|false|C0231218|Malaise|malaise
Finding|Idea or Concept|SIMPLE_SEGMENT|1176,1179|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|1176,1179|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|1184,1189|false|false|false|||fever
Finding|Finding|SIMPLE_SEGMENT|1184,1189|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|1184,1189|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Event|Event|SIMPLE_SEGMENT|1192,1198|false|false|false|||rigors
Finding|Sign or Symptom|SIMPLE_SEGMENT|1192,1198|false|false|false|C0424790|Rigor - Temperature-associated observation|rigors
Finding|Finding|SIMPLE_SEGMENT|1213,1220|false|false|false|C4534363|At home|at home
Finding|Idea or Concept|SIMPLE_SEGMENT|1216,1220|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|1216,1220|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|1216,1220|false|false|false|C1553498|home health encounter|home
Event|Event|SIMPLE_SEGMENT|1226,1231|false|false|false|||notes
Event|Event|SIMPLE_SEGMENT|1242,1250|false|false|false|||drainage
Finding|Body Substance|SIMPLE_SEGMENT|1242,1250|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Finding|Sign or Symptom|SIMPLE_SEGMENT|1242,1250|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1242,1250|false|false|false|C0013103|Drainage procedure|drainage
Finding|Functional Concept|SIMPLE_SEGMENT|1260,1275|false|false|false|C1512911|Intraabdominal Route of Administration|intra-abdominal
Drug|Substance|SIMPLE_SEGMENT|1276,1281|false|false|false|C1550628|Drain - SpecimenType|drain
Event|Event|SIMPLE_SEGMENT|1276,1281|false|false|false|||drain
Finding|Intellectual Product|SIMPLE_SEGMENT|1276,1281|false|false|false|C1546604|Drain Specimen Code|drain
Event|Event|SIMPLE_SEGMENT|1285,1291|false|false|false|||darker
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|1302,1310|false|false|false|C0559495|Urological stoma|urostomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1302,1310|false|false|false|C0856443|Urostomy procedure|urostomy
Event|Event|SIMPLE_SEGMENT|1311,1317|false|false|false|||output
Finding|Conceptual Entity|SIMPLE_SEGMENT|1311,1317|false|false|false|C1709366|system output|output
Procedure|Health Care Activity|SIMPLE_SEGMENT|1311,1317|false|false|false|C3251815|Measurement of fluid output|output
Event|Event|SIMPLE_SEGMENT|1327,1336|false|false|false|||unchanged
Finding|Finding|SIMPLE_SEGMENT|1327,1336|false|false|false|C0442739||unchanged
Event|Event|SIMPLE_SEGMENT|1342,1347|false|false|false|||notes
Finding|Intellectual Product|SIMPLE_SEGMENT|1365,1369|false|false|false|C1547225|Mild Severity of Illness Code|mild
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1370,1373|false|false|false|C0230180|Structure of left lower quadrant of abdomen|LLQ
Finding|Sign or Symptom|SIMPLE_SEGMENT|1370,1378|false|false|false|C0238551|Left lower quadrant pain|LLQ pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1374,1378|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|1374,1378|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|1374,1378|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1374,1378|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|1384,1390|false|false|false|||denies
Event|Event|SIMPLE_SEGMENT|1391,1399|true|false|false|||diarrhea
Finding|Finding|SIMPLE_SEGMENT|1391,1399|true|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|SIMPLE_SEGMENT|1391,1399|true|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1401,1406|true|false|false|C0018932|Hematochezia|BRBPR
Event|Event|SIMPLE_SEGMENT|1401,1406|true|false|false|||BRBPR
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1408,1412|true|false|false|C5779629|Eruption of skin (disorder)|rash
Event|Event|SIMPLE_SEGMENT|1408,1412|true|false|false|||rash
Finding|Pathologic Function|SIMPLE_SEGMENT|1408,1412|true|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Sign or Symptom|SIMPLE_SEGMENT|1408,1412|true|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Drug|Organic Chemical|SIMPLE_SEGMENT|1414,1419|true|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1414,1419|true|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|SIMPLE_SEGMENT|1414,1419|true|false|false|||cough
Finding|Sign or Symptom|SIMPLE_SEGMENT|1414,1419|true|false|false|C0010200|Coughing|cough
Event|Event|SIMPLE_SEGMENT|1422,1430|false|false|false|||headache
Finding|Sign or Symptom|SIMPLE_SEGMENT|1422,1430|false|false|false|C0018681|Headache|headache
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1432,1436|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|SIMPLE_SEGMENT|1432,1436|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|SIMPLE_SEGMENT|1432,1436|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Finding|Sign or Symptom|SIMPLE_SEGMENT|1432,1446|false|false|false|C0151315|Neck stiffness|neck stiffness
Event|Event|SIMPLE_SEGMENT|1437,1446|false|false|false|||stiffness
Finding|Sign or Symptom|SIMPLE_SEGMENT|1437,1446|false|false|false|C0427008|Stiffness|stiffness
Event|Event|SIMPLE_SEGMENT|1452,1461|false|false|false|||presented
Event|Event|SIMPLE_SEGMENT|1495,1504|false|false|false|||evaluated
Drug|Substance|SIMPLE_SEGMENT|1518,1523|false|false|false|C1550628|Drain - SpecimenType|drain
Event|Event|SIMPLE_SEGMENT|1518,1523|false|false|false|||drain
Finding|Intellectual Product|SIMPLE_SEGMENT|1518,1523|false|false|false|C1546604|Drain Specimen Code|drain
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|1524,1531|false|false|false|C1706355|Culture Dose Form|culture
Event|Event|SIMPLE_SEGMENT|1524,1531|false|false|false|||culture
Finding|Functional Concept|SIMPLE_SEGMENT|1524,1531|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Finding|Idea or Concept|SIMPLE_SEGMENT|1524,1531|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1524,1531|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|culture
Event|Event|SIMPLE_SEGMENT|1540,1547|false|false|false|||started
Drug|Antibiotic|SIMPLE_SEGMENT|1552,1557|false|false|false|C0250482|Zosyn|zosyn
Drug|Organic Chemical|SIMPLE_SEGMENT|1552,1557|false|false|false|C0250482|Zosyn|zosyn
Event|Event|SIMPLE_SEGMENT|1552,1557|false|false|false|||zosyn
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1562,1572|false|false|false|C0042313|vancomycin|vancomycin
Drug|Antibiotic|SIMPLE_SEGMENT|1562,1572|false|false|false|C0042313|vancomycin|vancomycin
Event|Event|SIMPLE_SEGMENT|1562,1572|false|false|false|||vancomycin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1562,1572|false|false|false|C0489941|Vancomycin measurement|vancomycin
Drug|Organic Chemical|SIMPLE_SEGMENT|1589,1602|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1589,1602|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Event|Event|SIMPLE_SEGMENT|1589,1602|false|false|false|||acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1589,1602|false|false|false|C0373527|Acetaminophen measurement|acetaminophen
Event|Event|SIMPLE_SEGMENT|1613,1624|false|false|false|||transferred
Event|Event|SIMPLE_SEGMENT|1644,1654|false|false|false|||management
Event|Occupational Activity|SIMPLE_SEGMENT|1644,1654|false|false|false|C0001554;C1273870|Administration occupational activities;Management procedure|management
Procedure|Health Care Activity|SIMPLE_SEGMENT|1644,1654|false|false|false|C0376636|Disease Management|management
Finding|Finding|SIMPLE_SEGMENT|1661,1681|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Event|Event|SIMPLE_SEGMENT|1666,1673|false|false|false|||Medical
Finding|Functional Concept|SIMPLE_SEGMENT|1666,1673|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|1666,1673|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|1666,1673|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|1666,1673|false|false|false|C0199168|Medical service|Medical
Finding|Finding|SIMPLE_SEGMENT|1666,1681|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1674,1681|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1674,1681|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|1674,1681|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1685,1697|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|SIMPLE_SEGMENT|1685,1697|false|false|false|||Hypertension
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1707,1710|false|false|false|C0396060|Congenital laryngeal adductor palsy|lap
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1707,1710|false|false|false|C1870042|ACP2 protein, human|lap
Drug|Enzyme|SIMPLE_SEGMENT|1707,1710|false|false|false|C1870042|ACP2 protein, human|lap
Event|Event|SIMPLE_SEGMENT|1707,1710|false|false|false|||lap
Finding|Finding|SIMPLE_SEGMENT|1707,1710|false|false|false|C0456170;C1412132;C1413323;C1423544;C1424863;C1425522;C2827449;C3540509;C5575443;C5890955|ACP2 gene;ACP2 wt Allele;CEBPB gene;CEBPB wt Allele;CENPJ gene;LAP3 gene;LAP3 wt Allele;Left atrial pressure;PICALM gene;PICALM wt Allele|lap
Finding|Gene or Genome|SIMPLE_SEGMENT|1707,1710|false|false|false|C0456170;C1412132;C1413323;C1423544;C1424863;C1425522;C2827449;C3540509;C5575443;C5890955|ACP2 gene;ACP2 wt Allele;CEBPB gene;CEBPB wt Allele;CENPJ gene;LAP3 gene;LAP3 wt Allele;Left atrial pressure;PICALM gene;PICALM wt Allele|lap
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1707,1710|false|false|false|C0031150|Laparoscopy|lap
Event|Event|SIMPLE_SEGMENT|1711,1716|false|false|false|||chole
Finding|Functional Concept|SIMPLE_SEGMENT|1726,1730|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1726,1735|false|false|false|C0230432;C4281599|Structure of left knee;Structure of left knee region|left knee
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1726,1735|false|false|false|C0230432;C4281599|Structure of left knee;Structure of left knee region|left knee
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1731,1735|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1731,1735|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|1731,1735|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1731,1735|false|false|false|C0562271|Examination of knee joint|knee
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1731,1747|false|false|false|C5575606||knee replacement
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1731,1747|false|false|false|C0086511|Knee Replacement Arthroplasty|knee replacement
Event|Event|SIMPLE_SEGMENT|1736,1747|false|false|false|||replacement
Finding|Functional Concept|SIMPLE_SEGMENT|1736,1747|false|false|false|C0559956|Replacement|replacement
Procedure|Health Care Activity|SIMPLE_SEGMENT|1736,1747|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|replacement
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1736,1747|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|replacement
Event|Event|SIMPLE_SEGMENT|1757,1768|false|false|false|||laminectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1757,1768|false|false|false|C0022983|Laminectomy|laminectomy
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1781,1784|false|false|false|C1114365||age
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1781,1784|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|SIMPLE_SEGMENT|1781,1784|false|false|false|C0162574|Glycation End Products, Advanced|age
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1794,1801|false|false|false|C0005682|Urinary Bladder|Bladder
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1794,1801|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|Bladder
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1794,1801|false|false|false|C0872388|Procedures on bladder|Bladder
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1794,1808|false|false|false|C0005684;C0005695;C0699885|Bladder Neoplasm;Carcinoma of bladder;Malignant neoplasm of urinary bladder|Bladder Cancer
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1802,1808|false|false|false|C0006826|Malignant Neoplasms|Cancer
Event|Event|SIMPLE_SEGMENT|1802,1808|false|false|false|||Cancer
Finding|Finding|SIMPLE_SEGMENT|1809,1813|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|SIMPLE_SEGMENT|1809,1813|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|SIMPLE_SEGMENT|1809,1813|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Finding|SIMPLE_SEGMENT|1809,1819|false|false|false|C0205082;C4554016|Enneking High Surgical Grade;Severe (severity modifier)|high grade
Finding|Intellectual Product|SIMPLE_SEGMENT|1809,1819|false|false|false|C0205082;C4554016|Enneking High Surgical Grade;Severe (severity modifier)|high grade
Finding|Classification|SIMPLE_SEGMENT|1814,1819|false|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|grade
Finding|Finding|SIMPLE_SEGMENT|1814,1819|false|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|grade
Anatomy|Cell Component|SIMPLE_SEGMENT|1820,1823|false|false|false|C1167383|membrane attack complex location|TCC
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1820,1823|false|false|false|C1861305|TARSAL-CARPAL COALITION SYNDROME|TCC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1820,1823|false|false|false|C0077072;C5552697|Membrane Attack Complex;triclocarban|TCC
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1820,1823|false|false|false|C0077072;C5552697|Membrane Attack Complex;triclocarban|TCC
Drug|Organic Chemical|SIMPLE_SEGMENT|1820,1823|false|false|false|C0077072;C5552697|Membrane Attack Complex;triclocarban|TCC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1820,1823|false|false|false|C0077072;C5552697|Membrane Attack Complex;triclocarban|TCC
Event|Event|SIMPLE_SEGMENT|1820,1823|false|false|false|||TCC
Event|Event|SIMPLE_SEGMENT|1828,1837|false|false|false|||diagnosed
Finding|Intellectual Product|SIMPLE_SEGMENT|1846,1850|false|false|false|C1720594|Then - dosing instruction fragment|then
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1856,1862|false|false|false|C0030797|Pelvis|pelvic
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1856,1866|false|false|false|C0203201|Magnetic Resonance Imaging (MRI) of Pelvis|pelvic MRI
Event|Event|SIMPLE_SEGMENT|1863,1866|false|false|false|||MRI
Finding|Gene or Genome|SIMPLE_SEGMENT|1863,1866|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1863,1866|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|SIMPLE_SEGMENT|1863,1866|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1869,1877|false|false|false|C1269955|Tumor Cell Invasion|invasion
Event|Event|SIMPLE_SEGMENT|1869,1877|false|false|false|||invasion
Finding|Pathologic Function|SIMPLE_SEGMENT|1869,1877|false|false|false|C2699153|Cell Invasion|invasion
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1883,1890|false|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1883,1890|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1883,1890|false|false|false|C0872388|Procedures on bladder|bladder
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1883,1895|false|false|false|C0458421|Wall of bladder|bladder wall
Event|Event|SIMPLE_SEGMENT|1897,1908|false|false|false|||perivesical
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1910,1914|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1910,1921|false|false|false|C0225317;C4532079|Neck+Chest>Soft tissue;soft tissue|soft tissue
Anatomy|Tissue|SIMPLE_SEGMENT|1910,1921|false|false|false|C0225317;C4532079|Neck+Chest>Soft tissue;soft tissue|soft tissue
Anatomy|Tissue|SIMPLE_SEGMENT|1915,1921|false|false|false|C0040300|Body tissue|tissue
Finding|Intellectual Product|SIMPLE_SEGMENT|1915,1921|false|false|false|C1547928|Tissue Specimen Code|tissue
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1926,1934|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1935,1942|false|false|false|C0042232|Vagina|vaginal
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|1935,1942|false|false|false|C1272941|Vaginal Dosage Form|vaginal
Finding|Finding|SIMPLE_SEGMENT|1935,1942|false|false|false|C1522570;C4521343|Vaginal (intended site);Vaginal Route of Administration|vaginal
Finding|Functional Concept|SIMPLE_SEGMENT|1935,1942|false|false|false|C1522570;C4521343|Vaginal (intended site);Vaginal Route of Administration|vaginal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1935,1947|false|false|false|C0447612|Vaginal wall|vaginal wall
Event|Event|SIMPLE_SEGMENT|1949,1950|false|false|false|||/
Event|Event|SIMPLE_SEGMENT|1955,1962|false|false|false|||staging
Finding|Functional Concept|SIMPLE_SEGMENT|1955,1962|false|false|false|C0332305|With staging|staging
Event|Event|SIMPLE_SEGMENT|1972,1984|false|false|false|||hysterectomy
Finding|Finding|SIMPLE_SEGMENT|1972,1984|false|false|false|C1548863|Consent Type - Hysterectomy|hysterectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1972,1984|false|false|false|C0020699|Hysterectomy|hysterectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1989,2011|false|false|false|C0278321|Bilateral oophorectomy|bilateral oophorectomy
Event|Event|SIMPLE_SEGMENT|1999,2011|false|false|false|||oophorectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1999,2011|false|false|false|C0029936|Ovariectomy|oophorectomy
Finding|Gene or Genome|SIMPLE_SEGMENT|2016,2021|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Finding|Finding|SIMPLE_SEGMENT|2016,2028|false|false|false|C0151994|Enlarged uterus|large uterus
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2022,2028|false|false|false|C0042149;C1519876;C4266525|Mouse Uterus;Pelvis>Uterus;Uterus|uterus
Anatomy|Tissue|SIMPLE_SEGMENT|2022,2028|false|false|false|C0042149;C1519876;C4266525|Mouse Uterus;Pelvis>Uterus;Uterus|uterus
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2022,2028|false|false|false|C0042131;C0496919|Neoplasm of uncertain or unknown behavior of uterus;Uterine Diseases|uterus
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2022,2028|false|false|false|C0042131;C0496919|Neoplasm of uncertain or unknown behavior of uterus;Uterine Diseases|uterus
Event|Event|SIMPLE_SEGMENT|2022,2028|false|false|false|||uterus
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2022,2028|false|false|false|C0869889|examination of uterus|uterus
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2032,2039|false|false|false|C0023267|Fibroid Tumor|fibroid
Event|Event|SIMPLE_SEGMENT|2032,2039|false|false|false|||fibroid
Event|Event|SIMPLE_SEGMENT|2058,2059|false|false|false|||b
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2062,2068|false|false|false|C0030797|Pelvis|pelvic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2062,2079|false|false|false|C0729595|Pelvic lymph node group|pelvic lymph node
Finding|Body Substance|SIMPLE_SEGMENT|2069,2074|false|false|false|C0024202|Lymph|lymph
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2069,2079|false|false|false|C0024204|lymph nodes|lymph node
Event|Event|SIMPLE_SEGMENT|2080,2089|false|false|false|||resection
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2080,2089|false|false|false|C0015252;C0728940|Excision;removal technique|resection
Drug|Chemical Viewed Structurally|SIMPLE_SEGMENT|2096,2103|false|false|false|C0302912|Radicals (chemistry)|radical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2096,2114|false|false|false|C0194401|Complete cystectomy|radical cystectomy
Event|Event|SIMPLE_SEGMENT|2104,2114|false|false|false|||cystectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2104,2114|false|false|false|C0010651|Cystectomy|cystectomy
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2119,2127|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Event|Event|SIMPLE_SEGMENT|2128,2139|false|false|false|||vaginectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2128,2139|false|false|false|C0195130|Vaginectomy|vaginectomy
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2145,2152|false|false|false|C0042232|Vagina|vaginal
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|2145,2152|false|false|false|C1272941|Vaginal Dosage Form|vaginal
Finding|Finding|SIMPLE_SEGMENT|2145,2152|false|false|false|C1522570;C4521343|Vaginal (intended site);Vaginal Route of Administration|vaginal
Finding|Functional Concept|SIMPLE_SEGMENT|2145,2152|false|false|false|C1522570;C4521343|Vaginal (intended site);Vaginal Route of Administration|vaginal
Event|Event|SIMPLE_SEGMENT|2154,2168|false|false|false|||reconstruction
Procedure|Machine Activity|SIMPLE_SEGMENT|2154,2168|false|false|false|C0020912;C0524865|Optical Image Reconstruction;Reconstructive Surgical Procedures|reconstruction
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2154,2168|false|false|false|C0020912;C0524865|Optical Image Reconstruction;Reconstructive Surgical Procedures|reconstruction
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2174,2179|false|false|false|C0020885|ileum|ileal
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|2174,2187|false|false|false|C0441253|Structure of ileal conduit|ileal conduit
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2174,2187|false|false|false|C0348002|Ileal conduit procedure|ileal conduit
Event|Activity|SIMPLE_SEGMENT|2188,2196|false|false|false|C1706214|Creation|creation
Event|Event|SIMPLE_SEGMENT|2188,2196|false|false|false|||creation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2188,2196|false|false|false|C0441513|Surgical construction|creation
Event|Event|SIMPLE_SEGMENT|2210,2221|false|false|false|||complicated
Event|Event|SIMPLE_SEGMENT|2225,2235|false|false|false|||bacteremia
Finding|Finding|SIMPLE_SEGMENT|2225,2235|false|false|false|C0004610|Bacteremia|bacteremia
Event|Event|SIMPLE_SEGMENT|2240,2251|true|false|false|||development
Finding|Functional Concept|SIMPLE_SEGMENT|2240,2251|true|false|false|C0018271;C0243107;C0678723;C1527148|Development;Growth and Development function;biological development;development aspects|development
Finding|Organism Function|SIMPLE_SEGMENT|2240,2251|true|false|false|C0018271;C0243107;C0678723;C1527148|Development;Growth and Development function;biological development;development aspects|development
Event|Event|SIMPLE_SEGMENT|2255,2270|true|false|false|||intra-abdominal
Finding|Functional Concept|SIMPLE_SEGMENT|2255,2270|true|false|false|C1512911|Intraabdominal Route of Administration|intra-abdominal
Drug|Substance|SIMPLE_SEGMENT|2272,2277|true|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|2272,2277|true|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|2278,2288|true|false|false|||collection
Finding|Conceptual Entity|SIMPLE_SEGMENT|2278,2288|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|SIMPLE_SEGMENT|2278,2288|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|SIMPLE_SEGMENT|2278,2288|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|SIMPLE_SEGMENT|2278,2288|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Drug|Substance|SIMPLE_SEGMENT|2297,2302|true|false|false|C1550628|Drain - SpecimenType|drain
Finding|Intellectual Product|SIMPLE_SEGMENT|2297,2302|true|false|false|C1546604|Drain Specimen Code|drain
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2297,2312|true|false|false|C3495845|Drain placement|drain placement
Event|Event|SIMPLE_SEGMENT|2303,2312|true|false|false|||placement
Procedure|Health Care Activity|SIMPLE_SEGMENT|2303,2312|true|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2303,2312|true|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Event|Event|SIMPLE_SEGMENT|2330,2331|false|false|false|||/
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2337,2340|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2337,2340|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2337,2340|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Event|Event|SIMPLE_SEGMENT|2337,2340|false|false|false|||DVT
Event|Event|SIMPLE_SEGMENT|2345,2347|false|false|false|||PE
Drug|Organic Chemical|SIMPLE_SEGMENT|2351,2358|false|false|false|C0728963|Lovenox|lovenox
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2351,2358|false|false|false|C0728963|Lovenox|lovenox
Event|Event|SIMPLE_SEGMENT|2351,2358|false|false|false|||lovenox
Finding|Functional Concept|SIMPLE_SEGMENT|2364,2370|false|false|false|C0728831|Social|Social
Finding|Finding|SIMPLE_SEGMENT|2364,2378|false|false|false|C0424945;C3714536|Social History;Social and personal history|Social History
Event|Event|SIMPLE_SEGMENT|2371,2378|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2371,2378|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2371,2378|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2371,2378|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Classification|SIMPLE_SEGMENT|2384,2390|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|SIMPLE_SEGMENT|2384,2390|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|SIMPLE_SEGMENT|2384,2390|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|SIMPLE_SEGMENT|2384,2390|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Finding|SIMPLE_SEGMENT|2384,2398|false|false|false|C0241889|Family Medical History|Family History
Event|Event|SIMPLE_SEGMENT|2391,2398|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2391,2398|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2391,2398|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2391,2398|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Event|Event|SIMPLE_SEGMENT|2400,2408|false|false|false|||Negative
Finding|Classification|SIMPLE_SEGMENT|2400,2408|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|Negative
Finding|Finding|SIMPLE_SEGMENT|2400,2408|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|Negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2400,2408|false|false|false|C5237010|Expression Negative|Negative
Finding|Finding|SIMPLE_SEGMENT|2400,2412|false|false|false|C0205160|Negative|Negative for
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2413,2420|true|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2413,2420|true|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Event|Event|SIMPLE_SEGMENT|2413,2420|true|false|false|||bladder
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2413,2420|true|false|false|C0872388|Procedures on bladder|bladder
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2413,2423|true|true|false|C0005684|Malignant neoplasm of urinary bladder|bladder CA
Event|Event|SIMPLE_SEGMENT|2428,2436|false|false|false|||Physical
Finding|Finding|SIMPLE_SEGMENT|2428,2436|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|2428,2436|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|2428,2436|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|2428,2441|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2428,2441|false|false|false|C0031809|Physical Examination|Physical Exam
Event|Event|SIMPLE_SEGMENT|2437,2441|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|2437,2441|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2437,2441|false|false|false|C0582103|Medical Examination|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2443,2452|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|SIMPLE_SEGMENT|2453,2457|false|false|false|||EXAM
Finding|Functional Concept|SIMPLE_SEGMENT|2453,2457|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|SIMPLE_SEGMENT|2453,2457|false|false|false|C0582103|Medical Examination|EXAM
Drug|Food|SIMPLE_SEGMENT|2476,2481|false|false|false|C1875856|Vital High Nitrogen Enteral Nutrition|Vital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2476,2487|false|false|false|C0488614;C0518766|Vital signs|Vital Signs
Procedure|Health Care Activity|SIMPLE_SEGMENT|2476,2487|false|false|false|C0150404|Taking vital signs|Vital Signs
Event|Event|SIMPLE_SEGMENT|2482,2487|false|false|false|||Signs
Finding|Finding|SIMPLE_SEGMENT|2482,2487|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|Signs
Finding|Functional Concept|SIMPLE_SEGMENT|2482,2487|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|Signs
Event|Event|SIMPLE_SEGMENT|2509,2514|false|false|false|||Lying
Finding|Individual Behavior|SIMPLE_SEGMENT|2509,2514|false|false|false|C0600261|Telling untruths|Lying
Event|Event|SIMPLE_SEGMENT|2530,2537|false|false|false|||General
Finding|Classification|SIMPLE_SEGMENT|2530,2537|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|SIMPLE_SEGMENT|2530,2537|false|false|false|C3812897|General medical service|General
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2539,2544|true|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|2539,2544|true|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2539,2544|true|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|SIMPLE_SEGMENT|2539,2544|true|false|false|||Alert
Finding|Finding|SIMPLE_SEGMENT|2539,2544|true|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|2539,2544|true|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|2539,2544|true|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|SIMPLE_SEGMENT|2546,2554|true|false|false|||oriented
Finding|Intellectual Product|SIMPLE_SEGMENT|2559,2564|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|SIMPLE_SEGMENT|2565,2573|true|false|false|||distress
Finding|Finding|SIMPLE_SEGMENT|2565,2573|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|SIMPLE_SEGMENT|2565,2573|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2577,2582|true|false|false|C1512338|HEENT|HEENT
Event|Event|SIMPLE_SEGMENT|2592,2601|false|false|false|||anicteric
Finding|Finding|SIMPLE_SEGMENT|2592,2601|false|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2603,2606|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2603,2606|false|false|false|C0026987|Myelofibrosis|MMM
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2608,2618|false|false|false|C0521367|Oropharyngeal|oropharynx
Event|Event|SIMPLE_SEGMENT|2619,2624|false|false|false|||clear
Finding|Idea or Concept|SIMPLE_SEGMENT|2619,2624|false|false|false|C1550016|Remote control command - Clear|clear
Event|Event|SIMPLE_SEGMENT|2632,2635|false|false|false|||RRR
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|2651,2659|true|false|false|C0039155|Systole|systolic
Finding|Finding|SIMPLE_SEGMENT|2651,2666|true|false|false|C0232257|Systolic Murmurs|systolic murmur
Finding|Finding|SIMPLE_SEGMENT|2660,2666|true|false|false|C0018808|Heart murmur|murmur
Event|Event|SIMPLE_SEGMENT|2667,2671|true|false|false|||RUBS
Finding|Finding|SIMPLE_SEGMENT|2667,2671|true|false|false|C0232267|Pericardial friction rub|RUBS
Event|Event|SIMPLE_SEGMENT|2676,2680|true|false|false|||rubs
Finding|Finding|SIMPLE_SEGMENT|2676,2680|true|false|false|C0232267|Pericardial friction rub|rubs
Event|Event|SIMPLE_SEGMENT|2682,2689|true|false|false|||gallops
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2693,2698|true|false|false|C0024109|Lung|Lungs
Event|Event|SIMPLE_SEGMENT|2700,2705|true|false|false|||Clear
Finding|Idea or Concept|SIMPLE_SEGMENT|2700,2705|true|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|SIMPLE_SEGMENT|2709,2721|true|false|false|||auscultation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2709,2721|true|false|false|C0004339|Auscultation|auscultation
Event|Event|SIMPLE_SEGMENT|2738,2745|true|false|false|||wheezes
Finding|Sign or Symptom|SIMPLE_SEGMENT|2738,2745|true|false|false|C0043144|Wheezing|wheezes
Event|Event|SIMPLE_SEGMENT|2747,2752|true|false|false|||rales
Finding|Finding|SIMPLE_SEGMENT|2747,2752|true|false|false|C0034642;C0240859|Basilar Rales;Rales|rales
Event|Event|SIMPLE_SEGMENT|2755,2762|true|false|false|||rhonchi
Finding|Finding|SIMPLE_SEGMENT|2755,2762|true|false|false|C0035508|Rhonchi|rhonchi
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2766,2773|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2766,2773|false|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Event|Event|SIMPLE_SEGMENT|2766,2773|false|false|false|||Abdomen
Finding|Finding|SIMPLE_SEGMENT|2766,2773|false|false|false|C0941288|Abdomen problem|Abdomen
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2775,2779|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Event|Event|SIMPLE_SEGMENT|2775,2779|false|false|false|||Soft
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2808,2813|false|false|false|C0021853|Intestines|bowel
Finding|Finding|SIMPLE_SEGMENT|2808,2820|false|false|false|C0232693|Bowel sounds|bowel sounds
Event|Event|SIMPLE_SEGMENT|2814,2820|false|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|2814,2820|false|false|false|C0037709||sounds
Finding|Finding|SIMPLE_SEGMENT|2821,2828|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|SIMPLE_SEGMENT|2821,2828|false|false|false|C0150312;C0449450|Present;Presentation|present
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2832,2837|false|false|false|C0020885|ileum|ileal
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|2832,2845|false|false|false|C0441253|Structure of ileal conduit|ileal conduit
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2832,2845|false|false|false|C0348002|Ileal conduit procedure|ileal conduit
Event|Event|SIMPLE_SEGMENT|2838,2845|false|false|false|||conduit
Drug|Substance|SIMPLE_SEGMENT|2846,2851|false|false|false|C1550628|Drain - SpecimenType|drain
Event|Event|SIMPLE_SEGMENT|2846,2851|false|false|false|||drain
Finding|Intellectual Product|SIMPLE_SEGMENT|2846,2851|false|false|false|C1546604|Drain Specimen Code|drain
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2855,2858|false|false|false|C0230178|Structure of right lower quadrant of abdomen|RLQ
Drug|Substance|SIMPLE_SEGMENT|2873,2878|false|false|false|C1550628|Drain - SpecimenType|drain
Event|Event|SIMPLE_SEGMENT|2873,2878|false|false|false|||drain
Finding|Intellectual Product|SIMPLE_SEGMENT|2873,2878|false|false|false|C1546604|Drain Specimen Code|drain
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2882,2885|false|false|false|C0230180|Structure of left lower quadrant of abdomen|LLQ
Finding|Gene or Genome|SIMPLE_SEGMENT|2901,2905|false|false|false|C1864650|GNAS-AS1 gene|sang
Drug|Substance|SIMPLE_SEGMENT|2906,2911|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|2906,2911|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|2906,2911|false|false|false|C1546638|Fluid Specimen Code|fluid
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|2931,2934|true|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Event|Event|SIMPLE_SEGMENT|2931,2934|true|false|false|||Ext
Finding|Gene or Genome|SIMPLE_SEGMENT|2931,2934|true|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Event|Event|SIMPLE_SEGMENT|2936,2940|false|false|false|||Warm
Finding|Finding|SIMPLE_SEGMENT|2936,2940|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|2936,2940|false|false|false|C0687712|warming process|Warm
Finding|Finding|SIMPLE_SEGMENT|2942,2946|false|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|2947,2955|false|false|false|||perfused
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2971,2976|false|false|false|C1717255||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|2971,2976|false|false|false|C0013604|Edema|edema
Event|Event|SIMPLE_SEGMENT|2977,2980|false|false|false|||LLE
Finding|Gene or Genome|SIMPLE_SEGMENT|2991,2994|false|false|false|C1539110|CNDP2 gene|CN2
Event|Event|SIMPLE_SEGMENT|3006,3012|false|false|false|||intact
Finding|Finding|SIMPLE_SEGMENT|3006,3012|false|false|false|C1554187|Gender Status - Intact|intact
Event|Event|SIMPLE_SEGMENT|3014,3020|false|false|false|||moving
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3021,3036|false|false|false|C0278454|All extremities|all extremities
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3025,3036|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Finding|Body Substance|SIMPLE_SEGMENT|3053,3062|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|3053,3062|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|3053,3062|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|3053,3062|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|SIMPLE_SEGMENT|3063,3067|false|false|false|||EXAM
Finding|Functional Concept|SIMPLE_SEGMENT|3063,3067|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|SIMPLE_SEGMENT|3063,3067|false|false|false|C0582103|Medical Examination|EXAM
Drug|Food|SIMPLE_SEGMENT|3087,3092|false|false|false|C1875856|Vital High Nitrogen Enteral Nutrition|Vital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3087,3098|false|false|false|C0488614;C0518766|Vital signs|Vital signs
Procedure|Health Care Activity|SIMPLE_SEGMENT|3087,3098|false|false|false|C0150404|Taking vital signs|Vital signs
Event|Event|SIMPLE_SEGMENT|3093,3098|false|false|false|||signs
Finding|Finding|SIMPLE_SEGMENT|3093,3098|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|SIMPLE_SEGMENT|3093,3098|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Event|Event|SIMPLE_SEGMENT|3130,3137|false|false|false|||General
Finding|Classification|SIMPLE_SEGMENT|3130,3137|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|SIMPLE_SEGMENT|3130,3137|false|false|false|C3812897|General medical service|General
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3147,3152|false|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3154,3160|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3154,3160|false|false|false|C0036412|Scleral Diseases|Sclera
Event|Event|SIMPLE_SEGMENT|3154,3160|false|false|false|||Sclera
Procedure|Health Care Activity|SIMPLE_SEGMENT|3154,3160|false|false|false|C2228481|examination of sclera|Sclera
Event|Event|SIMPLE_SEGMENT|3161,3170|false|false|false|||anicteric
Finding|Finding|SIMPLE_SEGMENT|3161,3170|false|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3172,3176|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Anatomy|Cell Component|SIMPLE_SEGMENT|3172,3176|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Finding|Finding|SIMPLE_SEGMENT|3172,3176|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|Neck
Finding|Functional Concept|SIMPLE_SEGMENT|3178,3184|false|false|false|C0332254|Supple|supple
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3187,3192|false|false|false|C0024109|Lung|Lungs
Event|Event|SIMPLE_SEGMENT|3194,3199|true|false|false|||Clear
Finding|Idea or Concept|SIMPLE_SEGMENT|3194,3199|true|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|SIMPLE_SEGMENT|3203,3215|true|false|false|||auscultation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3203,3215|true|false|false|C0004339|Auscultation|auscultation
Event|Event|SIMPLE_SEGMENT|3232,3239|true|false|false|||wheezes
Finding|Sign or Symptom|SIMPLE_SEGMENT|3232,3239|true|false|false|C0043144|Wheezing|wheezes
Event|Event|SIMPLE_SEGMENT|3241,3246|true|false|false|||rales
Finding|Finding|SIMPLE_SEGMENT|3241,3246|true|false|false|C0034642;C0240859|Basilar Rales;Rales|rales
Event|Event|SIMPLE_SEGMENT|3249,3256|true|false|false|||rhonchi
Finding|Finding|SIMPLE_SEGMENT|3249,3256|true|false|false|C0035508|Rhonchi|rhonchi
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3260,3268|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Event|Event|SIMPLE_SEGMENT|3269,3281|false|false|false|||auscultation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3269,3281|false|false|false|C0004339|Auscultation|auscultation
Event|Activity|SIMPLE_SEGMENT|3296,3300|false|false|false|C0871208|Rating (action)|rate
Event|Event|SIMPLE_SEGMENT|3296,3300|false|false|false|||rate
Finding|Idea or Concept|SIMPLE_SEGMENT|3296,3300|false|false|false|C1549480|Amount type - Rate|rate
Event|Event|SIMPLE_SEGMENT|3305,3311|false|false|false|||rhythm
Finding|Finding|SIMPLE_SEGMENT|3305,3311|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|SIMPLE_SEGMENT|3305,3311|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Event|Event|SIMPLE_SEGMENT|3336,3339|false|false|false|||SEM
Finding|Finding|SIMPLE_SEGMENT|3336,3339|false|false|false|C0694547|SYSTOLIC EJECTION MURMUR|SEM
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3341,3348|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3341,3348|false|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Event|Event|SIMPLE_SEGMENT|3341,3348|false|false|false|||Abdomen
Finding|Finding|SIMPLE_SEGMENT|3341,3348|false|false|false|C0941288|Abdomen problem|Abdomen
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3355,3360|false|false|false|C0020885|ileum|ileal
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|3355,3368|false|false|false|C0441253|Structure of ileal conduit|ileal conduit
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3355,3368|false|false|false|C0348002|Ileal conduit procedure|ileal conduit
Event|Event|SIMPLE_SEGMENT|3378,3383|false|false|false|||clear
Finding|Idea or Concept|SIMPLE_SEGMENT|3378,3383|false|false|false|C1550016|Remote control command - Clear|clear
Event|Event|SIMPLE_SEGMENT|3391,3396|false|false|false|||urine
Finding|Body Substance|SIMPLE_SEGMENT|3391,3396|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Functional Concept|SIMPLE_SEGMENT|3391,3396|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Intellectual Product|SIMPLE_SEGMENT|3391,3396|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3408,3411|false|false|false|C0230180|Structure of left lower quadrant of abdomen|LLQ
Drug|Substance|SIMPLE_SEGMENT|3412,3417|false|false|false|C1550628|Drain - SpecimenType|drain
Event|Event|SIMPLE_SEGMENT|3412,3417|false|false|false|||drain
Finding|Intellectual Product|SIMPLE_SEGMENT|3412,3417|false|false|false|C1546604|Drain Specimen Code|drain
Event|Activity|SIMPLE_SEGMENT|3421,3426|false|false|false|C1882509|put - instruction imperative|place
Finding|Functional Concept|SIMPLE_SEGMENT|3421,3426|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|SIMPLE_SEGMENT|3421,3426|false|false|false|C1533810||place
Finding|Body Substance|SIMPLE_SEGMENT|3436,3456|false|false|false|C4518404|Serosanguinous fluid|serosanguinous fluid
Drug|Substance|SIMPLE_SEGMENT|3451,3456|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|3451,3456|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|3451,3456|false|false|false|C1546638|Fluid Specimen Code|fluid
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|3460,3463|false|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Event|Event|SIMPLE_SEGMENT|3460,3463|false|false|false|||Ext
Finding|Gene or Genome|SIMPLE_SEGMENT|3460,3463|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Event|Event|SIMPLE_SEGMENT|3465,3469|false|false|false|||Warm
Finding|Finding|SIMPLE_SEGMENT|3465,3469|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3465,3469|false|false|false|C0687712|warming process|Warm
Finding|Finding|SIMPLE_SEGMENT|3471,3475|true|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|3476,3484|true|false|false|||perfused
Drug|Food|SIMPLE_SEGMENT|3489,3495|true|false|false|C5890763||pulses
Event|Event|SIMPLE_SEGMENT|3489,3495|true|false|false|||pulses
Finding|Physiologic Function|SIMPLE_SEGMENT|3489,3495|true|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|SIMPLE_SEGMENT|3489,3495|true|false|false|C0034107|Pulse taking|pulses
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|3500,3508|true|false|false|C0149651|Clubbing|clubbing
Event|Event|SIMPLE_SEGMENT|3500,3508|true|false|false|||clubbing
Event|Event|SIMPLE_SEGMENT|3510,3518|true|false|false|||cyanosis
Finding|Sign or Symptom|SIMPLE_SEGMENT|3510,3518|true|false|false|C0010520|Cyanosis|cyanosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3523,3528|true|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|3523,3528|true|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|3523,3528|true|false|false|C0013604|Edema|edema
Procedure|Health Care Activity|SIMPLE_SEGMENT|3552,3561|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|SIMPLE_SEGMENT|3562,3566|false|false|false|||LABS
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3562,3566|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3596,3601|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3596,3601|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3596,3601|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|3602,3605|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|3613,3616|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3613,3616|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3613,3616|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3623,3626|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3623,3626|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|3623,3626|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3623,3626|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3632,3635|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3632,3635|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|3643,3646|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|3643,3646|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3643,3646|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3643,3646|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3643,3646|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|3650,3653|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3650,3653|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|3650,3653|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|3650,3653|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|3650,3653|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3650,3653|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|SIMPLE_SEGMENT|3659,3663|false|false|false|||MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3659,3663|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3691,3694|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3711,3716|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3711,3716|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3711,3716|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3729,3735|false|false|false|C0024202|Lymph|Lymphs
Drug|Antibiotic|SIMPLE_SEGMENT|3741,3746|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3741,3746|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|SIMPLE_SEGMENT|3741,3746|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3752,3755|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|Eos
Event|Event|SIMPLE_SEGMENT|3752,3755|false|false|false|||Eos
Finding|Gene or Genome|SIMPLE_SEGMENT|3752,3755|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|Eos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3859,3864|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3859,3864|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3859,3864|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3869,3872|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|SIMPLE_SEGMENT|3869,3872|false|false|false|||PTT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3869,3872|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3894,3899|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3894,3899|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3894,3899|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3900,3903|false|false|false|C0389252|RET protein, human|Ret
Finding|Gene or Genome|SIMPLE_SEGMENT|3900,3903|false|false|false|C0389252;C0694890;C0813143;C1704885|Oncogene RET;RET gene;RET protein, human;RET wt Allele|Ret
Finding|Receptor|SIMPLE_SEGMENT|3900,3903|false|false|false|C0389252;C0694890;C0813143;C1704885|Oncogene RET;RET gene;RET protein, human;RET wt Allele|Ret
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|3913,3916|false|false|false|C0002636;C0220724|Amniotic Band Syndrome;CONSTRICTING BANDS, CONGENITAL|Abs
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3913,3916|false|false|false|C0002636;C0220724|Amniotic Band Syndrome;CONSTRICTING BANDS, CONGENITAL|Abs
Finding|Gene or Genome|SIMPLE_SEGMENT|3913,3916|false|false|false|C1425698;C4723885|DDX41 gene;DDX41 wt Allele|Abs
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3917,3920|false|false|false|C0389252|RET protein, human|Ret
Finding|Gene or Genome|SIMPLE_SEGMENT|3917,3920|false|false|false|C0389252;C0694890;C0813143;C1704885|Oncogene RET;RET gene;RET protein, human;RET wt Allele|Ret
Finding|Receptor|SIMPLE_SEGMENT|3917,3920|false|false|false|C0389252;C0694890;C0813143;C1704885|Oncogene RET;RET gene;RET protein, human;RET wt Allele|Ret
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3938,3943|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3938,3943|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3938,3943|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|3938,3951|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3938,3951|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3938,3951|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3944,3951|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|3944,3951|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3944,3951|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|3944,3951|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3944,3951|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3944,3951|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|SIMPLE_SEGMENT|3997,4001|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3997,4001|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3997,4001|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4026,4031|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4026,4031|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4026,4031|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4032,4035|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4032,4035|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|SIMPLE_SEGMENT|4032,4035|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|SIMPLE_SEGMENT|4032,4035|false|false|false|||ALT
Finding|Gene or Genome|SIMPLE_SEGMENT|4032,4035|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|SIMPLE_SEGMENT|4032,4035|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|SIMPLE_SEGMENT|4032,4035|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4032,4035|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4038,4041|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4038,4041|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4038,4041|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4038,4041|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|SIMPLE_SEGMENT|4038,4041|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|SIMPLE_SEGMENT|4038,4041|false|false|false|||AST
Finding|Gene or Genome|SIMPLE_SEGMENT|4038,4041|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4044,4051|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|SIMPLE_SEGMENT|4044,4051|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Event|Event|SIMPLE_SEGMENT|4044,4051|false|false|false|||AlkPhos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4079,4084|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4079,4084|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4079,4084|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4085,4091|false|false|false|C0023764|lipase|Lipase
Drug|Enzyme|SIMPLE_SEGMENT|4085,4091|false|false|false|C0023764|lipase|Lipase
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4085,4091|false|false|false|C0023764|lipase|Lipase
Event|Event|SIMPLE_SEGMENT|4085,4091|false|false|false|||Lipase
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4085,4091|false|false|false|C0373670|Lipase measurement|Lipase
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4106,4111|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4106,4111|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4106,4111|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4106,4119|false|false|false|C0853248|Blood albumin|BLOOD Albumin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4112,4119|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4112,4119|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4112,4119|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Event|Event|SIMPLE_SEGMENT|4112,4119|false|false|false|||Albumin
Finding|Gene or Genome|SIMPLE_SEGMENT|4112,4119|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Finding|Physiologic Function|SIMPLE_SEGMENT|4112,4119|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4112,4119|false|false|false|C0201838|Albumin measurement|Albumin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4125,4129|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4125,4129|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4125,4129|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4125,4129|false|false|false|C0337439|Iron measurement|Iron
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4145,4150|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4145,4150|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4145,4150|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4189,4192|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4189,4192|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Drug|Hormone|SIMPLE_SEGMENT|4189,4192|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4189,4192|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Event|Event|SIMPLE_SEGMENT|4189,4192|false|false|false|||TRF
Finding|Gene or Genome|SIMPLE_SEGMENT|4189,4192|false|false|false|C1334121;C1336604;C1705002|IL5 gene;TERF1 gene;TERF1 wt Allele|TRF
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4210,4215|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4210,4215|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4210,4215|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4210,4223|false|false|false|C3824990|lactate in blood (lab test)|BLOOD Lactate
Drug|Organic Chemical|SIMPLE_SEGMENT|4216,4223|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4216,4223|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Event|Event|SIMPLE_SEGMENT|4216,4223|false|false|false|||Lactate
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4216,4223|false|false|false|C0202115|Lactic acid measurement|Lactate
Finding|Body Substance|SIMPLE_SEGMENT|4229,4238|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|4229,4238|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|4229,4238|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|4229,4238|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|SIMPLE_SEGMENT|4239,4243|false|false|false|||LABS
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4239,4243|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4273,4278|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4273,4278|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4273,4278|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|4279,4282|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|4287,4290|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4287,4290|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4287,4290|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4297,4300|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4297,4300|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|4297,4300|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4297,4300|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4306,4309|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4306,4309|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|4317,4320|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|4317,4320|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4317,4320|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4317,4320|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4317,4320|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|4324,4327|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4324,4327|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|4324,4327|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|4324,4327|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|4324,4327|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4324,4327|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|SIMPLE_SEGMENT|4333,4337|false|false|false|||MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4333,4337|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4365,4368|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4385,4390|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4385,4390|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4385,4390|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4395,4398|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|SIMPLE_SEGMENT|4395,4398|false|false|false|||PTT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4395,4398|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4420,4425|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4420,4425|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4426,4429|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4446,4451|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4446,4451|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4446,4451|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|4446,4459|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4446,4459|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4446,4459|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4452,4459|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|4452,4459|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4452,4459|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|4452,4459|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4452,4459|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4452,4459|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4502,4506|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4502,4506|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4502,4506|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4531,4536|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4531,4536|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4531,4536|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4531,4544|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4537,4544|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4537,4544|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4537,4544|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4537,4544|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|4537,4544|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|SIMPLE_SEGMENT|4537,4544|false|false|false|||Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|4537,4544|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4537,4544|false|false|false|C0201925|Calcium measurement|Calcium
Event|Event|SIMPLE_SEGMENT|4547,4548|false|false|false|||5
Event|Event|SIMPLE_SEGMENT|4567,4579|false|false|false|||MICROBIOLOGY
Finding|Functional Concept|SIMPLE_SEGMENT|4567,4579|false|false|false|C0025953;C1571921;C4049106|Microbiological;Microbiology - Laboratory Class;Microbiology Diagnostic Service Section ID|MICROBIOLOGY
Finding|Intellectual Product|SIMPLE_SEGMENT|4567,4579|false|false|false|C0025953;C1571921;C4049106|Microbiological;Microbiology - Laboratory Class;Microbiology Diagnostic Service Section ID|MICROBIOLOGY
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4567,4579|false|false|false|C0085672|Microbiology procedure|MICROBIOLOGY
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4595,4600|false|false|false|C0851353|Blood and lymphatic system disorders|Blood
Event|Event|SIMPLE_SEGMENT|4595,4600|false|false|false|||Blood
Finding|Body Substance|SIMPLE_SEGMENT|4595,4600|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4595,4609|false|true|false|C0200949|Blood culture|Blood cultures
Event|Event|SIMPLE_SEGMENT|4601,4609|false|false|false|||cultures
Finding|Idea or Concept|SIMPLE_SEGMENT|4601,4609|false|false|false|C0010453|Culture (Anthropological)|cultures
Event|Event|SIMPLE_SEGMENT|4613,4620|false|false|false|||pending
Finding|Idea or Concept|SIMPLE_SEGMENT|4613,4620|false|false|false|C1691786;C1704475|Pending - Allergy Clinical Status;Pending - referral status|pending
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4634,4640|false|false|false|C0030797|Pelvis|pelvic
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|4641,4651|false|false|false|C1720922|Respiratory Aspiration|aspiration
Event|Event|SIMPLE_SEGMENT|4641,4651|false|false|false|||aspiration
Finding|Finding|SIMPLE_SEGMENT|4641,4651|false|false|false|C0220787;C0700198;C2712334|Aspiration into respiratory tract;Endotracheal aspiration;Pulmonary aspiration|aspiration
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|4641,4651|false|false|false|C0220787;C0700198;C2712334|Aspiration into respiratory tract;Endotracheal aspiration;Pulmonary aspiration|aspiration
Finding|Pathologic Function|SIMPLE_SEGMENT|4641,4651|false|false|false|C0220787;C0700198;C2712334|Aspiration into respiratory tract;Endotracheal aspiration;Pulmonary aspiration|aspiration
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4641,4651|false|false|false|C0349707||aspiration
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|4655,4665|false|false|false|C0061856|Gram's stain|GRAM STAIN
Drug|Organic Chemical|SIMPLE_SEGMENT|4655,4665|false|false|false|C0061856|Gram's stain|GRAM STAIN
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4655,4665|false|false|false|C0200966|Bacterial stain, routine|GRAM STAIN
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|4660,4665|false|false|false|C0038128|Stains|STAIN
Event|Event|SIMPLE_SEGMENT|4660,4665|false|false|false|||STAIN
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4660,4665|false|false|false|C0487602|Staining method|STAIN
Finding|Idea or Concept|SIMPLE_SEGMENT|4667,4672|false|false|false|C1546485|Diagnosis Type - Final|Final
Event|Event|SIMPLE_SEGMENT|4705,4710|false|false|false|||FIELD
Finding|Conceptual Entity|SIMPLE_SEGMENT|4705,4710|false|false|false|C1521738;C2346620;C2349184|Field;Force Field;Knowledge Field|FIELD
Procedure|Health Care Activity|SIMPLE_SEGMENT|4705,4710|false|false|false|C1553496|field - patient encounter|FIELD
Event|Event|SIMPLE_SEGMENT|4715,4732|false|false|false|||POLYMORPHONUCLEAR
Anatomy|Cell|SIMPLE_SEGMENT|4734,4744|false|false|false|C0023516|Leukocytes|LEUKOCYTES
Event|Event|SIMPLE_SEGMENT|4734,4744|false|false|false|||LEUKOCYTES
Finding|Body Substance|SIMPLE_SEGMENT|4734,4744|false|false|false|C1547962;C1550647|Specimen Type - Leukocytes|LEUKOCYTES
Finding|Intellectual Product|SIMPLE_SEGMENT|4734,4744|false|false|false|C1547962;C1550647|Specimen Type - Leukocytes|LEUKOCYTES
Finding|Finding|SIMPLE_SEGMENT|4756,4775|true|false|false|C2924473|Microorganisms seen|MICROORGANISMS SEEN
Event|Event|SIMPLE_SEGMENT|4771,4775|true|false|false|||SEEN
Drug|Substance|SIMPLE_SEGMENT|4781,4786|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|FLUID
Event|Event|SIMPLE_SEGMENT|4781,4786|false|false|false|||FLUID
Finding|Intellectual Product|SIMPLE_SEGMENT|4781,4786|false|false|false|C1546638|Fluid Specimen Code|FLUID
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4787,4794|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|SIMPLE_SEGMENT|4787,4794|false|false|false|||CULTURE
Finding|Functional Concept|SIMPLE_SEGMENT|4787,4794|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|SIMPLE_SEGMENT|4787,4794|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4787,4794|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Event|Event|SIMPLE_SEGMENT|4796,4801|false|false|false|||Final
Finding|Idea or Concept|SIMPLE_SEGMENT|4796,4801|false|false|false|C1546485|Diagnosis Type - Final|Final
Event|Event|SIMPLE_SEGMENT|4813,4819|true|false|false|||GROWTH
Finding|Finding|SIMPLE_SEGMENT|4813,4819|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|4813,4819|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organism Function|SIMPLE_SEGMENT|4813,4819|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Physiologic Function|SIMPLE_SEGMENT|4813,4819|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|4813,4819|true|false|false|C2911660|Growth action|GROWTH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4825,4842|false|false|false|C1273935|Anaerobic microbial culture|ANAEROBIC CULTURE
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4835,4842|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|SIMPLE_SEGMENT|4835,4842|false|false|false|||CULTURE
Finding|Functional Concept|SIMPLE_SEGMENT|4835,4842|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|SIMPLE_SEGMENT|4835,4842|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4835,4842|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Event|Event|SIMPLE_SEGMENT|4864,4870|true|false|false|||GROWTH
Finding|Finding|SIMPLE_SEGMENT|4864,4870|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|4864,4870|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organism Function|SIMPLE_SEGMENT|4864,4870|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Physiologic Function|SIMPLE_SEGMENT|4864,4870|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|4864,4870|true|false|false|C2911660|Growth action|GROWTH
Event|Event|SIMPLE_SEGMENT|4884,4891|false|false|false|||IMAGING
Finding|Finding|SIMPLE_SEGMENT|4884,4891|false|false|false|C0740845|Imaging problem|IMAGING
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4884,4891|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|IMAGING
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4912,4918|false|false|false|C1644645||CT ABD
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4915,4918|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|ABD
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|4915,4918|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|ABD
Event|Event|SIMPLE_SEGMENT|4915,4918|false|false|false|||ABD
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4919,4922|false|false|false|C0449203|PEL (body structure)|PEL
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4919,4922|false|false|false|C1292753;C1394210;C4520841|Pel crisis;Primary Effusion Lymphoma;Pure Erythroid Leukemia|PEL
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4919,4922|false|false|false|C1292753;C1394210;C4520841|Pel crisis;Primary Effusion Lymphoma;Pure Erythroid Leukemia|PEL
Event|Event|SIMPLE_SEGMENT|4923,4924|false|false|false|||W
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|4926,4934|false|false|false|C0009924|Contrast Media|CONTRAST
Event|Event|SIMPLE_SEGMENT|4926,4934|false|false|false|||CONTRAST
Finding|Intellectual Product|SIMPLE_SEGMENT|4943,4951|false|false|false|C1552654|Parameterized Data Type - Interval|Interval
Event|Event|SIMPLE_SEGMENT|4952,4960|false|false|false|||decrease
Finding|Finding|SIMPLE_SEGMENT|4952,4960|false|false|false|C0392756|Reduced|decrease
Finding|Functional Concept|SIMPLE_SEGMENT|4976,4981|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Drug|Substance|SIMPLE_SEGMENT|4993,4998|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|4993,4998|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|4993,4998|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|5000,5010|false|false|false|||collection
Finding|Conceptual Entity|SIMPLE_SEGMENT|5000,5010|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|SIMPLE_SEGMENT|5000,5010|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|SIMPLE_SEGMENT|5000,5010|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|SIMPLE_SEGMENT|5000,5010|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5077,5085|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Finding|Functional Concept|SIMPLE_SEGMENT|5086,5094|false|false|false|C5445118|Approach (contact)|approach
Event|Event|SIMPLE_SEGMENT|5103,5111|false|false|false|||catheter
Finding|Intellectual Product|SIMPLE_SEGMENT|5103,5111|false|false|false|C1546572||catheter
Finding|Finding|SIMPLE_SEGMENT|5112,5121|false|false|false|C0442739||unchanged
Event|Event|SIMPLE_SEGMENT|5126,5134|false|false|false|||position
Event|Event|SIMPLE_SEGMENT|5158,5165|false|false|false|||located
Event|Event|SIMPLE_SEGMENT|5185,5195|false|false|false|||collection
Finding|Conceptual Entity|SIMPLE_SEGMENT|5185,5195|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|SIMPLE_SEGMENT|5185,5195|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|SIMPLE_SEGMENT|5185,5195|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|SIMPLE_SEGMENT|5185,5195|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|SIMPLE_SEGMENT|5229,5237|false|false|false|C1552654|Parameterized Data Type - Interval|Interval
Event|Event|SIMPLE_SEGMENT|5238,5246|false|false|false|||increase
Finding|Functional Concept|SIMPLE_SEGMENT|5238,5246|false|false|false|C0442805|Increase|increase
Finding|Finding|SIMPLE_SEGMENT|5238,5254|false|false|false|C1268652|increase in size|increase in size
Finding|Functional Concept|SIMPLE_SEGMENT|5262,5266|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5267,5273|false|false|false|C0030797|Pelvis|pelvic
Drug|Substance|SIMPLE_SEGMENT|5274,5279|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|5274,5279|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|5274,5279|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|5281,5291|false|false|false|||collection
Finding|Conceptual Entity|SIMPLE_SEGMENT|5281,5291|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|SIMPLE_SEGMENT|5281,5291|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|SIMPLE_SEGMENT|5281,5291|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|SIMPLE_SEGMENT|5281,5291|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Event|Event|SIMPLE_SEGMENT|5298,5307|false|false|false|||measuring
Event|Event|SIMPLE_SEGMENT|5367,5376|false|false|false|||Increased
Event|Activity|SIMPLE_SEGMENT|5388,5399|false|false|false|C2349975|Enhance (action)|enhancement
Event|Event|SIMPLE_SEGMENT|5388,5399|false|false|false|||enhancement
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5388,5399|false|false|false|C1627358|Refractive surgery enhancement|enhancement
Event|Event|SIMPLE_SEGMENT|5404,5411|false|false|false|||suggest
Event|Event|SIMPLE_SEGMENT|5412,5424|false|false|false|||superimposed
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5426,5435|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|SIMPLE_SEGMENT|5426,5435|false|false|false|||infection
Finding|Pathologic Function|SIMPLE_SEGMENT|5426,5435|false|false|false|C3714514|Infection|infection
Finding|Finding|SIMPLE_SEGMENT|5444,5447|true|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|5444,5447|true|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Drug|Substance|SIMPLE_SEGMENT|5448,5453|true|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|5448,5453|true|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|5448,5453|true|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|5454,5464|true|false|false|||collection
Finding|Conceptual Entity|SIMPLE_SEGMENT|5454,5464|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|SIMPLE_SEGMENT|5454,5464|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|SIMPLE_SEGMENT|5454,5464|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|SIMPLE_SEGMENT|5454,5464|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Event|Event|SIMPLE_SEGMENT|5465,5475|true|false|false|||identified
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5481,5484|false|false|false|C3813556|Cancer/Testis Antigen|CTA
Event|Event|SIMPLE_SEGMENT|5481,5484|false|false|false|||CTA
Finding|Gene or Genome|SIMPLE_SEGMENT|5481,5484|false|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5481,5484|false|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5485,5488|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|ABD
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|5485,5488|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|ABD
Event|Event|SIMPLE_SEGMENT|5485,5488|false|false|false|||ABD
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5491,5497|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|PELVIS
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5491,5497|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|PELVIS
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5491,5497|false|false|false|C0153663|Malignant neoplasm of pelvis|PELVIS
Event|Event|SIMPLE_SEGMENT|5491,5497|false|false|false|||PELVIS
Finding|Finding|SIMPLE_SEGMENT|5491,5497|false|false|false|C0812455|Pelvis problem|PELVIS
Event|Event|SIMPLE_SEGMENT|5505,5513|false|false|false|||Decrease
Finding|Finding|SIMPLE_SEGMENT|5505,5513|false|false|false|C0392756|Reduced|Decrease
Finding|Functional Concept|SIMPLE_SEGMENT|5525,5530|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5525,5545|false|false|false|C0230178|Structure of right lower quadrant of abdomen|right lower quadrant
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5531,5536|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|5531,5536|false|false|false|C2003888|Lower (action)|lower
Drug|Substance|SIMPLE_SEGMENT|5546,5551|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|5546,5551|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|5552,5562|false|false|false|||collection
Finding|Conceptual Entity|SIMPLE_SEGMENT|5552,5562|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|SIMPLE_SEGMENT|5552,5562|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|SIMPLE_SEGMENT|5552,5562|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|SIMPLE_SEGMENT|5552,5562|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|SIMPLE_SEGMENT|5574,5586|false|false|false|C1522243|Percutaneous Route of Drug Administration|percutaneous
Drug|Substance|SIMPLE_SEGMENT|5587,5592|false|false|false|C1550628|Drain - SpecimenType|drain
Event|Event|SIMPLE_SEGMENT|5587,5592|false|false|false|||drain
Finding|Intellectual Product|SIMPLE_SEGMENT|5587,5592|false|false|false|C1546604|Drain Specimen Code|drain
Finding|Finding|SIMPLE_SEGMENT|5618,5622|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|SIMPLE_SEGMENT|5618,5622|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|SIMPLE_SEGMENT|5618,5622|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Event|Activity|SIMPLE_SEGMENT|5623,5634|false|false|false|C0599946|Attenuation|attenuation
Event|Event|SIMPLE_SEGMENT|5651,5655|false|false|false|||exam
Finding|Functional Concept|SIMPLE_SEGMENT|5651,5655|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|5651,5655|false|false|false|C0582103|Medical Examination|exam
Event|Event|SIMPLE_SEGMENT|5656,5666|false|false|false|||consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|5656,5666|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|5656,5671|false|false|false|C0332290|Consistent with|consistent with
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5672,5677|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|5672,5677|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|5672,5677|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5672,5686|false|false|false|C0456388|Blood product|blood products
Event|Event|SIMPLE_SEGMENT|5678,5686|false|false|false|||products
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5704,5713|false|false|false|C0020452|Hyperemia|hyperemia
Event|Event|SIMPLE_SEGMENT|5704,5713|false|false|false|||hyperemia
Finding|Finding|SIMPLE_SEGMENT|5723,5729|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|5723,5729|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Finding|SIMPLE_SEGMENT|5723,5742|false|false|false|C4050249|Likely Inflammatory Activity|likely inflammatory
Event|Event|SIMPLE_SEGMENT|5730,5742|false|false|false|||inflammatory
Finding|Functional Concept|SIMPLE_SEGMENT|5730,5742|false|true|false|C0333348|Inflammatory|inflammatory
Event|Event|SIMPLE_SEGMENT|5756,5764|true|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|5756,5764|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|5756,5767|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|5769,5777|true|false|false|C0009924|Contrast Media|contrast
Event|Event|SIMPLE_SEGMENT|5769,5777|true|false|false|||contrast
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|5778,5791|true|false|false|C0015379|Extravasation of Diagnostic and Therapeutic Materials|extravasation
Event|Event|SIMPLE_SEGMENT|5778,5791|true|false|false|||extravasation
Finding|Pathologic Function|SIMPLE_SEGMENT|5778,5791|true|false|false|C0015376|Extravasation|extravasation
Finding|Gene or Genome|SIMPLE_SEGMENT|5806,5811|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Finding|Intellectual Product|SIMPLE_SEGMENT|5812,5818|false|false|false|C1547311|Patient Condition Code - Stable|stable
Drug|Substance|SIMPLE_SEGMENT|5819,5824|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|5819,5824|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|5819,5824|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|5825,5835|false|false|false|||collection
Finding|Conceptual Entity|SIMPLE_SEGMENT|5825,5835|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|SIMPLE_SEGMENT|5825,5835|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|SIMPLE_SEGMENT|5825,5835|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|SIMPLE_SEGMENT|5825,5835|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Finding|SIMPLE_SEGMENT|5843,5846|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|SIMPLE_SEGMENT|5843,5846|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Functional Concept|SIMPLE_SEGMENT|5847,5851|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5853,5860|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|abdomen
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5853,5860|false|false|false|C0153662|Malignant neoplasm of abdomen|abdomen
Finding|Finding|SIMPLE_SEGMENT|5853,5860|false|false|false|C0941288|Abdomen problem|abdomen
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5862,5868|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5862,5868|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5862,5868|false|false|false|C0153663|Malignant neoplasm of pelvis|pelvis
Event|Event|SIMPLE_SEGMENT|5862,5868|false|false|false|||pelvis
Finding|Finding|SIMPLE_SEGMENT|5862,5868|false|false|false|C0812455|Pelvis problem|pelvis
Finding|Intellectual Product|SIMPLE_SEGMENT|5874,5878|false|false|false|C1547225|Mild Severity of Illness Code|mild
Event|Activity|SIMPLE_SEGMENT|5897,5908|true|false|false|C2349975|Enhance (action)|enhancement
Event|Event|SIMPLE_SEGMENT|5897,5908|true|false|false|||enhancement
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5897,5908|true|false|false|C1627358|Refractive surgery enhancement|enhancement
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5911,5920|true|true|false|C0009450|Communicable Diseases|infection
Event|Event|SIMPLE_SEGMENT|5911,5920|true|false|false|||infection
Finding|Pathologic Function|SIMPLE_SEGMENT|5911,5920|true|true|false|C3714514|Infection|infection
Event|Event|SIMPLE_SEGMENT|5931,5939|true|false|false|||excluded
Finding|Finding|SIMPLE_SEGMENT|5954,5960|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|SIMPLE_SEGMENT|5954,5960|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Event|Event|SIMPLE_SEGMENT|5961,5965|false|false|false|||left
Finding|Functional Concept|SIMPLE_SEGMENT|5961,5965|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Event|Event|SIMPLE_SEGMENT|5971,5979|false|false|false|||moderate
Finding|Finding|SIMPLE_SEGMENT|5971,5979|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|SIMPLE_SEGMENT|5971,5979|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Finding|SIMPLE_SEGMENT|5983,5989|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|SIMPLE_SEGMENT|5983,5989|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Event|Event|SIMPLE_SEGMENT|5990,5995|false|false|false|||right
Finding|Functional Concept|SIMPLE_SEGMENT|5990,5995|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5997,6018|false|false|false|C0268804|Hydroureteronephrosis|hydroureteronephrosis
Event|Event|SIMPLE_SEGMENT|5997,6018|false|false|false|||hydroureteronephrosis
Finding|Functional Concept|SIMPLE_SEGMENT|6033,6037|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Event|Event|SIMPLE_SEGMENT|6038,6048|false|false|false|||nephrogram
Event|Event|SIMPLE_SEGMENT|6050,6056|false|false|false|||stable
Finding|Intellectual Product|SIMPLE_SEGMENT|6050,6056|false|false|false|C1547311|Patient Condition Code - Stable|stable
Finding|Finding|SIMPLE_SEGMENT|6071,6075|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|Mass
Finding|Gene or Genome|SIMPLE_SEGMENT|6071,6075|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|Mass
Finding|Intellectual Product|SIMPLE_SEGMENT|6071,6075|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|Mass
Finding|Finding|SIMPLE_SEGMENT|6071,6082|false|false|false|C4086564|Mass Effect|Mass effect
Event|Event|SIMPLE_SEGMENT|6076,6082|false|false|false|||effect
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|6089,6100|false|false|false|C0500470|Anatomical anastomosis|anastomosis
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|6089,6100|false|false|false|C0332853|Anastomosis|anastomosis
Event|Event|SIMPLE_SEGMENT|6089,6100|false|false|false|||anastomosis
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6089,6100|false|false|false|C0677554||anastomosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6109,6115|false|false|false|C4522154|Distal Resection Margin|distal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6116,6123|false|false|false|C0041951|Ureter|ureters
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|6129,6139|false|false|false|C3898148|Neobladder|neobladder
Event|Event|SIMPLE_SEGMENT|6144,6152|false|false|false|||resolved
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6179,6193|false|false|false|C0020295|Hydronephrosis|hydronephrosis
Event|Event|SIMPLE_SEGMENT|6179,6193|false|false|false|||hydronephrosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6215,6220|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|6215,6220|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|6215,6220|false|false|false|C0013604|Edema|edema
Event|Event|SIMPLE_SEGMENT|6240,6247|true|false|false|||resolve
Event|Event|SIMPLE_SEGMENT|6261,6271|true|false|false|||etiologies
Finding|Functional Concept|SIMPLE_SEGMENT|6261,6271|true|false|false|C0015127|Etiology aspects|etiologies
Event|Event|SIMPLE_SEGMENT|6282,6290|true|false|false|||stenosis
Finding|Pathologic Function|SIMPLE_SEGMENT|6282,6290|true|false|false|C1261287|Stenosis|stenosis
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6292,6297|false|false|false|C0027651|Neoplasms|tumor
Event|Event|SIMPLE_SEGMENT|6292,6297|false|false|false|||tumor
Finding|Finding|SIMPLE_SEGMENT|6292,6297|false|false|false|C1578706;C3273930|Tumor Mass|tumor
Finding|Intellectual Product|SIMPLE_SEGMENT|6292,6297|false|false|false|C1578706;C3273930|Tumor Mass|tumor
Event|Event|SIMPLE_SEGMENT|6299,6311|false|false|false|||infiltration
Finding|Functional Concept|SIMPLE_SEGMENT|6299,6311|false|false|false|C0332448;C1523986;C3669041|Infiltration;Infiltration Route of Administration;Spread by direct extension|infiltration
Finding|Pathologic Function|SIMPLE_SEGMENT|6299,6311|false|false|false|C0332448;C1523986;C3669041|Infiltration;Infiltration Route of Administration;Spread by direct extension|infiltration
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6299,6311|false|false|false|C0702249|Infiltration (procedure)|infiltration
Event|Event|SIMPLE_SEGMENT|6322,6330|false|false|false|||excluded
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6341,6348|false|false|false|C0205054|Hepatic|hepatic
Finding|Finding|SIMPLE_SEGMENT|6341,6355|false|false|false|C0577053|Lesion of liver|hepatic lesion
Event|Event|SIMPLE_SEGMENT|6349,6355|false|false|false|||lesion
Finding|Finding|SIMPLE_SEGMENT|6349,6355|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|SIMPLE_SEGMENT|6349,6355|false|false|false|C0221198;C1546698|Lesion|lesion
Event|Event|SIMPLE_SEGMENT|6369,6378|false|false|false|||attention
Finding|Intellectual Product|SIMPLE_SEGMENT|6369,6378|false|false|false|C0004268;C4281780|Attention;Attention - G-code|attention
Finding|Mental Process|SIMPLE_SEGMENT|6369,6378|false|false|false|C0004268;C4281780|Attention;Attention - G-code|attention
Event|Governmental or Regulatory Activity|SIMPLE_SEGMENT|6387,6391|false|false|false|C1510751|Academic Research Enhancement Awards|area
Event|Event|SIMPLE_SEGMENT|6408,6417|false|false|false|||followups
Event|Event|SIMPLE_SEGMENT|6418,6429|false|false|false|||recommended
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6436,6450|false|false|false|C0184661;C2183254|Interventional procedure;interventional (invasive) radiology|INTERVENTIONAL
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6436,6450|false|false|false|C0184661;C2183254|Interventional procedure;interventional (invasive) radiology|INTERVENTIONAL
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6436,6460|false|false|false|C0184661|Interventional procedure|INTERVENTIONAL PROCEDURE
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6451,6460|false|false|false|C0945766||PROCEDURE
Event|Event|SIMPLE_SEGMENT|6451,6460|false|false|false|||PROCEDURE
Event|Occupational Activity|SIMPLE_SEGMENT|6451,6460|false|false|false|C1546467|Act Class - procedure|PROCEDURE
Finding|Functional Concept|SIMPLE_SEGMENT|6451,6460|false|false|false|C2700391|Procedure (set of actions)|PROCEDURE
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6451,6460|false|false|false|C0184661|Interventional procedure|PROCEDURE
Drug|Organic Chemical|SIMPLE_SEGMENT|6470,6478|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|Complete
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6470,6478|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|Complete
Drug|Vitamin|SIMPLE_SEGMENT|6470,6478|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|Complete
Finding|Functional Concept|SIMPLE_SEGMENT|6470,6478|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|Complete
Finding|Idea or Concept|SIMPLE_SEGMENT|6470,6478|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|Complete
Event|Event|SIMPLE_SEGMENT|6479,6487|false|false|false|||collapse
Finding|Finding|SIMPLE_SEGMENT|6479,6487|false|false|false|C0036974;C0344329;C2210463|Collapse (finding);Shock|collapse
Finding|Pathologic Function|SIMPLE_SEGMENT|6479,6487|false|false|false|C0036974;C0344329;C2210463|Collapse (finding);Shock|collapse
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|6479,6487|false|false|false|C0332521|Collapse (morphologic abnormality)|collapse
Finding|Body Substance|SIMPLE_SEGMENT|6492,6499|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|6492,6499|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|6492,6499|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|SIMPLE_SEGMENT|6492,6503|false|false|false|C0332310|Has patient|patient has
Event|Event|SIMPLE_SEGMENT|6513,6520|false|false|false|||drained
Finding|Functional Concept|SIMPLE_SEGMENT|6521,6525|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6527,6532|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|6527,6532|false|false|false|C2003888|Lower (action)|lower
Event|Event|SIMPLE_SEGMENT|6543,6553|false|false|false|||collection
Finding|Conceptual Entity|SIMPLE_SEGMENT|6543,6553|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|SIMPLE_SEGMENT|6543,6553|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|SIMPLE_SEGMENT|6543,6553|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|SIMPLE_SEGMENT|6543,6553|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Event|Event|SIMPLE_SEGMENT|6560,6568|false|false|false|||catheter
Finding|Intellectual Product|SIMPLE_SEGMENT|6560,6568|false|false|false|C1546572||catheter
Event|Event|SIMPLE_SEGMENT|6579,6589|false|false|false|||collection
Finding|Conceptual Entity|SIMPLE_SEGMENT|6579,6589|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|SIMPLE_SEGMENT|6579,6589|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|SIMPLE_SEGMENT|6579,6589|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|SIMPLE_SEGMENT|6579,6589|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Event|Event|SIMPLE_SEGMENT|6594,6601|false|false|false|||removed
Finding|Finding|SIMPLE_SEGMENT|6608,6621|false|false|false|C4489118|Near complete|Near complete
Drug|Organic Chemical|SIMPLE_SEGMENT|6613,6621|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6613,6621|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|SIMPLE_SEGMENT|6613,6621|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|SIMPLE_SEGMENT|6613,6621|false|false|false|||complete
Finding|Functional Concept|SIMPLE_SEGMENT|6613,6621|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|SIMPLE_SEGMENT|6613,6621|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Event|Event|SIMPLE_SEGMENT|6622,6630|false|false|false|||collapse
Finding|Finding|SIMPLE_SEGMENT|6622,6630|false|false|false|C0036974;C0344329;C2210463|Collapse (finding);Shock|collapse
Finding|Pathologic Function|SIMPLE_SEGMENT|6622,6630|false|false|false|C0036974;C0344329;C2210463|Collapse (finding);Shock|collapse
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|6622,6630|false|false|false|C0332521|Collapse (morphologic abnormality)|collapse
Finding|Body Substance|SIMPLE_SEGMENT|6638,6645|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|6638,6645|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|6638,6645|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|6660,6667|false|false|false|||drained
Event|Event|SIMPLE_SEGMENT|6669,6679|false|false|false|||collection
Finding|Conceptual Entity|SIMPLE_SEGMENT|6669,6679|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|SIMPLE_SEGMENT|6669,6679|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|SIMPLE_SEGMENT|6669,6679|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|SIMPLE_SEGMENT|6669,6679|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6691,6697|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|6691,6697|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6691,6697|false|false|false|C0153663|Malignant neoplasm of pelvis|pelvis
Finding|Finding|SIMPLE_SEGMENT|6691,6697|false|false|false|C0812455|Pelvis problem|pelvis
Event|Event|SIMPLE_SEGMENT|6712,6720|false|false|false|||catheter
Finding|Intellectual Product|SIMPLE_SEGMENT|6712,6720|false|false|false|C1546572||catheter
Event|Activity|SIMPLE_SEGMENT|6724,6729|false|false|false|C1882509|put - instruction imperative|place
Event|Event|SIMPLE_SEGMENT|6724,6729|false|false|false|||place
Finding|Functional Concept|SIMPLE_SEGMENT|6724,6729|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|SIMPLE_SEGMENT|6724,6729|false|false|false|C1533810||place
Finding|Functional Concept|SIMPLE_SEGMENT|6736,6740|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6736,6755|false|false|false|C0230180|Structure of left lower quadrant of abdomen|Left lower quadrant
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6741,6746|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|6741,6746|false|false|false|C2003888|Lower (action)|lower
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6760,6764|false|false|false|C4318566|Deep Resection Margin|deep
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6765,6771|false|false|false|C0030797|Pelvis|pelvic
Event|Event|SIMPLE_SEGMENT|6772,6783|false|false|false|||collections
Finding|Idea or Concept|SIMPLE_SEGMENT|6787,6792|false|false|false|C1552828|Table Frame - above|above
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6802,6810|false|false|true|C2926606||findings
Event|Event|SIMPLE_SEGMENT|6802,6810|false|false|false|||findings
Finding|Functional Concept|SIMPLE_SEGMENT|6802,6810|false|false|true|C2607943|findings aspects|findings
Event|Event|SIMPLE_SEGMENT|6816,6825|false|false|false|||discussed
Event|Event|SIMPLE_SEGMENT|6842,6847|false|false|false|||Given
Finding|Body Substance|SIMPLE_SEGMENT|6853,6860|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|6853,6860|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|6853,6860|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|6863,6872|false|false|false|||improving
Finding|Intellectual Product|SIMPLE_SEGMENT|6873,6881|false|false|false|C1315013|Clinical NEC (not elsewhere classified in LNC)|clinical
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6873,6888|false|false|false|C0449440;C5890498|Clinical status|clinical status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6882,6888|false|false|false|C5889824||status
Event|Event|SIMPLE_SEGMENT|6882,6888|false|false|false|||status
Finding|Idea or Concept|SIMPLE_SEGMENT|6882,6888|false|false|false|C1546481|What subject filter - Status|status
Event|Event|SIMPLE_SEGMENT|6894,6902|true|false|false|||decision
Finding|Mental Process|SIMPLE_SEGMENT|6894,6902|true|false|false|C0679006|Decision|decision
Finding|Conceptual Entity|SIMPLE_SEGMENT|6934,6944|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|SIMPLE_SEGMENT|6934,6944|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|SIMPLE_SEGMENT|6934,6944|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|SIMPLE_SEGMENT|6934,6944|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Event|Event|SIMPLE_SEGMENT|6945,6953|true|false|false|||drainage
Finding|Body Substance|SIMPLE_SEGMENT|6945,6953|true|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Finding|Sign or Symptom|SIMPLE_SEGMENT|6945,6953|true|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6945,6953|true|false|false|C0013103|Drainage procedure|drainage
Finding|Finding|SIMPLE_SEGMENT|6962,6966|true|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|6962,6966|true|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|6962,6966|true|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Finding|SIMPLE_SEGMENT|6973,6979|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|Severe
Finding|Intellectual Product|SIMPLE_SEGMENT|6973,6979|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|Severe
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6980,7004|false|false|false|C0521622|Bilateral hydronephrosis|bilateral hydronephrosis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6990,7004|false|false|false|C0020295|Hydronephrosis|hydronephrosis
Event|Event|SIMPLE_SEGMENT|6990,7004|false|false|false|||hydronephrosis
Event|Event|SIMPLE_SEGMENT|7018,7030|false|false|false|||examinations
Procedure|Health Care Activity|SIMPLE_SEGMENT|7018,7030|false|false|false|C0031809|Physical Examination|examinations
Event|Event|SIMPLE_SEGMENT|7033,7047|false|false|false|||RECOMMENDATION
Finding|Idea or Concept|SIMPLE_SEGMENT|7033,7047|false|false|false|C0034866|Recommendation|RECOMMENDATION
Event|Event|SIMPLE_SEGMENT|7056,7067|false|false|false|||persistence
Finding|Mental Process|SIMPLE_SEGMENT|7056,7067|false|false|false|C0546816|Persistence|persistence
Finding|Finding|SIMPLE_SEGMENT|7071,7077|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|SIMPLE_SEGMENT|7071,7077|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7071,7092|false|false|false|C0237061|Severe hydronephrosis|severe hydronephrosis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7078,7092|false|false|false|C0020295|Hydronephrosis|hydronephrosis
Event|Event|SIMPLE_SEGMENT|7078,7092|false|false|false|||hydronephrosis
Event|Event|SIMPLE_SEGMENT|7095,7107|false|false|false|||percutaneous
Finding|Functional Concept|SIMPLE_SEGMENT|7095,7107|false|false|false|C1522243|Percutaneous Route of Drug Administration|percutaneous
Event|Event|SIMPLE_SEGMENT|7109,7120|false|false|false|||nephrostomy
Finding|Finding|SIMPLE_SEGMENT|7109,7120|false|false|false|C0481713|Has nephrostomy|nephrostomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7109,7120|false|false|false|C0278314|Nephrostomy (procedure)|nephrostomy
Event|Event|SIMPLE_SEGMENT|7121,7126|false|false|false|||tubes
Finding|Intellectual Product|SIMPLE_SEGMENT|7121,7126|false|false|false|C1547937||tubes
Event|Event|SIMPLE_SEGMENT|7137,7147|false|false|false|||considered
Finding|Intellectual Product|SIMPLE_SEGMENT|7153,7158|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|Brief
Finding|Idea or Concept|SIMPLE_SEGMENT|7159,7167|false|false|false|C1547192|Organization unit type - Hospital|Hospital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7159,7174|false|false|false|C0488549||Hospital Course
Finding|Finding|SIMPLE_SEGMENT|7159,7174|false|false|false|C0489547|Hospital course|Hospital Course
Finding|Intellectual Product|SIMPLE_SEGMENT|7176,7181|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|BRIEF
Event|Event|SIMPLE_SEGMENT|7182,7189|false|false|false|||SUMMARY
Finding|Intellectual Product|SIMPLE_SEGMENT|7182,7189|false|false|false|C1552616;C1706244|Summary (document);summary - ActRelationshipSubset|SUMMARY
Finding|Idea or Concept|SIMPLE_SEGMENT|7210,7214|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|SIMPLE_SEGMENT|7210,7214|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Event|Event|SIMPLE_SEGMENT|7219,7224|false|false|false|||women
Event|Event|SIMPLE_SEGMENT|7232,7239|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|7232,7239|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|7232,7239|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|7232,7239|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|7232,7242|false|false|false|C0262926|Medical History|history of
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7243,7250|false|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7243,7250|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7243,7250|false|false|false|C0872388|Procedures on bladder|bladder
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7243,7257|false|false|false|C0005684;C0005695;C0699885|Bladder Neoplasm;Carcinoma of bladder;Malignant neoplasm of urinary bladder|bladder cancer
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7251,7257|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|SIMPLE_SEGMENT|7251,7257|false|false|false|||cancer
Event|Event|SIMPLE_SEGMENT|7263,7273|false|false|false|||cystectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7263,7273|false|false|false|C0010651|Cystectomy|cystectomy
Event|Event|SIMPLE_SEGMENT|7275,7287|false|false|false|||hysterectomy
Finding|Finding|SIMPLE_SEGMENT|7275,7287|false|false|false|C1548863|Consent Type - Hysterectomy|hysterectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7275,7287|false|false|false|C0020699|Hysterectomy|hysterectomy
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7293,7296|false|false|false|C0054252|Buthionine Sulfoximine|BSO
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|7293,7296|false|false|false|C0054252|Buthionine Sulfoximine|BSO
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7293,7296|false|false|false|C0054252|Buthionine Sulfoximine|BSO
Event|Event|SIMPLE_SEGMENT|7293,7296|false|false|false|||BSO
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7306,7311|false|false|false|C0020885|ileum|ileal
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|7306,7319|false|false|false|C0441253|Structure of ileal conduit|ileal conduit
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7306,7319|false|false|false|C0348002|Ileal conduit procedure|ileal conduit
Event|Event|SIMPLE_SEGMENT|7312,7319|false|false|false|||conduit
Finding|Finding|SIMPLE_SEGMENT|7328,7342|false|false|false|C0241311|post operative (finding)|post operative
Event|Event|SIMPLE_SEGMENT|7343,7349|false|false|false|||course
Event|Event|SIMPLE_SEGMENT|7359,7370|false|false|false|||complicated
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7374,7377|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7374,7377|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7374,7377|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7382,7387|false|false|false|C1258215;C4019039|Ileus;Intestinal obstruction co-occurrent and due to decreased peristalsis|ileus
Event|Event|SIMPLE_SEGMENT|7382,7387|false|false|false|||ileus
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7394,7400|false|false|false|C0030797|Pelvis|pelvic
Drug|Substance|SIMPLE_SEGMENT|7401,7406|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|7401,7406|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|7401,7406|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|7407,7418|false|false|false|||collections
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7426,7429|false|false|false|C0230180|Structure of left lower quadrant of abdomen|LLQ
Drug|Substance|SIMPLE_SEGMENT|7430,7435|false|false|false|C1550628|Drain - SpecimenType|drain
Event|Event|SIMPLE_SEGMENT|7430,7435|false|false|false|||drain
Finding|Intellectual Product|SIMPLE_SEGMENT|7430,7435|false|false|false|C1546604|Drain Specimen Code|drain
Event|Event|SIMPLE_SEGMENT|7436,7445|false|false|false|||presented
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7452,7462|false|false|false|C2979880||subjective
Finding|Finding|SIMPLE_SEGMENT|7452,7462|false|false|false|C2266644|subjective (symptom)|subjective
Event|Event|SIMPLE_SEGMENT|7463,7469|false|false|false|||fevers
Finding|Sign or Symptom|SIMPLE_SEGMENT|7463,7469|false|false|false|C0015967|Fever|fevers
Event|Event|SIMPLE_SEGMENT|7471,7479|false|false|false|||lethargy
Finding|Sign or Symptom|SIMPLE_SEGMENT|7471,7479|false|false|false|C0023380|Lethargy|lethargy
Finding|Finding|SIMPLE_SEGMENT|7485,7491|false|false|false|C4554530|Bloody|bloody
Drug|Substance|SIMPLE_SEGMENT|7492,7497|false|false|false|C1550628|Drain - SpecimenType|drain
Event|Event|SIMPLE_SEGMENT|7492,7497|false|false|false|||drain
Finding|Intellectual Product|SIMPLE_SEGMENT|7492,7497|false|false|false|C1546604|Drain Specimen Code|drain
Event|Event|SIMPLE_SEGMENT|7498,7504|false|false|false|||output
Finding|Conceptual Entity|SIMPLE_SEGMENT|7498,7504|false|false|false|C1709366|system output|output
Procedure|Health Care Activity|SIMPLE_SEGMENT|7498,7504|false|false|false|C3251815|Measurement of fluid output|output
Event|Event|SIMPLE_SEGMENT|7515,7520|false|false|false|||found
Finding|Idea or Concept|SIMPLE_SEGMENT|7529,7538|false|false|false|C1546960|Patient Outcome - Worsening|worsening
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7539,7545|false|false|false|C0002871|Anemia|anemia
Event|Event|SIMPLE_SEGMENT|7539,7545|false|false|false|||anemia
Event|Event|SIMPLE_SEGMENT|7554,7559|false|false|false|||given
Event|Event|SIMPLE_SEGMENT|7562,7567|false|false|false|||units
Event|Event|SIMPLE_SEGMENT|7594,7602|false|false|false|||increase
Finding|Functional Concept|SIMPLE_SEGMENT|7594,7602|false|false|false|C0442805|Increase|increase
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7606,7616|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7606,7616|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Organic Chemical|SIMPLE_SEGMENT|7606,7616|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7606,7616|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Event|Event|SIMPLE_SEGMENT|7606,7616|false|false|false|||hemoglobin
Finding|Finding|SIMPLE_SEGMENT|7606,7616|false|false|false|C1561562|Hemoglobin finding|hemoglobin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7606,7616|false|false|false|C0518015|Hemoglobin measurement|hemoglobin
Event|Event|SIMPLE_SEGMENT|7617,7622|false|false|false|||noted
Event|Event|SIMPLE_SEGMENT|7638,7643|false|false|false|||found
Event|Event|SIMPLE_SEGMENT|7650,7657|false|false|false|||imaging
Finding|Finding|SIMPLE_SEGMENT|7650,7657|false|false|false|C0740845|Imaging problem|imaging
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7650,7657|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|imaging
Finding|Intellectual Product|SIMPLE_SEGMENT|7669,7677|false|false|false|C1552654|Parameterized Data Type - Interval|interval
Event|Event|SIMPLE_SEGMENT|7678,7686|false|false|false|||increase
Finding|Functional Concept|SIMPLE_SEGMENT|7678,7686|false|false|false|C0442805|Increase|increase
Finding|Finding|SIMPLE_SEGMENT|7678,7694|false|false|false|C1268652|increase in size|increase in size
Finding|Functional Concept|SIMPLE_SEGMENT|7701,7705|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7706,7715|false|false|false|C0000726|Abdomen|abdominal
Finding|Body Substance|SIMPLE_SEGMENT|7706,7721|false|false|false|C2699330|Abdominal Fluid|abdominal fluid
Drug|Substance|SIMPLE_SEGMENT|7716,7721|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|7716,7721|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|7716,7721|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|7722,7732|false|false|false|||collection
Finding|Conceptual Entity|SIMPLE_SEGMENT|7722,7732|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|SIMPLE_SEGMENT|7722,7732|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|SIMPLE_SEGMENT|7722,7732|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|SIMPLE_SEGMENT|7722,7732|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Event|Event|SIMPLE_SEGMENT|7734,7742|false|false|false|||Decision
Finding|Mental Process|SIMPLE_SEGMENT|7734,7742|false|false|false|C0679006|Decision|Decision
Event|Activity|SIMPLE_SEGMENT|7755,7760|false|false|false|C1882509|put - instruction imperative|place
Finding|Functional Concept|SIMPLE_SEGMENT|7755,7760|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|SIMPLE_SEGMENT|7755,7760|false|false|false|C1533810||place
Drug|Substance|SIMPLE_SEGMENT|7764,7769|false|false|false|C1550628|Drain - SpecimenType|drain
Event|Event|SIMPLE_SEGMENT|7764,7769|false|false|false|||drain
Finding|Intellectual Product|SIMPLE_SEGMENT|7764,7769|false|false|false|C1546604|Drain Specimen Code|drain
Drug|Substance|SIMPLE_SEGMENT|7778,7783|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|Fluid
Event|Event|SIMPLE_SEGMENT|7778,7783|false|false|false|||Fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|7778,7783|false|false|false|C1546638|Fluid Specimen Code|Fluid
Event|Event|SIMPLE_SEGMENT|7788,7792|false|false|false|||sent
Event|Event|SIMPLE_SEGMENT|7797,7805|false|false|false|||revealed
Finding|Classification|SIMPLE_SEGMENT|7807,7815|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|7807,7815|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|7807,7815|false|false|false|C5237010|Expression Negative|negative
Event|Event|SIMPLE_SEGMENT|7816,7824|true|false|false|||cultures
Finding|Idea or Concept|SIMPLE_SEGMENT|7816,7824|true|true|false|C0010453|Culture (Anthropological)|cultures
Event|Event|SIMPLE_SEGMENT|7827,7835|true|false|false|||negative
Finding|Classification|SIMPLE_SEGMENT|7827,7835|true|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|7827,7835|true|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|7827,7835|true|false|false|C5237010|Expression Negative|negative
Anatomy|Cell|SIMPLE_SEGMENT|7836,7851|true|false|false|C0334227|Tumor cells, malignant|malignant cells
Anatomy|Cell|SIMPLE_SEGMENT|7846,7851|true|false|false|C0007634|Cells|cells
Event|Event|SIMPLE_SEGMENT|7856,7864|true|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|7856,7864|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|7856,7867|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7868,7877|true|false|false|C0229889|Lymphatic vessel|lymphatic
Finding|Finding|SIMPLE_SEGMENT|7868,7877|true|false|false|C0740775|Lymphatic problem|lymphatic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7881,7888|true|false|false|C0042027|Urinary tract|urinary
Drug|Substance|SIMPLE_SEGMENT|7890,7895|true|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|7890,7895|true|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|7890,7895|true|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Finding|SIMPLE_SEGMENT|7902,7905|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|7902,7905|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Drug|Substance|SIMPLE_SEGMENT|7906,7911|false|false|false|C1550628|Drain - SpecimenType|drain
Event|Event|SIMPLE_SEGMENT|7906,7911|false|false|false|||drain
Finding|Intellectual Product|SIMPLE_SEGMENT|7906,7911|false|false|false|C1546604|Drain Specimen Code|drain
Event|Event|SIMPLE_SEGMENT|7929,7936|false|false|false|||removed
Drug|Substance|SIMPLE_SEGMENT|7948,7953|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|7948,7953|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|7948,7953|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|7955,7965|false|false|false|||collection
Finding|Conceptual Entity|SIMPLE_SEGMENT|7955,7965|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|SIMPLE_SEGMENT|7955,7965|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|SIMPLE_SEGMENT|7955,7965|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|SIMPLE_SEGMENT|7955,7965|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|SIMPLE_SEGMENT|7970,7980|false|false|false|C4554154|Completely - dosing instruction fragment|completely
Event|Event|SIMPLE_SEGMENT|7981,7988|false|false|false|||drained
Drug|Substance|SIMPLE_SEGMENT|8000,8005|false|false|false|C1550628|Drain - SpecimenType|drain
Event|Event|SIMPLE_SEGMENT|8000,8005|false|false|false|||drain
Finding|Intellectual Product|SIMPLE_SEGMENT|8000,8005|false|false|false|C1546604|Drain Specimen Code|drain
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8010,8015|false|false|false|C1410088|Still|still
Event|Event|SIMPLE_SEGMENT|8017,8025|false|false|false|||draining
Finding|Body Substance|SIMPLE_SEGMENT|8026,8046|false|false|false|C4518404|Serosanguinous fluid|serosanguinous fluid
Drug|Substance|SIMPLE_SEGMENT|8041,8046|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|8041,8046|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|8041,8046|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|8055,8059|false|false|false|||kept
Event|Event|SIMPLE_SEGMENT|8067,8079|false|false|false|||repositioned
Event|Event|SIMPLE_SEGMENT|8089,8098|false|false|false|||consulted
Event|Event|SIMPLE_SEGMENT|8107,8113|false|false|false|||fevers
Finding|Sign or Symptom|SIMPLE_SEGMENT|8107,8113|false|false|false|C0015967|Fever|fevers
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8115,8127|false|false|false|C0023518|Leukocytosis|leukocytosis
Event|Event|SIMPLE_SEGMENT|8115,8127|false|false|false|||leukocytosis
Finding|Finding|SIMPLE_SEGMENT|8115,8127|false|false|false|C0750426|Blood leukocyte number above reference range|leukocytosis
Drug|Substance|SIMPLE_SEGMENT|8132,8137|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|8132,8137|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|8132,8137|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|8139,8150|false|false|false|||collections
Event|Event|SIMPLE_SEGMENT|8159,8165|false|false|false|||deemed
Drug|Antibiotic|SIMPLE_SEGMENT|8174,8185|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|SIMPLE_SEGMENT|8174,8185|false|false|false|||antibiotics
Event|Event|SIMPLE_SEGMENT|8216,8224|false|false|false|||spectrum
Finding|Conceptual Entity|SIMPLE_SEGMENT|8216,8224|false|false|false|C2827424|Spectrum|spectrum
Drug|Antibiotic|SIMPLE_SEGMENT|8231,8240|false|false|false|C1120106|ertapenem|ertapenem
Drug|Organic Chemical|SIMPLE_SEGMENT|8231,8240|false|false|false|C1120106|ertapenem|ertapenem
Event|Event|SIMPLE_SEGMENT|8231,8240|false|false|false|||ertapenem
Event|Event|SIMPLE_SEGMENT|8244,8253|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|8244,8253|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|8244,8253|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|8244,8253|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|8244,8253|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|SIMPLE_SEGMENT|8260,8267|false|false|false|||require
Finding|Functional Concept|SIMPLE_SEGMENT|8278,8284|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|SIMPLE_SEGMENT|8278,8284|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Disorder|Neoplastic Process|SIMPLE_SEGMENT|8285,8288|false|false|false|C0334463|Malignant Fibrous Histiocytoma|ups
Event|Event|SIMPLE_SEGMENT|8285,8288|false|false|false|||ups
Finding|Gene or Genome|SIMPLE_SEGMENT|8285,8288|false|false|false|C1415597|HMBS gene|ups
Event|Event|SIMPLE_SEGMENT|8293,8300|false|false|false|||imaging
Finding|Finding|SIMPLE_SEGMENT|8293,8300|false|false|false|C0740845|Imaging problem|imaging
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8293,8300|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|imaging
Event|Event|SIMPLE_SEGMENT|8304,8313|false|false|false|||specified
Finding|Idea or Concept|SIMPLE_SEGMENT|8321,8333|false|false|false|C1548597|Marketing basis - Transitional|transitional
Event|Event|SIMPLE_SEGMENT|8335,8341|false|false|false|||issues
Finding|Intellectual Product|SIMPLE_SEGMENT|8346,8351|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|ACUTE
Event|Event|SIMPLE_SEGMENT|8352,8358|false|false|false|||ISSUES
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8375,8381|false|false|false|C0030797|Pelvis|Pelvic
Drug|Substance|SIMPLE_SEGMENT|8382,8387|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|8382,8387|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|8382,8387|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|8388,8399|false|false|false|||collections
Finding|Body Substance|SIMPLE_SEGMENT|8401,8408|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|8401,8408|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|8401,8408|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|8409,8416|false|false|false|||arrived
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8426,8434|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Drug|Substance|SIMPLE_SEGMENT|8436,8441|false|false|false|C1550628|Drain - SpecimenType|drain
Event|Event|SIMPLE_SEGMENT|8436,8441|false|false|false|||drain
Finding|Intellectual Product|SIMPLE_SEGMENT|8436,8441|false|false|false|C1546604|Drain Specimen Code|drain
Event|Event|SIMPLE_SEGMENT|8442,8449|false|false|false|||putting
Finding|Body Substance|SIMPLE_SEGMENT|8454,8474|false|false|false|C4518404|Serosanguinous fluid|serosanguinous fluid
Drug|Substance|SIMPLE_SEGMENT|8469,8474|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|8469,8474|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|8469,8474|false|false|false|C1546638|Fluid Specimen Code|fluid
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8476,8486|false|false|false|C1644645||CT abdomen
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8476,8486|false|false|false|C0412620|CT of abdomen|CT abdomen
Anatomy|Body Location or Region|SIMPLE_SEGMENT|8479,8486|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|abdomen
Disorder|Neoplastic Process|SIMPLE_SEGMENT|8479,8486|false|false|false|C0153662|Malignant neoplasm of abdomen|abdomen
Event|Event|SIMPLE_SEGMENT|8479,8486|false|false|false|||abdomen
Finding|Finding|SIMPLE_SEGMENT|8479,8486|false|false|false|C0941288|Abdomen problem|abdomen
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8487,8493|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|8487,8493|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Disorder|Neoplastic Process|SIMPLE_SEGMENT|8487,8493|false|false|false|C0153663|Malignant neoplasm of pelvis|pelvis
Finding|Finding|SIMPLE_SEGMENT|8487,8493|false|false|false|C0812455|Pelvis problem|pelvis
Event|Event|SIMPLE_SEGMENT|8495,8503|false|false|false|||revealed
Finding|Functional Concept|SIMPLE_SEGMENT|8514,8518|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Drug|Substance|SIMPLE_SEGMENT|8519,8524|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|8519,8524|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|8525,8535|false|false|false|||collection
Finding|Conceptual Entity|SIMPLE_SEGMENT|8525,8535|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|SIMPLE_SEGMENT|8525,8535|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|SIMPLE_SEGMENT|8525,8535|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|SIMPLE_SEGMENT|8525,8535|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Event|Event|SIMPLE_SEGMENT|8541,8549|false|false|false|||decision
Finding|Mental Process|SIMPLE_SEGMENT|8541,8549|false|false|false|C0679006|Decision|decision
Event|Event|SIMPLE_SEGMENT|8554,8558|false|false|false|||made
Event|Activity|SIMPLE_SEGMENT|8563,8568|false|false|false|C1882509|put - instruction imperative|place
Event|Event|SIMPLE_SEGMENT|8563,8568|false|false|false|||place
Finding|Functional Concept|SIMPLE_SEGMENT|8563,8568|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|SIMPLE_SEGMENT|8563,8568|false|false|false|C1533810||place
Drug|Substance|SIMPLE_SEGMENT|8571,8576|false|false|false|C1550628|Drain - SpecimenType|drain
Event|Event|SIMPLE_SEGMENT|8571,8576|false|false|false|||drain
Finding|Intellectual Product|SIMPLE_SEGMENT|8571,8576|false|false|false|C1546604|Drain Specimen Code|drain
Drug|Substance|SIMPLE_SEGMENT|8590,8595|true|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|8590,8595|true|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|8590,8595|true|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|8600,8608|false|false|false|||negative
Finding|Classification|SIMPLE_SEGMENT|8600,8608|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|8600,8608|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|8600,8608|false|false|false|C5237010|Expression Negative|negative
Finding|Finding|SIMPLE_SEGMENT|8600,8612|false|false|false|C0205160|Negative|negative for
Event|Event|SIMPLE_SEGMENT|8613,8622|true|false|false|||malignant
Anatomy|Cell|SIMPLE_SEGMENT|8624,8629|true|false|false|C0007634|Cells|cells
Drug|Substance|SIMPLE_SEGMENT|8635,8640|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|8635,8640|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|8635,8640|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|8645,8647|false|false|false|||Cr
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8654,8667|false|false|false|C0041004|Triglycerides|triglycerides
Drug|Organic Chemical|SIMPLE_SEGMENT|8654,8667|false|false|false|C0041004|Triglycerides|triglycerides
Event|Event|SIMPLE_SEGMENT|8654,8667|false|false|false|||triglycerides
Finding|Physiologic Function|SIMPLE_SEGMENT|8654,8667|false|false|false|C4554056|Triglycerides metabolic function|triglycerides
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8654,8667|false|false|false|C0202236|Triglycerides measurement|triglycerides
Drug|Substance|SIMPLE_SEGMENT|8688,8693|true|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|8688,8693|true|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|8688,8693|true|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|8694,8704|true|false|false|||collection
Finding|Conceptual Entity|SIMPLE_SEGMENT|8694,8704|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|SIMPLE_SEGMENT|8694,8704|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|SIMPLE_SEGMENT|8694,8704|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|SIMPLE_SEGMENT|8694,8704|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Event|Event|SIMPLE_SEGMENT|8716,8721|true|false|false|||urine
Finding|Body Substance|SIMPLE_SEGMENT|8716,8721|true|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Functional Concept|SIMPLE_SEGMENT|8716,8721|true|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Intellectual Product|SIMPLE_SEGMENT|8716,8721|true|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8726,8735|true|false|false|C0229889|Lymphatic vessel|lymphatic
Finding|Finding|SIMPLE_SEGMENT|8726,8735|true|false|false|C0740775|Lymphatic problem|lymphatic
Drug|Substance|SIMPLE_SEGMENT|8736,8741|true|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|8736,8741|true|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|8736,8741|true|false|false|C1546638|Fluid Specimen Code|fluid
Drug|Substance|SIMPLE_SEGMENT|8743,8748|true|false|false|C0302908;C1704353|Liquid substance;fluid - substance|Fluid
Event|Event|SIMPLE_SEGMENT|8743,8748|true|false|false|||Fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|8743,8748|true|false|false|C1546638|Fluid Specimen Code|Fluid
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8750,8757|true|false|false|C1706355|Culture Dose Form|culture
Event|Event|SIMPLE_SEGMENT|8750,8757|true|false|false|||culture
Finding|Functional Concept|SIMPLE_SEGMENT|8750,8757|true|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Finding|Idea or Concept|SIMPLE_SEGMENT|8750,8757|true|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8750,8757|true|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|culture
Event|Event|SIMPLE_SEGMENT|8762,8770|false|false|false|||negative
Finding|Classification|SIMPLE_SEGMENT|8762,8770|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|8762,8770|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|8762,8770|false|false|false|C5237010|Expression Negative|negative
Finding|Finding|SIMPLE_SEGMENT|8762,8774|false|false|false|C0205160|Negative|negative for
Event|Event|SIMPLE_SEGMENT|8775,8783|true|false|false|||bacteria
Finding|Functional Concept|SIMPLE_SEGMENT|8775,8783|true|false|false|C1510439|bacteria aspects|bacteria
Finding|Intellectual Product|SIMPLE_SEGMENT|8788,8796|false|false|false|C1552654|Parameterized Data Type - Interval|interval
Event|Event|SIMPLE_SEGMENT|8797,8804|false|false|false|||imaging
Finding|Finding|SIMPLE_SEGMENT|8797,8804|false|false|false|C0740845|Imaging problem|imaging
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8797,8804|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|imaging
Finding|Finding|SIMPLE_SEGMENT|8810,8813|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|8810,8813|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Drug|Substance|SIMPLE_SEGMENT|8825,8830|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|8825,8830|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|8825,8830|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|8831,8841|false|false|false|||collection
Finding|Conceptual Entity|SIMPLE_SEGMENT|8831,8841|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|SIMPLE_SEGMENT|8831,8841|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|SIMPLE_SEGMENT|8831,8841|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|SIMPLE_SEGMENT|8831,8841|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|SIMPLE_SEGMENT|8846,8856|false|false|false|C4554154|Completely - dosing instruction fragment|completely
Event|Event|SIMPLE_SEGMENT|8857,8866|false|false|false|||collapsed
Drug|Substance|SIMPLE_SEGMENT|8876,8881|false|false|false|C1550628|Drain - SpecimenType|drain
Event|Event|SIMPLE_SEGMENT|8876,8881|false|false|false|||drain
Finding|Intellectual Product|SIMPLE_SEGMENT|8876,8881|false|false|false|C1546604|Drain Specimen Code|drain
Event|Event|SIMPLE_SEGMENT|8886,8893|false|false|false|||removed
Drug|Substance|SIMPLE_SEGMENT|8912,8917|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|8912,8917|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|8912,8917|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|8918,8928|false|false|false|||collection
Finding|Conceptual Entity|SIMPLE_SEGMENT|8918,8928|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|SIMPLE_SEGMENT|8918,8928|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|SIMPLE_SEGMENT|8918,8928|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|SIMPLE_SEGMENT|8918,8928|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Drug|Substance|SIMPLE_SEGMENT|8949,8954|false|false|false|C1550628|Drain - SpecimenType|drain
Event|Event|SIMPLE_SEGMENT|8949,8954|false|false|false|||drain
Finding|Intellectual Product|SIMPLE_SEGMENT|8949,8954|false|false|false|C1546604|Drain Specimen Code|drain
Event|Event|SIMPLE_SEGMENT|8955,8962|false|false|false|||putting
Finding|Body Substance|SIMPLE_SEGMENT|8967,8987|false|false|false|C4518404|Serosanguinous fluid|serosanguinous fluid
Drug|Substance|SIMPLE_SEGMENT|8982,8987|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|8982,8987|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|8982,8987|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|8993,9002|false|false|false|||continued
Event|Event|SIMPLE_SEGMENT|9006,9011|false|false|false|||drain
Finding|Body Substance|SIMPLE_SEGMENT|9012,9032|false|false|false|C4518404|Serosanguinous fluid|serosanguinous fluid
Drug|Substance|SIMPLE_SEGMENT|9027,9032|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|9027,9032|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|9027,9032|false|false|false|C1546638|Fluid Specimen Code|fluid
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9042,9047|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|9042,9047|false|false|false|C2003888|Lower (action)|lower
Event|Activity|SIMPLE_SEGMENT|9048,9052|false|false|false|C0871208|Rating (action)|rate
Finding|Idea or Concept|SIMPLE_SEGMENT|9048,9052|false|false|false|C1549480|Amount type - Rate|rate
Event|Event|SIMPLE_SEGMENT|9068,9077|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|9068,9077|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Drug|Substance|SIMPLE_SEGMENT|9083,9088|false|false|false|C1550628|Drain - SpecimenType|drain
Event|Event|SIMPLE_SEGMENT|9083,9088|false|false|false|||drain
Finding|Intellectual Product|SIMPLE_SEGMENT|9083,9088|false|false|false|C1546604|Drain Specimen Code|drain
Event|Event|SIMPLE_SEGMENT|9093,9097|false|false|false|||left
Finding|Functional Concept|SIMPLE_SEGMENT|9093,9097|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Event|Activity|SIMPLE_SEGMENT|9101,9106|false|false|false|C1882509|put - instruction imperative|place
Event|Event|SIMPLE_SEGMENT|9101,9106|false|false|false|||place
Finding|Functional Concept|SIMPLE_SEGMENT|9101,9106|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|SIMPLE_SEGMENT|9101,9106|false|false|false|C1533810||place
Drug|Substance|SIMPLE_SEGMENT|9114,9119|true|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|9114,9119|true|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|9114,9119|true|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|9121,9131|true|false|false|||collection
Finding|Conceptual Entity|SIMPLE_SEGMENT|9121,9131|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|SIMPLE_SEGMENT|9121,9131|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|SIMPLE_SEGMENT|9121,9131|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|SIMPLE_SEGMENT|9121,9131|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Event|Event|SIMPLE_SEGMENT|9135,9142|true|false|false|||imaging
Finding|Finding|SIMPLE_SEGMENT|9135,9142|true|false|false|C0740845|Imaging problem|imaging
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|9135,9142|true|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|imaging
Finding|Intellectual Product|SIMPLE_SEGMENT|9151,9161|true|false|false|C4554154|Completely - dosing instruction fragment|completely
Event|Event|SIMPLE_SEGMENT|9162,9171|true|false|false|||collapsed
Finding|Finding|SIMPLE_SEGMENT|9162,9171|true|true|false|C0344329;C0392748|Collapse (finding);Collapsed|collapsed
Finding|Functional Concept|SIMPLE_SEGMENT|9162,9171|true|true|false|C0344329;C0392748|Collapse (finding);Collapsed|collapsed
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|9173,9176|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9173,9176|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9173,9176|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|9173,9176|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|9173,9176|false|false|false|C1332410|BID gene|BID
Event|Event|SIMPLE_SEGMENT|9182,9190|false|false|false|||cultures
Finding|Idea or Concept|SIMPLE_SEGMENT|9182,9190|false|true|false|C0010453|Culture (Anthropological)|cultures
Drug|Substance|SIMPLE_SEGMENT|9214,9219|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|9214,9219|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|9220,9230|false|false|false|||collection
Finding|Conceptual Entity|SIMPLE_SEGMENT|9220,9230|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|SIMPLE_SEGMENT|9220,9230|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|SIMPLE_SEGMENT|9220,9230|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|SIMPLE_SEGMENT|9220,9230|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Event|Event|SIMPLE_SEGMENT|9231,9235|false|false|false|||came
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|9242,9250|false|false|false|C4727483|BRAF Gene Rearrangement|positive
Event|Event|SIMPLE_SEGMENT|9242,9250|false|false|false|||positive
Finding|Classification|SIMPLE_SEGMENT|9242,9250|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|SIMPLE_SEGMENT|9242,9250|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|SIMPLE_SEGMENT|9242,9254|false|false|false|C1446409|Positive|positive for
Event|Event|SIMPLE_SEGMENT|9255,9259|false|false|false|||MSSA
Finding|Finding|SIMPLE_SEGMENT|9255,9259|false|false|false|C2355591|Encounter due to being carrier or suspected carrier of Methicillin susceptible Staphylococcus aureus|MSSA
Event|Event|SIMPLE_SEGMENT|9281,9288|true|false|false|||reflect
Drug|Organic Chemical|SIMPLE_SEGMENT|9289,9292|true|true|false|C0939812|Ruta graveolens preparation|rue
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9289,9292|true|true|false|C0939812|Ruta graveolens preparation|rue
Event|Event|SIMPLE_SEGMENT|9289,9292|true|false|false|||rue
Finding|Functional Concept|SIMPLE_SEGMENT|9294,9309|true|false|false|C1512911|Intraabdominal Route of Administration|intra-abdominal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9294,9319|true|false|false|C1112209|Abdominal Infection|intra-abdominal infection
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9310,9319|true|false|false|C0009450|Communicable Diseases|infection
Event|Event|SIMPLE_SEGMENT|9310,9319|true|false|false|||infection
Finding|Pathologic Function|SIMPLE_SEGMENT|9310,9319|true|false|false|C3714514|Infection|infection
Event|Event|SIMPLE_SEGMENT|9321,9326|false|false|false|||Given
Finding|Body Substance|SIMPLE_SEGMENT|9332,9339|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|9332,9339|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|9332,9339|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|9346,9351|false|false|false|||fever
Finding|Finding|SIMPLE_SEGMENT|9346,9351|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|9346,9351|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9366,9378|false|false|false|C0023518|Leukocytosis|leukocytosis
Event|Event|SIMPLE_SEGMENT|9366,9378|false|false|false|||leukocytosis
Finding|Finding|SIMPLE_SEGMENT|9366,9378|false|false|false|C0750426|Blood leukocyte number above reference range|leukocytosis
Event|Event|SIMPLE_SEGMENT|9388,9394|false|false|false|||placed
Finding|Conceptual Entity|SIMPLE_SEGMENT|9404,9412|false|false|false|C2827424|Spectrum|spectrum
Drug|Antibiotic|SIMPLE_SEGMENT|9413,9424|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|SIMPLE_SEGMENT|9413,9424|false|false|false|||antibiotics
Event|Event|SIMPLE_SEGMENT|9437,9443|false|false|false|||ceftaz
Drug|Organic Chemical|SIMPLE_SEGMENT|9448,9454|false|false|false|C0699678|Flagyl|flagyl
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9448,9454|false|false|false|C0699678|Flagyl|flagyl
Event|Event|SIMPLE_SEGMENT|9448,9454|false|false|false|||flagyl
Event|Event|SIMPLE_SEGMENT|9465,9472|false|false|false|||tapered
Event|Event|SIMPLE_SEGMENT|9480,9484|false|false|false|||team
Drug|Antibiotic|SIMPLE_SEGMENT|9492,9497|false|false|false|C0250482|Zosyn|zosyn
Drug|Organic Chemical|SIMPLE_SEGMENT|9492,9497|false|false|false|C0250482|Zosyn|zosyn
Event|Event|SIMPLE_SEGMENT|9492,9497|false|false|false|||zosyn
Event|Event|SIMPLE_SEGMENT|9502,9511|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|9502,9511|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|9502,9511|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|9502,9511|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|9502,9511|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|SIMPLE_SEGMENT|9516,9527|false|false|false|||recommended
Drug|Antibiotic|SIMPLE_SEGMENT|9528,9537|false|false|false|C1120106|ertapenem|ertapenem
Drug|Organic Chemical|SIMPLE_SEGMENT|9528,9537|false|false|false|C1120106|ertapenem|ertapenem
Event|Event|SIMPLE_SEGMENT|9528,9537|false|false|false|||ertapenem
Finding|Idea or Concept|SIMPLE_SEGMENT|9570,9575|false|false|false|C1546485|Diagnosis Type - Final|final
Event|Event|SIMPLE_SEGMENT|9586,9595|false|false|false|||treatment
Finding|Conceptual Entity|SIMPLE_SEGMENT|9586,9595|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|SIMPLE_SEGMENT|9586,9595|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|SIMPLE_SEGMENT|9586,9595|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9586,9595|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Event|Event|SIMPLE_SEGMENT|9602,9612|false|false|false|||determined
Drug|Substance|SIMPLE_SEGMENT|9616,9621|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|9616,9621|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|9616,9621|false|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Conceptual Entity|SIMPLE_SEGMENT|9623,9633|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|SIMPLE_SEGMENT|9623,9633|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|SIMPLE_SEGMENT|9623,9633|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|SIMPLE_SEGMENT|9623,9633|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Event|Event|SIMPLE_SEGMENT|9634,9641|false|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|9634,9641|false|false|false|C0392747|Changing|changes
Finding|Functional Concept|SIMPLE_SEGMENT|9645,9651|false|false|false|C0205341;C1705914|Repeat;Repeat Object|repeat
Event|Event|SIMPLE_SEGMENT|9652,9659|false|false|false|||imaging
Finding|Finding|SIMPLE_SEGMENT|9652,9659|false|false|false|C0740845|Imaging problem|imaging
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|9652,9659|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|imaging
Finding|Classification|SIMPLE_SEGMENT|9663,9673|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|9663,9673|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9674,9679|false|false|false|C1874451|Basis|basis
Event|Event|SIMPLE_SEGMENT|9674,9679|false|false|false|||basis
Finding|Functional Concept|SIMPLE_SEGMENT|9674,9679|false|false|false|C1527178|Basis - conceptual entity|basis
Event|Event|SIMPLE_SEGMENT|9691,9699|false|false|false|||remained
Event|Event|SIMPLE_SEGMENT|9700,9708|false|false|false|||afebrile
Finding|Finding|SIMPLE_SEGMENT|9700,9708|false|false|false|C0277797|Apyrexial|afebrile
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9714,9726|false|false|false|C0023518|Leukocytosis|leukocytosis
Event|Event|SIMPLE_SEGMENT|9714,9726|false|false|false|||leukocytosis
Finding|Finding|SIMPLE_SEGMENT|9714,9726|false|false|false|C0750426|Blood leukocyte number above reference range|leukocytosis
Event|Event|SIMPLE_SEGMENT|9727,9735|false|false|false|||resolved
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9740,9749|false|false|false|C0024109|Lung|Pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9740,9749|false|false|false|C2707265||Pulmonary
Finding|Finding|SIMPLE_SEGMENT|9740,9749|false|false|false|C4522268|Pulmonary (intended site)|Pulmonary
Finding|Pathologic Function|SIMPLE_SEGMENT|9740,9758|false|false|false|C0034065|Pulmonary Embolism|Pulmonary embolism
Event|Event|SIMPLE_SEGMENT|9750,9758|false|false|false|||embolism
Finding|Finding|SIMPLE_SEGMENT|9750,9758|false|false|false|C0013922;C1704212|Embolism;Embolus|embolism
Finding|Pathologic Function|SIMPLE_SEGMENT|9750,9758|false|false|false|C0013922;C1704212|Embolism;Embolus|embolism
Finding|Finding|SIMPLE_SEGMENT|9760,9766|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Finding|Idea or Concept|SIMPLE_SEGMENT|9760,9766|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Event|Event|SIMPLE_SEGMENT|9767,9776|false|false|false|||developed
Finding|Mental Process|SIMPLE_SEGMENT|9784,9791|false|false|false|C0542559|contextual factors|setting
Event|Event|SIMPLE_SEGMENT|9802,9811|false|false|false|||diagnosed
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9827,9830|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9827,9830|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9827,9830|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Event|Event|SIMPLE_SEGMENT|9827,9830|false|false|false|||DVT
Event|Event|SIMPLE_SEGMENT|9840,9846|false|false|false|||placed
Drug|Organic Chemical|SIMPLE_SEGMENT|9850,9857|false|false|false|C0728963|Lovenox|lovenox
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9850,9857|false|false|false|C0728963|Lovenox|lovenox
Event|Event|SIMPLE_SEGMENT|9850,9857|false|false|false|||lovenox
Event|Event|SIMPLE_SEGMENT|9869,9881|false|false|false|||transitioned
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9885,9892|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Organic Chemical|SIMPLE_SEGMENT|9885,9892|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9885,9892|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9893,9896|false|false|false|C0017040|Gamma-glutamyl transferase|ggt
Drug|Enzyme|SIMPLE_SEGMENT|9893,9896|false|false|false|C0017040|Gamma-glutamyl transferase|ggt
Event|Event|SIMPLE_SEGMENT|9893,9896|false|false|false|||ggt
Finding|Gene or Genome|SIMPLE_SEGMENT|9893,9896|false|false|false|C1415053;C1415054|GGT1 gene;GGT2P gene|ggt
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9893,9896|false|false|false|C0202035|Gamma glutamyl transferase measurement|ggt
Event|Event|SIMPLE_SEGMENT|9904,9910|false|false|false|||needed
Event|Event|SIMPLE_SEGMENT|9915,9925|false|false|false|||procedures
Finding|Functional Concept|SIMPLE_SEGMENT|9915,9925|false|false|false|C0025664;C2700391|Methods aspects;Procedure (set of actions)|procedures
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9915,9925|false|false|false|C0184661|Interventional procedure|procedures
Event|Event|SIMPLE_SEGMENT|9935,9947|false|false|false|||transitioned
Drug|Organic Chemical|SIMPLE_SEGMENT|9956,9963|false|false|false|C0728963|Lovenox|lovenox
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9956,9963|false|false|false|C0728963|Lovenox|lovenox
Event|Event|SIMPLE_SEGMENT|9956,9963|false|false|false|||lovenox
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9973,9978|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|9973,9978|false|false|false|C2003888|Lower (action)|lower
Event|Event|SIMPLE_SEGMENT|9979,9983|false|false|false|||dose
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9988,9994|false|false|false|C0944911||weight
Event|Event|SIMPLE_SEGMENT|9988,9994|false|false|false|||weight
Finding|Finding|SIMPLE_SEGMENT|9988,9994|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|SIMPLE_SEGMENT|9988,9994|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|SIMPLE_SEGMENT|9988,9994|false|false|false|C1305866|Weighing patient|weight
Event|Event|SIMPLE_SEGMENT|9996,10002|false|false|false|||dosing
Event|Event|SIMPLE_SEGMENT|10021,10030|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|10021,10030|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|10021,10030|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|10021,10030|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|10021,10030|false|false|false|C0030685|Patient Discharge|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|10035,10040|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|Acute
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|10035,10053|false|false|false|C2609414|Acute kidney injury|Acute renal injury
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10041,10046|false|false|false|C0022646|Kidney|renal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10041,10046|false|false|false|C0042075|Urologic Diseases|renal
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|10041,10053|false|false|false|C0160420|Injury of kidney|renal injury
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|10047,10053|false|false|false|C3263722;C3263723|Traumatic AND/OR non-traumatic injury;Traumatic injury|injury
Event|Event|SIMPLE_SEGMENT|10047,10053|false|false|false|||injury
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10055,10058|false|false|false|C5239292|Solitary Cutaneous Reticulohistiocytosis|SCr
Event|Event|SIMPLE_SEGMENT|10055,10058|false|false|false|||SCr
Finding|Finding|SIMPLE_SEGMENT|10055,10058|false|false|false|C1539487;C4050416|FBXL20 gene;Stringent Complete Response|SCr
Finding|Gene or Genome|SIMPLE_SEGMENT|10055,10058|false|false|false|C1539487;C4050416|FBXL20 gene;Stringent Complete Response|SCr
Event|Event|SIMPLE_SEGMENT|10077,10083|false|false|false|||rising
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10092,10100|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|SIMPLE_SEGMENT|10092,10100|false|false|false|||baseline
Finding|Idea or Concept|SIMPLE_SEGMENT|10092,10100|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Event|Event|SIMPLE_SEGMENT|10136,10142|false|false|false|||likely
Finding|Finding|SIMPLE_SEGMENT|10136,10142|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|10136,10142|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10159,10167|false|false|false|C0042075|Urologic Diseases|uropathy
Event|Event|SIMPLE_SEGMENT|10159,10167|false|false|false|||uropathy
Finding|Gene or Genome|SIMPLE_SEGMENT|10172,10177|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Drug|Substance|SIMPLE_SEGMENT|10185,10190|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|10185,10190|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|10191,10202|false|false|false|||collections
Event|Event|SIMPLE_SEGMENT|10209,10217|false|false|false|||resolved
Finding|Idea or Concept|SIMPLE_SEGMENT|10241,10249|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|SIMPLE_SEGMENT|10250,10254|false|false|false|||stay
Finding|Idea or Concept|SIMPLE_SEGMENT|10260,10265|false|false|false|C1546485|Diagnosis Type - Final|final
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10278,10292|false|false|false|C0020295|Hydronephrosis|Hydronephrosis
Event|Event|SIMPLE_SEGMENT|10278,10292|false|false|false|||Hydronephrosis
Event|Event|SIMPLE_SEGMENT|10308,10317|false|false|false|||worsening
Finding|Intellectual Product|SIMPLE_SEGMENT|10321,10329|false|false|false|C1552654|Parameterized Data Type - Interval|interval
Event|Event|SIMPLE_SEGMENT|10330,10337|false|false|false|||imaging
Finding|Finding|SIMPLE_SEGMENT|10330,10337|false|false|false|C0740845|Imaging problem|imaging
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10330,10337|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|imaging
Event|Event|SIMPLE_SEGMENT|10350,10357|false|false|false|||studies
Procedure|Research Activity|SIMPLE_SEGMENT|10350,10357|false|false|false|C0947630|Scientific Study|studies
Finding|Body Substance|SIMPLE_SEGMENT|10365,10372|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|10365,10372|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|10365,10372|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10375,10378|false|false|false|C1114365||age
Drug|Biologically Active Substance|SIMPLE_SEGMENT|10375,10378|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|SIMPLE_SEGMENT|10375,10378|false|false|false|C0162574|Glycation End Products, Advanced|age
Event|Event|SIMPLE_SEGMENT|10375,10378|false|false|false|||age
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10389,10396|false|false|false|C0042027|Urinary tract|urinary
Event|Event|SIMPLE_SEGMENT|10398,10404|true|false|false|||output
Finding|Conceptual Entity|SIMPLE_SEGMENT|10398,10404|true|false|false|C1709366|system output|output
Procedure|Health Care Activity|SIMPLE_SEGMENT|10398,10404|true|false|false|C3251815|Measurement of fluid output|output
Drug|Biologically Active Substance|SIMPLE_SEGMENT|10415,10425|true|false|false|C0010294|creatinine|creatinine
Drug|Organic Chemical|SIMPLE_SEGMENT|10415,10425|true|false|false|C0010294|creatinine|creatinine
Event|Event|SIMPLE_SEGMENT|10415,10425|true|false|false|||creatinine
Finding|Physiologic Function|SIMPLE_SEGMENT|10415,10425|true|false|false|C4551889|Creatinine metabolic function|creatinine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10415,10425|true|false|false|C0201975|Creatinine measurement|creatinine
Phenomenon|Biologic Function|SIMPLE_SEGMENT|10415,10435|true|false|false|C0812399|Creatinine clearance|creatinine clearance
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10415,10435|true|false|false|C0373595|Creatinine renal clearance measurement|creatinine clearance
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10426,10435|true|false|false|C1382187|Clearance of substance|clearance
Event|Event|SIMPLE_SEGMENT|10426,10435|true|false|false|||clearance
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|10426,10435|true|false|false|C2825073|Clearance [PK]|clearance
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10426,10435|true|false|false|C4554548|Clearance procedure|clearance
Event|Event|SIMPLE_SEGMENT|10444,10455|true|false|false|||significant
Finding|Idea or Concept|SIMPLE_SEGMENT|10444,10455|true|false|false|C0750502|Significant|significant
Drug|Inorganic Chemical|SIMPLE_SEGMENT|10457,10468|true|false|false|C0013832;C3536863|Electrolyte [EPC];Electrolytes|electrolyte
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10457,10468|true|false|false|C0013832;C3536863|Electrolyte [EPC];Electrolytes|electrolyte
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|10469,10482|true|false|false|C0000768|Congenital Abnormality|abnormalities
Event|Event|SIMPLE_SEGMENT|10469,10482|true|false|false|||abnormalities
Finding|Functional Concept|SIMPLE_SEGMENT|10469,10482|true|false|false|C0000769|teratologic|abnormalities
Finding|Body Substance|SIMPLE_SEGMENT|10484,10491|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|10484,10491|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|10484,10491|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Finding|SIMPLE_SEGMENT|10492,10498|true|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|10492,10498|true|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|SIMPLE_SEGMENT|10524,10531|true|false|false|||benefit
Event|Event|SIMPLE_SEGMENT|10537,10549|true|false|false|||intervention
Procedure|Health Care Activity|SIMPLE_SEGMENT|10537,10549|true|false|false|C0184661;C0886296;C1273869|Intervention regimes;Interventional procedure;Nursing interventions|intervention
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10537,10549|true|false|false|C0184661;C0886296;C1273869|Intervention regimes;Interventional procedure;Nursing interventions|intervention
Finding|Finding|SIMPLE_SEGMENT|10558,10562|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|10558,10562|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|10558,10562|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Anatomy|Body Location or Region|SIMPLE_SEGMENT|10564,10567|false|false|false|C0449201|PER (body structure)|Per
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10564,10567|false|false|false|C1861457|PROGRESSIVE ENCEPHALOMYELITIS WITH RIGIDITY|Per
Event|Event|SIMPLE_SEGMENT|10564,10567|false|false|false|||Per
Finding|Functional Concept|SIMPLE_SEGMENT|10564,10567|false|false|false|C1418464;C1704764;C3273590;C4281991|Follow;PER1 gene;PER1 wt Allele;Per - dosing instruction fragment|Per
Finding|Gene or Genome|SIMPLE_SEGMENT|10564,10567|false|false|false|C1418464;C1704764;C3273590;C4281991|Follow;PER1 gene;PER1 wt Allele;Per - dosing instruction fragment|Per
Finding|Intellectual Product|SIMPLE_SEGMENT|10564,10567|false|false|false|C1418464;C1704764;C3273590;C4281991|Follow;PER1 gene;PER1 wt Allele;Per - dosing instruction fragment|Per
Event|Event|SIMPLE_SEGMENT|10577,10584|false|false|false|||consult
Procedure|Health Care Activity|SIMPLE_SEGMENT|10577,10584|false|false|false|C0009818|Consultation|consult
Event|Event|SIMPLE_SEGMENT|10586,10592|false|false|false|||deemed
Event|Event|SIMPLE_SEGMENT|10593,10599|false|false|false|||stable
Finding|Intellectual Product|SIMPLE_SEGMENT|10593,10599|false|false|false|C1547311|Patient Condition Code - Stable|stable
Event|Event|SIMPLE_SEGMENT|10604,10613|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|10604,10613|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|10604,10613|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|10604,10613|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|10604,10613|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|SIMPLE_SEGMENT|10618,10629|false|false|false|||recommended
Finding|Idea or Concept|SIMPLE_SEGMENT|10618,10629|false|false|false|C0034866|Recommendation|recommended
Finding|Classification|SIMPLE_SEGMENT|10631,10641|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|10631,10641|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|SIMPLE_SEGMENT|10650,10658|false|false|false|||followup
Procedure|Health Care Activity|SIMPLE_SEGMENT|10650,10658|false|false|false|C1522577|follow-up|followup
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10663,10669|false|false|false|C0002871|Anemia|Anemia
Event|Event|SIMPLE_SEGMENT|10663,10669|false|false|false|||Anemia
Finding|Finding|SIMPLE_SEGMENT|10671,10677|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|10671,10677|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|SIMPLE_SEGMENT|10680,10691|false|false|false|||combination
Finding|Finding|SIMPLE_SEGMENT|10680,10691|false|true|false|C3811910|combination - answer to question|combination
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10695,10701|false|false|false|C0002871|Anemia|anemia
Event|Event|SIMPLE_SEGMENT|10695,10701|false|false|false|||anemia
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10695,10725|false|false|false|C0002873|Anemia of chronic disease|anemia of chronic inflammation
Finding|Intellectual Product|SIMPLE_SEGMENT|10705,10712|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|10705,10712|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Finding|Pathologic Function|SIMPLE_SEGMENT|10705,10725|false|false|false|C0021376|Chronic inflammation|chronic inflammation
Event|Event|SIMPLE_SEGMENT|10713,10725|false|false|false|||inflammation
Finding|Pathologic Function|SIMPLE_SEGMENT|10713,10725|false|false|false|C0021368|Inflammation|inflammation
Finding|Intellectual Product|SIMPLE_SEGMENT|10731,10736|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Pathologic Function|SIMPLE_SEGMENT|10731,10747|false|false|false|C0333276|Acute hemorrhage|acute blood loss
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10737,10742|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|10737,10742|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|10737,10742|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Finding|SIMPLE_SEGMENT|10737,10747|false|false|false|C0019080;C3163616|Blood Loss;Hemorrhage|blood loss
Finding|Pathologic Function|SIMPLE_SEGMENT|10737,10747|false|false|false|C0019080;C3163616|Blood Loss;Hemorrhage|blood loss
Event|Event|SIMPLE_SEGMENT|10743,10747|false|false|false|||loss
Finding|Finding|SIMPLE_SEGMENT|10743,10747|false|false|false|C5890125|Loss (adaptation)|loss
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10755,10763|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Anatomy|Body Location or Region|SIMPLE_SEGMENT|10764,10773|false|false|false|C0000726|Abdomen|abdominal
Finding|Finding|SIMPLE_SEGMENT|10764,10779|false|false|false|C2266645|abdominal drain in place|abdominal drain
Drug|Substance|SIMPLE_SEGMENT|10774,10779|false|false|false|C1550628|Drain - SpecimenType|drain
Event|Event|SIMPLE_SEGMENT|10774,10779|false|false|false|||drain
Finding|Intellectual Product|SIMPLE_SEGMENT|10774,10779|false|false|false|C1546604|Drain Specimen Code|drain
Event|Event|SIMPLE_SEGMENT|10780,10787|false|false|false|||showing
Finding|Body Substance|SIMPLE_SEGMENT|10789,10809|false|false|false|C4518404|Serosanguinous fluid|serosanguinous fluid
Drug|Substance|SIMPLE_SEGMENT|10804,10809|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|10804,10809|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|10804,10809|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|10811,10815|true|false|false|||Labs
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|10811,10815|true|false|false|C0587081|Laboratory test finding|Labs
Event|Event|SIMPLE_SEGMENT|10820,10830|true|false|false|||consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|10820,10830|true|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|10820,10835|true|false|false|C0332290|Consistent with|consistent with
Event|Event|SIMPLE_SEGMENT|10836,10845|true|false|false|||hemolysis
Finding|Cell Function|SIMPLE_SEGMENT|10836,10845|true|true|false|C0019054;C1553188;C2937287;C2945560|Hemolysis (biological function);Hemolysis (disorder);Hemolysis (finding)|hemolysis
Finding|Finding|SIMPLE_SEGMENT|10836,10845|true|true|false|C0019054;C1553188;C2937287;C2945560|Hemolysis (biological function);Hemolysis (disorder);Hemolysis (finding)|hemolysis
Finding|Pathologic Function|SIMPLE_SEGMENT|10836,10845|true|true|false|C0019054;C1553188;C2937287;C2945560|Hemolysis (biological function);Hemolysis (disorder);Hemolysis (finding)|hemolysis
Event|Event|SIMPLE_SEGMENT|10848,10856|false|false|false|||Received
Event|Event|SIMPLE_SEGMENT|10890,10898|false|false|false|||response
Finding|Finding|SIMPLE_SEGMENT|10890,10898|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Intellectual Product|SIMPLE_SEGMENT|10890,10898|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Mental Process|SIMPLE_SEGMENT|10890,10898|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Body Substance|SIMPLE_SEGMENT|10900,10907|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|10900,10907|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|10900,10907|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|10913,10923|false|false|false|||discharged
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10929,10932|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|10929,10932|false|false|false|C0019046|Hemoglobin|Hgb
Event|Event|SIMPLE_SEGMENT|10929,10932|false|false|false|||Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|10929,10932|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|10929,10932|false|false|false|C0019029|Hemoglobin concentration|Hgb
Event|Event|SIMPLE_SEGMENT|10944,10947|false|false|false|||hem
Finding|Pathologic Function|SIMPLE_SEGMENT|10944,10947|false|false|false|C0019080|Hemorrhage|hem
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10944,10947|false|false|false|C0280599|altretamine/etoposide/methotrexate protocol|hem
Event|Event|SIMPLE_SEGMENT|10952,10966|false|false|false|||recommendation
Finding|Idea or Concept|SIMPLE_SEGMENT|10952,10966|false|false|false|C0034866|Recommendation|recommendation
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10982,10985|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|10982,10985|false|false|false|C0019046|Hemoglobin|Hgb
Event|Event|SIMPLE_SEGMENT|10982,10985|false|false|false|||Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|10982,10985|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|10982,10985|false|false|false|C0019029|Hemoglobin concentration|Hgb
Finding|Body Substance|SIMPLE_SEGMENT|10991,10998|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|10991,10998|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|10991,10998|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|10999,11004|false|false|false|||feels
Event|Event|SIMPLE_SEGMENT|11022,11030|false|false|false|||performs
Event|Event|SIMPLE_SEGMENT|11032,11038|false|false|false|||better
Finding|Idea or Concept|SIMPLE_SEGMENT|11032,11038|false|false|false|C1550462|Observation Interpretation - better|better
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11051,11056|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|11051,11056|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|11051,11056|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Event|Event|SIMPLE_SEGMENT|11057,11063|false|false|false|||counts
Event|Event|SIMPLE_SEGMENT|11068,11079|false|false|false|||Hypokalemia
Finding|Finding|SIMPLE_SEGMENT|11068,11079|false|false|false|C0020621|Hypokalemia|Hypokalemia
Event|Event|SIMPLE_SEGMENT|11085,11096|false|false|false|||hypokalemic
Event|Event|SIMPLE_SEGMENT|11105,11113|false|false|false|||repleted
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|11119,11123|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|11119,11123|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|11119,11123|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|11119,11123|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Drug|Inorganic Chemical|SIMPLE_SEGMENT|11124,11127|false|false|false|C0032825|potassium chloride|KCl
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11124,11127|false|false|false|C0032825|potassium chloride|KCl
Event|Event|SIMPLE_SEGMENT|11124,11127|false|false|false|||KCl
Event|Event|SIMPLE_SEGMENT|11129,11132|false|false|false|||PRN
Finding|Gene or Genome|SIMPLE_SEGMENT|11129,11132|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|SIMPLE_SEGMENT|11136,11143|false|false|false|||CHRONIC
Finding|Intellectual Product|SIMPLE_SEGMENT|11136,11143|false|false|false|C1547296|Chronic - Admission Level of Care Code|CHRONIC
Procedure|Health Care Activity|SIMPLE_SEGMENT|11136,11143|false|false|false|C1555457|Provision of recurring care for chronic illness|CHRONIC
Finding|Finding|SIMPLE_SEGMENT|11178,11182|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|SIMPLE_SEGMENT|11178,11182|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|SIMPLE_SEGMENT|11178,11182|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Disorder|Neoplastic Process|SIMPLE_SEGMENT|11178,11209|false|false|false|C5556496|Urothelial Carcinoma, High Grade|high-grade urothelial carcinoma
Finding|Classification|SIMPLE_SEGMENT|11183,11188|false|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|grade
Finding|Finding|SIMPLE_SEGMENT|11183,11188|false|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|grade
Disorder|Neoplastic Process|SIMPLE_SEGMENT|11189,11209|false|false|false|C0007138;C2145472|Carcinoma, Transitional Cell;Urothelial Carcinoma|urothelial carcinoma
Disorder|Neoplastic Process|SIMPLE_SEGMENT|11200,11209|false|false|false|C0007097|Carcinoma|carcinoma
Event|Event|SIMPLE_SEGMENT|11200,11209|false|false|false|||carcinoma
Event|Event|SIMPLE_SEGMENT|11211,11220|false|false|false|||involving
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11225,11229|false|false|false|C4318566|Deep Resection Margin|deep
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11231,11241|false|false|false|C0225358;C4551532|Bladder Detrusor Muscle;Muscle layer|muscularis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11231,11249|false|false|false|C0225358|Bladder Detrusor Muscle|muscularis propria
Event|Event|SIMPLE_SEGMENT|11254,11264|false|false|false|||cystectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11254,11264|false|false|false|C0010651|Cystectomy|cystectomy
Event|Event|SIMPLE_SEGMENT|11266,11278|false|false|false|||hysterectomy
Finding|Finding|SIMPLE_SEGMENT|11266,11278|false|false|false|C1548863|Consent Type - Hysterectomy|hysterectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11266,11278|false|false|false|C0020699|Hysterectomy|hysterectomy
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|11284,11287|false|false|false|C0054252|Buthionine Sulfoximine|BSO
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|11284,11287|false|false|false|C0054252|Buthionine Sulfoximine|BSO
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11284,11287|false|false|false|C0054252|Buthionine Sulfoximine|BSO
Event|Event|SIMPLE_SEGMENT|11284,11287|false|false|false|||BSO
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11297,11302|false|false|false|C0020885|ileum|ileal
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|11297,11310|false|false|false|C0441253|Structure of ileal conduit|ileal conduit
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11297,11310|false|false|false|C0348002|Ileal conduit procedure|ileal conduit
Event|Event|SIMPLE_SEGMENT|11303,11310|false|false|false|||conduit
Finding|Finding|SIMPLE_SEGMENT|11319,11333|false|false|false|C0241311|post operative (finding)|post operative
Event|Event|SIMPLE_SEGMENT|11334,11340|false|false|false|||course
Event|Event|SIMPLE_SEGMENT|11350,11361|false|false|false|||complicated
Anatomy|Body Location or Region|SIMPLE_SEGMENT|11365,11368|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11365,11368|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11365,11368|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11374,11379|false|false|false|C1258215;C4019039|Ileus;Intestinal obstruction co-occurrent and due to decreased peristalsis|ileus
Event|Event|SIMPLE_SEGMENT|11374,11379|false|false|false|||ileus
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11385,11391|false|false|false|C0030797|Pelvis|pelvic
Drug|Substance|SIMPLE_SEGMENT|11392,11397|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|11392,11397|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|11398,11409|false|false|false|||collections
Finding|Body Substance|SIMPLE_SEGMENT|11412,11419|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|11412,11419|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|11412,11419|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|11420,11427|true|false|false|||stating
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11446,11450|true|false|false|C0270724|Infantile Neuroaxonal Dystrophy|plan
Event|Event|SIMPLE_SEGMENT|11446,11450|true|false|false|||plan
Finding|Functional Concept|SIMPLE_SEGMENT|11446,11450|true|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Intellectual Product|SIMPLE_SEGMENT|11446,11450|true|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Mental Process|SIMPLE_SEGMENT|11446,11450|true|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Event|Event|SIMPLE_SEGMENT|11455,11460|true|false|false|||chemo
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11455,11460|true|false|false|C0392920;C3665472|Chemotherapy;Chemotherapy Regimen|chemo
Event|Event|SIMPLE_SEGMENT|11465,11474|true|false|false|||radiation
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|11465,11474|true|false|false|C0034519;C0851346|Electromagnetic Radiation;Radiation|radiation
Procedure|Research Activity|SIMPLE_SEGMENT|11465,11474|true|false|false|C1522449;C1524020;C1524021|Radiation Ionizing Radiotherapy;Radiation therapy (procedure);Radiotherapy Research|radiation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11465,11474|true|false|false|C1522449;C1524020;C1524021|Radiation Ionizing Radiotherapy;Radiation therapy (procedure);Radiotherapy Research|radiation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|11480,11483|false|false|false|C0032743;C0040398|Positron-Emission Tomography;Tomography, Emission-Computed|PET
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|11480,11488|false|false|false|C0032743|Positron-Emission Tomography|PET scan
Event|Event|SIMPLE_SEGMENT|11484,11488|false|false|false|||scan
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|11484,11488|false|false|false|C0034606;C0441633|Radionuclide Imaging;Scanning|scan
Event|Event|SIMPLE_SEGMENT|11494,11498|false|false|false|||show
Event|Event|SIMPLE_SEGMENT|11511,11515|false|false|false|||foci
Finding|Finding|SIMPLE_SEGMENT|11511,11515|false|false|false|C4321394|Foci|foci
Finding|Functional Concept|SIMPLE_SEGMENT|11519,11529|false|false|false|C0036525;C1522484|Metastatic to;metastatic qualifier|metastatic
Disorder|Neoplastic Process|SIMPLE_SEGMENT|11519,11537|false|false|false|C0027627;C2939419;C2939420|Metastatic Neoplasm;Metastatic malignant neoplasm;Neoplasm Metastasis|metastatic disease
Finding|Finding|SIMPLE_SEGMENT|11519,11537|false|false|false|C1513183|Metastatic Lesion|metastatic disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11530,11537|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|11530,11537|false|false|false|||disease
Anatomy|Body Location or Region|SIMPLE_SEGMENT|11545,11549|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11545,11549|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11545,11549|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|SIMPLE_SEGMENT|11545,11549|false|false|false|C0740941|Lung Problem|lung
Anatomy|Tissue|SIMPLE_SEGMENT|11555,11565|false|false|false|C0031153;C0230198;C4482223|Abdomen>Peritoneum;Peritoneum;Serous layer of peritoneum|peritoneum
Disorder|Neoplastic Process|SIMPLE_SEGMENT|11555,11565|false|false|false|C0496874;C0496954|Benign neoplasm of peritoneum;Neoplasm of uncertain or unknown behavior of peritoneum|peritoneum
Event|Event|SIMPLE_SEGMENT|11555,11565|false|false|false|||peritoneum
Finding|Body Substance|SIMPLE_SEGMENT|11571,11578|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|11571,11578|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|11571,11578|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Gene or Genome|SIMPLE_SEGMENT|11581,11584|false|false|false|C1420310|SON gene|son
Event|Event|SIMPLE_SEGMENT|11599,11603|false|false|false|||seen
Event|Event|SIMPLE_SEGMENT|11606,11612|false|false|false|||doctor
Finding|Intellectual Product|SIMPLE_SEGMENT|11606,11612|false|false|false|C2348314|Doctor - Title|doctor
Event|Event|SIMPLE_SEGMENT|11617,11621|false|false|false|||work
Event|Occupational Activity|SIMPLE_SEGMENT|11617,11621|false|false|false|C0043227|Work|work
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|11617,11624|false|false|false|C0750430|Work-up|work up
Anatomy|Body Location or Region|SIMPLE_SEGMENT|11629,11633|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11629,11633|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11629,11633|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|SIMPLE_SEGMENT|11629,11633|false|false|false|C0740941|Lung Problem|lung
Finding|Finding|SIMPLE_SEGMENT|11629,11638|false|false|false|C0149726|Lung mass|lung mass
Event|Event|SIMPLE_SEGMENT|11634,11638|false|false|false|||mass
Finding|Finding|SIMPLE_SEGMENT|11634,11638|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|SIMPLE_SEGMENT|11634,11638|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|SIMPLE_SEGMENT|11634,11638|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Idea or Concept|SIMPLE_SEGMENT|11650,11657|false|false|false|C0549178|Continuous|ongoing
Event|Event|SIMPLE_SEGMENT|11658,11668|false|false|false|||discussion
Finding|Social Behavior|SIMPLE_SEGMENT|11658,11668|false|false|false|C2584313|Discussion (communication)|discussion
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11658,11668|false|false|false|C0557061|Discussion (procedure)|discussion
Finding|Classification|SIMPLE_SEGMENT|11675,11685|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|11675,11685|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|SIMPLE_SEGMENT|11686,11689|false|false|false|||hem
Finding|Pathologic Function|SIMPLE_SEGMENT|11686,11689|false|false|false|C0019080|Hemorrhage|hem
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11686,11689|false|false|false|C0280599|altretamine/etoposide/methotrexate protocol|hem
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11711,11715|false|false|false|C0339510|Vitelliform Macular Dystrophy|best
Finding|Gene or Genome|SIMPLE_SEGMENT|11711,11715|false|false|false|C1826421;C5781213|BEST1 gene;BEST1 wt Allele|best
Event|Event|SIMPLE_SEGMENT|11716,11722|false|false|false|||manage
Event|Event|SIMPLE_SEGMENT|11723,11733|false|false|false|||concerning
Event|Event|SIMPLE_SEGMENT|11735,11742|false|false|false|||lesions
Finding|Finding|SIMPLE_SEGMENT|11735,11742|false|false|false|C0221198|Lesion|lesions
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11747,11753|false|false|false|C0006141|Breast|Breast
Disorder|Neoplastic Process|SIMPLE_SEGMENT|11747,11753|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|Breast
Event|Event|SIMPLE_SEGMENT|11747,11753|false|false|false|||Breast
Finding|Finding|SIMPLE_SEGMENT|11747,11753|false|false|false|C0567499|Breast problem|Breast
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11747,11753|false|false|false|C0191838|Procedures on breast|Breast
Finding|Finding|SIMPLE_SEGMENT|11747,11758|false|false|false|C0024103|Mass in breast|Breast mass
Event|Event|SIMPLE_SEGMENT|11754,11758|false|false|false|||mass
Finding|Finding|SIMPLE_SEGMENT|11754,11758|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|SIMPLE_SEGMENT|11754,11758|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|SIMPLE_SEGMENT|11754,11758|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Event|Event|SIMPLE_SEGMENT|11763,11772|false|false|false|||mammogram
Finding|Finding|SIMPLE_SEGMENT|11763,11772|false|false|false|C0260913|Encounter due to Screening for malignant neoplasm of breast|mammogram
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|11763,11772|false|false|false|C0024671|Mammography|mammogram
Event|Event|SIMPLE_SEGMENT|11773,11780|false|false|false|||showing
Finding|Intellectual Product|SIMPLE_SEGMENT|11781,11788|false|false|false|C1511314|Breast Imaging Reporting and Data System|BI-RADS
Finding|Intellectual Product|SIMPLE_SEGMENT|11781,11790|false|false|false|C5960924|Breast Imaging-Reporting and Data System Assessment Category 5|BI-RADS 5
Event|Event|SIMPLE_SEGMENT|11789,11790|false|false|false|||5
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|11792,11797|false|false|false|C0302909;C1378566|Solid Dose Form;solid substance|Solid
Drug|Substance|SIMPLE_SEGMENT|11792,11797|false|false|false|C0302909;C1378566|Solid Dose Form;solid substance|Solid
Event|Event|SIMPLE_SEGMENT|11798,11802|false|false|false|||mass
Finding|Finding|SIMPLE_SEGMENT|11798,11802|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|SIMPLE_SEGMENT|11798,11802|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|SIMPLE_SEGMENT|11798,11802|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|11815,11820|false|false|false|C1743089|CLOCK protein, human|clock
Drug|Enzyme|SIMPLE_SEGMENT|11815,11820|false|false|false|C1743089|CLOCK protein, human|clock
Finding|Gene or Genome|SIMPLE_SEGMENT|11815,11820|false|false|false|C1413503|CLOCK gene|clock
Finding|Functional Concept|SIMPLE_SEGMENT|11821,11825|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11821,11832|false|false|false|C0222601|Left breast|left breast
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11826,11832|false|false|false|C0006141|Breast|breast
Disorder|Neoplastic Process|SIMPLE_SEGMENT|11826,11832|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|breast
Event|Event|SIMPLE_SEGMENT|11826,11832|false|false|false|||breast
Finding|Finding|SIMPLE_SEGMENT|11826,11832|false|false|false|C0567499|Breast problem|breast
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11826,11832|false|false|false|C0191838|Procedures on breast|breast
Event|Event|SIMPLE_SEGMENT|11838,11846|false|false|false|||features
Finding|Finding|SIMPLE_SEGMENT|11860,11885|false|false|false|C4050405|Suspicious for Malignancy|suspicious for malignancy
Disorder|Neoplastic Process|SIMPLE_SEGMENT|11875,11885|false|true|false|C0006826;C1306459|Malignant Neoplasms;Primary malignant neoplasm|malignancy
Event|Event|SIMPLE_SEGMENT|11875,11885|false|false|false|||malignancy
Finding|Body Substance|SIMPLE_SEGMENT|11891,11898|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|11891,11898|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|11891,11898|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Gene or Genome|SIMPLE_SEGMENT|11901,11904|false|false|false|C1420310|SON gene|son
Event|Event|SIMPLE_SEGMENT|11914,11918|false|false|false|||seen
Event|Event|SIMPLE_SEGMENT|11922,11928|false|false|false|||doctor
Finding|Intellectual Product|SIMPLE_SEGMENT|11922,11928|false|false|false|C2348314|Doctor - Title|doctor
Event|Event|SIMPLE_SEGMENT|11933,11943|false|false|false|||evaluating
Finding|Finding|SIMPLE_SEGMENT|11948,11951|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|11948,11951|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11952,11958|false|false|false|C0006141|Breast|breast
Disorder|Neoplastic Process|SIMPLE_SEGMENT|11952,11958|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|breast
Finding|Finding|SIMPLE_SEGMENT|11952,11958|false|false|false|C0567499|Breast problem|breast
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11952,11958|false|false|false|C0191838|Procedures on breast|breast
Finding|Finding|SIMPLE_SEGMENT|11952,11963|false|false|false|C0024103|Mass in breast|breast mass
Event|Event|SIMPLE_SEGMENT|11959,11963|false|false|false|||mass
Finding|Finding|SIMPLE_SEGMENT|11959,11963|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|SIMPLE_SEGMENT|11959,11963|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|SIMPLE_SEGMENT|11959,11963|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Event|Event|SIMPLE_SEGMENT|11971,11980|false|false|false|||recommend
Finding|Idea or Concept|SIMPLE_SEGMENT|11982,11989|false|false|false|C0549178|Continuous|ongoing
Event|Event|SIMPLE_SEGMENT|11990,12000|false|false|false|||discussion
Finding|Social Behavior|SIMPLE_SEGMENT|11990,12000|false|false|false|C2584313|Discussion (communication)|discussion
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11990,12000|false|false|false|C0557061|Discussion (procedure)|discussion
Event|Event|SIMPLE_SEGMENT|12021,12027|false|false|false|||doctor
Finding|Intellectual Product|SIMPLE_SEGMENT|12021,12027|false|false|true|C2348314|Doctor - Title|doctor
Event|Event|SIMPLE_SEGMENT|12032,12042|false|false|false|||outpatient
Finding|Classification|SIMPLE_SEGMENT|12032,12042|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|12032,12042|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12058,12062|false|false|false|C0270724|Infantile Neuroaxonal Dystrophy|plan
Event|Event|SIMPLE_SEGMENT|12058,12062|false|false|false|||plan
Finding|Functional Concept|SIMPLE_SEGMENT|12058,12062|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Intellectual Product|SIMPLE_SEGMENT|12058,12062|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Mental Process|SIMPLE_SEGMENT|12058,12062|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Event|Event|SIMPLE_SEGMENT|12066,12072|false|false|false|||manage
Event|Event|SIMPLE_SEGMENT|12077,12080|false|false|false|||HLD
Event|Event|SIMPLE_SEGMENT|12082,12091|true|false|false|||continued
Drug|Organic Chemical|SIMPLE_SEGMENT|12092,12104|true|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12092,12104|true|false|false|C0286651|atorvastatin|atorvastatin
Event|Event|SIMPLE_SEGMENT|12092,12104|true|false|false|||atorvastatin
Event|Event|SIMPLE_SEGMENT|12113,12120|true|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|12113,12120|true|false|false|C0392747|Changing|changes
Finding|Idea or Concept|SIMPLE_SEGMENT|12122,12130|false|false|false|C0750591|consider|Consider
Event|Event|SIMPLE_SEGMENT|12132,12142|false|false|false|||evaluation
Finding|Idea or Concept|SIMPLE_SEGMENT|12132,12142|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|SIMPLE_SEGMENT|12132,12142|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Drug|Inorganic Chemical|SIMPLE_SEGMENT|12153,12161|false|false|false|C0723457|Stop brand of fluoride|stopping
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12153,12161|false|false|false|C0723457|Stop brand of fluoride|stopping
Event|Event|SIMPLE_SEGMENT|12153,12161|false|false|false|||stopping
Drug|Organic Chemical|SIMPLE_SEGMENT|12162,12174|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12162,12174|false|false|false|C0286651|atorvastatin|atorvastatin
Event|Event|SIMPLE_SEGMENT|12162,12174|false|false|false|||atorvastatin
Finding|Classification|SIMPLE_SEGMENT|12178,12188|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|12178,12188|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12189,12194|false|false|false|C1874451|Basis|basis
Event|Event|SIMPLE_SEGMENT|12189,12194|false|false|false|||basis
Finding|Functional Concept|SIMPLE_SEGMENT|12189,12194|false|false|false|C1527178|Basis - conceptual entity|basis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12200,12214|false|false|false|C0020676|Hypothyroidism|Hypothyroidism
Event|Event|SIMPLE_SEGMENT|12200,12214|false|false|false|||Hypothyroidism
Event|Event|SIMPLE_SEGMENT|12216,12225|true|false|false|||continued
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|12226,12239|true|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Hormone|SIMPLE_SEGMENT|12226,12239|true|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Organic Chemical|SIMPLE_SEGMENT|12226,12239|true|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12226,12239|true|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Event|Event|SIMPLE_SEGMENT|12226,12239|true|false|false|||levothyroxine
Event|Event|SIMPLE_SEGMENT|12248,12255|true|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|12248,12255|true|false|false|C0392747|Changing|changes
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12264,12267|false|false|false|C0162531|Hereditary Coproporphyria|HCP
Event|Event|SIMPLE_SEGMENT|12264,12267|false|false|false|||HCP
Finding|Gene or Genome|SIMPLE_SEGMENT|12264,12267|false|false|false|C1335283;C1412376;C1413681;C1705637;C5780748|AMBP gene;AMBP wt Allele;CPOX gene;PTPN6 gene;PTPN6 wt Allele|HCP
Finding|Gene or Genome|SIMPLE_SEGMENT|12279,12282|false|false|false|C1420310|SON gene|son
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12288,12297|false|false|false|C0804815||physician
Event|Occupational Activity|SIMPLE_SEGMENT|12304,12308|false|false|false|C0009219|Coding|Code
Finding|Intellectual Product|SIMPLE_SEGMENT|12304,12308|false|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|Code
Procedure|Health Care Activity|SIMPLE_SEGMENT|12304,12315|false|false|false|C0742531|CODE STATUS|Code status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12309,12315|false|false|false|C5889824||status
Event|Event|SIMPLE_SEGMENT|12309,12315|false|false|false|||status
Finding|Idea or Concept|SIMPLE_SEGMENT|12309,12315|false|false|false|C1546481|What subject filter - Status|status
Event|Event|SIMPLE_SEGMENT|12322,12326|false|false|false|||code
Event|Occupational Activity|SIMPLE_SEGMENT|12322,12326|false|false|false|C0009219|Coding|code
Finding|Intellectual Product|SIMPLE_SEGMENT|12322,12326|false|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|code
Event|Event|SIMPLE_SEGMENT|12328,12337|false|false|false|||confirmed
Finding|Body Substance|SIMPLE_SEGMENT|12343,12350|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|12343,12350|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|12343,12350|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|12360,12372|false|false|false|C1548597|Marketing basis - Transitional|TRANSITIONAL
Event|Event|SIMPLE_SEGMENT|12373,12379|false|false|false|||ISSUES
Event|Event|SIMPLE_SEGMENT|12411,12415|false|false|false|||need
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12416,12426|false|false|false|C0009450|Communicable Diseases|infectious
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12416,12434|false|false|false|C0009450|Communicable Diseases|infectious disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12427,12434|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|12427,12434|false|false|false|||disease
Event|Event|SIMPLE_SEGMENT|12435,12441|false|false|false|||follow
Finding|Functional Concept|SIMPLE_SEGMENT|12435,12441|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|SIMPLE_SEGMENT|12435,12441|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|SIMPLE_SEGMENT|12435,12444|false|false|false|C0589120|Follow-up status|follow up
Procedure|Health Care Activity|SIMPLE_SEGMENT|12435,12444|false|false|false|C1522577|follow-up|follow up
Event|Event|SIMPLE_SEGMENT|12442,12444|false|false|false|||up
Event|Event|SIMPLE_SEGMENT|12498,12502|false|false|false|||call
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|12511,12514|false|false|false|C1137947|SET protein, human|set
Drug|Biologically Active Substance|SIMPLE_SEGMENT|12511,12514|false|false|false|C1137947|SET protein, human|set
Event|Event|SIMPLE_SEGMENT|12511,12514|false|false|false|||set
Finding|Conceptual Entity|SIMPLE_SEGMENT|12511,12514|false|false|false|C0036849;C1366517;C1442518;C1552652;C1705195|Parameterized Data Type - Set;SET gene;Set (Psychology);Set scale;set (group)|set
Finding|Functional Concept|SIMPLE_SEGMENT|12511,12514|false|false|false|C0036849;C1366517;C1442518;C1552652;C1705195|Parameterized Data Type - Set;SET gene;Set (Psychology);Set scale;set (group)|set
Finding|Gene or Genome|SIMPLE_SEGMENT|12511,12514|false|false|false|C0036849;C1366517;C1442518;C1552652;C1705195|Parameterized Data Type - Set;SET gene;Set (Psychology);Set scale;set (group)|set
Finding|Idea or Concept|SIMPLE_SEGMENT|12511,12514|false|false|false|C0036849;C1366517;C1442518;C1552652;C1705195|Parameterized Data Type - Set;SET gene;Set (Psychology);Set scale;set (group)|set
Finding|Mental Process|SIMPLE_SEGMENT|12511,12514|false|false|false|C0036849;C1366517;C1442518;C1552652;C1705195|Parameterized Data Type - Set;SET gene;Set (Psychology);Set scale;set (group)|set
Event|Activity|SIMPLE_SEGMENT|12511,12517|false|false|false|C1521827|Preparation|set up
Event|Activity|SIMPLE_SEGMENT|12521,12532|false|false|false|C0003629|Appointments|appointment
Event|Event|SIMPLE_SEGMENT|12521,12532|false|false|false|||appointment
Event|Activity|SIMPLE_SEGMENT|12541,12552|false|false|false|C0003629|Appointments|appointment
Event|Event|SIMPLE_SEGMENT|12541,12552|false|false|false|||appointment
Event|Event|SIMPLE_SEGMENT|12576,12578|false|false|false|||CT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12576,12586|false|false|false|C1644645||CT abdomen
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|12576,12586|false|false|false|C0412620|CT of abdomen|CT abdomen
Anatomy|Body Location or Region|SIMPLE_SEGMENT|12579,12586|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|abdomen
Disorder|Neoplastic Process|SIMPLE_SEGMENT|12579,12586|false|false|false|C0153662|Malignant neoplasm of abdomen|abdomen
Finding|Finding|SIMPLE_SEGMENT|12579,12586|false|false|false|C0941288|Abdomen problem|abdomen
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|12587,12593|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|12587,12593|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Disorder|Neoplastic Process|SIMPLE_SEGMENT|12587,12593|false|false|false|C0153663|Malignant neoplasm of pelvis|pelvis
Finding|Finding|SIMPLE_SEGMENT|12587,12593|false|false|false|C0812455|Pelvis problem|pelvis
Event|Event|SIMPLE_SEGMENT|12621,12627|false|false|false|||Assure
Event|Event|SIMPLE_SEGMENT|12649,12651|false|false|false|||CT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12649,12659|false|false|false|C1644645||CT abdomen
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|12649,12659|false|false|false|C0412620|CT of abdomen|CT abdomen
Anatomy|Body Location or Region|SIMPLE_SEGMENT|12652,12659|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|abdomen
Disorder|Neoplastic Process|SIMPLE_SEGMENT|12652,12659|false|false|false|C0153662|Malignant neoplasm of abdomen|abdomen
Event|Event|SIMPLE_SEGMENT|12652,12659|false|false|false|||abdomen
Finding|Finding|SIMPLE_SEGMENT|12652,12659|false|false|false|C0941288|Abdomen problem|abdomen
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|12662,12668|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|12662,12668|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Disorder|Neoplastic Process|SIMPLE_SEGMENT|12662,12668|false|false|false|C0153663|Malignant neoplasm of pelvis|pelvis
Finding|Finding|SIMPLE_SEGMENT|12662,12668|false|false|false|C0812455|Pelvis problem|pelvis
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|12675,12683|false|false|false|C0009924|Contrast Media|contrast
Event|Event|SIMPLE_SEGMENT|12675,12683|false|false|false|||contrast
Finding|Intellectual Product|SIMPLE_SEGMENT|12691,12695|false|false|false|C1561540|Transaction counts and value totals - week|week
Finding|Gene or Genome|SIMPLE_SEGMENT|12729,12732|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|lab
Finding|Intellectual Product|SIMPLE_SEGMENT|12729,12732|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|lab
Event|Event|SIMPLE_SEGMENT|12733,12738|false|false|false|||draws
Anatomy|Cell Component|SIMPLE_SEGMENT|12757,12760|false|false|false|C2263086|Nuclear cap binding complex location|CBC
Event|Event|SIMPLE_SEGMENT|12757,12760|false|false|false|||CBC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|12757,12760|false|false|false|C0009555|Complete Blood Count|CBC
Event|Event|SIMPLE_SEGMENT|12767,12779|false|false|false|||differential
Finding|Idea or Concept|SIMPLE_SEGMENT|12767,12779|false|false|false|C1549478|Amount type - Differential|differential
Drug|Biologically Active Substance|SIMPLE_SEGMENT|12781,12784|false|false|false|C0600137|Blood Urea Nitrogen|BUN
Drug|Inorganic Chemical|SIMPLE_SEGMENT|12781,12784|false|false|false|C0600137|Blood Urea Nitrogen|BUN
Event|Event|SIMPLE_SEGMENT|12781,12784|false|false|false|||BUN
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|12781,12784|false|false|false|C0005845|Blood urea nitrogen measurement|BUN
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|12790,12793|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|SIMPLE_SEGMENT|12790,12793|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|12790,12793|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|SIMPLE_SEGMENT|12790,12793|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|SIMPLE_SEGMENT|12790,12793|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|SIMPLE_SEGMENT|12790,12793|false|false|false|||AST
Finding|Gene or Genome|SIMPLE_SEGMENT|12790,12793|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Disorder|Neoplastic Process|SIMPLE_SEGMENT|12795,12798|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|12795,12798|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|SIMPLE_SEGMENT|12795,12798|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|SIMPLE_SEGMENT|12795,12798|false|false|false|||ALT
Finding|Gene or Genome|SIMPLE_SEGMENT|12795,12798|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|SIMPLE_SEGMENT|12795,12798|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|SIMPLE_SEGMENT|12795,12798|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|12795,12798|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Event|Event|SIMPLE_SEGMENT|12800,12802|false|false|false|||TB
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|12804,12807|false|false|false|C1663627|ALK protein, human|ALK
Drug|Enzyme|SIMPLE_SEGMENT|12804,12807|false|false|false|C1663627|ALK protein, human|ALK
Event|Event|SIMPLE_SEGMENT|12804,12807|false|false|false|||ALK
Finding|Gene or Genome|SIMPLE_SEGMENT|12804,12807|false|false|false|C1332080;C1663627;C1704943|ALK gene;ALK protein, human;ALK wt Allele|ALK
Finding|Receptor|SIMPLE_SEGMENT|12804,12807|false|false|false|C1332080;C1663627;C1704943|ALK gene;ALK protein, human;ALK wt Allele|ALK
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|12804,12812|false|false|false|C0002059|Alkaline Phosphatase|ALK PHOS
Drug|Enzyme|SIMPLE_SEGMENT|12804,12812|false|false|false|C0002059|Alkaline Phosphatase|ALK PHOS
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|12804,12812|false|false|false|C0201850|Alkaline phosphatase measurement|ALK PHOS
Event|Event|SIMPLE_SEGMENT|12808,12812|false|false|false|||PHOS
Finding|Gene or Genome|SIMPLE_SEGMENT|12818,12821|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|LAB
Finding|Intellectual Product|SIMPLE_SEGMENT|12818,12821|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|LAB
Event|Activity|SIMPLE_SEGMENT|12822,12830|false|false|false|C1272683||REQUESTS
Finding|Idea or Concept|SIMPLE_SEGMENT|12842,12851|false|false|false|C1552657|Annotated - ParameterizedDataType|ANNOTATED
Event|Event|SIMPLE_SEGMENT|12879,12882|false|false|false|||FAX
Finding|Idea or Concept|SIMPLE_SEGMENT|12879,12882|false|false|false|C1547563;C1549619|Authorization Mode - Fax;Fax Number|FAX
Finding|Intellectual Product|SIMPLE_SEGMENT|12879,12882|false|false|false|C1547563;C1549619|Authorization Mode - Fax;Fax Number|FAX
Finding|Finding|SIMPLE_SEGMENT|12896,12904|false|false|false|C0332149|Possible|possible
Event|Event|SIMPLE_SEGMENT|12906,12912|false|false|false|||please
Drug|Antibiotic|SIMPLE_SEGMENT|12918,12927|false|false|false|C1120106|ertapenem|ertapenem
Drug|Organic Chemical|SIMPLE_SEGMENT|12918,12927|false|false|false|C1120106|ertapenem|ertapenem
Event|Event|SIMPLE_SEGMENT|12918,12927|false|false|false|||ertapenem
Finding|Finding|SIMPLE_SEGMENT|12937,12941|true|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|12937,12941|true|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|12937,12941|true|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|SIMPLE_SEGMENT|12958,12967|true|false|false|||interfere
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|12977,12993|true|false|false|C0871707|daily activities|daily activities
Event|Activity|SIMPLE_SEGMENT|12983,12993|true|false|false|C0441655|Activities|activities
Event|Event|SIMPLE_SEGMENT|12983,12993|true|false|false|||activities
Finding|Finding|SIMPLE_SEGMENT|12983,12993|true|false|false|C2239122|activities (history)|activities
Drug|Antibiotic|SIMPLE_SEGMENT|13031,13040|false|false|false|C1120106|ertapenem|ertapenem
Drug|Organic Chemical|SIMPLE_SEGMENT|13031,13040|false|false|false|C1120106|ertapenem|ertapenem
Event|Event|SIMPLE_SEGMENT|13031,13040|false|false|false|||ertapenem
Finding|Idea or Concept|SIMPLE_SEGMENT|13064,13069|false|false|false|C1546485|Diagnosis Type - Final|final
Event|Event|SIMPLE_SEGMENT|13070,13079|false|false|false|||treatment
Finding|Conceptual Entity|SIMPLE_SEGMENT|13070,13079|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|SIMPLE_SEGMENT|13070,13079|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|SIMPLE_SEGMENT|13070,13079|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|13070,13079|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Event|Event|SIMPLE_SEGMENT|13088,13098|false|false|false|||determined
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13106,13116|false|false|false|C0009450|Communicable Diseases|infectious
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13106,13124|false|false|false|C0009450|Communicable Diseases|infectious disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13117,13124|false|false|false|C0012634|Disease|disease
Finding|Idea or Concept|SIMPLE_SEGMENT|13146,13153|false|false|false|C0549178|Continuous|ongoing
Event|Event|SIMPLE_SEGMENT|13154,13164|false|false|false|||discussion
Finding|Social Behavior|SIMPLE_SEGMENT|13154,13164|false|false|false|C2584313|Discussion (communication)|discussion
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|13154,13164|false|false|false|C0557061|Discussion (procedure)|discussion
Finding|Classification|SIMPLE_SEGMENT|13170,13180|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|13170,13180|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13181,13184|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|13181,13184|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|13181,13184|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|13181,13184|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|SIMPLE_SEGMENT|13181,13184|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|13181,13184|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|SIMPLE_SEGMENT|13181,13184|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13181,13184|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|SIMPLE_SEGMENT|13181,13184|false|false|false|||PCP
Finding|Gene or Genome|SIMPLE_SEGMENT|13181,13184|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|SIMPLE_SEGMENT|13181,13184|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Event|SIMPLE_SEGMENT|13189,13192|false|false|false|||hem
Finding|Pathologic Function|SIMPLE_SEGMENT|13189,13192|false|false|false|C0019080|Hemorrhage|hem
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|13189,13192|false|false|false|C0280599|altretamine/etoposide/methotrexate protocol|hem
Finding|Finding|SIMPLE_SEGMENT|13222,13225|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|13222,13225|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|13226,13232|false|false|false|C0006141|Breast|breast
Disorder|Neoplastic Process|SIMPLE_SEGMENT|13226,13232|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|breast
Finding|Finding|SIMPLE_SEGMENT|13226,13232|false|false|false|C0567499|Breast problem|breast
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|13226,13232|false|false|false|C0191838|Procedures on breast|breast
Finding|Finding|SIMPLE_SEGMENT|13226,13239|false|false|false|C0567489|Lesion of breast|breast lesion
Event|Event|SIMPLE_SEGMENT|13233,13239|false|false|false|||lesion
Finding|Finding|SIMPLE_SEGMENT|13233,13239|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|SIMPLE_SEGMENT|13233,13239|false|false|false|C0221198;C1546698|Lesion|lesion
Anatomy|Body Location or Region|SIMPLE_SEGMENT|13244,13248|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|13244,13248|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13244,13248|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|SIMPLE_SEGMENT|13244,13248|false|false|false|C0740941|Lung Problem|lung
Anatomy|Tissue|SIMPLE_SEGMENT|13249,13259|false|false|false|C0031153;C0230198;C4482223|Abdomen>Peritoneum;Peritoneum;Serous layer of peritoneum|peritoneum
Disorder|Neoplastic Process|SIMPLE_SEGMENT|13249,13259|false|false|false|C0496874;C0496954|Benign neoplasm of peritoneum;Neoplasm of uncertain or unknown behavior of peritoneum|peritoneum
Event|Event|SIMPLE_SEGMENT|13261,13268|false|false|false|||lesions
Finding|Finding|SIMPLE_SEGMENT|13261,13268|false|false|false|C0221198|Lesion|lesions
Event|Event|SIMPLE_SEGMENT|13275,13285|false|false|false|||Reevaluate
Event|Event|SIMPLE_SEGMENT|13286,13290|false|false|false|||need
Finding|Functional Concept|SIMPLE_SEGMENT|13286,13290|false|false|false|C0686904|Patient need for (contextual qualifier)|need
Finding|Functional Concept|SIMPLE_SEGMENT|13286,13294|false|false|false|C0686904|Patient need for (contextual qualifier)|need for
Drug|Organic Chemical|SIMPLE_SEGMENT|13295,13307|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13295,13307|false|false|false|C0286651|atorvastatin|atorvastatin
Event|Event|SIMPLE_SEGMENT|13295,13307|false|false|false|||atorvastatin
Event|Event|SIMPLE_SEGMENT|13317,13321|false|false|false|||need
Event|Event|SIMPLE_SEGMENT|13322,13332|false|false|false|||outpatient
Finding|Classification|SIMPLE_SEGMENT|13322,13332|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|13322,13332|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|SIMPLE_SEGMENT|13333,13339|false|false|false|||follow
Finding|Idea or Concept|SIMPLE_SEGMENT|13385,13394|false|false|false|C1546960|Patient Outcome - Worsening|worsening
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13395,13409|false|false|false|C0020295|Hydronephrosis|hydronephrosis
Event|Event|SIMPLE_SEGMENT|13395,13409|false|false|false|||hydronephrosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13413,13424|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13413,13424|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|13413,13424|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|13413,13424|false|false|false|C4284232|Medications|Medications
Finding|Finding|SIMPLE_SEGMENT|13413,13437|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|SIMPLE_SEGMENT|13428,13437|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|13428,13437|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13456,13466|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|13456,13466|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|13456,13471|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|SIMPLE_SEGMENT|13467,13471|false|false|false|||list
Finding|Intellectual Product|SIMPLE_SEGMENT|13467,13471|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|SIMPLE_SEGMENT|13475,13483|false|false|false|||accurate
Drug|Organic Chemical|SIMPLE_SEGMENT|13488,13496|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13488,13496|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|SIMPLE_SEGMENT|13488,13496|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|SIMPLE_SEGMENT|13488,13496|false|false|false|||complete
Finding|Functional Concept|SIMPLE_SEGMENT|13488,13496|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|SIMPLE_SEGMENT|13488,13496|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Organic Chemical|SIMPLE_SEGMENT|13501,13514|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13501,13514|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|SIMPLE_SEGMENT|13501,13514|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|13501,13514|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Drug|Organic Chemical|SIMPLE_SEGMENT|13533,13545|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13533,13545|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|SIMPLE_SEGMENT|13563,13573|false|false|false|C0206460|enoxaparin|Enoxaparin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13563,13573|false|false|false|C0206460|enoxaparin|Enoxaparin
Drug|Organic Chemical|SIMPLE_SEGMENT|13563,13580|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13563,13580|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|13574,13580|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|13574,13580|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13574,13580|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|SIMPLE_SEGMENT|13574,13580|false|false|false|||Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|13574,13580|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|13574,13580|false|false|false|C0337443|Sodium measurement|Sodium
Event|Event|SIMPLE_SEGMENT|13596,13601|false|false|false|||Start
Finding|Idea or Concept|SIMPLE_SEGMENT|13620,13624|false|false|false|C1552851|next - HtmlLinkType|Next
Event|Event|SIMPLE_SEGMENT|13625,13632|false|false|false|||Routine
Finding|Idea or Concept|SIMPLE_SEGMENT|13625,13632|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|Routine
Finding|Intellectual Product|SIMPLE_SEGMENT|13625,13632|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|Routine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|13625,13632|false|false|false|C1979801|Routine coag|Routine
Event|Occupational Activity|SIMPLE_SEGMENT|13633,13647|false|false|false|C0001554|Administration occupational activities|Administration
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|13633,13647|false|false|false|C1533734|Administration (procedure)|Administration
Finding|Finding|SIMPLE_SEGMENT|13648,13652|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Finding|Idea or Concept|SIMPLE_SEGMENT|13648,13652|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Finding|Intellectual Product|SIMPLE_SEGMENT|13648,13652|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|13657,13670|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Hormone|SIMPLE_SEGMENT|13657,13670|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Organic Chemical|SIMPLE_SEGMENT|13657,13670|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13657,13670|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Event|Event|SIMPLE_SEGMENT|13657,13670|false|false|false|||Levothyroxine
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|13657,13677|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Hormone|SIMPLE_SEGMENT|13657,13677|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13657,13677|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|13671,13677|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|13671,13677|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13671,13677|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|SIMPLE_SEGMENT|13671,13677|false|false|false|||Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|13671,13677|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|13671,13677|false|false|false|C0337443|Sodium measurement|Sodium
Drug|Organic Chemical|SIMPLE_SEGMENT|13699,13708|false|false|false|C0024002|lorazepam|LORazepam
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13699,13708|false|false|false|C0024002|lorazepam|LORazepam
Finding|Gene or Genome|SIMPLE_SEGMENT|13730,13733|false|false|false|C1422467|CIAO3 gene|PRN
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|13734,13741|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Event|Event|SIMPLE_SEGMENT|13734,13741|false|false|false|||anxiety
Finding|Sign or Symptom|SIMPLE_SEGMENT|13734,13741|false|false|false|C0860603|Anxiety symptoms|anxiety
Event|Event|SIMPLE_SEGMENT|13746,13755|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|13746,13755|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|13746,13755|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|13746,13755|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|13746,13755|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|13746,13767|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13756,13767|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13756,13767|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|13756,13767|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|13756,13767|false|false|false|C4284232|Medications|Medications
Drug|Antibiotic|SIMPLE_SEGMENT|13773,13782|false|false|false|C1120106|ertapenem|Ertapenem
Drug|Organic Chemical|SIMPLE_SEGMENT|13773,13782|false|false|false|C1120106|ertapenem|Ertapenem
Event|Event|SIMPLE_SEGMENT|13773,13782|false|false|false|||Ertapenem
Drug|Organic Chemical|SIMPLE_SEGMENT|13773,13789|false|false|false|C1170745|ertapenem sodium|Ertapenem Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13773,13789|false|false|false|C1170745|ertapenem sodium|Ertapenem Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|13783,13789|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|13783,13789|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13783,13789|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|SIMPLE_SEGMENT|13783,13789|false|false|false|||Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|13783,13789|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|13783,13789|false|false|false|C0337443|Sodium measurement|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13800,13808|false|false|false|C0720099|Duration brand of oxymetazoline|Duration
Event|Event|SIMPLE_SEGMENT|13800,13808|false|false|false|||Duration
Event|Event|SIMPLE_SEGMENT|13812,13816|false|false|false|||Dose
Drug|Antibiotic|SIMPLE_SEGMENT|13830,13839|true|false|false|C1120106|ertapenem|ertapenem
Drug|Organic Chemical|SIMPLE_SEGMENT|13830,13839|true|false|false|C1120106|ertapenem|ertapenem
Event|Event|SIMPLE_SEGMENT|13830,13839|true|false|false|||ertapenem
Event|Event|SIMPLE_SEGMENT|13879,13888|true|false|false|||interfere
Finding|Functional Concept|SIMPLE_SEGMENT|13879,13888|true|false|false|C0521102|Interferes with|interfere
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|13898,13914|true|false|false|C0871707|daily activities|daily activities
Event|Activity|SIMPLE_SEGMENT|13904,13914|true|false|false|C0441655|Activities|activities
Event|Event|SIMPLE_SEGMENT|13904,13914|true|false|false|||activities
Finding|Finding|SIMPLE_SEGMENT|13904,13914|true|false|false|C2239122|activities (history)|activities
Drug|Food|SIMPLE_SEGMENT|13921,13925|false|false|false|C0349374;C0444318;C1446647;C2702362;C2825079;C5551141;C5552693|Cow's milk;Milk Beverage;Milk Specimen;Milk antigen;Plant-Based Milk;cow milk allergenic extract|Milk
Drug|Immunologic Factor|SIMPLE_SEGMENT|13921,13925|false|false|false|C0349374;C0444318;C1446647;C2702362;C2825079;C5551141;C5552693|Cow's milk;Milk Beverage;Milk Specimen;Milk antigen;Plant-Based Milk;cow milk allergenic extract|Milk
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13921,13925|false|false|false|C0349374;C0444318;C1446647;C2702362;C2825079;C5551141;C5552693|Cow's milk;Milk Beverage;Milk Specimen;Milk antigen;Plant-Based Milk;cow milk allergenic extract|Milk
Drug|Substance|SIMPLE_SEGMENT|13921,13925|false|false|false|C0349374;C0444318;C1446647;C2702362;C2825079;C5551141;C5552693|Cow's milk;Milk Beverage;Milk Specimen;Milk antigen;Plant-Based Milk;cow milk allergenic extract|Milk
Event|Event|SIMPLE_SEGMENT|13921,13925|false|false|false|||Milk
Finding|Body Substance|SIMPLE_SEGMENT|13921,13925|false|false|false|C0026131;C1546713|Milk (body substance);Milk Specimen Code|Milk
Finding|Intellectual Product|SIMPLE_SEGMENT|13921,13925|false|false|false|C0026131;C1546713|Milk (body substance);Milk Specimen Code|Milk
Drug|Clinical Drug|SIMPLE_SEGMENT|13921,13937|false|false|false|C0591789;C0782828|Milk of Magnesia (Brand Name);magnesium hydroxide Oral Suspension|Milk of Magnesia
Drug|Inorganic Chemical|SIMPLE_SEGMENT|13921,13937|false|false|false|C0591789;C0782828|Milk of Magnesia (Brand Name);magnesium hydroxide Oral Suspension|Milk of Magnesia
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13921,13937|false|false|false|C0591789;C0782828|Milk of Magnesia (Brand Name);magnesium hydroxide Oral Suspension|Milk of Magnesia
Drug|Inorganic Chemical|SIMPLE_SEGMENT|13929,13937|false|false|false|C0024477|magnesium oxide|Magnesia
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13929,13937|false|false|false|C0024477|magnesium oxide|Magnesia
Event|Event|SIMPLE_SEGMENT|13929,13937|false|false|false|||Magnesia
Finding|Gene or Genome|SIMPLE_SEGMENT|13951,13954|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|SIMPLE_SEGMENT|13955,13967|false|false|false|||constipation
Finding|Sign or Symptom|SIMPLE_SEGMENT|13955,13967|false|false|false|C0009806|Constipation|constipation
Drug|Organic Chemical|SIMPLE_SEGMENT|13974,13984|false|false|false|C0206460|enoxaparin|Enoxaparin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13974,13984|false|false|false|C0206460|enoxaparin|Enoxaparin
Event|Event|SIMPLE_SEGMENT|13974,13984|false|false|false|||Enoxaparin
Drug|Organic Chemical|SIMPLE_SEGMENT|13974,13991|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13974,13991|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|13985,13991|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|13985,13991|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13985,13991|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|SIMPLE_SEGMENT|13985,13991|false|false|false|||Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|13985,13991|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|13985,13991|false|false|false|C0337443|Sodium measurement|Sodium
Event|Event|SIMPLE_SEGMENT|14007,14012|false|false|false|||Start
Finding|Idea or Concept|SIMPLE_SEGMENT|14039,14043|false|false|false|C1552851|next - HtmlLinkType|Next
Finding|Idea or Concept|SIMPLE_SEGMENT|14044,14051|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|Routine
Finding|Intellectual Product|SIMPLE_SEGMENT|14044,14051|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|Routine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|14044,14051|false|false|false|C1979801|Routine coag|Routine
Event|Event|SIMPLE_SEGMENT|14052,14066|false|false|false|||Administration
Event|Occupational Activity|SIMPLE_SEGMENT|14052,14066|false|false|false|C0001554|Administration occupational activities|Administration
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|14052,14066|false|false|false|C1533734|Administration (procedure)|Administration
Finding|Finding|SIMPLE_SEGMENT|14068,14072|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Finding|Idea or Concept|SIMPLE_SEGMENT|14068,14072|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Finding|Intellectual Product|SIMPLE_SEGMENT|14068,14072|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Drug|Organic Chemical|SIMPLE_SEGMENT|14079,14092|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14079,14092|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|SIMPLE_SEGMENT|14079,14092|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|14079,14092|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Drug|Organic Chemical|SIMPLE_SEGMENT|14113,14125|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14113,14125|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|14145,14158|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Hormone|SIMPLE_SEGMENT|14145,14158|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Organic Chemical|SIMPLE_SEGMENT|14145,14158|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14145,14158|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|14145,14165|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Hormone|SIMPLE_SEGMENT|14145,14165|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14145,14165|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|14159,14165|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|14159,14165|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14159,14165|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|SIMPLE_SEGMENT|14159,14165|false|false|false|||Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|14159,14165|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|14159,14165|false|false|false|C0337443|Sodium measurement|Sodium
Drug|Organic Chemical|SIMPLE_SEGMENT|14189,14198|false|false|false|C0024002|lorazepam|LORazepam
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14189,14198|false|false|false|C0024002|lorazepam|LORazepam
Finding|Gene or Genome|SIMPLE_SEGMENT|14220,14223|false|false|false|C1422467|CIAO3 gene|PRN
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|14224,14231|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Event|Event|SIMPLE_SEGMENT|14224,14231|false|false|false|||anxiety
Finding|Sign or Symptom|SIMPLE_SEGMENT|14224,14231|false|false|false|C0860603|Anxiety symptoms|anxiety
Event|Event|SIMPLE_SEGMENT|14237,14246|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|14237,14246|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|14237,14246|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|14237,14246|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|14237,14246|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14237,14258|false|false|false|C4019243||Discharge Disposition
Finding|Finding|SIMPLE_SEGMENT|14237,14258|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14247,14258|false|false|false|C2926604||Disposition
Event|Event|SIMPLE_SEGMENT|14247,14258|false|false|false|||Disposition
Procedure|Health Care Activity|SIMPLE_SEGMENT|14247,14258|false|false|false|C0184758|Patient disposition|Disposition
Finding|Finding|SIMPLE_SEGMENT|14260,14268|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|SIMPLE_SEGMENT|14260,14268|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Procedure|Health Care Activity|SIMPLE_SEGMENT|14260,14273|false|false|false|C0023977|long-term care|Extended Care
Event|Activity|SIMPLE_SEGMENT|14269,14273|false|false|false|C1947933|care activity|Care
Event|Event|SIMPLE_SEGMENT|14269,14273|false|false|false|||Care
Finding|Finding|SIMPLE_SEGMENT|14269,14273|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|SIMPLE_SEGMENT|14269,14273|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Event|Event|SIMPLE_SEGMENT|14276,14284|false|false|false|||Facility
Finding|Intellectual Product|SIMPLE_SEGMENT|14276,14284|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|SIMPLE_SEGMENT|14292,14301|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|14292,14301|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|14292,14301|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|14292,14301|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|14292,14301|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|14292,14311|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14302,14311|false|false|false|C0945731||Diagnosis
Event|Event|SIMPLE_SEGMENT|14302,14311|false|false|false|||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|14302,14311|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|14302,14311|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|14302,14311|false|false|false|C0011900|Diagnosis|Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14313,14330|false|false|false|C0801658||Primary diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14321,14330|false|false|false|C0945731||diagnosis
Event|Event|SIMPLE_SEGMENT|14321,14330|false|false|false|||diagnosis
Finding|Classification|SIMPLE_SEGMENT|14321,14330|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|14321,14330|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|14321,14330|false|false|false|C0011900|Diagnosis|diagnosis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|14332,14338|false|false|false|C0030797|Pelvis|Pelvic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14332,14355|false|false|false|C1697454|Pelvic fluid collection|Pelvic fluid collection
Drug|Substance|SIMPLE_SEGMENT|14339,14344|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|14339,14344|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|14345,14355|false|false|false|||collection
Finding|Conceptual Entity|SIMPLE_SEGMENT|14345,14355|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|SIMPLE_SEGMENT|14345,14355|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|SIMPLE_SEGMENT|14345,14355|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|SIMPLE_SEGMENT|14345,14355|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14356,14365|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|SIMPLE_SEGMENT|14356,14365|false|false|false|||infection
Finding|Pathologic Function|SIMPLE_SEGMENT|14356,14365|false|false|false|C3714514|Infection|infection
Event|Event|SIMPLE_SEGMENT|14372,14377|false|false|false|||acute
Finding|Intellectual Product|SIMPLE_SEGMENT|14372,14377|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14379,14384|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|14379,14384|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|14379,14384|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Finding|SIMPLE_SEGMENT|14379,14389|false|false|false|C0019080;C3163616|Blood Loss;Hemorrhage|blood loss
Finding|Pathologic Function|SIMPLE_SEGMENT|14379,14389|false|false|false|C0019080;C3163616|Blood Loss;Hemorrhage|blood loss
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14379,14396|false|false|false|C0154286;C0154298;C0948824|Acute posthaemorrhagic anaemia;Anemia due to blood loss;Iron deficiency anemia secondary to chronic blood loss|blood loss anemia
Finding|Finding|SIMPLE_SEGMENT|14385,14389|false|false|false|C5890125|Loss (adaptation)|loss
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14390,14396|false|false|false|C0002871|Anemia|anemia
Event|Event|SIMPLE_SEGMENT|14390,14396|false|false|false|||anemia
Disorder|Neoplastic Process|SIMPLE_SEGMENT|14398,14407|false|false|false|C0027627|Neoplasm Metastasis|Secondary
Event|Event|SIMPLE_SEGMENT|14398,14407|false|false|false|||Secondary
Finding|Functional Concept|SIMPLE_SEGMENT|14398,14407|false|false|false|C1522484|metastatic qualifier|Secondary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14398,14417|false|false|false|C4255018||Secondary diagnosis
Finding|Finding|SIMPLE_SEGMENT|14398,14417|false|false|false|C0332138|Secondary diagnosis|Secondary diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14408,14417|false|false|false|C0945731||diagnosis
Event|Event|SIMPLE_SEGMENT|14408,14417|false|false|false|||diagnosis
Finding|Classification|SIMPLE_SEGMENT|14408,14417|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|14408,14417|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|14408,14417|false|false|false|C0011900|Diagnosis|diagnosis
Finding|Intellectual Product|SIMPLE_SEGMENT|14419,14424|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14419,14438|false|false|false|C0022660|Kidney Failure, Acute|acute renal failure
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|14425,14430|false|false|false|C0022646|Kidney|renal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14425,14430|false|false|false|C0042075|Urologic Diseases|renal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14425,14438|false|false|false|C0035078|Kidney Failure|renal failure
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14425,14445|false|false|false|C0022660|Kidney Failure, Acute|renal failure, acute
Event|Event|SIMPLE_SEGMENT|14431,14438|false|false|false|||failure
Finding|Functional Concept|SIMPLE_SEGMENT|14431,14438|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|SIMPLE_SEGMENT|14431,14438|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|SIMPLE_SEGMENT|14431,14438|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Event|Event|SIMPLE_SEGMENT|14440,14445|false|false|false|||acute
Finding|Intellectual Product|SIMPLE_SEGMENT|14440,14445|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|SIMPLE_SEGMENT|14449,14456|false|false|false|||chronic
Finding|Intellectual Product|SIMPLE_SEGMENT|14449,14456|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|14449,14456|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14458,14464|false|false|false|C0002871|Anemia|anemia
Event|Event|SIMPLE_SEGMENT|14458,14464|false|false|false|||anemia
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|14473,14482|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14473,14482|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|14473,14482|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|SIMPLE_SEGMENT|14473,14491|false|false|false|C0034065|Pulmonary Embolism|pulmonary embolism
Event|Event|SIMPLE_SEGMENT|14483,14491|false|false|false|||embolism
Finding|Finding|SIMPLE_SEGMENT|14483,14491|false|false|false|C0013922;C1704212|Embolism;Embolus|embolism
Finding|Pathologic Function|SIMPLE_SEGMENT|14483,14491|false|false|false|C0013922;C1704212|Embolism;Embolus|embolism
Finding|Finding|SIMPLE_SEGMENT|14502,14506|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|SIMPLE_SEGMENT|14502,14506|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|SIMPLE_SEGMENT|14502,14506|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Classification|SIMPLE_SEGMENT|14507,14512|false|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|grade
Finding|Finding|SIMPLE_SEGMENT|14507,14512|false|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|grade
Disorder|Neoplastic Process|SIMPLE_SEGMENT|14514,14534|false|false|false|C0007138;C2145472|Carcinoma, Transitional Cell;Urothelial Carcinoma|urothelial carcinoma
Disorder|Neoplastic Process|SIMPLE_SEGMENT|14525,14534|false|false|false|C0007097|Carcinoma|carcinoma
Event|Event|SIMPLE_SEGMENT|14525,14534|false|false|false|||carcinoma
Finding|Functional Concept|SIMPLE_SEGMENT|14536,14540|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|14536,14547|false|false|false|C0222601|Left breast|left breast
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|14541,14547|false|false|false|C0006141|Breast|breast
Disorder|Neoplastic Process|SIMPLE_SEGMENT|14541,14547|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|breast
Finding|Finding|SIMPLE_SEGMENT|14541,14547|false|false|false|C0567499|Breast problem|breast
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|14541,14547|false|false|false|C0191838|Procedures on breast|breast
Finding|Finding|SIMPLE_SEGMENT|14541,14552|false|false|false|C0024103|Mass in breast|breast mass
Event|Event|SIMPLE_SEGMENT|14548,14552|false|false|false|||mass
Finding|Finding|SIMPLE_SEGMENT|14548,14552|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|SIMPLE_SEGMENT|14548,14552|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|SIMPLE_SEGMENT|14548,14552|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|SIMPLE_SEGMENT|14554,14560|false|false|false|C1511314|Breast Imaging Reporting and Data System|BIRADS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14566,14580|false|false|false|C0020676|Hypothyroidism|hypothyroidism
Event|Event|SIMPLE_SEGMENT|14566,14580|false|false|false|||hypothyroidism
Event|Event|SIMPLE_SEGMENT|14586,14595|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|14586,14595|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|14586,14595|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|14586,14595|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|14586,14595|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14596,14605|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14596,14605|false|false|false|C0012634|Disease|Condition
Event|Event|SIMPLE_SEGMENT|14596,14605|false|false|false|||Condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|14596,14605|false|false|false|C1705253|Logical Condition|Condition
Finding|Mental Process|SIMPLE_SEGMENT|14607,14613|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14607,14620|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|SIMPLE_SEGMENT|14607,14620|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14614,14620|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|14614,14620|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|14622,14627|false|false|false|||Clear
Finding|Idea or Concept|SIMPLE_SEGMENT|14622,14627|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|SIMPLE_SEGMENT|14632,14640|false|false|false|||coherent
Finding|Finding|SIMPLE_SEGMENT|14632,14640|false|false|false|C4068804|Coherent|coherent
Event|Event|SIMPLE_SEGMENT|14642,14647|false|false|false|||Level
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14642,14664|false|false|false|C4050479||Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|14642,14664|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|SIMPLE_SEGMENT|14651,14664|false|false|false|||Consciousness
Finding|Finding|SIMPLE_SEGMENT|14651,14664|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|SIMPLE_SEGMENT|14651,14664|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14666,14671|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|14666,14671|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14666,14671|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|SIMPLE_SEGMENT|14666,14671|false|false|false|||Alert
Finding|Finding|SIMPLE_SEGMENT|14666,14671|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|14666,14671|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|14666,14671|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|SIMPLE_SEGMENT|14676,14687|false|false|false|||interactive
Finding|Functional Concept|SIMPLE_SEGMENT|14676,14687|false|false|false|C1704675|Interaction|interactive
Event|Activity|SIMPLE_SEGMENT|14689,14697|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|14689,14697|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|SIMPLE_SEGMENT|14689,14697|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14698,14704|false|false|false|C5889824||Status
Event|Event|SIMPLE_SEGMENT|14698,14704|false|false|false|||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|14698,14704|false|false|false|C1546481|What subject filter - Status|Status
Finding|Functional Concept|SIMPLE_SEGMENT|14706,14716|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|SIMPLE_SEGMENT|14706,14716|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|SIMPLE_SEGMENT|14706,14716|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|SIMPLE_SEGMENT|14706,14716|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|SIMPLE_SEGMENT|14719,14727|false|false|false|||requires
Event|Event|SIMPLE_SEGMENT|14728,14738|false|false|false|||assistance
Finding|Social Behavior|SIMPLE_SEGMENT|14728,14738|false|false|false|C0018896|Helping Behavior|assistance
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|14742,14745|false|false|false|C1454018|AICDA protein, human|aid
Drug|Enzyme|SIMPLE_SEGMENT|14742,14745|false|false|false|C1454018|AICDA protein, human|aid
Event|Event|SIMPLE_SEGMENT|14742,14745|false|false|false|||aid
Finding|Gene or Genome|SIMPLE_SEGMENT|14742,14745|false|false|false|C1421876;C3540469|AICDA gene;AICDA wt Allele|aid
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|14742,14745|false|false|false|C0021588;C0280108|AID - Artificial insemination by donor;dacarbazine/doxorubicin/ifosfamide protocol|aid
Event|Event|SIMPLE_SEGMENT|14747,14753|false|false|false|||walker
Event|Event|SIMPLE_SEGMENT|14768,14777|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|14768,14777|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|14768,14777|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|14768,14777|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|14768,14777|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14768,14790|false|false|false|C3669312||Discharge Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|14768,14790|false|false|false|C4282220|Discharge instructions|Discharge Instructions
Procedure|Health Care Activity|SIMPLE_SEGMENT|14768,14790|false|false|false|C2266673|hospital discharge instructions (treatment)|Discharge Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14778,14790|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|14778,14790|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|14778,14790|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Finding|Gene or Genome|SIMPLE_SEGMENT|14792,14796|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Event|Event|SIMPLE_SEGMENT|14815,14819|false|false|false|||come
Finding|Idea or Concept|SIMPLE_SEGMENT|14827,14835|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|SIMPLE_SEGMENT|14848,14855|false|false|false|||feeling
Finding|Finding|SIMPLE_SEGMENT|14848,14861|false|false|false|C0849970|Feeling tired|feeling tired
Event|Event|SIMPLE_SEGMENT|14856,14861|false|false|false|||tired
Finding|Finding|SIMPLE_SEGMENT|14856,14861|false|false|false|C0015672;C0849970;C3539029|Fatigue;Feel Tired question;Feeling tired|tired
Finding|Intellectual Product|SIMPLE_SEGMENT|14856,14861|false|false|false|C0015672;C0849970;C3539029|Fatigue;Feel Tired question;Feeling tired|tired
Finding|Sign or Symptom|SIMPLE_SEGMENT|14856,14861|false|false|false|C0015672;C0849970;C3539029|Fatigue;Feel Tired question;Feeling tired|tired
Drug|Substance|SIMPLE_SEGMENT|14871,14876|false|false|false|C1550628|Drain - SpecimenType|drain
Finding|Intellectual Product|SIMPLE_SEGMENT|14871,14876|false|false|false|C1546604|Drain Specimen Code|drain
Event|Event|SIMPLE_SEGMENT|14877,14883|false|false|false|||output
Finding|Conceptual Entity|SIMPLE_SEGMENT|14877,14883|false|false|false|C1709366|system output|output
Procedure|Health Care Activity|SIMPLE_SEGMENT|14877,14883|false|false|false|C3251815|Measurement of fluid output|output
Event|Event|SIMPLE_SEGMENT|14888,14894|false|false|false|||bloody
Finding|Finding|SIMPLE_SEGMENT|14888,14894|false|false|false|C4554530|Bloody|bloody
Event|Event|SIMPLE_SEGMENT|14903,14911|false|false|false|||happened
Finding|Idea or Concept|SIMPLE_SEGMENT|14919,14927|false|false|false|C1547192|Organization unit type - Hospital|hospital
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|14933,14940|false|false|false|C0040405|X-Ray Computed Tomography|CT scan
Event|Event|SIMPLE_SEGMENT|14936,14940|false|false|false|||scan
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|14936,14940|false|false|false|C0034606;C0441633|Radionuclide Imaging;Scanning|scan
Event|Event|SIMPLE_SEGMENT|14941,14947|false|false|false|||showed
Finding|Finding|SIMPLE_SEGMENT|14948,14958|false|false|false|C0450093|Very large|very large
Finding|Gene or Genome|SIMPLE_SEGMENT|14953,14958|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Drug|Substance|SIMPLE_SEGMENT|14959,14964|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|14959,14964|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|14965,14976|false|false|false|||collections
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|14985,14991|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|14985,14991|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Disorder|Neoplastic Process|SIMPLE_SEGMENT|14985,14991|false|false|false|C0153663|Malignant neoplasm of pelvis|pelvis
Finding|Finding|SIMPLE_SEGMENT|14985,14991|false|false|false|C0812455|Pelvis problem|pelvis
Event|Event|SIMPLE_SEGMENT|14999,15011|false|false|false|||radiologists
Event|Event|SIMPLE_SEGMENT|15012,15018|false|false|false|||placed
Drug|Substance|SIMPLE_SEGMENT|15027,15032|false|false|false|C1550628|Drain - SpecimenType|drain
Event|Event|SIMPLE_SEGMENT|15027,15032|false|false|false|||drain
Finding|Intellectual Product|SIMPLE_SEGMENT|15027,15032|false|false|false|C1546604|Drain Specimen Code|drain
Event|Event|SIMPLE_SEGMENT|15037,15044|false|false|false|||removed
Finding|Intellectual Product|SIMPLE_SEGMENT|15048,15052|false|false|false|C1720092|Once - dosing instruction fragment|once
Event|Event|SIMPLE_SEGMENT|15057,15065|false|false|false|||appeared
Finding|Gene or Genome|SIMPLE_SEGMENT|15075,15080|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Drug|Substance|SIMPLE_SEGMENT|15081,15086|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|15081,15086|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|15087,15097|false|false|false|||collection
Finding|Conceptual Entity|SIMPLE_SEGMENT|15087,15097|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|SIMPLE_SEGMENT|15087,15097|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|SIMPLE_SEGMENT|15087,15097|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|SIMPLE_SEGMENT|15087,15097|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Event|Event|SIMPLE_SEGMENT|15102,15106|false|false|false|||gone
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15126,15131|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|SIMPLE_SEGMENT|15126,15131|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|15126,15143|false|false|false|C0005841|Blood Transfusion|blood transfusion
Event|Event|SIMPLE_SEGMENT|15132,15143|false|false|false|||transfusion
Finding|Functional Concept|SIMPLE_SEGMENT|15132,15143|false|false|false|C0199960||transfusion
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|15132,15143|false|false|false|C0005841;C1879316|Blood Transfusion;Transfusion (procedure)|transfusion
Event|Event|SIMPLE_SEGMENT|15149,15155|false|false|false|||placed
Event|Event|SIMPLE_SEGMENT|15158,15162|false|false|false|||PICC
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|15158,15162|false|false|false|C2049629|Peripherally Inserted Central Catheter Line Insertion|PICC
Drug|Antibiotic|SIMPLE_SEGMENT|15200,15211|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|SIMPLE_SEGMENT|15200,15211|false|false|false|||antibiotics
Event|Event|SIMPLE_SEGMENT|15226,15236|false|false|false|||discharged
Finding|Idea or Concept|SIMPLE_SEGMENT|15246,15254|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|SIMPLE_SEGMENT|15261,15266|false|false|false|||needs
Event|Event|SIMPLE_SEGMENT|15270,15276|false|false|false|||happen
Event|Event|SIMPLE_SEGMENT|15286,15291|false|false|false|||leave
Finding|Idea or Concept|SIMPLE_SEGMENT|15296,15304|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|SIMPLE_SEGMENT|15315,15323|false|false|false|||continue
Event|Event|SIMPLE_SEGMENT|15324,15330|false|false|false|||seeing
Anatomy|Body Location or Region|SIMPLE_SEGMENT|15362,15366|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|15362,15366|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15362,15366|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|SIMPLE_SEGMENT|15362,15366|false|false|false|C0740941|Lung Problem|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|15371,15377|false|false|false|C0006141|Breast|breast
Disorder|Neoplastic Process|SIMPLE_SEGMENT|15371,15377|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|breast
Finding|Finding|SIMPLE_SEGMENT|15371,15377|false|false|false|C0567499|Breast problem|breast
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|15371,15377|false|false|false|C0191838|Procedures on breast|breast
Finding|Finding|SIMPLE_SEGMENT|15371,15385|false|false|false|C0567489|Lesion of breast|breast lesions
Event|Event|SIMPLE_SEGMENT|15378,15385|false|false|false|||lesions
Finding|Finding|SIMPLE_SEGMENT|15378,15385|false|false|false|C0221198|Lesion|lesions
Event|Event|SIMPLE_SEGMENT|15390,15396|false|false|false|||follow
Event|Event|SIMPLE_SEGMENT|15403,15418|false|false|false|||recommendations
Finding|Idea or Concept|SIMPLE_SEGMENT|15403,15418|false|false|false|C0034866|Recommendation|recommendations
Event|Event|SIMPLE_SEGMENT|15423,15431|false|false|false|||Continue
Finding|Idea or Concept|SIMPLE_SEGMENT|15423,15431|false|false|false|C0549178|Continuous|Continue
Event|Event|SIMPLE_SEGMENT|15432,15438|false|false|false|||taking
Drug|Organic Chemical|SIMPLE_SEGMENT|15439,15446|false|false|false|C0728963|Lovenox|Lovenox
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|15439,15446|false|false|false|C0728963|Lovenox|Lovenox
Finding|Idea or Concept|SIMPLE_SEGMENT|15453,15456|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|15453,15456|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|15460,15465|false|false|false|||treat
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15470,15475|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|15470,15475|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|15470,15475|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Pathologic Function|SIMPLE_SEGMENT|15470,15480|false|false|false|C0087086;C0302148|Blood Clot;Thrombus|blood clot
Drug|Organic Chemical|SIMPLE_SEGMENT|15476,15480|false|false|false|C0009074|clotrimazole|clot
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|15476,15480|false|false|false|C0009074|clotrimazole|clot
Finding|Pathologic Function|SIMPLE_SEGMENT|15476,15480|false|false|false|C0302148|Blood Clot|clot
Event|Event|SIMPLE_SEGMENT|15481,15483|false|false|false|||in
Anatomy|Body Location or Region|SIMPLE_SEGMENT|15490,15494|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|15490,15494|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15490,15494|false|false|false|C0024115|Lung diseases|lung
Event|Event|SIMPLE_SEGMENT|15490,15494|false|false|false|||lung
Finding|Finding|SIMPLE_SEGMENT|15490,15494|false|false|false|C0740941|Lung Problem|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15506,15516|true|false|false|C0009450|Communicable Diseases|infectious
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15506,15524|true|false|false|C0009450|Communicable Diseases|infectious disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15517,15524|true|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|15517,15524|true|false|false|||disease
Event|Event|SIMPLE_SEGMENT|15525,15531|true|false|false|||doctor
Finding|Intellectual Product|SIMPLE_SEGMENT|15525,15531|true|false|false|C2348314|Doctor - Title|doctor
Event|Event|SIMPLE_SEGMENT|15540,15549|true|false|false|||contacted
Event|Event|SIMPLE_SEGMENT|15569,15573|false|false|false|||call
Event|Event|SIMPLE_SEGMENT|15588,15594|false|false|false|||number
Finding|Idea or Concept|SIMPLE_SEGMENT|15588,15594|false|false|false|C1554106|MDF AttributeType - Number|number
Event|Activity|SIMPLE_SEGMENT|15608,15619|false|false|false|C0003629|Appointments|appointment
Event|Event|SIMPLE_SEGMENT|15608,15619|false|false|false|||appointment
Event|Event|SIMPLE_SEGMENT|15642,15646|false|false|false|||sure
Finding|Intellectual Product|SIMPLE_SEGMENT|15642,15646|false|false|false|C4724437|SURE Test|sure
Finding|Functional Concept|SIMPLE_SEGMENT|15658,15664|false|false|false|C0205341;C1705914|Repeat;Repeat Object|repeat
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|15665,15672|false|false|false|C0040405|X-Ray Computed Tomography|CT scan
Event|Event|SIMPLE_SEGMENT|15668,15672|false|false|false|||scan
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|15668,15672|false|false|false|C0034606;C0441633|Radionuclide Imaging;Scanning|scan
Event|Activity|SIMPLE_SEGMENT|15691,15702|false|false|false|C0003629|Appointments|appointment
Event|Event|SIMPLE_SEGMENT|15691,15702|false|false|false|||appointment
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15712,15722|false|false|false|C0009450|Communicable Diseases|infectious
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15712,15730|false|false|false|C0009450|Communicable Diseases|infectious disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15723,15730|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|15731,15737|false|false|false|||doctor
Finding|Intellectual Product|SIMPLE_SEGMENT|15731,15737|false|false|false|C2348314|Doctor - Title|doctor
Drug|Antibiotic|SIMPLE_SEGMENT|15763,15774|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|SIMPLE_SEGMENT|15763,15774|false|false|false|||antibiotics
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15799,15809|false|false|false|C0009450|Communicable Diseases|infectious
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15799,15817|false|false|false|C0009450|Communicable Diseases|infectious disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15810,15817|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|15810,15817|false|false|false|||disease
Event|Event|SIMPLE_SEGMENT|15818,15824|false|false|false|||doctor
Finding|Intellectual Product|SIMPLE_SEGMENT|15818,15824|false|false|false|C2348314|Doctor - Title|doctor
Event|Event|SIMPLE_SEGMENT|15829,15838|false|false|false|||determine
Event|Event|SIMPLE_SEGMENT|15857,15861|false|false|false|||need
Event|Event|SIMPLE_SEGMENT|15887,15895|false|false|false|||pleasure
Finding|Intellectual Product|SIMPLE_SEGMENT|15887,15895|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|SIMPLE_SEGMENT|15887,15895|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|SIMPLE_SEGMENT|15903,15907|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|15903,15907|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|15903,15907|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|15903,15907|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|15903,15910|false|false|false|C1555558|care of - AddressPartType|care of
Procedure|Health Care Activity|SIMPLE_SEGMENT|15934,15942|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|15943,15955|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|15943,15955|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|15943,15955|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

