CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Pharmaceutical Preparations|Drug|false|false||MEDICINEnull|Medicine|Title|false|false||MEDICINEnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|amoxicillin|Drug|false|false||amoxicillin
null|amoxicillin|Drug|false|false||amoxicillinnull|Iron Drug Class|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|Ferrum metallicum, Homeopathic preparation|Drug|false|false||ironnull|Iron measurement|Procedure|false|false||ironnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Claims attachment|Finding|false|false||attach
null|HIPAA attachments|Finding|false|false||attachnull|Fix|Phenomenon|false|false||attachnull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|Laboratory test finding|Lab|false|false||LABSnull|Primed lymphocyte test|Procedure|false|false||PLTnull|Count Dosing Unit|LabModifier|false|false||COUNT
null|Count|LabModifier|false|false||COUNTnull|Monos|Drug|false|false||MONOS
null|Mono-S|Drug|false|false||MONOS
null|Monos|Drug|false|false||MONOSnull|SARCOIDOSIS, EARLY-ONSET|Disorder|false|false||EOS
null|Familial eosinophilia|Disorder|false|false||EOSnull|PRSS33 gene|Finding|false|false||EOS
null|IKZF4 gene|Finding|false|false||EOSnull|Eos <Loriini>|Entity|false|false||EOSnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C0014792;C1114281|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||HGB
null|Hemoglobin|Drug|false|false||HGBnull|CYGB gene|Finding|false|false||HGBnull|Hemoglobin concentration|Lab|false|false||HGBnull|Hemopoietic stem cell transplant|Procedure|false|false||HCT
null|Hematocrit Measurement|Procedure|false|false||HCTnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Arylsulfatase A, human|Drug|false|false||ASA
null|Arylsulfatase A, human|Drug|false|false||ASA
null|aspirin|Drug|false|false||ASA
null|aspirin|Drug|false|false||ASAnull|ARSA gene|Finding|false|false||ASAnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|CNS depressants ethanol|Drug|false|false||ETHANOL
null|CNS depressants ethanol|Drug|false|false||ETHANOL
null|antiseptics ethanol|Drug|false|false||ETHANOL
null|antiseptics ethanol|Drug|false|false||ETHANOL
null|ethanol|Drug|false|false||ETHANOL
null|ethanol|Drug|false|false||ETHANOLnull|Toxic effect of ethyl alcohol|Disorder|false|false||ETHANOLnull|Ethanol measurement|Procedure|false|false||ETHANOLnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Albumin|Drug|false|false||ALBUMIN
null|Albumins|Drug|false|false||ALBUMIN
null|Albumins|Drug|false|false||ALBUMIN
null|Albumin|Drug|false|false||ALBUMINnull|Albumin metabolic function|Finding|false|false||ALBUMIN
null|ALB gene|Finding|false|false||ALBUMINnull|Albumin measurement|Procedure|false|false||ALBUMINnull|CALCIUM SUPPLEMENTS|Drug|false|false||CALCIUM
null|calcium|Drug|false|false||CALCIUM
null|calcium|Drug|false|false||CALCIUM
null|calcium|Drug|false|false||CALCIUM
null|CALCIUM SUPPLEMENTS|Drug|false|false||CALCIUM
null|Calcium, Dietary|Drug|false|false||CALCIUM
null|Calcium [EPC]|Drug|false|false||CALCIUM
null|Calcium Drug Class|Drug|false|false||CALCIUMnull|Calcium metabolic function|Finding|false|false||CALCIUMnull|Calcium measurement|Procedure|false|false||CALCIUMnull|phosphate ion|Drug|false|false||PHOSPHATE
null|Phosphates|Drug|false|false||PHOSPHATE
null|phosphate ion|Drug|false|false||PHOSPHATEnull|Phosphate measurement|Procedure|false|false||PHOSPHATEnull|Magnesium supplements, alimentary tract and metabolism|Drug|false|false||MAGNESIUM
null|magnesium|Drug|false|false||MAGNESIUM
null|magnesium|Drug|false|false||MAGNESIUM
null|Magnesium Drug Class|Drug|false|false||MAGNESIUM
null|Magnesium supplements, alimentary tract and metabolism|Drug|false|false||MAGNESIUMnull|Magnesium measurement|Procedure|false|false||MAGNESIUMnull|lipase|Drug|false|false||LIPASE
null|lipase|Drug|false|false||LIPASE
null|lipase|Drug|false|false||LIPASEnull|Lipase measurement|Procedure|false|false||LIPASEnull|Alanine Transaminase|Drug|false|false||ALT
null|Alanine Transaminase|Drug|false|false||ALTnull|Liposarcoma, well differentiated|Disorder|false|false||ALT
null|Atypical Lipoma|Disorder|false|false||ALTnull|null|Finding|false|false||ALT
null|Alternative Billing Concepts|Finding|false|false||ALT
null|GPT gene|Finding|false|false||ALTnull|Antibiotic Lock Therapy|Procedure|false|false||ALTnull|Southern Altai Language|Entity|false|false||ALTnull|SGPT - Glutamate pyruvate transaminase|Drug|false|false||SGPT
null|SGPT - Glutamate pyruvate transaminase|Drug|false|false||SGPTnull|GPT gene|Finding|false|false||SGPTnull|Serum Alanine Transaminase Test|Procedure|false|false||SGPTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false|C1185650|AST
null|Aspartate Transaminase|Drug|false|false|C1185650|AST
null|Aspartate Transaminase|Drug|false|false|C1185650|AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false|C1185650|AST
null|SLC17A5 protein, human|Drug|false|false|C1185650|AST
null|SLC17A5 protein, human|Drug|false|false|C1185650|ASTnull|Atypical Spitz Nevus|Disorder|false|false|C1185650|ASTnull|SLC17A5 wt Allele|Finding|false|false|C1185650|AST
null|SLC17A5 gene|Finding|false|false|C1185650|AST
null|GOT1 gene|Finding|false|false|C1185650|ASTnull|Asterion|Anatomy|false|false|C4522245;C0004002;C0242192;C1121182;C0201899;C1415181;C1420113;C5960784;C1415181|ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||SGOT
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||SGOTnull|GOT1 gene|Finding|false|false|C1185650|SGOTnull|Aspartate aminotransferase measurement|Procedure|false|false|C1185650|SGOTnull|Alkaline Phosphatase|Drug|false|false||ALK PHOS
null|Alkaline Phosphatase|Drug|false|false||ALK PHOSnull|Alkaline phosphatase measurement|Procedure|false|false||ALK PHOSnull|ALK protein, human|Drug|false|false||ALK
null|ALK protein, human|Drug|false|false||ALKnull|ALK protein, human|Finding|false|false||ALK
null|ALK gene|Finding|false|false||ALK
null|ALK wt Allele|Finding|false|false||ALKnull|Phos <Photinae>|Entity|false|false||PHOSnull|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSEnull|Glucose measurement|Procedure|false|false||GLUCOSEnull|Glucose^1.5H post dose glucagon|Lab|false|false||GLUCOSEnull|urea|Drug|false|false||UREA
null|urea|Drug|false|false||UREA
null|urea|Drug|false|false||UREAnull|Urea measurement|Procedure|false|false||UREAnull|Sodium supplements|Drug|false|false||SODIUM
null|sodium|Drug|false|false||SODIUM
null|sodium|Drug|false|false||SODIUM
null|Sodium Drug Class|Drug|false|false||SODIUMnull|Sodium metabolic function|Finding|false|false||SODIUMnull|Sodium measurement|Procedure|false|false||SODIUMnull|Potassium Drug Class|Drug|false|false||POTASSIUM
null|Dietary Potassium|Drug|false|false||POTASSIUM
null|potassium|Drug|false|false||POTASSIUM
null|potassium|Drug|false|false||POTASSIUM
null|potassium|Drug|false|false||POTASSIUM
null|Potassium supplement|Drug|false|false||POTASSIUM
null|Potassium supplement|Drug|false|false||POTASSIUMnull|Potassium metabolic function|Finding|false|false||POTASSIUMnull|Potassium measurement|Procedure|false|false||POTASSIUMnull|chloride ion|Drug|false|false||CHLORIDE
null|Chlorides|Drug|false|false||CHLORIDEnull|Chloride metabolic function|Finding|false|false||CHLORIDEnull|Chloride measurement|Procedure|false|false||CHLORIDEnull|Total|Modifier|false|false||TOTALnull|carbon dioxide|Drug|false|false||CO2
null|carbon dioxide|Drug|false|false||CO2null|MT-CO2 gene|Finding|false|false||CO2
null|null|Finding|false|false||CO2
null|C2 wt Allele|Finding|false|false||CO2null|blood anion gap (lab test)|Procedure|false|false||ANION GAP
null|Anion gap measurement|Procedure|false|false||ANION GAPnull|Anion Gap|Attribute|false|false||ANION GAPnull|Anion gap result|Lab|false|false||ANION GAPnull|Anions|Drug|false|false||ANIONnull|Ras GTPase-Activating Protein 1, Human|Drug|false|false||GAP
null|Ras GTPase-Activating Protein 1, Human|Drug|false|false||GAP
null|GTPase-Activating Proteins|Drug|false|false||GAP
null|GTPase-Activating Proteins|Drug|false|false||GAPnull|RASA1 wt Allele|Finding|false|false||GAP
null|RASA1 gene|Finding|false|false||GAPnull|Gap (space)|Modifier|false|false||GAPnull|Mandibular left third molar abutment mesial hemisection|Device|false|false||17AMnull|Hematuria|Disorder|false|false||URINE  BLOODnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|nitrite ion|Drug|false|false||NITRITE
null|Nitrites|Drug|false|false||NITRITE
null|Nitrites|Drug|false|false||NITRITE
null|Nitrites|Drug|false|false||NITRITE
null|nitrite ion|Drug|false|false||NITRITE
null|nitrite ion|Drug|false|false||NITRITEnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Proteins|Drug|false|false||PROTEIN
null|Proteins|Drug|false|false||PROTEINnull|Protein Info|Finding|false|false||PROTEINnull|Protein measurement|Procedure|false|false||PROTEINnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSEnull|Glucose measurement|Procedure|false|false||GLUCOSEnull|Glucose^1.5H post dose glucagon|Lab|false|false||GLUCOSEnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Ketones|Drug|false|false||KETONEnull|bilirubin preparation|Drug|false|false||BILIRUBIN
null|bilirubin preparation|Drug|false|false||BILIRUBIN
null|Bilirubin|Drug|false|false||BILIRUBIN
null|Bilirubin|Drug|false|false||BILIRUBINnull|Bilirubin, total measurement|Procedure|false|false||BILIRUBIN
null|blood bilirubin level test|Procedure|false|false||BILIRUBINnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Mandibular left third molar abutment mesial hemisection|Device|false|false||17AMnull|Color of urine|Finding|false|false||URINE  COLORnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|color additive|Drug|false|false||COLOR
null|Coloring Excipient|Drug|false|false||COLORnull|color - solid dosage form|Modifier|false|false||COLOR
null|Color|Modifier|false|false||COLORnull|Color quantity|LabModifier|false|false||COLORnull|Cereal plant straw|Drug|false|false||Strawnull|Straw package type|Device|false|false||Strawnull|Straw Color|Modifier|false|false||Strawnull|Straw (unit of presentation)|LabModifier|false|false||Strawnull|Remote control command - Clear|Finding|false|false||CLEARnull|Clear|Modifier|false|false||CLEAR
null|Transparent (qualitative concept)|Modifier|false|false||CLEARnull|Mandibular left third molar abutment mesial hemisection|Device|false|false||17AMnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Opiates|Drug|false|false||opiates
null|Opiates|Drug|false|false||opiates
null|Opiates|Drug|false|false||opiates
null|Opiate Alkaloids|Drug|false|false||opiates
null|Opiate Alkaloids|Drug|false|false||opiates
null|Opiate Alkaloids|Drug|false|false||opiatesnull|Opiate Measurement|Procedure|false|false||opiatesnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|cocaine|Drug|false|false||cocaine
null|cocaine|Drug|false|false||cocaine
null|cocaine|Drug|false|false||cocaine
null|cocaine|Drug|false|false||cocainenull|Poisoning by cocaine|Disorder|false|false||cocainenull|Cocaine measurement|Procedure|false|false||cocainenull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Mandibular left third molar abutment mesial hemisection|Device|false|false||17AMnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Rh Negative Blood Group|Finding|false|false||NEGATIVE
null|Negative|Finding|false|false||NEGATIVE
null|Negative Finding|Finding|false|false||NEGATIVEnull|Expression Negative|Lab|false|false||NEGATIVEnull|Negative - qualifier|Modifier|false|false||NEGATIVE
null|Negative Charge|Modifier|false|false||NEGATIVEnull|Negative Number|LabModifier|false|false||NEGATIVEnull|Mandibular left third molar abutment mesial hemisection|Device|false|false||17AMnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Hour|Time|false|false||HOURSnull|Random|Modifier|false|false||RANDOMnull|Laboratory test finding|Lab|false|false||LABSnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|thyrotropin|Drug|false|false||TSH
null|thyrotropin|Drug|false|false||TSH
null|thyrotropin|Drug|false|false||TSHnull|Thyroid stimulating hormone measurement|Procedure|false|false||TSHnull|null|Attribute|false|false||TSHnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|T4 free measurement|Procedure|false|false||Free T4null|Free of (attribute)|Finding|false|false||Freenull|Empty (qualifier)|Modifier|false|false||Freenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|thiamine|Drug|false|false||VITAMIN B1
null|thiamine|Drug|false|false||VITAMIN B1
null|thiamine|Drug|false|false||VITAMIN B1null|Thiamine measurement|Procedure|false|false||VITAMIN B1null|Vitamins|Drug|false|false||VITAMIN
null|Vitamins|Drug|false|false||VITAMIN
null|Vitamins|Drug|false|false||VITAMINnull|whole blood specimen|Finding|false|false||WHOLE BLOOD
null|whole blood|Finding|false|false||WHOLE BLOOD
null|null|Finding|false|false||WHOLE BLOODnull|null|LabModifier|false|false||WHOLEnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Paroxysmal nocturnal dyspnea|Disorder|false|false||PNDnull|NPPA wt Allele|Finding|false|false||PND
null|NPPA gene|Finding|false|false||PNDnull|Micro (prefix)|Finding|false|false||MICRO
null|Microbiology - Laboratory Class|Finding|false|false||MICROnull|Microbiology procedure|Procedure|false|false||MICROnull|Unit Of Measure Prefix - micro|LabModifier|false|false||MICROnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Final report|Finding|false|false||FINAL REPORTnull|Diagnosis Type - Final|Finding|false|false||FINALnull|Final|Time|false|false||FINALnull|End-stage|Modifier|false|false||FINALnull|Report (document)|Finding|false|false||REPORTnull|Reporting|Procedure|false|false||REPORTnull|null|Attribute|false|false||REPORTnull|Urine culture|Procedure|false|false||URINE CULTUREnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Culture Dose Form|Drug|false|false||CULTUREnull|Culture (Anthropological)|Finding|false|false||CULTURE
null|Cultural aspects|Finding|false|false||CULTUREnull|Microbial culture (procedure)|Procedure|false|false||CULTURE
null|Laboratory culture|Procedure|false|false||CULTUREnull|Diagnosis Type - Final|Finding|false|false||Finalnull|Final|Time|false|false||Finalnull|End-stage|Modifier|false|false||Finalnull|Bacterial|Modifier|false|false||BACTERIALnull|Colony (cells or organisms)|Anatomy|false|false||COLONYnull|colonies (qualifier value)|LabModifier|false|false||COLONYnull|null|Modifier|false|false||TYPESnull|Consistent with|Finding|false|false||CONSISTENTnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false|C1123023;C4520765|SKIN
null|Skin and subcutaneous tissue disorders|Disorder|false|false|C1123023;C4520765|SKINnull|Skin Specimen Source Code|Finding|false|false|C1123023;C4520765|SKIN
null|Skin Specimen|Finding|false|false|C1123023;C4520765|SKINnull|Skin, Human|Anatomy|false|false|C1546781;C0444099;C0178298;C0496955|SKIN
null|Skin|Anatomy|false|false|C1546781;C0444099;C0178298;C0496955|SKINnull|Specimen Type - Genital|Finding|false|false|C0017420;C0559522|GENITAL
null|null|Finding|false|false|C0017420;C0559522|GENITALnull|Genital system|Anatomy|false|false|C1550642;C1546649;C0259846;C2349974|GENITAL
null|Genitalia|Anatomy|false|false|C1550642;C1546649;C0259846;C2349974|GENITALnull|Contamination|Finding|false|false|C0017420;C0559522|CONTAMINATIONnull|adulteration|Phenomenon|false|false|C0017420;C0559522|CONTAMINATIONnull|Specimen Reject Reason - Contamination|Modifier|false|false||CONTAMINATIONnull|Imaging problem|Finding|false|false||IMAGINGnull|Diagnostic Imaging|Procedure|false|false||IMAGING
null|Imaging Techniques|Procedure|false|false||IMAGINGnull|Imaging Technology|Title|false|false||IMAGINGnull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|Laboratory test finding|Lab|false|false||LABSnull|Laboratory test finding|Lab|true|false||labsnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|physical examination (physical finding)|Finding|false|false||PHYSICAL EXAMnull|Physical Examination|Procedure|false|false||PHYSICAL EXAMnull|physical examination (physical finding)|Finding|false|false||PHYSICAL
null|Physical|Finding|false|false||PHYSICALnull|Physical Examination|Procedure|false|false||PHYSICALnull|Exam|Finding|false|false||EXAMnull|Medical Examination|Procedure|false|false||EXAMnull|C1orf210 gene|Finding|false|false||Tempnull|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Procedure|false|false||Tempnull|Temperature|LabModifier|false|false||Tempnull|delivery (history)|Finding|false|false||delivery
null|Transfer Technique|Finding|false|false||delivery
null|null|Finding|false|false||deliverynull|Obstetric Delivery|Procedure|false|false||deliverynull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||GENERALnull|General medical service|Procedure|false|false||GENERALnull|Generalized|Modifier|false|false||GENERALnull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|Chairs|Device|false|false||chairnull|Chairperson|Subject|false|false||chairnull|Smiling|Finding|false|false||smilingnull|Problems with head|Disorder|false|false|C0018670;C0152336|headnull|Procedure on head|Procedure|false|false|C0018670;C0152336|headnull|Structure of head of caudate nucleus|Anatomy|false|false|C0362076;C0876917|head
null|Head|Anatomy|false|false|C0362076;C0876917|headnull|Head Device|Device|false|false||headnull|Eye|Anatomy|false|false|C5848506|EYESnull|null|Attribute|false|false|C0015392|EYESnull|Scleral Diseases|Disorder|false|false|C0036410|Scleranull|examination of sclera|Procedure|false|false|C0036410|Scleranull|Sclera|Anatomy|false|false|C0205180;C0036412;C2228481;C1828121|Scleranull|Anicteric|Finding|false|false|C0036410|anictericnull|Injection|Drug|true|false||injectionnull|Injection Route of Administration|Finding|true|false|C0036410|injectionnull|Injection of therapeutic agent|Procedure|true|false||injection
null|Injection procedure|Procedure|true|false||injectionnull|Cardiac attachment|Finding|false|false|C0018787|CARDIACnull|Heart|Anatomy|false|false|C1314974|CARDIACnull|Cardiac - anatomy qualifier|Modifier|false|false||CARDIACnull|Heart murmur|Finding|true|false||murmursnull|Pericardial friction rub|Finding|true|false||rubsnull|Respiratory, thoracic and mediastinal disorders|Disorder|false|false||RESPnull|Respiratory rate|Attribute|false|false||RESPnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Auscultation|Procedure|false|false||auscultationnull|Wheezing|Finding|true|false||wheezesnull|Rhonchi|Finding|true|false||rhonchinull|Basilar Rales|Finding|false|false||rales
null|Rales|Finding|false|false||ralesnull|Increased work of breathing|Finding|true|false||increased work of breathingnull|Increased (finding)|Finding|true|false||increased
null|Increase|Finding|true|false||increasednull|Increased|LabModifier|false|false||increasednull|Work of Breathing|Finding|true|false||work of breathingnull|Work|Event|true|false||worknull|outcomes otolaryngology breathing|Finding|false|false||breathing
null|Inspiration (function)|Finding|false|false||breathing
null|Respiration|Finding|false|false||breathingnull|null|Attribute|false|false||breathingnull|respiratory system process|Phenomenon|false|false||breathingnull|Malignant neoplasm of abdomen|Disorder|false|false|C0230168;C0000726|ABDOMENnull|Abdomen problem|Finding|false|false|C0230168;C0000726|ABDOMENnull|Abdomen|Anatomy|false|false|C0153662;C0941288|ABDOMEN
null|Abdominal Cavity|Anatomy|false|false|C0153662;C0941288|ABDOMENnull|Intestines|Anatomy|false|false||bowelsnull|null|Device|false|false||soundsnull|null|Phenomenon|false|false||soundsnull|Dilated|Finding|false|false||distendednull|Distended|Modifier|false|false||distendednull|All extremities|Anatomy|false|false||EXTREMITIES
null|Limb structure|Anatomy|false|false||EXTREMITIESnull|null|Drug|false|false||Pulsesnull|Physiologic pulse|Finding|false|false||Pulsesnull|Pulse taking|Procedure|false|false||Pulsesnull|Radial|Finding|false|false||Radial
null|Circumpennate|Finding|false|false||Radialnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false|C1123023;C4520765|SKIN
null|Skin and subcutaneous tissue disorders|Disorder|false|false|C1123023;C4520765|SKINnull|Skin Specimen Source Code|Finding|false|false|C1123023;C4520765|SKIN
null|Skin Specimen|Finding|false|false|C1123023;C4520765|SKINnull|Skin, Human|Anatomy|false|false|C1546781;C0444099;C0178298;C0496955|SKIN
null|Skin|Anatomy|false|false|C1546781;C0444099;C0178298;C0496955|SKINnull|Feels warm|Finding|false|false||Warmnull|warming process|Phenomenon|false|false||Warmnull|capsule (pharmacologic)|Drug|false|false||Capnull|CATARACT, ANTERIOR POLAR|Disorder|false|false||Capnull|BRD4 wt Allele|Finding|false|false||Cap
null|HACD1 gene|Finding|false|false||Cap
null|SERPINB6 gene|Finding|false|false||Cap
null|BRD4 gene|Finding|false|false||Cap
null|CAP1 gene|Finding|false|false||Cap
null|SORBS1 gene|Finding|false|false||Cap
null|LNPEP gene|Finding|false|false||Capnull|CAP Regimen|Procedure|false|false||Cap
null|cisplatin/cyclophosphamide/doxorubicin protocol|Procedure|false|false||Cap
null|cyclophosphamide/doxorubicin/prednisone protocol|Procedure|false|false||Capnull|Cap (physical object)|Device|false|false||Cap
null|Syringe Caps|Device|false|false||Cap
null|Cap device|Device|false|false||Capnull|College of American Pathologists|Subject|false|false||Capnull|Controlled Attenuation Parameter|Modifier|false|false||Capnull|Capsule Dosing Unit|LabModifier|false|false||Capnull|refill|Finding|false|false||refillnull|Eruption of skin (disorder)|Disorder|true|false||rashnull|Skin rash|Finding|true|false||rash
null|Eruptions|Finding|true|false||rash
null|Exanthema|Finding|true|false||rashnull|Neurologic (qualifier value)|Modifier|false|false||NEUROLOGICnull|Speech|Finding|false|false||Speechnull|Speech assessment|Procedure|false|false||Speechnull|Slow|Modifier|false|false||slownull|Massive|Modifier|false|false||markedlynull|Admission Level of Care Code - Improved|Finding|false|false||improved
null|Improved - answer to question|Finding|false|false||improved
null|Improved|Finding|false|false||improvednull|Better|Modifier|false|false||improvednull|Does speak|Finding|false|false||speaksnull|LITAF gene|Finding|false|false||simplenull|Simple|Modifier|false|false||simplenull|Sentence|Finding|false|false||sentencesnull|Sitting position|Finding|false|false|C0278454;C0278454;C0015385|Sitting
null|Sitting Function|Finding|false|false|C0278454;C0278454;C0015385|Sittingnull|Chairs|Device|false|false||chairnull|Chairperson|Subject|false|false||chairnull|Able (qualifier value)|Finding|false|false||ablenull|Ability|Subject|false|false||ablenull|All extremities|Anatomy|false|false|C2584297;C0277814|all extremitiesnull|All extremities|Anatomy|false|false|C2584297;C0277814|extremities
null|Limb structure|Anatomy|false|false|C2584297;C0277814|extremitiesnull|Fingers|Anatomy|false|false||fingersnull|Fingers, unit of measurement|LabModifier|false|false||fingersnull|Lower extremity>Toes|Anatomy|false|false||toes
null|Toes|Anatomy|false|false||toesnull|Thumb structure|Anatomy|false|false||thumbnull|Psychiatric problem|Disorder|false|false||PSYCH
null|Mental disorders|Disorder|false|false||PSYCHnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Awake (finding)|Finding|false|false||awakenull|Awakening (time frame)|Time|false|false||awakenull|Pleasant|Finding|false|false||pleasantnull|Smiling|Finding|false|false||smilingnull|BRIEF Health Literacy Screening Tool|Finding|false|false||Brief
null|Behavior Rating Inventory of Executive Function|Finding|false|false||Briefnull|Brief|Time|false|false||Briefnull|Shortened|Modifier|false|false||Briefnull|Hospital course|Finding|false|false||Hospital Coursenull|null|Attribute|false|false||Hospital Coursenull|Organization unit type - Hospital|Finding|false|false||Hospitalnull|Hospitals|Device|false|false||Hospitalnull|Hospitals|Entity|false|false||Hospitalnull|Hospital environment|Modifier|false|false||Hospitalnull|Course|Time|false|false||Coursenull|BRIEF Health Literacy Screening Tool|Finding|false|false||BRIEF
null|Behavior Rating Inventory of Executive Function|Finding|false|false||BRIEFnull|Brief|Time|false|false||BRIEFnull|Shortened|Modifier|false|false||BRIEFnull|Organization unit type - Hospital|Finding|false|false||HOSPITALnull|Hospitals|Device|false|false||HOSPITALnull|Hospitals|Entity|false|false||HOSPITALnull|Hospital environment|Modifier|false|false||HOSPITALnull|summary - ActRelationshipSubset|Finding|false|false||SUMMARY
null|Summary (document)|Finding|false|false||SUMMARYnull|Females|Subject|false|false||female
null|Woman|Subject|false|false||femalenull|Female, Self-Report|Modifier|false|false||female
null|Female Phenotype|Modifier|false|false||femalenull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Eating disorder symptom|Disorder|false|false||disordered eatingnull|Eating|Finding|false|false||eatingnull|6-pyruvoyl-tetrahydropterin synthase deficiency|Disorder|false|false||PTSD
null|Post-Traumatic Stress Disorder|Disorder|false|false||PTSDnull|Glutamate Decarboxylase|Drug|false|false||GAD
null|Glutamate Decarboxylase|Drug|false|false||GADnull|Generalized Anxiety Disorder|Disorder|false|false||GADnull|GAD1 wt Allele|Finding|false|false||GAD
null|GAD1 gene|Finding|false|false||GADnull|Panic Disorder|Disorder|false|false||panic disordernull|Panic|Finding|false|false||panicnull|Disease|Disorder|false|false||disordernull|Cancer patients and suicide and depression|Disorder|false|false||depression
null|Mental Depression|Disorder|false|false||depression
null|Depressive disorder|Disorder|false|false||depression
null|Depressed mood|Disorder|false|false||depressionnull|Depression - motion|Finding|false|false||depression
null|null|Finding|false|false||depressionnull|Depression - recess|Modifier|false|false||depressionnull|Functional Relationship|Finding|false|false||functional
null|Function (attribute)|Finding|false|false||functional
null|Functional|Finding|false|false||functionalnull|Neurologic (qualifier value)|Modifier|false|false||neurologicalnull|Disease|Disorder|false|false||disordernull|Therapy Object (animal model)|Finding|false|false||therapy
null|therapeutic aspects|Finding|false|false||therapynull|Therapeutic procedure|Procedure|false|false||therapynull|Session|Finding|false|false||sessionnull|Activity Session|Event|false|false||sessionnull|Weakness|Finding|false|false||weakness
null|Asthenia|Finding|false|false||weaknessnull|Dyskinetic syndrome|Disorder|false|false||abnormal movementnull|Abnormal movement|Finding|false|false||abnormal movementnull|Observation Interpretation - Abnormal|Finding|false|false||abnormal
null|Abnormal|Finding|false|false||abnormalnull|Movement|Finding|false|false||movementnull|Aphasia|Disorder|false|false||aphasianull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Functional Relationship|Finding|false|false||functional
null|Function (attribute)|Finding|false|false||functional
null|Functional|Finding|false|false||functionalnull|Neurologic (qualifier value)|Modifier|false|false||neurologicalnull|Episode of|Time|false|false||episodenull|Neurology speciality|Title|false|false||neurologynull|psychology qualifier|Finding|false|false||psychologynull|Psychology|Title|false|false||psychologynull|Consistent with|Finding|false|false||consistent withnull|Compatible|Modifier|false|false||consistent withnull|Consistent with|Finding|false|false||consistentnull|Functional Relationship|Finding|false|false||functional
null|Function (attribute)|Finding|false|false||functional
null|Functional|Finding|false|false||functionalnull|nervous system disorder|Disorder|false|false||neurological disordernull|Neurologic (qualifier value)|Modifier|false|false||neurologicalnull|Disease|Disorder|false|false||disordernull|Similarity|Modifier|false|false||similarnull|null|Time|false|false||priornull|Presentation|Finding|false|false||presentationnull|RXFP2 gene|Finding|false|false||greatnull|Greater|LabModifier|false|false||great
null|Large|LabModifier|false|false||greatnull|Improvement|Finding|false|false||improvementnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Rehabilitation therapy|Procedure|false|false||rehabnull|Marketing basis - Transitional|Finding|false|false||TRANSITIONALnull|Transitional cell morphology|Modifier|false|false||TRANSITIONALnull|Rehabilitation therapy|Procedure|false|false||rehabnull|Precaution Code - Aggressive|Finding|false|false||aggressive
null|Aggressive behavior|Finding|false|false||aggressive
null|Risk Codes - Aggressive|Finding|false|false||aggressivenull|Aggressive course|Time|false|false||aggressivenull|Entity Risk - aggressive|Modifier|false|false||aggressivenull|Further|Modifier|false|false||furthernull|Improvement|Finding|false|false||improvementnull|functional status (history)|Finding|false|false||functional status
null|Functional Status|Finding|false|false||functional statusnull|null|Attribute|false|false||functional statusnull|Functional Relationship|Finding|false|false||functional
null|Function (attribute)|Finding|false|false||functional
null|Functional|Finding|false|false||functionalnull|What subject filter - Status|Finding|false|false||statusnull|null|Attribute|false|false||statusnull|Social status|Modifier|false|false||status
null|Status|Modifier|false|false||statusnull|On discharge|Time|false|false||On dischargenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Has patient|Finding|false|false||patient hasnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|therapist|Subject|false|false||therapistnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Intermittent|Time|false|false||intermittentnull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|Desire for food|Finding|false|false||appetitenull|Zofran|Drug|false|false||Zofran
null|Zofran|Drug|false|false||Zofrannull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|CIAO3 gene|Finding|false|false||prnnull|As required|Time|false|false||prn
null|Pro Re Nata|Time|false|false||prnnull|Corrected QT Interval|LabModifier|false|false||QTcnull|Electrocardiogram image|Finding|false|false||EKG
null|Electrocardiogram|Finding|false|false||EKGnull|Electrocardiography|Procedure|false|false||EKGnull|Zofran|Drug|false|false||Zofran
null|Zofran|Drug|false|false||Zofrannull|Use - dosing instruction imperative|Finding|false|false||use
null|utilization qualifier|Finding|false|false||use
null|Usage|Finding|false|false||usenull|1 Week|Time|false|false||1 weeknull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|Corrected QT Interval|LabModifier|false|false||QTcnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Has patient|Finding|false|false||Patient hasnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Restrained eating behavior|Finding|false|false||restrictive eatingnull|Eating|Finding|false|false||eatingnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|encouragement|Finding|false|false||encouragementnull|Evidence of (contextual qualifier)|Finding|false|false||evidence ofnull|Evidence|Finding|false|false||evidencenull|Disease|Disorder|false|false||disordernull|Referral category - Inpatient|Finding|false|false||inpatient
null|Patient Class - Inpatient|Finding|false|false||inpatientnull|inpatient encounter|Procedure|false|false||inpatientnull|inpatient|Subject|false|false||inpatientnull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|With meals|Time|false|false||with mealsnull|Meal (occasion for eating)|Finding|false|false||mealsnull|With meals|Time|false|false||mealsnull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|therapist|Subject|false|false||therapistnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Psychiatrist|Subject|false|false||psychiatristnull|Further|Modifier|false|false||furthernull|Titration Method|Procedure|false|false||titrationnull|Referral type - Psychiatric|Finding|false|false||psychiatric
null|Psychiatric|Finding|false|false||psychiatricnull|Psychiatric service|Procedure|false|false||psychiatricnull|Psychiatry Specialty|Title|false|false||psychiatricnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Report (document)|Finding|false|false||reportnull|Reporting|Procedure|false|false||reportnull|null|Attribute|false|false||reportnull|Act Relationship Subset - previous|Time|false|false||previous
null|Previous|Time|false|false||previousnull|Sensitivity (Personality)|Finding|false|false||sensitivity
null|Hypersensitivity|Finding|false|false||sensitivity
null|Antimicrobial susceptibility|Finding|false|false||sensitivitynull|stimulus sensitivity|Modifier|false|false||sensitivity
null|Signal Sensitivity|Modifier|false|false||sensitivitynull|Statistical sensitivity|LabModifier|false|false||sensitivity
null|Diagnostic Sensitivity|LabModifier|false|false||sensitivitynull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Concern|Finding|false|false||concernnull|Possible|Finding|false|false||possiblenull|Possible diagnosis|Modifier|false|false||possible
null|Possibly Related to Intervention|Modifier|false|false||possiblenull|Bipolar Disorder|Disorder|false|false||bipolar disordernull|Bipolar|Modifier|false|false||bipolarnull|Disease|Disorder|false|false||disordernull|Diagnosis Classification - Diagnosis|Finding|false|false||diagnosis
null|diagnosis aspects|Finding|false|false||diagnosisnull|Diagnosis|Procedure|false|false||diagnosisnull|null|Attribute|false|false||diagnosisnull|Pending - Allergy Clinical Status|Finding|false|false||pending
null|Pending - referral status|Finding|false|false||pendingnull|Pending - status|Time|false|false||pendingnull|pending - ManagedParticipationStatus|Modifier|false|false||pending
null|pending - RoleStatus|Modifier|false|false||pending
null|Pending - Day type|Modifier|false|false||pendingnull|Thiamine Drug Class|Drug|false|false||thiamine
null|thiamine|Drug|false|false||thiamine
null|thiamine|Drug|false|false||thiamine
null|thiamine|Drug|false|false||thiamine
null|Thiamine Drug Class|Drug|false|false||thiaminenull|Thiamine measurement|Procedure|false|false||thiaminenull|Admission Level of Care Code - Acute|Finding|false|false||ACUTE
null|Acute - Triage Code|Finding|false|false||ACUTEnull|acute|Time|false|false||ACUTEnull|Glutamate Decarboxylase|Drug|false|false||GAD
null|Glutamate Decarboxylase|Drug|false|false||GADnull|Generalized Anxiety Disorder|Disorder|false|false||GADnull|GAD1 wt Allele|Finding|false|false||GAD
null|GAD1 gene|Finding|false|false||GADnull|Panic Disorder|Disorder|false|false||Panic disordernull|Panic|Finding|false|false||Panicnull|Disease|Disorder|false|false||disordernull|Cancer patients and suicide and depression|Disorder|false|false||Depression
null|Mental Depression|Disorder|false|false||Depression
null|Depressive disorder|Disorder|false|false||Depression
null|Depressed mood|Disorder|false|false||Depressionnull|Depression - motion|Finding|false|false||Depression
null|null|Finding|false|false||Depressionnull|Depression - recess|Modifier|false|false||Depressionnull|6-pyruvoyl-tetrahydropterin synthase deficiency|Disorder|false|false||PTSD
null|Post-Traumatic Stress Disorder|Disorder|false|false||PTSDnull|Dissociative neurological symptom disorder (disorder)|Disorder|false|false||Functional neurological disorder
null|Conversion disorder|Disorder|false|false||Functional neurological disordernull|Functional Relationship|Finding|false|false||Functional
null|Function (attribute)|Finding|false|false||Functional
null|Functional|Finding|false|false||Functionalnull|nervous system disorder|Disorder|false|false||neurological disordernull|Neurologic (qualifier value)|Modifier|false|false||neurologicalnull|Disease|Disorder|false|false||disordernull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Therapy Object (animal model)|Finding|false|false||therapy
null|therapeutic aspects|Finding|false|false||therapynull|Therapeutic procedure|Procedure|false|false||therapynull|Session|Finding|false|false||sessionnull|Activity Session|Event|false|false||sessionnull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Onset of (contextual qualifier)|Modifier|false|false||onset ofnull|Onset of (contextual qualifier)|Modifier|false|false||onsetnull|Age of Onset|LabModifier|false|false||onsetnull|Weakness|Finding|false|false||weakness
null|Asthenia|Finding|false|false||weaknessnull|Dyskinetic syndrome|Disorder|false|false||abnormal movementnull|Abnormal movement|Finding|false|false||abnormal movementnull|Observation Interpretation - Abnormal|Finding|false|false||abnormal
null|Abnormal|Finding|false|false||abnormalnull|Movement|Finding|false|false||movementnull|Aphasia|Disorder|false|false||aphasianull|contextual factors|Finding|false|false||settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|Potential|Modifier|false|false||potentialnull|Precipitating Factors|Attribute|false|false||triggernull|Triggered by|Modifier|false|false||triggernull|Shadow|Finding|false|false||shadowsnull|Door (physical object)|Device|false|false||doornull|therapist|Subject|false|false||therapistnull|Several|LabModifier|false|false||severalnull|week|Time|false|false||weeksnull|More|LabModifier|false|false||morenull|Stress|Finding|false|false||stressednull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Holidays|Event|false|false||holidaysnull|mycolate outer membrane|Anatomy|false|false|C0878676;C0038436|momnull|Multiple of the median|LabModifier|false|false||momnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||majornull|Major <Sympycninae>|Entity|false|false||majornull|Major|Modifier|false|false||majornull|Precipitating Factors|Attribute|false|false||triggernull|Triggered by|Modifier|false|false||triggernull|6-pyruvoyl-tetrahydropterin synthase deficiency|Disorder|false|false|C3811401|PTSD
null|Post-Traumatic Stress Disorder|Disorder|false|false|C3811401|PTSDnull|therapist|Subject|false|false||therapistnull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Sex Behavior|Finding|false|false||sexualnull|physical examination (physical finding)|Finding|false|false||physical
null|Physical|Finding|false|false||physicalnull|Physical Examination|Procedure|false|false||physicalnull|Participation Mode - verbal|Finding|false|false||verbalnull|Consent Mode - Verbal|Procedure|false|false||verbalnull|Verbal|Modifier|false|false||verbalnull|Drug abuse|Disorder|false|false||abusenull|Victim of abuse (finding)|Finding|false|false||abusenull|Abuse|Event|false|false||abusenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Very|Modifier|false|false||verynull|Presentation|Finding|false|false||presentationnull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Functional Relationship|Finding|false|false||functional
null|Function (attribute)|Finding|false|false||functional
null|Functional|Finding|false|false||functionalnull|Neurologic Symptoms|Finding|false|false||neurological symptomsnull|Neurologic (qualifier value)|Modifier|false|false||neurologicalnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Weakness|Finding|false|false||weakness
null|Asthenia|Finding|false|false||weaknessnull|Observation Interpretation - Abnormal|Finding|false|false||abnormal
null|Abnormal|Finding|false|false||abnormalnull|Movement|Finding|false|false||movementnull|Aphasia|Disorder|false|false||aphasianull|Impaired|Finding|false|false||impairednull|Function (attribute)|Finding|false|false||functioning
null|Functional|Finding|false|false||functioningnull|Concern|Finding|false|false||concernnull|Catatonia|Disorder|false|false||catatonianull|Ativan|Drug|false|false||ativan
null|Ativan|Drug|false|false||ativannull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|Anxiety Disorders|Disorder|false|false||anxiety
null|Anxiety|Disorder|false|false||anxietynull|Anxiety symptoms|Finding|false|false||anxietynull|Psychiatry Specialty|Title|false|false||Psychiatrynull|criteria|Finding|false|false||criterianull|Similarity|Modifier|false|false||similarnull|Episode of|Time|false|false||episodenull|ferryl iron|Drug|false|false||IV ironnull|Iron Drug Class|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|Ferrum metallicum, Homeopathic preparation|Drug|false|false||ironnull|Iron measurement|Procedure|false|false||ironnull|Infusion route|Finding|false|false||infusionnull|Infusion procedures|Procedure|false|false||infusionnull|neurology services (treatment)|Procedure|false|false||neurology servicenull|Neurology service|Entity|false|false||neurology servicenull|Neurology speciality|Title|false|false||neurologynull|ActInformationPrivacyReason - service|Finding|false|false||servicenull|Software Service|Device|false|false||servicenull|Services|Event|false|false||servicenull|Dissociative neurological symptom disorder (disorder)|Disorder|false|false||functional neurological disorder
null|Conversion disorder|Disorder|false|false||functional neurological disordernull|Functional Relationship|Finding|false|false||functional
null|Function (attribute)|Finding|false|false||functional
null|Functional|Finding|false|false||functionalnull|nervous system disorder|Disorder|false|false||neurological disordernull|Neurologic (qualifier value)|Modifier|false|false||neurologicalnull|Disease|Disorder|false|false||disordernull|Rehabilitation therapy|Procedure|false|false||rehabnull|Once a day, at bedtime|Time|false|false||QHSnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|therapist|Subject|false|false||therapistnull|Sensitive|Finding|false|false||is sensitive tonull|Sensitive|Finding|false|false||sensitive tonull|Sensitive|Finding|false|false||sensitivenull|stimulus sensitivity|Modifier|false|false||sensitivenull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Selective Serotonin Reuptake Inhibitors|Drug|false|false||SSRIsnull|Manic|Disorder|false|false||manicnull|Manic mood|Finding|false|false||manicnull|Bipolar Disorder|Disorder|false|false||bipolar disordernull|Bipolar|Modifier|false|false||bipolarnull|Disease|Disorder|false|false||disordernull|Neurology speciality|Title|false|false||neuronull|Neurologic (qualifier value)|Modifier|false|false||neuronull|Psychiatry Specialty|Title|false|false||psychiatrynull|Consistent with|Finding|false|false||consistent withnull|Compatible|Modifier|false|false||consistent withnull|Consistent with|Finding|false|false||consistentnull|Catatonia|Disorder|false|false||catatonianull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Dissociative neurological symptom disorder (disorder)|Disorder|false|false||functional neurological disorder
null|Conversion disorder|Disorder|false|false||functional neurological disordernull|Functional Relationship|Finding|false|false||functional
null|Function (attribute)|Finding|false|false||functional
null|Functional|Finding|false|false||functionalnull|nervous system disorder|Disorder|false|false||neurological disordernull|Neurologic (qualifier value)|Modifier|false|false||neurologicalnull|Disease|Disorder|false|false||disordernull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Rehabilitation therapy|Procedure|false|false||rehabnull|Precaution Code - Aggressive|Finding|false|false||aggressive
null|Aggressive behavior|Finding|false|false||aggressive
null|Risk Codes - Aggressive|Finding|false|false||aggressivenull|Aggressive course|Time|false|false||aggressivenull|Entity Risk - aggressive|Modifier|false|false||aggressivenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Once a day, at bedtime|Time|false|false||qhsnull|Eating|Finding|false|false||eatingnull|Restrained eating behavior|Finding|false|false||Restrictive eatingnull|Eating|Finding|false|false||eatingnull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Restrained eating behavior|Finding|false|false||restrictive eatingnull|Eating|Finding|false|false||eatingnull|Bradycardia by ECG Finding|Finding|false|false||bradycardia
null|Bradycardia|Finding|false|false||bradycardianull|Electrolyte [EPC]|Drug|false|false||electrolyte
null|Electrolytes|Drug|false|false||electrolyte
null|Electrolytes|Drug|false|false||electrolytenull|Congenital Abnormality|Disorder|false|false||abnormalitiesnull|teratologic|Finding|false|false||abnormalitiesnull|therapist|Subject|false|false||therapistnull|Eating disorder symptom|Disorder|false|false||disordered eatingnull|Eating|Finding|false|false||eatingnull|Much worse|Finding|false|false||much worsenull|Much|Finding|false|false||muchnull|Observation Interpretation - worse|Finding|false|false||worse
null|Worse|Finding|false|false||worsenull|Worsening (qualifier value)|Modifier|false|false||worsenull|month|Time|false|false||monthsnull|contextual factors|Finding|false|false||settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|travel|Finding|false|false|C0175218;C0162435|travelingnull|Very Much|Finding|false|false|C0175218;C0162435|a lotnull|Stock (in-store merchandise)|Finding|false|false|C0175218;C0162435|lotnull|nucleus of the lateral olfactory tract|Anatomy|false|false|C2984081;C0040802;C1710198;C0043227|lot
null|Olfactory tract|Anatomy|false|false|C2984081;C0040802;C1710198;C0043227|lotnull|Lot (entire collection)|Modifier|false|false||lotnull|Work|Event|false|false|C0175218;C0162435|worknull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|Program|Drug|false|false||program
null|Program|Drug|false|false||programnull|Program - framework of goals|Finding|false|false||program
null|Programs - Publication Format|Finding|false|false||program
null|Programs|Finding|false|false||programnull|therapist|Subject|false|false||therapistnull|Nutrition, Calories|LabModifier|false|false||calories
null|calorie unit of energy|LabModifier|false|false||caloriesnull|Smaller|Modifier|false|false||lessnull|Less Than|LabModifier|false|false||lessnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Language Ability Proficiency - Good|Finding|false|false||good
null|Language Proficiency - Good|Finding|false|false||goodnull|Specimen Quality - Good|Modifier|false|false||good
null|Good|Modifier|false|false||goodnull|Persons|Subject|false|false||peoplenull|Review of|Finding|false|false||review ofnull|Review (Publication Type)|Finding|false|false||review
null|Act Class - review|Finding|false|false||reviewnull|ATP5F1A gene|Finding|false|false||OMRnull|Finding of body mass index|Finding|false|false||BMInull|null|Attribute|false|false||BMI
null|Body mass index|Attribute|false|false||BMInull|Current (present time)|Time|false|false||currentlynull|Electrolyte [EPC]|Drug|true|false||electrolyte
null|Electrolytes|Drug|true|false||electrolyte
null|Electrolytes|Drug|true|false||electrolytenull|Congenital Abnormality|Disorder|true|false||abnormalitiesnull|teratologic|Finding|true|false||abnormalitiesnull|Desire for food|Finding|false|false||appetitenull|Neurologic Symptoms|Finding|false|false||neurological symptomsnull|Neurologic (qualifier value)|Modifier|false|false||neurologicalnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Nutrition (function)|Finding|false|false||nutrition
null|Nutritional status|Finding|false|false||nutrition
null|Nutrition outcomes|Finding|false|false||nutritionnull|Feeding and dietary regimes|Procedure|false|false||nutrition
null|Nutritional Study|Procedure|false|false||nutritionnull|Science of nutrition|Title|false|false||nutritionnull|Processing type - Evaluation|Finding|false|false||evaluationnull|Evaluation procedure|Procedure|false|false||evaluation
null|Evaluation|Procedure|false|false||evaluationnull|Patient need for (contextual qualifier)|Finding|true|false||need fornull|Patient need for (contextual qualifier)|Finding|true|false||neednull|Needs|Modifier|false|false||neednull|Eating Disorders|Disorder|false|false||eating disordernull|Eating|Finding|false|false||eatingnull|Disease|Disorder|false|false||disordernull|Clinical trial protocol document|Finding|false|false||protocol
null|Study Protocol|Finding|false|false||protocol
null|Protocols documentation|Finding|false|false||protocol
null|Protocol - answer to question|Finding|false|false||protocol
null|Library Protocol|Finding|false|false||protocolnull|Referral category - Inpatient|Finding|false|false||inpatient
null|Patient Class - Inpatient|Finding|false|false||inpatientnull|inpatient encounter|Procedure|false|false||inpatientnull|inpatient|Subject|false|false||inpatientnull|Ensure (product)|Drug|false|false||Ensurenull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787|Heart
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787|Heartnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|Heartnull|Chest>Heart|Anatomy|false|false|C0153957;C0153500;C0795691|Heart
null|Heart|Anatomy|false|false|C0153957;C0153500;C0795691|Heartnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Electrolytes|Drug|false|false||Electrolytes
null|Electrolytes|Drug|false|false||Electrolytes
null|Electrolyte [EPC]|Drug|false|false||Electrolytesnull|thyrotropin|Drug|false|false||TSH
null|thyrotropin|Drug|false|false||TSH
null|thyrotropin|Drug|false|false||TSHnull|Thyroid stimulating hormone measurement|Procedure|false|false||TSHnull|null|Attribute|false|false||TSHnull|TNFAIP1 wt Allele|Finding|false|false||B12
null|NDUFB3 gene|Finding|false|false||B12
null|TNFAIP1 gene|Finding|false|false||B12null|Levels (qualifier value)|Modifier|false|false||levelsnull|Thiamin supplementation|Procedure|false|false||thiamine supplementationnull|Thiamine Drug Class|Drug|false|false||thiamine
null|thiamine|Drug|false|false||thiamine
null|thiamine|Drug|false|false||thiamine
null|thiamine|Drug|false|false||thiamine
null|Thiamine Drug Class|Drug|false|false||thiaminenull|Thiamine measurement|Procedure|false|false||thiaminenull|Dietary Supplementation|Procedure|false|false||supplementationnull|Zofran|Drug|false|false||Zofran
null|Zofran|Drug|false|false||Zofrannull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|Corrected QT Interval|LabModifier|false|false||QTcnull|Core Specimen|Finding|false|false|C1167518|COREnull|viral nucleocapsid location|Anatomy|false|false|C1879489;C3274653|COREnull|Processor Core|Device|false|false||CORE
null|Core Device|Device|false|false||COREnull|Core|Modifier|false|false||COREnull|Measures (attribute)|Finding|false|false|C1167518|MEASURESnull|Measures|LabModifier|false|false||MEASURESnull|MDF Attribute Type - Code|Finding|false|false||CODE
null|A Codes|Finding|false|false||CODE
null|Code|Finding|false|false||CODEnull|Coding|Event|false|false||CODEnull|Full|Modifier|false|false||fullnull|MDF Attribute Type - Code|Finding|false|false||code
null|A Codes|Finding|false|false||code
null|Code|Finding|false|false||codenull|Coding|Event|false|false||codenull|Contact - HL7 Attribution|Finding|false|false||CONTACT
null|Contact with|Finding|false|false||CONTACT
null|Communication Contact|Finding|false|false||CONTACTnull|contact person|Subject|false|false||CONTACTnull|Physical contact|Phenomenon|false|false||CONTACTnull|Personal Contact|Event|false|false||CONTACTnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Request - ActReason|Finding|false|false||request
null|request - ActMood|Finding|false|false||request
null|Question (inquiry)|Finding|false|false||requestnull|null|Event|false|false||requestnull|Relationship - Mother|Finding|false|false||mothernull|Mother (person)|Subject|false|false||mothernull|Consent Non-Disclosure Reason - Emergency|Finding|false|false||Emergency
null|Admission Type - Emergency|Finding|false|false||Emergency
null|Referral category - Emergency|Finding|false|false||Emergency
null|Emergencies [Disease/Finding]|Finding|false|false||Emergency
null|Consent Bypass Reason - Emergency|Finding|false|false||Emergency
null|Level of Care - Emergency|Finding|false|false||Emergency
null|Certification patient type - Emergency|Finding|false|false||Emergency
null|Encounter Admission Source - emergency|Finding|false|false||Emergency
null|Patient Class - Emergency|Finding|false|false||Emergency
null|Visit Priority Code - Emergency|Finding|false|false||Emergencynull|emergency encounter|Procedure|false|false||Emergencynull|Specialty Type - Emergency|Title|false|false||Emergencynull|Emergency Situation|Phenomenon|false|false||Emergencynull|Bale out|Time|false|false||Emergencynull|Contacts|Procedure|false|false||Contactsnull|Uncle|Subject|false|false||Unclenull|therapist|Subject|false|false||Therapistnull|null|Finding|false|false||coordinates
null|Coordinated|Finding|false|false||coordinatesnull|Coordinate on an axis or a grid|Modifier|false|false||coordinatesnull|Continuity Assessment Record and Evaluation|Finding|false|false||care
null|In care (finding)|Finding|false|false||carenull|care activity|Event|false|false||carenull|Availability of|Finding|false|false||availablenull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|MEDICATION LIST|Finding|false|false||Medication listnull|Pharmaceutical Preparations|Drug|false|false||Medicationnull|medication - HL7 publishing domain|Finding|false|false||Medication
null|Medications|Finding|false|false||Medicationnull|List|Finding|false|false||list
null|Sequence Data Type|Finding|false|false||listnull|Accurate (qualifier value)|Modifier|false|false||accuratenull|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||completenull|Completion Status for valid values - Complete|Finding|false|false||complete
null|Data operation - complete|Finding|false|false||complete
null|Finish - dosing instruction imperative|Finding|false|false||completenull|Complete|Modifier|false|false||completenull|Once a day, at bedtime|Time|false|false||QHSnull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin Drug Class|Drug|false|false||Multivitamins
null|Multivitamin Drug Class|Drug|false|false||Multivitaminsnull|Minerals|Drug|false|false||mineralsnull|Tablet Dosage Form|Drug|false|false||TABnull|Tablet Dosing Unit|LabModifier|false|false||TABnull|Daily|Time|false|false||DAILYnull|ondansetron|Drug|false|false||Ondansetron
null|ondansetron|Drug|false|false||Ondansetronnull|Optical Doppler Tomography|Procedure|false|false||ODTnull|Every eight hours|Time|false|false||Q8Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Nausea and vomiting|Finding|false|false||Nausea/Vomitingnull|Nausea|Finding|false|false||Nauseanull|null|Attribute|false|false||Nauseanull|Vomiting|Finding|false|false||Vomitingnull|Firstly|Modifier|false|false||Firstnull|First (number)|LabModifier|false|false||Firstnull|Line Specimen|Drug|false|false||Line
null|Long Interspersed Elements|Drug|false|false||Line
null|Long Interspersed Elements|Drug|false|false||Linenull|line source specimen code|Finding|false|false||Linenull|Intravascular line|Device|false|false||Linenull|Linear|Modifier|false|false||Linenull|Line Unit of Length|LabModifier|false|false||Linenull|Thiamine Drug Class|Drug|false|false||Thiamine
null|thiamine|Drug|false|false||Thiamine
null|thiamine|Drug|false|false||Thiamine
null|thiamine|Drug|false|false||Thiamine
null|Thiamine Drug Class|Drug|false|false||Thiaminenull|Thiamine measurement|Procedure|false|false||Thiaminenull|Daily|Time|false|false||DAILYnull|Once a day, at bedtime|Time|false|false||QHSnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|long-term care|Procedure|false|false||Extended Carenull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|In care (finding)|Finding|false|false||Care
null|Continuity Assessment Record and Evaluation|Finding|false|false||Carenull|care activity|Event|false|false||Carenull|ADMIN.FACILITY|Finding|false|false||Facilitynull|Facility (object)|Device|false|false||Facilitynull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Dissociative neurological symptom disorder (disorder)|Disorder|false|false||Functional neurological disorder
null|Conversion disorder|Disorder|false|false||Functional neurological disordernull|Functional Relationship|Finding|false|false||Functional
null|Function (attribute)|Finding|false|false||Functional
null|Functional|Finding|false|false||Functionalnull|nervous system disorder|Disorder|false|false||neurological disordernull|Neurologic (qualifier value)|Modifier|false|false||neurologicalnull|Disease|Disorder|false|false||disordernull|Glutamate Decarboxylase|Drug|false|false||GAD
null|Glutamate Decarboxylase|Drug|false|false||GADnull|Generalized Anxiety Disorder|Disorder|false|false||GADnull|GAD1 wt Allele|Finding|false|false||GAD
null|GAD1 gene|Finding|false|false||GADnull|Cancer patients and suicide and depression|Disorder|false|false||depression
null|Mental Depression|Disorder|false|false||depression
null|Depressive disorder|Disorder|false|false||depression
null|Depressed mood|Disorder|false|false||depressionnull|Depression - motion|Finding|false|false||depression
null|null|Finding|false|false||depressionnull|Depression - recess|Modifier|false|false||depressionnull|6-pyruvoyl-tetrahydropterin synthase deficiency|Disorder|false|false||PTSD
null|Post-Traumatic Stress Disorder|Disorder|false|false||PTSDnull|Eating disorder symptom|Disorder|false|false||disordered eatingnull|Eating|Finding|false|false||eatingnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Disease|Disorder|false|false||Conditionnull|Logical Condition|Finding|false|false||Conditionnull|null|Attribute|false|false||Conditionnull|Condition|Modifier|false|false||Conditionnull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|BORNHOLM EYE DISEASE|Disorder|false|false||Bednull|Bachelor of Education|Finding|false|false||Bednull|Beds|Device|false|false||Bednull|Patient Location - Bed|Modifier|false|false||Bednull|Helping Behavior|Finding|false|false||assistancenull|Assisted (qualifier value)|Modifier|false|false||assistancenull|Chairs|Device|false|false||chairnull|Chairperson|Subject|false|false||chairnull|has wheelchair at home (history)|Finding|false|false||wheelchair
null|Wheelchair Usually Used|Finding|false|false||wheelchairnull|wheelchair|Device|false|false||wheelchairnull|Discharge instructions|Finding|false|false||Discharge Instructionsnull|hospital discharge instructions (treatment)|Procedure|false|false||Discharge Instructionsnull|null|Attribute|false|false||Discharge Instructionsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructionsnull|FBXW7-AS1 gene|Finding|false|false||Dearnull|Role Privilege|Finding|false|false||privilege
null|User Privilege|Finding|false|false||privilege
null|Privilege|Finding|false|false||privilegenull|care of - AddressPartType|Finding|false|false||care ofnull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Organization unit type - Hospital|Finding|false|false||HOSPITALnull|Hospitals|Device|false|false||HOSPITALnull|Hospitals|Entity|false|false||HOSPITALnull|Hospital environment|Modifier|false|false||HOSPITALnull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Speaking (function)|Finding|false|false||speakingnull|Occur (action)|Event|false|false||HAPPENEDnull|Organization unit type - Hospital|Finding|false|false||HOSPITALnull|Hospitals|Device|false|false||HOSPITALnull|Hospitals|Entity|false|false||HOSPITALnull|Hospital environment|Modifier|false|false||HOSPITALnull|Neurologists|Subject|false|false||neurologistsnull|Dissociative neurological symptom disorder (disorder)|Disorder|false|false||functional neurological disorder
null|Conversion disorder|Disorder|false|false||functional neurological disordernull|Functional Relationship|Finding|false|false||functional
null|Function (attribute)|Finding|false|false||functional
null|Functional|Finding|false|false||functionalnull|nervous system disorder|Disorder|false|false||neurological disordernull|Neurologic (qualifier value)|Modifier|false|false||neurologicalnull|Disease|Disorder|false|false||disordernull|physical examination (physical finding)|Finding|false|false||physical
null|Physical|Finding|false|false||physicalnull|Physical Examination|Procedure|false|false||physicalnull|Occupational therapist|Subject|false|false||occupational therapistsnull|Occupational|Finding|false|false||occupationalnull|therapist|Subject|false|false||therapistsnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Organization unit type - Hospital|Finding|false|false||HOSPITALnull|Hospitals|Device|false|false||HOSPITALnull|Hospitals|Entity|false|false||HOSPITALnull|Hospital environment|Modifier|false|false||HOSPITALnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Physicians|Subject|false|false||doctorsnull|Appointments|Event|false|false||appointmentsnull|physical examination (physical finding)|Finding|false|false||physical
null|Physical|Finding|false|false||physicalnull|Physical Examination|Procedure|false|false||physicalnull|Occupational|Finding|false|false||occupationalnull|therapist|Subject|false|false||therapistsnull|Vitelliform Macular Dystrophy|Disorder|false|false||bestnull|BEST1 wt Allele|Finding|false|false||best
null|BEST1 gene|Finding|false|false||bestnull|best (quality)|Modifier|false|false||bestnull|Care team|Finding|false|false||Care Teamnull|null|Attribute|false|false||Care Teamnull|In care (finding)|Finding|false|false||Care
null|Continuity Assessment Record and Evaluation|Finding|false|false||Carenull|care activity|Event|false|false||Carenull|Team|Subject|false|false||Teamnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions