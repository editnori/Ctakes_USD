 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|50,59|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|50,59|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|50,64|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|84,93|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|84,93|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|84,93|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|84,93|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|84,93|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|84,98|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|116,121|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|116,121|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|116,121|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|140,143|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|140,143|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|140,143|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|140,143|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|140,143|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|151,158|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|151,158|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|160,168|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|SIMPLE_SEGMENT|171,180|false|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|171,180|false|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|171,180|false|false|false|C0020517|Hypersensitivity|Allergies
Attribute|Clinical Attribute|SIMPLE_SEGMENT|192,201|false|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|192,201|false|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|192,201|false|false|false|C0020517|Hypersensitivity|Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|204,226|true|false|false|C0041755|Adverse reaction to drug|Adverse Drug Reactions
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|212,216|false|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|Drug
Finding|Finding|SIMPLE_SEGMENT|212,216|false|false|false|C0740721|Drug problem|Drug
Finding|Pathologic Function|SIMPLE_SEGMENT|212,226|true|false|false|C0041755|Adverse reaction to drug|Drug Reactions
Event|Event|SIMPLE_SEGMENT|217,226|false|false|false|||Reactions
Event|Event|SIMPLE_SEGMENT|229,238|false|false|false|||Attending
Finding|Functional Concept|SIMPLE_SEGMENT|229,238|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|SIMPLE_SEGMENT|246,261|false|false|false|C0277786|Chief complaint (finding)|Chief Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|252,261|false|false|false|C3864418||Complaint
Event|Event|SIMPLE_SEGMENT|252,261|false|false|false|||Complaint
Finding|Finding|SIMPLE_SEGMENT|252,261|false|false|false|C5441521|Complaint (finding)|Complaint
Finding|Idea or Concept|SIMPLE_SEGMENT|263,272|false|false|false|C1546960|Patient Outcome - Worsening|Worsening
Anatomy|Body Location or Region|SIMPLE_SEGMENT|273,276|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|ABD
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|273,276|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|ABD
Event|Event|SIMPLE_SEGMENT|277,287|false|false|false|||distension
Finding|Finding|SIMPLE_SEGMENT|277,287|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distension
Finding|Pathologic Function|SIMPLE_SEGMENT|277,287|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distension
Attribute|Clinical Attribute|SIMPLE_SEGMENT|292,296|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|292,296|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|292,296|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|292,296|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Classification|SIMPLE_SEGMENT|300,305|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|SIMPLE_SEGMENT|306,314|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|306,314|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|318,336|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|327,336|false|false|false|C0945766||Procedure
Event|Event|SIMPLE_SEGMENT|327,336|false|false|false|||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|327,336|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|327,336|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|327,336|false|false|false|C0184661|Interventional procedure|Procedure
Event|Event|SIMPLE_SEGMENT|338,350|false|false|false|||Paracentesis
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|338,350|false|false|false|C0034115|Paracentesis|Paracentesis
Event|Event|SIMPLE_SEGMENT|354,361|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|354,361|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|354,361|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|354,361|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|354,364|false|false|false|C0262926|Medical History|History of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|354,380|false|false|false|C0488508||History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|354,380|false|false|false|C0262512|History of present illness (finding)|History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|365,372|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Idea or Concept|SIMPLE_SEGMENT|365,372|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Finding|SIMPLE_SEGMENT|365,380|false|false|false|C4264312|Present illness|Present Illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|373,380|false|false|false|C0221423|Illness (finding)|Illness
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|386,389|false|false|false|C0019196;C0220847|Hepatitis C;hepatitis C virus|HCV
Disorder|Virus|SIMPLE_SEGMENT|386,389|false|false|false|C0019196;C0220847|Hepatitis C;hepatitis C virus|HCV
Event|Event|SIMPLE_SEGMENT|386,389|false|false|false|||HCV
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|390,399|false|false|false|C0023890;C1623038|Cirrhosis;Liver Cirrhosis|cirrhosis
Event|Event|SIMPLE_SEGMENT|390,399|false|false|false|||cirrhosis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|404,411|false|false|false|C0003962|Ascites|ascites
Event|Event|SIMPLE_SEGMENT|404,411|false|false|false|||ascites
Finding|Pathologic Function|SIMPLE_SEGMENT|404,411|false|false|false|C5441966|Peritoneal Effusion|ascites
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|413,416|false|false|false|C0019682;C0019693|HIV;HIV Infections|hiv
Disorder|Virus|SIMPLE_SEGMENT|413,416|false|false|false|C0019682;C0019693|HIV;HIV Infections|hiv
Drug|Immunologic Factor|SIMPLE_SEGMENT|413,416|false|false|false|C0086413|HIV Vaccine|hiv
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|413,416|false|false|false|C0086413|HIV Vaccine|hiv
Event|Event|SIMPLE_SEGMENT|413,416|false|false|false|||hiv
Drug|Organic Chemical|SIMPLE_SEGMENT|420,423|false|false|false|C0052432|artesunate|ART
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|420,423|false|false|false|C0052432|artesunate|ART
Event|Event|SIMPLE_SEGMENT|420,423|false|false|false|||ART
Finding|Gene or Genome|SIMPLE_SEGMENT|420,423|false|false|false|C1412286;C3890191|AGRP gene;AGRP wt Allele|ART
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|420,423|false|false|false|C0872104;C1963724|Antiretroviral therapy;Assisted Reproductive Technologies|ART
Event|Event|SIMPLE_SEGMENT|429,433|false|false|false|||IVDU
Finding|Individual Behavior|SIMPLE_SEGMENT|429,433|false|false|false|C0699778|intravenous drug use|IVDU
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|435,439|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|435,439|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|SIMPLE_SEGMENT|435,439|false|false|false|||COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|435,439|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|451,455|false|false|false|C0038436;C0878676|6-pyruvoyl-tetrahydropterin synthase deficiency;Post-Traumatic Stress Disorder|PTSD
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|451,455|false|false|false|C0038436;C0878676|6-pyruvoyl-tetrahydropterin synthase deficiency;Post-Traumatic Stress Disorder|PTSD
Event|Event|SIMPLE_SEGMENT|451,455|false|false|false|||PTSD
Event|Event|SIMPLE_SEGMENT|457,466|false|false|false|||presented
Finding|Idea or Concept|SIMPLE_SEGMENT|484,493|false|false|false|C1546960|Patient Outcome - Worsening|worsening
Anatomy|Body Location or Region|SIMPLE_SEGMENT|494,497|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|abd
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|494,497|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|abd
Event|Event|SIMPLE_SEGMENT|499,509|false|false|false|||distension
Finding|Finding|SIMPLE_SEGMENT|499,509|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distension
Finding|Pathologic Function|SIMPLE_SEGMENT|499,509|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distension
Finding|Intellectual Product|SIMPLE_SEGMENT|520,524|false|false|false|C1561540|Transaction counts and value totals - week|week
Event|Event|SIMPLE_SEGMENT|531,538|false|false|false|||reports
Finding|Idea or Concept|SIMPLE_SEGMENT|539,543|false|false|false|C0036588;C1551994|Self;subscriber - self|self
Finding|Intellectual Product|SIMPLE_SEGMENT|539,543|false|false|false|C0036588;C1551994|Self;subscriber - self|self
Drug|Organic Chemical|SIMPLE_SEGMENT|558,563|false|false|false|C0699992|Lasix|lasix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|558,563|false|false|false|C0699992|Lasix|lasix
Event|Event|SIMPLE_SEGMENT|558,563|false|false|false|||lasix
Event|Event|SIMPLE_SEGMENT|568,581|false|false|false|||spirnolactone
Finding|Gene or Genome|SIMPLE_SEGMENT|593,596|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Event|Event|SIMPLE_SEGMENT|616,620|false|false|false|||like
Drug|Chemical|SIMPLE_SEGMENT|686,695|false|false|false|C0220806|Chemicals|chemicals
Event|Event|SIMPLE_SEGMENT|686,695|false|false|false|||chemicals
Finding|Functional Concept|SIMPLE_SEGMENT|729,739|false|false|false|C0443288;C1548390;C1549594;C1610594|Confidentiality - restricted;Confidentiality code - Restricted;Document Confidentiality Status - Restricted;Restricted|restricted
Finding|Idea or Concept|SIMPLE_SEGMENT|729,739|false|false|false|C0443288;C1548390;C1549594;C1610594|Confidentiality - restricted;Confidentiality code - Restricted;Document Confidentiality Status - Restricted;Restricted|restricted
Finding|Intellectual Product|SIMPLE_SEGMENT|729,739|false|false|false|C0443288;C1548390;C1549594;C1610594|Confidentiality - restricted;Confidentiality code - Restricted;Document Confidentiality Status - Restricted;Restricted|restricted
Drug|Food|SIMPLE_SEGMENT|740,745|false|false|false|C0012155|Diet|diets
Event|Event|SIMPLE_SEGMENT|740,745|false|false|false|||diets
Finding|Intellectual Product|SIMPLE_SEGMENT|759,763|false|false|false|C1561540|Transaction counts and value totals - week|week
Event|Event|SIMPLE_SEGMENT|769,774|false|false|false|||notes
Finding|Idea or Concept|SIMPLE_SEGMENT|801,810|false|false|false|C1546960|Patient Outcome - Worsening|worsening
Anatomy|Body Location or Region|SIMPLE_SEGMENT|811,814|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|abd
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|811,814|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|abd
Event|Event|SIMPLE_SEGMENT|815,825|false|false|false|||distension
Finding|Finding|SIMPLE_SEGMENT|815,825|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distension
Finding|Pathologic Function|SIMPLE_SEGMENT|815,825|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distension
Event|Event|SIMPLE_SEGMENT|830,840|false|false|false|||discomfort
Finding|Sign or Symptom|SIMPLE_SEGMENT|830,840|false|false|false|C2364135|Discomfort|discomfort
Event|Event|SIMPLE_SEGMENT|847,853|false|false|false|||denies
Attribute|Clinical Attribute|SIMPLE_SEGMENT|858,863|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|858,863|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|858,863|false|false|false|C0013604|Edema|edema
Event|Event|SIMPLE_SEGMENT|868,871|false|false|false|||SOB
Finding|Sign or Symptom|SIMPLE_SEGMENT|868,871|false|false|false|C0013404|Dyspnea|SOB
Event|Event|SIMPLE_SEGMENT|876,885|false|false|false|||orthopnea
Finding|Finding|SIMPLE_SEGMENT|876,885|false|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|876,885|false|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Event|Event|SIMPLE_SEGMENT|891,897|false|false|false|||denies
Event|Event|SIMPLE_SEGMENT|913,920|false|false|false|||dysuria
Finding|Sign or Symptom|SIMPLE_SEGMENT|913,920|false|false|false|C0013428|Dysuria|dysuria
Drug|Food|SIMPLE_SEGMENT|930,934|false|false|false|C0016452;C3540798|Food;Food allergenic extracts|food
Drug|Immunologic Factor|SIMPLE_SEGMENT|930,934|false|false|false|C0016452;C3540798|Food;Food allergenic extracts|food
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|930,934|false|false|false|C0016452;C3540798|Food;Food allergenic extracts|food
Event|Event|SIMPLE_SEGMENT|930,934|false|false|false|||food
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|930,944|false|false|false|C0016479|Food Poisoning|food poisoning
Event|Event|SIMPLE_SEGMENT|935,944|false|false|false|||poisoning
Finding|Intellectual Product|SIMPLE_SEGMENT|947,951|false|false|false|C1561540|Transaction counts and value totals - week|week
Finding|Gene or Genome|SIMPLE_SEGMENT|952,955|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|968,973|false|false|false|C1838328|Lopes Gorlin syndrome|stale
Event|Event|SIMPLE_SEGMENT|968,973|false|false|false|||stale
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|975,979|false|false|false|C0452597;C0993597|Cake;Topical Cake|cake
Drug|Food|SIMPLE_SEGMENT|975,979|false|false|false|C0452597;C0993597|Cake;Topical Cake|cake
Event|Event|SIMPLE_SEGMENT|975,979|false|false|false|||cake
Drug|Food|SIMPLE_SEGMENT|998,1002|false|false|false|C0016452;C3540798|Food;Food allergenic extracts|food
Drug|Immunologic Factor|SIMPLE_SEGMENT|998,1002|false|false|false|C0016452;C3540798|Food;Food allergenic extracts|food
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|998,1002|false|false|false|C0016452;C3540798|Food;Food allergenic extracts|food
Event|Event|SIMPLE_SEGMENT|1003,1012|false|false|false|||ingestion
Phenomenon|Biologic Function|SIMPLE_SEGMENT|1003,1012|false|false|false|C0232478|Ingestion|ingestion
Event|Event|SIMPLE_SEGMENT|1021,1029|false|false|false|||resolved
Finding|Idea or Concept|SIMPLE_SEGMENT|1040,1043|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|1040,1043|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|1049,1055|false|false|false|||denies
Event|Event|SIMPLE_SEGMENT|1069,1076|false|false|false|||illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|1069,1076|false|false|false|C0221423|Illness (finding)|illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|1080,1084|false|false|false|C0221423|Illness (finding)|sick
Event|Event|SIMPLE_SEGMENT|1085,1093|false|false|false|||contacts
Procedure|Health Care Activity|SIMPLE_SEGMENT|1085,1093|false|false|false|C4036459|Contacts|contacts
Event|Event|SIMPLE_SEGMENT|1099,1104|false|false|false|||notes
Event|Event|SIMPLE_SEGMENT|1124,1132|false|false|false|||noticing
Anatomy|Tissue|SIMPLE_SEGMENT|1133,1136|false|false|false|C0017562|Gingiva|gum
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|1133,1136|false|false|false|C0812395;C1378701|Gum Dose Form;Gum as an ingredient|gum
Finding|Gene or Genome|SIMPLE_SEGMENT|1133,1136|false|false|false|C1825233;C5444202|OTULIN gene;OTULIN wt Allele|gum
Finding|Pathologic Function|SIMPLE_SEGMENT|1133,1145|false|false|false|C0017565|Gingival Hemorrhage|gum bleeding
Event|Event|SIMPLE_SEGMENT|1137,1145|false|false|false|||bleeding
Finding|Pathologic Function|SIMPLE_SEGMENT|1137,1145|false|false|false|C0019080|Hemorrhage|bleeding
Event|Event|SIMPLE_SEGMENT|1152,1160|false|false|false|||brushing
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1165,1170|false|false|false|C0040426;C4071855|Head>Teeth;Tooth structure|teeth
Procedure|Health Care Activity|SIMPLE_SEGMENT|1165,1170|false|false|false|C2239132|examination of teeth|teeth
Event|Event|SIMPLE_SEGMENT|1193,1199|false|false|false|||denies
Finding|Finding|SIMPLE_SEGMENT|1200,1204|false|false|false|C0332219|Easy|easy
Finding|Finding|SIMPLE_SEGMENT|1200,1213|true|false|false|C0423798|Increased tendency to bruise|easy bruising
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|1205,1213|true|false|false|C0009938|Contusions|bruising
Event|Event|SIMPLE_SEGMENT|1205,1213|false|false|false|||bruising
Finding|Finding|SIMPLE_SEGMENT|1205,1213|true|false|false|C2136686|reported bruising (history)|bruising
Event|Event|SIMPLE_SEGMENT|1215,1221|false|false|false|||melena
Finding|Pathologic Function|SIMPLE_SEGMENT|1215,1221|true|false|false|C0025222|Melena|melena
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1223,1228|true|false|false|C0018932|Hematochezia|BRBPR
Event|Event|SIMPLE_SEGMENT|1223,1228|false|false|false|||BRBPR
Event|Event|SIMPLE_SEGMENT|1231,1240|false|false|false|||hemetesis
Event|Event|SIMPLE_SEGMENT|1242,1252|false|false|false|||hemoptysis
Finding|Sign or Symptom|SIMPLE_SEGMENT|1242,1252|false|false|false|C0019079|Hemoptysis|hemoptysis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1257,1266|false|false|false|C0018965|Hematuria|hematuria
Event|Event|SIMPLE_SEGMENT|1257,1266|false|false|false|||hematuria
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1285,1288|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|abd
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|1285,1288|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|abd
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1289,1293|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|1289,1293|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|1289,1293|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1289,1293|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|1299,1303|false|false|false|||went
Event|Event|SIMPLE_SEGMENT|1322,1333|false|false|false|||transferred
Event|Activity|SIMPLE_SEGMENT|1354,1358|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|1354,1358|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|1354,1358|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|1354,1358|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1367,1373|false|false|false|C4255046||report
Event|Event|SIMPLE_SEGMENT|1367,1373|false|false|false|||report
Finding|Intellectual Product|SIMPLE_SEGMENT|1367,1373|false|false|false|C0684224|Report (document)|report
Procedure|Health Care Activity|SIMPLE_SEGMENT|1367,1373|false|false|false|C0700287|Reporting|report
Finding|Intellectual Product|SIMPLE_SEGMENT|1382,1387|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|brief
Event|Event|SIMPLE_SEGMENT|1388,1394|false|false|false|||period
Finding|Organism Function|SIMPLE_SEGMENT|1388,1394|false|false|false|C0025344|Menstruation|period
Procedure|Research Activity|SIMPLE_SEGMENT|1388,1394|false|false|false|C2347804|Clinical Trial Period|period
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|1399,1408|false|false|false|C0009676|Confusion|confusion
Event|Event|SIMPLE_SEGMENT|1399,1408|false|false|false|||confusion
Finding|Finding|SIMPLE_SEGMENT|1399,1408|false|false|false|C0683369|Clouded consciousness|confusion
Event|Event|SIMPLE_SEGMENT|1423,1429|false|false|false|||recall
Event|Event|SIMPLE_SEGMENT|1434,1444|false|false|false|||ultrasound
Finding|Functional Concept|SIMPLE_SEGMENT|1434,1444|true|true|false|C0220934|Ultrasonic|ultrasound
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|1434,1444|true|true|false|C0041621;C1456803|Ultrasonic Shockwave;Ultrasonics (sound)|ultrasound
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1434,1444|true|true|false|C0041618;C1315081|Ultrasonography;Urological ultrasound|ultrasound
Event|Event|SIMPLE_SEGMENT|1471,1477|false|false|false|||denies
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1485,1489|true|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|drug
Finding|Finding|SIMPLE_SEGMENT|1485,1489|true|false|false|C0740721|Drug problem|drug
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|1485,1493|true|false|false|C0242510|Drug usage|drug use
Finding|Finding|SIMPLE_SEGMENT|1485,1493|true|false|false|C0476643;C2239127|Drug use history;Encounter due to drug use|drug use
Event|Event|SIMPLE_SEGMENT|1490,1493|false|false|false|||use
Finding|Functional Concept|SIMPLE_SEGMENT|1490,1493|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|SIMPLE_SEGMENT|1490,1493|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Drug|Organic Chemical|SIMPLE_SEGMENT|1497,1504|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1497,1504|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Finding|Intellectual Product|SIMPLE_SEGMENT|1497,1504|false|false|false|C1547288|Alcohol - Recreational Drug Use Code|alcohol
Event|Event|SIMPLE_SEGMENT|1514,1520|false|false|false|||denies
Event|Event|SIMPLE_SEGMENT|1522,1529|false|false|false|||feeling
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|1530,1538|false|false|false|C0009676|Confusion|confused
Event|Event|SIMPLE_SEGMENT|1530,1538|false|false|false|||confused
Finding|Finding|SIMPLE_SEGMENT|1530,1538|false|false|false|C0683369;C1547301|Clouded consciousness;Precaution Code - Confused|confused
Finding|Intellectual Product|SIMPLE_SEGMENT|1530,1538|false|false|false|C0683369;C1547301|Clouded consciousness;Precaution Code - Confused|confused
Event|Event|SIMPLE_SEGMENT|1544,1551|false|false|false|||reports
Event|Event|SIMPLE_SEGMENT|1564,1573|false|false|false|||forgetful
Finding|Sign or Symptom|SIMPLE_SEGMENT|1564,1573|false|false|false|C0542476|Forgetful|forgetful
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1577,1582|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Event|Event|SIMPLE_SEGMENT|1577,1582|false|false|false|||times
Finding|Idea or Concept|SIMPLE_SEGMENT|1597,1604|false|false|false|C1555582|Initial (abbreviation)|initial
Event|Event|SIMPLE_SEGMENT|1605,1611|false|false|false|||vitals
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1643,1647|false|false|false|C0587081|Laboratory test finding|Labs
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1660,1663|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1660,1663|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|SIMPLE_SEGMENT|1660,1663|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|SIMPLE_SEGMENT|1660,1663|false|false|false|||ALT
Finding|Gene or Genome|SIMPLE_SEGMENT|1660,1663|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|SIMPLE_SEGMENT|1660,1663|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|SIMPLE_SEGMENT|1660,1663|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1660,1663|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|1664,1667|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1664,1667|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1664,1667|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1664,1667|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|SIMPLE_SEGMENT|1664,1667|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|SIMPLE_SEGMENT|1664,1667|false|false|false|||AST
Finding|Gene or Genome|SIMPLE_SEGMENT|1664,1667|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Event|Event|SIMPLE_SEGMENT|1686,1692|false|false|false|||Tbili1
Anatomy|Cell|SIMPLE_SEGMENT|1696,1699|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|1704,1712|false|false|false|C0005821|Blood Platelets|platelet
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1717,1720|false|false|false|C0368980|Coagulation tissue factor induced.INR|INR
Event|Event|SIMPLE_SEGMENT|1717,1720|false|false|false|||INR
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1717,1720|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1717,1720|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Finding|Finding|SIMPLE_SEGMENT|1730,1750|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Event|Event|SIMPLE_SEGMENT|1735,1742|false|false|false|||Medical
Finding|Functional Concept|SIMPLE_SEGMENT|1735,1742|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|1735,1742|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|1735,1742|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|1735,1742|false|false|false|C0199168|Medical service|Medical
Finding|Finding|SIMPLE_SEGMENT|1735,1750|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1743,1750|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1743,1750|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|1743,1750|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1755,1758|false|false|false|C0019196;C0220847|Hepatitis C;hepatitis C virus|HCV
Disorder|Virus|SIMPLE_SEGMENT|1755,1758|false|false|false|C0019196;C0220847|Hepatitis C;hepatitis C virus|HCV
Event|Event|SIMPLE_SEGMENT|1755,1758|false|false|false|||HCV
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1759,1768|false|false|false|C0023890;C1623038|Cirrhosis;Liver Cirrhosis|Cirrhosis
Event|Event|SIMPLE_SEGMENT|1759,1768|false|false|false|||Cirrhosis
Event|Event|SIMPLE_SEGMENT|1777,1784|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|1777,1784|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|1777,1784|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|1777,1784|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|1777,1787|true|false|false|C0262926|Medical History|history of
Finding|Finding|SIMPLE_SEGMENT|1788,1796|true|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Finding|Idea or Concept|SIMPLE_SEGMENT|1788,1796|true|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Finding|Finding|SIMPLE_SEGMENT|1788,1807|true|false|false|C0476427|Abnormal cervical smear|abnormal Pap smears
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1797,1800|false|false|false|C3496568|pars anterior of the paramedian lobule|Pap
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1797,1800|true|false|false|C0760170;C1740167|ACPP protein, human;alpha 2-plasmin inhibitor-plasmin complex|Pap
Drug|Enzyme|SIMPLE_SEGMENT|1797,1800|true|false|false|C0760170;C1740167|ACPP protein, human;alpha 2-plasmin inhibitor-plasmin complex|Pap
Drug|Immunologic Factor|SIMPLE_SEGMENT|1797,1800|true|false|false|C0760170;C1740167|ACPP protein, human;alpha 2-plasmin inhibitor-plasmin complex|Pap
Finding|Finding|SIMPLE_SEGMENT|1797,1800|true|false|false|C0428642;C1367456;C1413944;C1413945;C1418410;C1422804;C1423108;C1424700;C1538823;C1705529;C1705530;C1705531;C1863340;C2266415;C3538851;C3889402|ACP3 gene;ACP3 wt Allele;ASAP1 gene;ASAP1 wt Allele;ASAP2 gene;MRPS30 gene;PAPOLA gene;PAPOLA wt Allele;PDAP1 gene;PITUITARY ADENOMA PREDISPOSITION;Pulmonary artery pressure;REG3A gene;REG3A wt Allele;TUSC2 gene;TUSC2 wt Allele|Pap
Finding|Gene or Genome|SIMPLE_SEGMENT|1797,1800|true|false|false|C0428642;C1367456;C1413944;C1413945;C1418410;C1422804;C1423108;C1424700;C1538823;C1705529;C1705530;C1705531;C1863340;C2266415;C3538851;C3889402|ACP3 gene;ACP3 wt Allele;ASAP1 gene;ASAP1 wt Allele;ASAP2 gene;MRPS30 gene;PAPOLA gene;PAPOLA wt Allele;PDAP1 gene;PITUITARY ADENOMA PREDISPOSITION;Pulmonary artery pressure;REG3A gene;REG3A wt Allele;TUSC2 gene;TUSC2 wt Allele|Pap
Finding|Molecular Function|SIMPLE_SEGMENT|1797,1800|true|false|false|C0428642;C1367456;C1413944;C1413945;C1418410;C1422804;C1423108;C1424700;C1538823;C1705529;C1705530;C1705531;C1863340;C2266415;C3538851;C3889402|ACP3 gene;ACP3 wt Allele;ASAP1 gene;ASAP1 wt Allele;ASAP2 gene;MRPS30 gene;PAPOLA gene;PAPOLA wt Allele;PDAP1 gene;PITUITARY ADENOMA PREDISPOSITION;Pulmonary artery pressure;REG3A gene;REG3A wt Allele;TUSC2 gene;TUSC2 wt Allele|Pap
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1797,1807|true|false|false|C0079104|Pap smear|Pap smears
Event|Event|SIMPLE_SEGMENT|1801,1807|false|false|false|||smears
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1801,1807|true|false|false|C0444186|Smear test|smears
Event|Event|SIMPLE_SEGMENT|1822,1835|false|false|false|||calcification
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|1822,1835|false|false|false|C0006660;C0006663;C1533591|Calcification;Calcinosis;Physiologic calcification|calcification
Finding|Pathologic Function|SIMPLE_SEGMENT|1822,1835|false|false|false|C0006660;C0006663;C1533591|Calcification;Calcinosis;Physiologic calcification|calcification
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1843,1849|false|false|false|C0006141|Breast|breast
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1843,1849|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|breast
Event|Event|SIMPLE_SEGMENT|1843,1849|false|false|false|||breast
Finding|Finding|SIMPLE_SEGMENT|1843,1849|false|false|false|C0567499|Breast problem|breast
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1843,1849|false|false|false|C0191838|Procedures on breast|breast
Event|Event|SIMPLE_SEGMENT|1861,1868|false|false|false|||removed
Finding|Body Substance|SIMPLE_SEGMENT|1890,1897|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1890,1897|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1890,1897|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|1910,1916|false|false|false|||benign
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1927,1930|false|false|false|C0019682;C0019693|HIV;HIV Infections|HIV
Disorder|Virus|SIMPLE_SEGMENT|1927,1930|false|false|false|C0019682;C0019693|HIV;HIV Infections|HIV
Drug|Immunologic Factor|SIMPLE_SEGMENT|1927,1930|false|false|false|C0086413|HIV Vaccine|HIV
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1927,1930|false|false|false|C0086413|HIV Vaccine|HIV
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1927,1938|false|false|false|C0019693|HIV Infections|HIV disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1931,1938|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|1931,1938|false|false|false|||disease
Event|Event|SIMPLE_SEGMENT|1953,1961|false|false|false|||followed
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1989,1993|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1989,1993|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|SIMPLE_SEGMENT|1989,1993|false|false|false|||COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|1989,1993|false|false|false|C1412502|ARCN1 gene|COPD
Finding|Finding|SIMPLE_SEGMENT|1999,2011|false|false|false|C0332119|Past history of|Past history
Finding|Finding|SIMPLE_SEGMENT|1999,2014|false|false|false|C0332119|Past history of|Past history of
Event|Event|SIMPLE_SEGMENT|2004,2011|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|2004,2011|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|2004,2011|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|2004,2011|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|2004,2014|false|false|false|C0262926|Medical History|history of
Event|Event|SIMPLE_SEGMENT|2015,2022|false|false|false|||smoking
Finding|Individual Behavior|SIMPLE_SEGMENT|2015,2022|false|false|false|C0037369;C0453996;C1548578|Location characteristic ID - Smoking;Smoking;Tobacco smoking behavior|smoking
Finding|Intellectual Product|SIMPLE_SEGMENT|2015,2022|false|false|false|C0037369;C0453996;C1548578|Location characteristic ID - Smoking;Smoking;Tobacco smoking behavior|smoking
Anatomy|Body System|SIMPLE_SEGMENT|2044,2048|false|false|false|C1123023;C4520765|Skin;Skin, Human|skin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2044,2048|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2044,2048|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Finding|Body Substance|SIMPLE_SEGMENT|2044,2048|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Finding|Intellectual Product|SIMPLE_SEGMENT|2044,2048|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2044,2055|false|false|false|C0037284|Skin lesion|skin lesion
Event|Event|SIMPLE_SEGMENT|2049,2055|false|false|false|||lesion
Finding|Finding|SIMPLE_SEGMENT|2049,2055|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|SIMPLE_SEGMENT|2049,2055|false|false|false|C0221198;C1546698|Lesion|lesion
Event|Event|SIMPLE_SEGMENT|2067,2075|false|false|false|||biopsied
Event|Event|SIMPLE_SEGMENT|2080,2086|false|false|false|||showed
Anatomy|Body System|SIMPLE_SEGMENT|2089,2093|false|false|false|C1123023;C4520765|Skin;Skin, Human|skin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2089,2093|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2089,2093|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Finding|Body Substance|SIMPLE_SEGMENT|2089,2093|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Finding|Intellectual Product|SIMPLE_SEGMENT|2089,2093|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2089,2100|false|false|false|C0007114|Malignant neoplasm of skin|skin cancer
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2094,2100|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|SIMPLE_SEGMENT|2094,2100|false|false|false|||cancer
Finding|Body Substance|SIMPLE_SEGMENT|2105,2112|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|2105,2112|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|2105,2112|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|2105,2119|false|false|false|C0747307|Patient-Reported|patient report
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2113,2119|false|false|false|C4255046||report
Event|Event|SIMPLE_SEGMENT|2113,2119|false|false|false|||report
Finding|Intellectual Product|SIMPLE_SEGMENT|2113,2119|false|false|false|C0684224|Report (document)|report
Procedure|Health Care Activity|SIMPLE_SEGMENT|2113,2119|false|false|false|C0700287|Reporting|report
Event|Event|SIMPLE_SEGMENT|2127,2136|false|false|false|||scheduled
Drug|Organic Chemical|SIMPLE_SEGMENT|2143,2151|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2143,2151|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|SIMPLE_SEGMENT|2143,2151|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|SIMPLE_SEGMENT|2143,2151|false|false|false|||complete
Finding|Functional Concept|SIMPLE_SEGMENT|2143,2151|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|SIMPLE_SEGMENT|2143,2151|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Event|Activity|SIMPLE_SEGMENT|2154,2161|false|false|false|C1883720|Removing (action)|removal
Event|Event|SIMPLE_SEGMENT|2154,2161|false|false|false|||removal
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2154,2161|false|false|false|C0015252;C0185115;C0728940|Excision;Extraction;removal technique|removal
Anatomy|Body System|SIMPLE_SEGMENT|2169,2173|false|false|false|C1123023;C4520765|Skin;Skin, Human|skin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2169,2173|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2169,2173|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Finding|Body Substance|SIMPLE_SEGMENT|2169,2173|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Finding|Intellectual Product|SIMPLE_SEGMENT|2169,2173|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2169,2180|false|false|false|C0037284|Skin lesion|skin lesion
Event|Event|SIMPLE_SEGMENT|2174,2180|false|false|false|||lesion
Finding|Finding|SIMPLE_SEGMENT|2174,2180|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|SIMPLE_SEGMENT|2174,2180|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Idea or Concept|SIMPLE_SEGMENT|2196,2200|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|SIMPLE_SEGMENT|2196,2200|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Event|Event|SIMPLE_SEGMENT|2228,2234|false|false|false|||lesion
Finding|Finding|SIMPLE_SEGMENT|2228,2234|false|true|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|SIMPLE_SEGMENT|2228,2234|false|true|false|C0221198;C1546698|Lesion|lesion
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2242,2250|false|false|false|C0016540|Forehead|forehead
Event|Event|SIMPLE_SEGMENT|2265,2278|false|false|false|||discoloration
Finding|Finding|SIMPLE_SEGMENT|2265,2278|false|false|false|C0332572|Abnormal color|discoloration
Event|Event|SIMPLE_SEGMENT|2287,2295|false|false|false|||biopsied
Event|Event|SIMPLE_SEGMENT|2299,2306|false|false|false|||exclude
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2334,2341|false|false|false|C1261473;C4551686|Malignant neoplasm of soft tissue;Sarcoma|sarcoma
Event|Event|SIMPLE_SEGMENT|2334,2341|false|false|false|||sarcoma
Event|Event|SIMPLE_SEGMENT|2347,2354|false|false|false|||results
Event|Event|SIMPLE_SEGMENT|2358,2365|false|false|false|||pending
Finding|Idea or Concept|SIMPLE_SEGMENT|2358,2365|false|false|false|C1691786;C1704475|Pending - Allergy Clinical Status;Pending - referral status|pending
Finding|Finding|SIMPLE_SEGMENT|2380,2390|false|false|false|C5961011|Hypoechoic|hypoechoic
Event|Event|SIMPLE_SEGMENT|2391,2397|false|false|false|||lesion
Finding|Finding|SIMPLE_SEGMENT|2391,2397|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|SIMPLE_SEGMENT|2391,2397|false|false|false|C0221198;C1546698|Lesion|lesion
Event|Event|SIMPLE_SEGMENT|2405,2415|false|false|false|||ultrasound
Finding|Functional Concept|SIMPLE_SEGMENT|2405,2415|false|false|false|C0220934|Ultrasonic|ultrasound
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|2405,2415|false|false|false|C0041621;C1456803|Ultrasonic Shockwave;Ultrasonics (sound)|ultrasound
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2405,2415|false|false|false|C0041618;C1315081|Ultrasonography;Urological ultrasound|ultrasound
Event|Event|SIMPLE_SEGMENT|2438,2447|false|false|false|||monitored
Event|Event|SIMPLE_SEGMENT|2454,2457|false|false|false|||MRI
Finding|Gene or Genome|SIMPLE_SEGMENT|2454,2457|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2454,2457|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|SIMPLE_SEGMENT|2454,2457|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Event|Event|SIMPLE_SEGMENT|2465,2472|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2465,2472|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2465,2472|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2465,2472|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2465,2475|false|false|false|C0262926|Medical History|History of
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|2476,2485|false|false|false|C0334044|Dysplasia|dysplasia
Event|Event|SIMPLE_SEGMENT|2476,2485|false|false|false|||dysplasia
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2476,2493|false|false|false|C0347129|Dysplasia of anus|dysplasia of anus
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2489,2493|false|false|false|C0003461|Anus|anus
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2489,2493|false|false|false|C0003462|Anus Diseases|anus
Event|Event|SIMPLE_SEGMENT|2489,2493|false|false|false|||anus
Procedure|Health Care Activity|SIMPLE_SEGMENT|2489,2493|false|false|false|C0870072|Procedure on anus|anus
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|2508,2534|false|false|false|C0005586;C1839839;C1852197;C1970943;C1970945;C2700438;C2700439;C2700440|Bipolar Disorder;MAJOR AFFECTIVE DISORDER 1;MAJOR AFFECTIVE DISORDER 2;MAJOR AFFECTIVE DISORDER 4;MAJOR AFFECTIVE DISORDER 6;MAJOR AFFECTIVE DISORDER 7;MAJOR AFFECTIVE DISORDER 8;MAJOR AFFECTIVE DISORDER 9|Bipolar affective disorder
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|2508,2557|false|false|false|C0338875|Bipolar affective disorder, currently manic, mild|Bipolar affective disorder, currently manic, mild
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|2516,2534|false|false|false|C0525045|Mood Disorders|affective disorder
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2526,2534|false|false|false|C0012634|Disease|disorder
Event|Event|SIMPLE_SEGMENT|2526,2534|false|false|false|||disorder
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|2546,2551|false|false|false|C0338831|Manic|manic
Event|Event|SIMPLE_SEGMENT|2546,2551|false|false|false|||manic
Finding|Finding|SIMPLE_SEGMENT|2546,2551|false|false|false|C0564408|Manic mood|manic
Event|Event|SIMPLE_SEGMENT|2553,2557|false|false|false|||mild
Finding|Intellectual Product|SIMPLE_SEGMENT|2553,2557|false|false|false|C1547225|Mild Severity of Illness Code|mild
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2563,2567|false|false|false|C0038436;C0878676|6-pyruvoyl-tetrahydropterin synthase deficiency;Post-Traumatic Stress Disorder|PTSD
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|2563,2567|false|false|false|C0038436;C0878676|6-pyruvoyl-tetrahydropterin synthase deficiency;Post-Traumatic Stress Disorder|PTSD
Event|Event|SIMPLE_SEGMENT|2563,2567|false|false|false|||PTSD
Event|Event|SIMPLE_SEGMENT|2576,2583|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2576,2583|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2576,2583|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2576,2583|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2576,2586|false|false|false|C0262926|Medical History|History of
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|2587,2594|true|false|false|C0274659|Poisoning by cocaine|cocaine
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|2587,2594|true|false|false|C0009170|cocaine|cocaine
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|2587,2594|true|false|false|C0009170|cocaine|cocaine
Drug|Organic Chemical|SIMPLE_SEGMENT|2587,2594|true|false|false|C0009170|cocaine|cocaine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2587,2594|true|false|false|C0009170|cocaine|cocaine
Event|Event|SIMPLE_SEGMENT|2587,2594|false|false|false|||cocaine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2587,2594|true|false|false|C0202362|Cocaine measurement|cocaine
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|2599,2605|true|false|false|C0161541|Poisoning by heroin|heroin
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|2599,2605|true|false|false|C0011892|heroin|heroin
Drug|Organic Chemical|SIMPLE_SEGMENT|2599,2605|true|false|false|C0011892|heroin|heroin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2599,2605|true|false|false|C0011892|heroin|heroin
Event|Event|SIMPLE_SEGMENT|2599,2605|false|false|false|||heroin
Event|Event|SIMPLE_SEGMENT|2606,2609|false|false|false|||use
Finding|Functional Concept|SIMPLE_SEGMENT|2606,2609|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|SIMPLE_SEGMENT|2606,2609|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Functional Concept|SIMPLE_SEGMENT|2616,2622|false|false|false|C0728831|Social|Social
Finding|Finding|SIMPLE_SEGMENT|2616,2630|false|false|false|C0424945;C3714536|Social History;Social and personal history|Social History
Event|Event|SIMPLE_SEGMENT|2623,2630|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2623,2630|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2623,2630|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2623,2630|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Classification|SIMPLE_SEGMENT|2636,2642|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|SIMPLE_SEGMENT|2636,2642|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|SIMPLE_SEGMENT|2636,2642|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|SIMPLE_SEGMENT|2636,2642|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Finding|SIMPLE_SEGMENT|2636,2650|false|false|false|C0241889|Family Medical History|Family History
Event|Event|SIMPLE_SEGMENT|2643,2650|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2643,2650|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2643,2650|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2643,2650|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Event|Event|SIMPLE_SEGMENT|2699,2706|false|false|false|||talking
Finding|Conceptual Entity|SIMPLE_SEGMENT|2741,2748|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|brother
Finding|Idea or Concept|SIMPLE_SEGMENT|2741,2748|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|brother
Event|Event|SIMPLE_SEGMENT|2767,2772|false|false|false|||touch
Finding|Mental Process|SIMPLE_SEGMENT|2767,2772|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|2767,2772|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2767,2772|false|false|false|C0152054|Therapeutic Touch|touch
Event|Event|SIMPLE_SEGMENT|2782,2787|false|false|false|||lives
Event|Event|SIMPLE_SEGMENT|2807,2812|false|false|false|||aware
Finding|Mental Process|SIMPLE_SEGMENT|2807,2812|true|false|false|C0004448|Awareness|aware
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2834,2839|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2834,2839|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2834,2839|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|SIMPLE_SEGMENT|2834,2839|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2834,2839|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|SIMPLE_SEGMENT|2834,2839|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|SIMPLE_SEGMENT|2834,2839|false|false|false|||liver
Finding|Finding|SIMPLE_SEGMENT|2834,2839|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|SIMPLE_SEGMENT|2834,2839|false|false|false|C0872387|Procedures on liver|liver
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2834,2847|false|true|false|C0023895;C0267792|Hepatobiliary Disorder;Liver diseases|liver disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2840,2847|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|2840,2847|false|false|false|||disease
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2851,2861|false|false|false|C3812393|ErbB Receptors|her family
Drug|Enzyme|SIMPLE_SEGMENT|2851,2861|false|false|false|C3812393|ErbB Receptors|her family
Finding|Receptor|SIMPLE_SEGMENT|2851,2861|false|false|false|C3812393|ErbB Receptors|her family
Finding|Classification|SIMPLE_SEGMENT|2855,2861|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|2855,2861|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|2855,2861|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|2855,2861|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Drug|Organic Chemical|SIMPLE_SEGMENT|2874,2881|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2874,2881|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Finding|Intellectual Product|SIMPLE_SEGMENT|2874,2881|false|false|false|C1547288|Alcohol - Recreational Drug Use Code|alcohol
Finding|Finding|SIMPLE_SEGMENT|2874,2893|false|false|false|C0001948;C2215684|Alcohol consumption;alcohol consumption (history)|alcohol consumption
Finding|Individual Behavior|SIMPLE_SEGMENT|2874,2893|false|false|false|C0001948;C2215684|Alcohol consumption;alcohol consumption (history)|alcohol consumption
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2882,2893|false|false|false|C0220811|Consumption-archaic term for TB|consumption
Event|Activity|SIMPLE_SEGMENT|2882,2893|false|false|false|C0009830|Consumption of goods|consumption
Event|Event|SIMPLE_SEGMENT|2882,2893|false|false|false|||consumption
Finding|Physiologic Function|SIMPLE_SEGMENT|2882,2893|false|false|false|C1947907|biologic consumption|consumption
Drug|Food|SIMPLE_SEGMENT|2902,2907|false|false|false|C0452428|Drink (dietary substance)|drink
Event|Event|SIMPLE_SEGMENT|2902,2907|false|false|false|||drink
Finding|Gene or Genome|SIMPLE_SEGMENT|2919,2922|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Drug|Organic Chemical|SIMPLE_SEGMENT|2937,2944|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2937,2944|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Finding|Intellectual Product|SIMPLE_SEGMENT|2937,2944|false|false|false|C1547288|Alcohol - Recreational Drug Use Code|alcohol
Finding|Finding|SIMPLE_SEGMENT|2937,2956|false|false|false|C0001948;C2215684|Alcohol consumption;alcohol consumption (history)|alcohol consumption
Finding|Individual Behavior|SIMPLE_SEGMENT|2937,2956|false|false|false|C0001948;C2215684|Alcohol consumption;alcohol consumption (history)|alcohol consumption
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2945,2956|false|false|false|C0220811|Consumption-archaic term for TB|consumption
Event|Activity|SIMPLE_SEGMENT|2945,2956|false|false|false|C0009830|Consumption of goods|consumption
Event|Event|SIMPLE_SEGMENT|2945,2956|false|false|false|||consumption
Finding|Physiologic Function|SIMPLE_SEGMENT|2945,2956|false|false|false|C1947907|biologic consumption|consumption
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2963,2967|false|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|drug
Finding|Finding|SIMPLE_SEGMENT|2963,2967|false|false|false|C0740721|Drug problem|drug
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|2963,2971|false|false|false|C0242510|Drug usage|drug use
Finding|Finding|SIMPLE_SEGMENT|2963,2971|false|false|false|C0476643;C2239127|Drug use history;Encounter due to drug use|drug use
Event|Event|SIMPLE_SEGMENT|2968,2971|false|false|false|||use
Finding|Functional Concept|SIMPLE_SEGMENT|2968,2971|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|SIMPLE_SEGMENT|2968,2971|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Gene or Genome|SIMPLE_SEGMENT|2982,2985|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Event|Event|SIMPLE_SEGMENT|2993,2997|false|false|false|||quit
Event|Event|SIMPLE_SEGMENT|2998,3005|false|false|false|||smoking
Event|Event|SIMPLE_SEGMENT|3008,3014|false|false|false|||couple
Finding|Functional Concept|SIMPLE_SEGMENT|3008,3014|false|false|false|C1948027|Couple (action)|couple
Finding|Gene or Genome|SIMPLE_SEGMENT|3024,3027|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Event|Event|SIMPLE_SEGMENT|3034,3042|false|false|false|||Physical
Finding|Finding|SIMPLE_SEGMENT|3034,3042|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|3034,3042|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|3034,3042|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|3034,3047|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|3034,3047|false|false|false|C0031809|Physical Examination|Physical Exam
Event|Event|SIMPLE_SEGMENT|3043,3047|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|3043,3047|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|3043,3047|false|false|false|C0582103|Medical Examination|Exam
Event|Event|SIMPLE_SEGMENT|3078,3085|false|false|false|||General
Finding|Classification|SIMPLE_SEGMENT|3078,3085|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|SIMPLE_SEGMENT|3078,3085|false|false|false|C3812897|General medical service|General
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3090,3093|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3090,3093|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3090,3093|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|3090,3093|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3090,3093|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|SIMPLE_SEGMENT|3090,3093|false|false|false|||NAD
Finding|Finding|SIMPLE_SEGMENT|3090,3093|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3096,3101|false|false|false|C1512338|HEENT|HEENT
Drug|Organic Chemical|SIMPLE_SEGMENT|3103,3107|false|false|false|C0951233|cetrimonium bromide|CTAB
Event|Event|SIMPLE_SEGMENT|3103,3107|false|false|false|||CTAB
Finding|Finding|SIMPLE_SEGMENT|3109,3118|false|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3119,3125|false|false|false|C0036410|Sclera|sclera
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3119,3125|false|false|false|C0036412|Scleral Diseases|sclera
Event|Event|SIMPLE_SEGMENT|3119,3125|false|false|false|||sclera
Procedure|Health Care Activity|SIMPLE_SEGMENT|3119,3125|false|false|false|C2228481|examination of sclera|sclera
Event|Event|SIMPLE_SEGMENT|3130,3135|false|false|false|||clear
Finding|Idea or Concept|SIMPLE_SEGMENT|3130,3135|false|false|false|C1550016|Remote control command - Clear|clear
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3138,3142|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Anatomy|Cell Component|SIMPLE_SEGMENT|3138,3142|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Finding|Finding|SIMPLE_SEGMENT|3138,3142|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|Neck
Event|Event|SIMPLE_SEGMENT|3144,3150|false|false|false|||supple
Finding|Functional Concept|SIMPLE_SEGMENT|3144,3150|false|false|false|C0332254|Supple|supple
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3155,3158|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3155,3158|true|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|SIMPLE_SEGMENT|3155,3158|false|false|false|||LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|3155,3158|true|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Event|Event|SIMPLE_SEGMENT|3165,3168|false|false|false|||RRR
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3186,3191|false|false|false|C0024109|Lung|Lungs
Drug|Organic Chemical|SIMPLE_SEGMENT|3193,3197|false|false|false|C0951233|cetrimonium bromide|CTAb
Event|Event|SIMPLE_SEGMENT|3193,3197|false|false|false|||CTAb
Finding|Organism Function|SIMPLE_SEGMENT|3209,3219|false|false|false|C0231800|Expiration, Respiratory|expiratory
Event|Event|SIMPLE_SEGMENT|3220,3225|false|false|false|||phase
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3238,3245|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3238,3245|false|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Event|Event|SIMPLE_SEGMENT|3238,3245|false|false|false|||Abdomen
Finding|Finding|SIMPLE_SEGMENT|3238,3245|false|false|false|C0941288|Abdomen problem|Abdomen
Event|Event|SIMPLE_SEGMENT|3247,3256|false|false|false|||distended
Finding|Finding|SIMPLE_SEGMENT|3247,3256|false|false|false|C0700124|Dilated|distended
Finding|Intellectual Product|SIMPLE_SEGMENT|3258,3262|false|false|false|C1547225|Mild Severity of Illness Code|mild
Event|Event|SIMPLE_SEGMENT|3271,3281|false|false|false|||tenderness
Finding|Mental Process|SIMPLE_SEGMENT|3271,3281|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|SIMPLE_SEGMENT|3271,3281|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3284,3289|false|false|false|C0230171|Flank (surface region)|flank
Event|Event|SIMPLE_SEGMENT|3290,3298|false|false|false|||dullness
Finding|Finding|SIMPLE_SEGMENT|3290,3298|false|false|false|C0541911|Dullness|dullness
Event|Event|SIMPLE_SEGMENT|3308,3315|false|false|false|||percuss
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3316,3321|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3316,3321|false|true|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3316,3321|false|true|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|SIMPLE_SEGMENT|3316,3321|false|true|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3316,3321|false|true|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|SIMPLE_SEGMENT|3316,3321|false|true|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|SIMPLE_SEGMENT|3316,3321|false|false|false|||liver
Finding|Finding|SIMPLE_SEGMENT|3316,3321|false|true|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|SIMPLE_SEGMENT|3316,3321|false|true|false|C0872387|Procedures on liver|liver
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3322,3328|false|false|false|C0037993;C4037984|Abdomen>Spleen;Spleen|spleen
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3322,3328|false|false|false|C0153470|Malignant neoplasm of spleen|spleen
Finding|Finding|SIMPLE_SEGMENT|3322,3328|false|false|false|C0812414|Spleen problem|spleen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3322,3328|false|false|false|C0869677|Procedures on Spleen|spleen
Event|Event|SIMPLE_SEGMENT|3329,3333|false|false|false|||edge
Finding|Conceptual Entity|SIMPLE_SEGMENT|3329,3333|false|false|false|C2697523|Graph Edge|edge
Event|Event|SIMPLE_SEGMENT|3338,3348|false|false|false|||distension
Finding|Finding|SIMPLE_SEGMENT|3338,3348|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distension
Finding|Pathologic Function|SIMPLE_SEGMENT|3338,3348|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distension
Event|Event|SIMPLE_SEGMENT|3358,3363|false|false|false|||foley
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|3366,3369|false|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Event|Event|SIMPLE_SEGMENT|3366,3369|false|false|false|||Ext
Finding|Gene or Genome|SIMPLE_SEGMENT|3366,3369|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|3388,3396|false|false|false|C0149651|Clubbing|clubbing
Event|Event|SIMPLE_SEGMENT|3388,3396|false|false|false|||clubbing
Finding|Molecular Function|SIMPLE_SEGMENT|3406,3410|false|false|false|C1817552|abscisic aldehyde oxidase activity|AAO3
Event|Event|SIMPLE_SEGMENT|3431,3435|false|false|false|||able
Finding|Finding|SIMPLE_SEGMENT|3431,3435|false|false|false|C1299581|Able (qualifier value)|able
Event|Event|SIMPLE_SEGMENT|3439,3445|false|false|false|||recall
Event|Governmental or Regulatory Activity|SIMPLE_SEGMENT|3439,3445|false|false|false|C1705180|Recall (activity)|recall
Finding|Mental Process|SIMPLE_SEGMENT|3439,3445|false|false|false|C0034770|Mental Recall|recall
Finding|Finding|SIMPLE_SEGMENT|3446,3453|false|false|false|C4035626|3 times|3 times
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3448,3453|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Event|Event|SIMPLE_SEGMENT|3448,3453|false|false|false|||times
Event|Event|SIMPLE_SEGMENT|3482,3488|false|false|false|||intact
Finding|Finding|SIMPLE_SEGMENT|3482,3488|false|false|false|C1554187|Gender Status - Intact|intact
Event|Event|SIMPLE_SEGMENT|3492,3501|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|3492,3501|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|3492,3501|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|3492,3501|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|3492,3501|false|false|false|C0030685|Patient Discharge|Discharge
Event|Event|SIMPLE_SEGMENT|3504,3512|false|false|false|||PHYSICAL
Finding|Finding|SIMPLE_SEGMENT|3504,3512|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|SIMPLE_SEGMENT|3504,3512|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|3504,3512|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|SIMPLE_SEGMENT|3504,3524|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAMINATION
Procedure|Health Care Activity|SIMPLE_SEGMENT|3504,3524|false|false|false|C0031809|Physical Examination|PHYSICAL EXAMINATION
Event|Activity|SIMPLE_SEGMENT|3513,3524|false|false|false|C4321457|Examination|EXAMINATION
Event|Event|SIMPLE_SEGMENT|3513,3524|false|false|false|||EXAMINATION
Procedure|Health Care Activity|SIMPLE_SEGMENT|3513,3524|false|false|false|C0031809;C0582103|Medical Examination;Physical Examination|EXAMINATION
Event|Event|SIMPLE_SEGMENT|3545,3552|false|false|false|||General
Finding|Classification|SIMPLE_SEGMENT|3545,3552|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|SIMPLE_SEGMENT|3545,3552|false|false|false|C3812897|General medical service|General
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3557,3560|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3557,3560|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3557,3560|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|3557,3560|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3557,3560|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|SIMPLE_SEGMENT|3557,3560|false|false|false|||NAD
Finding|Finding|SIMPLE_SEGMENT|3557,3560|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3563,3568|false|false|false|C1512338|HEENT|HEENT
Finding|Finding|SIMPLE_SEGMENT|3570,3579|false|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3580,3586|false|false|false|C0036410|Sclera|sclera
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3580,3586|false|false|false|C0036412|Scleral Diseases|sclera
Event|Event|SIMPLE_SEGMENT|3580,3586|false|false|false|||sclera
Procedure|Health Care Activity|SIMPLE_SEGMENT|3580,3586|false|false|false|C2228481|examination of sclera|sclera
Event|Event|SIMPLE_SEGMENT|3591,3596|false|false|false|||clear
Finding|Idea or Concept|SIMPLE_SEGMENT|3591,3596|false|false|false|C1550016|Remote control command - Clear|clear
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3599,3603|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Anatomy|Cell Component|SIMPLE_SEGMENT|3599,3603|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Finding|Finding|SIMPLE_SEGMENT|3599,3603|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|Neck
Event|Event|SIMPLE_SEGMENT|3605,3611|false|false|false|||supple
Finding|Functional Concept|SIMPLE_SEGMENT|3605,3611|false|false|false|C0332254|Supple|supple
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3616,3619|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3616,3619|true|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|SIMPLE_SEGMENT|3616,3619|false|false|false|||LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|3616,3619|true|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Event|Event|SIMPLE_SEGMENT|3626,3629|false|false|false|||RRR
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3647,3652|false|false|false|C0024109|Lung|Lungs
Drug|Organic Chemical|SIMPLE_SEGMENT|3654,3658|false|false|false|C0951233|cetrimonium bromide|CTAb
Event|Event|SIMPLE_SEGMENT|3654,3658|false|false|false|||CTAb
Finding|Organism Function|SIMPLE_SEGMENT|3670,3680|false|false|false|C0231800|Expiration, Respiratory|expiratory
Event|Event|SIMPLE_SEGMENT|3681,3686|false|false|false|||phase
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3699,3706|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3699,3706|false|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Event|Event|SIMPLE_SEGMENT|3699,3706|false|false|false|||Abdomen
Finding|Finding|SIMPLE_SEGMENT|3699,3706|false|false|false|C0941288|Abdomen problem|Abdomen
Event|Event|SIMPLE_SEGMENT|3708,3717|false|false|false|||distended
Finding|Finding|SIMPLE_SEGMENT|3708,3717|false|false|false|C0700124|Dilated|distended
Event|Event|SIMPLE_SEGMENT|3722,3730|false|false|false|||improved
Finding|Finding|SIMPLE_SEGMENT|3722,3730|false|false|false|C0184511;C1561611;C4084203|Admission Level of Care Code - Improved;Improved;Improved - answer to question|improved
Finding|Intellectual Product|SIMPLE_SEGMENT|3722,3730|false|false|false|C0184511;C1561611;C4084203|Admission Level of Care Code - Improved;Improved;Improved - answer to question|improved
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3732,3735|false|false|false|C0034155;C1268935|Congenital Thrombotic Thrombocytopenic Purpura;Purpura, Thrombotic Thrombocytopenic|TTP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3732,3735|false|false|false|C1506603;C4723973|ZFP36 protein, human;thiamine triphosphorate|TTP
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3732,3735|false|false|false|C1506603;C4723973|ZFP36 protein, human;thiamine triphosphorate|TTP
Drug|Organic Chemical|SIMPLE_SEGMENT|3732,3735|false|false|false|C1506603;C4723973|ZFP36 protein, human;thiamine triphosphorate|TTP
Drug|Vitamin|SIMPLE_SEGMENT|3732,3735|false|false|false|C1506603;C4723973|ZFP36 protein, human;thiamine triphosphorate|TTP
Event|Event|SIMPLE_SEGMENT|3732,3735|false|false|false|||TTP
Finding|Gene or Genome|SIMPLE_SEGMENT|3732,3735|false|false|false|C1413036;C1421571;C3539814|ADAMTS13 gene;ZFP36 gene;ZFP36 wt Allele|TTP
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3739,3742|false|false|false|C0230177|Structure of right upper quadrant of abdomen|RUQ
Event|Event|SIMPLE_SEGMENT|3752,3757|false|false|false|||foley
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|3760,3763|false|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Event|Event|SIMPLE_SEGMENT|3760,3763|false|false|false|||Ext
Finding|Gene or Genome|SIMPLE_SEGMENT|3760,3763|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|3782,3790|false|false|false|C0149651|Clubbing|clubbing
Event|Event|SIMPLE_SEGMENT|3782,3790|false|false|false|||clubbing
Finding|Molecular Function|SIMPLE_SEGMENT|3800,3804|false|false|false|C1817552|abscisic aldehyde oxidase activity|AAO3
Event|Event|SIMPLE_SEGMENT|3817,3823|false|false|false|||intact
Finding|Finding|SIMPLE_SEGMENT|3817,3823|false|false|false|C1554187|Gender Status - Intact|intact
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3862,3869|false|false|false|C0017725|glucose|GLUCOSE
Drug|Organic Chemical|SIMPLE_SEGMENT|3862,3869|false|false|false|C0017725|glucose|GLUCOSE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3862,3869|false|false|false|C0017725|glucose|GLUCOSE
Event|Event|SIMPLE_SEGMENT|3862,3869|false|false|false|||GLUCOSE
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3862,3869|false|false|false|C5781949|Glucose^1.5H post dose glucagon|GLUCOSE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3862,3869|false|false|false|C0337438|Glucose measurement|GLUCOSE
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3875,3879|false|false|false|C0041942|urea|UREA
Drug|Organic Chemical|SIMPLE_SEGMENT|3875,3879|false|false|false|C0041942|urea|UREA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3875,3879|false|false|false|C0041942|urea|UREA
Event|Event|SIMPLE_SEGMENT|3875,3879|false|false|false|||UREA
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3875,3879|false|false|false|C0523961|Urea measurement|UREA
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3897,3903|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|3897,3903|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3897,3903|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Event|Event|SIMPLE_SEGMENT|3897,3903|false|false|false|||SODIUM
Finding|Physiologic Function|SIMPLE_SEGMENT|3897,3903|false|false|false|C4553025|Sodium metabolic function|SODIUM
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3897,3903|false|false|false|C0337443|Sodium measurement|SODIUM
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3909,3918|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|3909,3918|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Food|SIMPLE_SEGMENT|3909,3918|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Inorganic Chemical|SIMPLE_SEGMENT|3909,3918|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3909,3918|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Event|Event|SIMPLE_SEGMENT|3909,3918|false|false|false|||POTASSIUM
Finding|Physiologic Function|SIMPLE_SEGMENT|3909,3918|false|false|false|C4553027|Potassium metabolic function|POTASSIUM
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3909,3918|false|false|false|C0202194|Potassium measurement|POTASSIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|3923,3931|false|false|false|C0008203;C0596019|Chlorides;chloride ion|CHLORIDE
Event|Event|SIMPLE_SEGMENT|3923,3931|false|false|false|||CHLORIDE
Finding|Physiologic Function|SIMPLE_SEGMENT|3923,3931|false|false|false|C4553021|Chloride metabolic function|CHLORIDE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3923,3931|false|false|false|C0201952|Chloride measurement|CHLORIDE
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3942,3945|false|false|false|C0007012|carbon dioxide|CO2
Drug|Inorganic Chemical|SIMPLE_SEGMENT|3942,3945|false|false|false|C0007012|carbon dioxide|CO2
Event|Event|SIMPLE_SEGMENT|3942,3945|false|false|false|||CO2
Finding|Finding|SIMPLE_SEGMENT|3942,3945|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Finding|Gene or Genome|SIMPLE_SEGMENT|3942,3945|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|3949,3954|false|false|false|C0003075|Anions|ANION
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3949,3958|false|false|false|C0003074|Anion Gap|ANION GAP
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3949,3958|false|false|false|C1509129|Anion gap result|ANION GAP
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3949,3958|false|false|false|C0201889;C2189246|Anion gap measurement;blood anion gap (lab test)|ANION GAP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3955,3958|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3955,3958|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Event|Event|SIMPLE_SEGMENT|3955,3958|false|false|false|||GAP
Finding|Gene or Genome|SIMPLE_SEGMENT|3955,3958|false|false|false|C1419277;C2984552|RASA1 gene;RASA1 wt Allele|GAP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4007,4010|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4007,4010|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|SIMPLE_SEGMENT|4007,4010|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|SIMPLE_SEGMENT|4007,4010|false|false|false|||ALT
Finding|Gene or Genome|SIMPLE_SEGMENT|4007,4010|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|SIMPLE_SEGMENT|4007,4010|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|SIMPLE_SEGMENT|4007,4010|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4007,4010|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4011,4015|false|false|false|C0376147|SGPT - Glutamate pyruvate transaminase|SGPT
Drug|Enzyme|SIMPLE_SEGMENT|4011,4015|false|false|false|C0376147|SGPT - Glutamate pyruvate transaminase|SGPT
Event|Event|SIMPLE_SEGMENT|4011,4015|false|false|false|||SGPT
Finding|Gene or Genome|SIMPLE_SEGMENT|4011,4015|false|false|false|C1415274|GPT gene|SGPT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4011,4015|false|false|false|C0036828|Serum Alanine Transaminase Test|SGPT
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4022,4025|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4022,4025|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4022,4025|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4022,4025|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|SIMPLE_SEGMENT|4022,4025|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|SIMPLE_SEGMENT|4022,4025|false|false|false|||AST
Finding|Gene or Genome|SIMPLE_SEGMENT|4022,4025|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4026,4030|false|false|false|C0242192|SGOT - Glutamate oxaloacetate transaminase|SGOT
Drug|Enzyme|SIMPLE_SEGMENT|4026,4030|false|false|false|C0242192|SGOT - Glutamate oxaloacetate transaminase|SGOT
Event|Event|SIMPLE_SEGMENT|4026,4030|false|false|false|||SGOT
Finding|Gene or Genome|SIMPLE_SEGMENT|4026,4030|false|false|false|C1415181|GOT1 gene|SGOT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4026,4030|false|false|false|C0201899|Aspartate aminotransferase measurement|SGOT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4037,4040|false|false|false|C1663627|ALK protein, human|ALK
Drug|Enzyme|SIMPLE_SEGMENT|4037,4040|false|false|false|C1663627|ALK protein, human|ALK
Event|Event|SIMPLE_SEGMENT|4037,4040|false|false|false|||ALK
Finding|Gene or Genome|SIMPLE_SEGMENT|4037,4040|false|false|false|C1332080;C1663627;C1704943|ALK gene;ALK protein, human;ALK wt Allele|ALK
Finding|Receptor|SIMPLE_SEGMENT|4037,4040|false|false|false|C1332080;C1663627;C1704943|ALK gene;ALK protein, human;ALK wt Allele|ALK
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4037,4045|false|false|false|C0002059|Alkaline Phosphatase|ALK PHOS
Drug|Enzyme|SIMPLE_SEGMENT|4037,4045|false|false|false|C0002059|Alkaline Phosphatase|ALK PHOS
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4037,4045|false|false|false|C0201850|Alkaline phosphatase measurement|ALK PHOS
Event|Event|SIMPLE_SEGMENT|4041,4045|false|false|false|||PHOS
Event|Event|SIMPLE_SEGMENT|4052,4055|false|false|false|||TOT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4080,4086|false|false|false|C0023764|lipase|LIPASE
Drug|Enzyme|SIMPLE_SEGMENT|4080,4086|false|false|false|C0023764|lipase|LIPASE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4080,4086|false|false|false|C0023764|lipase|LIPASE
Event|Event|SIMPLE_SEGMENT|4080,4086|false|false|false|||LIPASE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4080,4086|false|false|false|C0373670|Lipase measurement|LIPASE
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4105,4112|false|false|false|C0001924;C5966160|Albumin;Albumins|ALBUMIN
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4105,4112|false|false|false|C0001924;C5966160|Albumin;Albumins|ALBUMIN
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4105,4112|false|false|false|C0001924;C5966160|Albumin;Albumins|ALBUMIN
Event|Event|SIMPLE_SEGMENT|4105,4112|false|false|false|||ALBUMIN
Finding|Gene or Genome|SIMPLE_SEGMENT|4105,4112|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|ALBUMIN
Finding|Physiologic Function|SIMPLE_SEGMENT|4105,4112|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|ALBUMIN
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4105,4112|false|false|false|C0201838|Albumin measurement|ALBUMIN
Anatomy|Cell|SIMPLE_SEGMENT|4132,4135|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|4141,4144|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4141,4144|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4141,4144|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4150,4153|false|false|false|C0019046|Hemoglobin|HGB
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4150,4153|false|false|false|C0019046|Hemoglobin|HGB
Event|Event|SIMPLE_SEGMENT|4150,4153|false|false|false|||HGB
Finding|Gene or Genome|SIMPLE_SEGMENT|4150,4153|false|false|false|C1424337|CYGB gene|HGB
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4150,4153|false|false|false|C0019029|Hemoglobin concentration|HGB
Event|Event|SIMPLE_SEGMENT|4159,4162|false|false|false|||HCT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4159,4162|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4159,4162|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Disorder|Virus|SIMPLE_SEGMENT|4168,4171|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|4168,4171|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4168,4171|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4168,4171|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4168,4171|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|4177,4180|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4177,4180|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|4177,4180|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|4177,4180|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|4177,4180|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4177,4180|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4187,4191|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Event|Event|SIMPLE_SEGMENT|4197,4200|false|false|false|||RDW
Finding|Body Substance|SIMPLE_SEGMENT|4233,4239|false|false|false|C0024202|Lymph|LYMPHS
Event|Event|SIMPLE_SEGMENT|4243,4244|false|false|false|||5
Drug|Antibiotic|SIMPLE_SEGMENT|4246,4251|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4246,4251|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Organic Chemical|SIMPLE_SEGMENT|4246,4251|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4256,4259|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|EOS
Event|Event|SIMPLE_SEGMENT|4256,4259|false|false|false|||EOS
Finding|Gene or Genome|SIMPLE_SEGMENT|4256,4259|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|EOS
Event|Event|SIMPLE_SEGMENT|4290,4293|false|false|false|||PLT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4290,4293|false|false|false|C0201617|Primed lymphocyte test|PLT
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4322,4325|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|SIMPLE_SEGMENT|4322,4325|false|false|false|||PTT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4322,4325|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Event|Event|SIMPLE_SEGMENT|4356,4359|false|false|false|||CXR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4356,4359|false|false|false|C0039985|Plain chest X-ray|CXR
Finding|Intellectual Product|SIMPLE_SEGMENT|4364,4369|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4370,4385|false|false|false|C0553534|Cardiopulmonary|cardiopulmonary
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4370,4385|false|false|false|C4072686|Cardiovascular disease+Pulmonary disease|cardiopulmonary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4386,4393|false|false|false|C1184743|bony process|process
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4386,4393|true|false|false|C1951340|Process Pharmacologic Substance|process
Event|Event|SIMPLE_SEGMENT|4386,4393|false|false|false|||process
Finding|Functional Concept|SIMPLE_SEGMENT|4386,4393|true|false|false|C4521054|Process (qualifier value)|process
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|4386,4393|true|false|false|C1522240|Process|process
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4415,4425|false|false|false|C0550215||appearance
Event|Event|SIMPLE_SEGMENT|4415,4425|false|false|false|||appearance
Procedure|Health Care Activity|SIMPLE_SEGMENT|4415,4425|false|false|false|C2051406|patient appearance regarding mental status exam|appearance
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4433,4438|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4433,4438|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4433,4438|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|SIMPLE_SEGMENT|4433,4438|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4433,4438|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|SIMPLE_SEGMENT|4433,4438|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|SIMPLE_SEGMENT|4433,4438|false|false|false|||liver
Finding|Finding|SIMPLE_SEGMENT|4433,4438|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|SIMPLE_SEGMENT|4433,4438|false|false|false|C0872387|Procedures on liver|liver
Event|Event|SIMPLE_SEGMENT|4439,4449|false|false|false|||compatible
Finding|Idea or Concept|SIMPLE_SEGMENT|4439,4449|false|false|false|C0332290|Consistent with|compatible
Finding|Idea or Concept|SIMPLE_SEGMENT|4439,4454|false|false|false|C0332290|Consistent with|compatible with
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4455,4464|false|false|false|C0023890;C1623038|Cirrhosis;Liver Cirrhosis|cirrhosis
Event|Event|SIMPLE_SEGMENT|4455,4464|false|false|false|||cirrhosis
Event|Event|SIMPLE_SEGMENT|4467,4472|false|false|false|||Signs
Finding|Finding|SIMPLE_SEGMENT|4467,4472|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|Signs
Finding|Functional Concept|SIMPLE_SEGMENT|4467,4472|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|Signs
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4476,4482|false|false|false|C0205054|Hepatic|portal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4485,4497|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|SIMPLE_SEGMENT|4485,4497|false|false|false|||hypertension
Event|Event|SIMPLE_SEGMENT|4514,4520|false|false|false|||amount
Finding|Intellectual Product|SIMPLE_SEGMENT|4514,4520|false|false|false|C1561574|Amount class - Amount|amount
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4524,4531|false|false|false|C0003962|Ascites|ascites
Event|Event|SIMPLE_SEGMENT|4524,4531|false|false|false|||ascites
Finding|Pathologic Function|SIMPLE_SEGMENT|4524,4531|false|false|false|C5441966|Peritoneal Effusion|ascites
Event|Event|SIMPLE_SEGMENT|4536,4548|false|false|false|||splenomegaly
Finding|Finding|SIMPLE_SEGMENT|4536,4548|false|false|false|C0038002|Splenomegaly|splenomegaly
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4556,4570|false|false|false|C0008350|Cholelithiasis|Cholelithiasis
Event|Event|SIMPLE_SEGMENT|4556,4570|false|false|false|||Cholelithiasis
Finding|Intellectual Product|SIMPLE_SEGMENT|4577,4583|false|false|false|C0030650|Legal patent|Patent
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4584,4590|false|false|false|C0205054|Hepatic|portal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4584,4596|false|false|false|C0032718|Portal vein structure|portal veins
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4591,4596|false|false|false|C0042449|Veins|veins
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4591,4596|false|false|false|C0398102|Procedure on vein|veins
Event|Event|SIMPLE_SEGMENT|4621,4625|false|false|false|||flow
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|4621,4625|false|false|false|C0806140|Flow|flow
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|4629,4639|false|false|false|C0358514|Diagnostic agents|Diagnostic
Event|Event|SIMPLE_SEGMENT|4629,4639|false|false|false|||Diagnostic
Finding|Functional Concept|SIMPLE_SEGMENT|4629,4639|false|false|false|C0348026;C1547424|Diagnostic;Location Service Code - Diagnostic|Diagnostic
Finding|Intellectual Product|SIMPLE_SEGMENT|4629,4639|false|false|false|C0348026;C1547424|Diagnostic;Location Service Code - Diagnostic|Diagnostic
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4629,4639|false|false|false|C0011900;C0430533|Diagnosis;Diagnostic dental procedure|Diagnostic
Event|Event|SIMPLE_SEGMENT|4640,4644|false|false|false|||para
Finding|Finding|SIMPLE_SEGMENT|4640,4644|false|false|false|C0030563|Parity|para
Event|Event|SIMPLE_SEGMENT|4645,4654|false|false|false|||attempted
Event|Event|SIMPLE_SEGMENT|4666,4678|false|false|false|||unsuccessful
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|4689,4694|false|false|false|C3714591|Floor (anatomic)|floor
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4703,4706|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|abd
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|4703,4706|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|abd
Event|Event|SIMPLE_SEGMENT|4707,4717|false|false|false|||distension
Finding|Finding|SIMPLE_SEGMENT|4707,4717|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distension
Finding|Pathologic Function|SIMPLE_SEGMENT|4707,4717|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distension
Event|Event|SIMPLE_SEGMENT|4722,4732|false|false|false|||discomfort
Finding|Sign or Symptom|SIMPLE_SEGMENT|4722,4732|false|false|false|C2364135|Discomfort|discomfort
Finding|Intellectual Product|SIMPLE_SEGMENT|4736,4741|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|Brief
Finding|Idea or Concept|SIMPLE_SEGMENT|4742,4750|false|false|false|C1547192|Organization unit type - Hospital|Hospital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4742,4757|false|false|false|C0488549||Hospital Course
Finding|Finding|SIMPLE_SEGMENT|4742,4757|false|false|false|C0489547|Hospital course|Hospital Course
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4763,4766|false|false|false|C0019196;C0220847|Hepatitis C;hepatitis C virus|HCV
Disorder|Virus|SIMPLE_SEGMENT|4763,4766|false|false|false|C0019196;C0220847|Hepatitis C;hepatitis C virus|HCV
Event|Event|SIMPLE_SEGMENT|4763,4766|false|false|false|||HCV
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4767,4776|false|false|false|C0023890;C1623038|Cirrhosis;Liver Cirrhosis|cirrhosis
Event|Event|SIMPLE_SEGMENT|4767,4776|false|false|false|||cirrhosis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4781,4788|false|false|false|C0003962|Ascites|ascites
Event|Event|SIMPLE_SEGMENT|4781,4788|false|false|false|||ascites
Finding|Pathologic Function|SIMPLE_SEGMENT|4781,4788|false|false|false|C5441966|Peritoneal Effusion|ascites
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4790,4793|false|false|false|C0019682;C0019693|HIV;HIV Infections|hiv
Disorder|Virus|SIMPLE_SEGMENT|4790,4793|false|false|false|C0019682;C0019693|HIV;HIV Infections|hiv
Drug|Immunologic Factor|SIMPLE_SEGMENT|4790,4793|false|false|false|C0086413|HIV Vaccine|hiv
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4790,4793|false|false|false|C0086413|HIV Vaccine|hiv
Event|Event|SIMPLE_SEGMENT|4790,4793|false|false|false|||hiv
Drug|Organic Chemical|SIMPLE_SEGMENT|4797,4800|false|false|false|C0052432|artesunate|ART
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4797,4800|false|false|false|C0052432|artesunate|ART
Event|Event|SIMPLE_SEGMENT|4797,4800|false|false|false|||ART
Finding|Gene or Genome|SIMPLE_SEGMENT|4797,4800|false|false|false|C1412286;C3890191|AGRP gene;AGRP wt Allele|ART
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4797,4800|false|false|false|C0872104;C1963724|Antiretroviral therapy;Assisted Reproductive Technologies|ART
Event|Event|SIMPLE_SEGMENT|4806,4810|false|false|false|||IVDU
Finding|Individual Behavior|SIMPLE_SEGMENT|4806,4810|false|false|false|C0699778|intravenous drug use|IVDU
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4812,4816|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4812,4816|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|SIMPLE_SEGMENT|4812,4816|false|false|false|||COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|4812,4816|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4828,4832|false|false|false|C0038436;C0878676|6-pyruvoyl-tetrahydropterin synthase deficiency;Post-Traumatic Stress Disorder|PTSD
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|4828,4832|false|false|false|C0038436;C0878676|6-pyruvoyl-tetrahydropterin synthase deficiency;Post-Traumatic Stress Disorder|PTSD
Event|Event|SIMPLE_SEGMENT|4828,4832|false|false|false|||PTSD
Event|Event|SIMPLE_SEGMENT|4834,4843|false|false|false|||presented
Finding|Idea or Concept|SIMPLE_SEGMENT|4861,4870|false|false|false|C1546960|Patient Outcome - Worsening|worsening
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4871,4874|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|abd
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|4871,4874|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|abd
Event|Event|SIMPLE_SEGMENT|4876,4886|false|false|false|||distension
Finding|Finding|SIMPLE_SEGMENT|4876,4886|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distension
Finding|Pathologic Function|SIMPLE_SEGMENT|4876,4886|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distension
Finding|Intellectual Product|SIMPLE_SEGMENT|4897,4901|false|false|false|C1561540|Transaction counts and value totals - week|week
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|4906,4915|false|false|false|C0009676|Confusion|confusion
Event|Event|SIMPLE_SEGMENT|4906,4915|false|false|false|||confusion
Finding|Finding|SIMPLE_SEGMENT|4906,4915|false|false|false|C0683369|Clouded consciousness|confusion
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4922,4929|false|false|false|C0003962|Ascites|Ascites
Finding|Pathologic Function|SIMPLE_SEGMENT|4922,4929|false|false|false|C5441966|Peritoneal Effusion|Ascites
Event|Event|SIMPLE_SEGMENT|4922,4931|false|false|false|||Ascites -
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4946,4949|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|abd
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|4946,4949|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|abd
Event|Event|SIMPLE_SEGMENT|4950,4960|false|false|false|||distension
Finding|Finding|SIMPLE_SEGMENT|4950,4960|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distension
Finding|Pathologic Function|SIMPLE_SEGMENT|4950,4960|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distension
Event|Event|SIMPLE_SEGMENT|4965,4975|false|false|false|||discomfort
Finding|Sign or Symptom|SIMPLE_SEGMENT|4965,4975|false|false|false|C2364135|Discomfort|discomfort
Event|Event|SIMPLE_SEGMENT|4986,4990|false|false|false|||week
Finding|Intellectual Product|SIMPLE_SEGMENT|4986,4990|false|false|false|C1561540|Transaction counts and value totals - week|week
Finding|Finding|SIMPLE_SEGMENT|4992,4998|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|4992,4998|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5003,5009|false|false|false|C0205054|Hepatic|portal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5010,5013|false|true|false|C0020538|Hypertensive disease|HTN
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5031,5036|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5031,5036|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5031,5036|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|SIMPLE_SEGMENT|5031,5036|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5031,5036|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|SIMPLE_SEGMENT|5031,5036|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Finding|Finding|SIMPLE_SEGMENT|5031,5036|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|SIMPLE_SEGMENT|5031,5036|false|false|false|C0872387|Procedures on liver|liver
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5031,5044|false|false|false|C0023895;C0267792|Hepatobiliary Disorder;Liver diseases|liver disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5037,5044|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|5037,5044|false|false|false|||disease
Finding|Body Substance|SIMPLE_SEGMENT|5057,5070|false|false|false|C5441965|Ascitic Fluid|ascitic fluid
Drug|Substance|SIMPLE_SEGMENT|5065,5070|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|5065,5070|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|5065,5070|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|5071,5080|false|false|false|||available
Finding|Functional Concept|SIMPLE_SEGMENT|5071,5080|false|false|false|C0470187|Availability of|available
Event|Event|SIMPLE_SEGMENT|5093,5102|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|5093,5102|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|SIMPLE_SEGMENT|5108,5113|false|false|false|||signs
Finding|Finding|SIMPLE_SEGMENT|5108,5113|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|SIMPLE_SEGMENT|5108,5113|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5117,5122|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5117,5122|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|5117,5122|false|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5117,5130|false|false|false|C0018801;C0018802|Congestive heart failure;Heart failure|heart failure
Event|Event|SIMPLE_SEGMENT|5123,5130|false|false|false|||failure
Finding|Functional Concept|SIMPLE_SEGMENT|5123,5130|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|SIMPLE_SEGMENT|5123,5130|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|SIMPLE_SEGMENT|5123,5130|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Event|Event|SIMPLE_SEGMENT|5131,5136|false|false|false|||noted
Event|Event|SIMPLE_SEGMENT|5140,5144|false|false|false|||exam
Finding|Functional Concept|SIMPLE_SEGMENT|5140,5144|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|5140,5144|false|false|false|C0582103|Medical Examination|exam
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|5162,5165|false|false|false|C0026760|Multiple Epiphyseal Dysplasia|med
Finding|Gene or Genome|SIMPLE_SEGMENT|5162,5165|false|false|false|C1413596;C1413597;C1419866;C1456376;C1549978;C4321267;C5781216|COL9A2 gene;COL9A3 gene;COMP gene;COMP wt Allele;Master of Education;SCN8A gene;SCN8A wt Allele|med
Finding|Intellectual Product|SIMPLE_SEGMENT|5162,5165|false|false|false|C1413596;C1413597;C1419866;C1456376;C1549978;C4321267;C5781216|COL9A2 gene;COL9A3 gene;COMP gene;COMP wt Allele;Master of Education;SCN8A gene;SCN8A wt Allele|med
Drug|Food|SIMPLE_SEGMENT|5194,5198|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|SIMPLE_SEGMENT|5194,5198|false|false|false|||diet
Finding|Functional Concept|SIMPLE_SEGMENT|5194,5198|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|SIMPLE_SEGMENT|5194,5198|false|false|false|C0012159|Diet therapy|diet
Event|Event|SIMPLE_SEGMENT|5199,5210|false|false|false|||restriction
Finding|Functional Concept|SIMPLE_SEGMENT|5199,5210|false|false|false|C0443288|Restricted|restriction
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5212,5215|true|false|false|C0871470|Systolic Pressure|SBP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5212,5215|true|false|false|C0085805|Androgen Binding Protein|SBP
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5212,5215|true|false|false|C0085805|Androgen Binding Protein|SBP
Event|Event|SIMPLE_SEGMENT|5212,5215|false|false|false|||SBP
Finding|Gene or Genome|SIMPLE_SEGMENT|5212,5215|true|false|false|C1705296;C3274833|CCHCR1 wt Allele;SHBG wt Allele|SBP
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5212,5215|true|false|false|C1306620|Systolic blood pressure measurement|SBP
Event|Event|SIMPLE_SEGMENT|5216,5224|false|false|false|||negative
Finding|Classification|SIMPLE_SEGMENT|5216,5224|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|5216,5224|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5216,5224|false|false|false|C5237010|Expression Negative|negative
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5225,5234|false|false|false|C0012798|Diuretics|diuretics
Event|Event|SIMPLE_SEGMENT|5225,5234|false|false|false|||diuretics
Drug|Organic Chemical|SIMPLE_SEGMENT|5240,5250|false|false|false|C0016860|furosemide|Furosemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5240,5250|false|false|false|C0016860|furosemide|Furosemide
Drug|Organic Chemical|SIMPLE_SEGMENT|5270,5284|false|false|false|C0037982|spironolactone|Spironolactone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5270,5284|false|false|false|C0037982|spironolactone|Spironolactone
Event|Event|SIMPLE_SEGMENT|5301,5307|false|false|false|||chosen
Event|Event|SIMPLE_SEGMENT|5330,5334|false|false|false|||dose
Event|Event|SIMPLE_SEGMENT|5336,5337|false|false|false|||/
Event|Event|SIMPLE_SEGMENT|5354,5357|false|false|false|||CXR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5354,5357|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|SIMPLE_SEGMENT|5370,5378|false|false|false|||negative
Finding|Classification|SIMPLE_SEGMENT|5370,5378|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|5370,5378|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5370,5378|false|false|false|C5237010|Expression Negative|negative
Finding|Body Substance|SIMPLE_SEGMENT|5380,5385|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Finding|Functional Concept|SIMPLE_SEGMENT|5380,5385|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Finding|Intellectual Product|SIMPLE_SEGMENT|5380,5385|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5380,5393|true|false|false|C0430404|Urine culture|Urine culture
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5386,5393|false|false|false|C1706355|Culture Dose Form|culture
Event|Event|SIMPLE_SEGMENT|5386,5393|false|false|false|||culture
Finding|Functional Concept|SIMPLE_SEGMENT|5386,5393|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Finding|Idea or Concept|SIMPLE_SEGMENT|5386,5393|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5386,5393|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|culture
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5386,5399|false|false|false|C0200949|Blood culture|culture blood
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5394,5399|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|5394,5399|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|5394,5399|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5394,5407|false|false|false|C0200949|Blood culture|blood culture
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5394,5416|false|false|false|C0852859|Blood culture negative|blood culture negative
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5400,5407|false|false|false|C1706355|Culture Dose Form|culture
Event|Event|SIMPLE_SEGMENT|5400,5407|false|false|false|||culture
Finding|Functional Concept|SIMPLE_SEGMENT|5400,5407|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Finding|Idea or Concept|SIMPLE_SEGMENT|5400,5407|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5400,5407|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|culture
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5400,5416|false|false|false|C0855652|Culture negative|culture negative
Event|Event|SIMPLE_SEGMENT|5408,5416|false|false|false|||negative
Finding|Classification|SIMPLE_SEGMENT|5408,5416|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|5408,5416|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5408,5416|false|false|false|C5237010|Expression Negative|negative
Event|Event|SIMPLE_SEGMENT|5428,5434|false|false|false|||losing
Finding|Pathologic Function|SIMPLE_SEGMENT|5435,5447|false|false|false|C0013604;C0546817|Edema;Hypervolemia (finding)|excess fluid
Drug|Substance|SIMPLE_SEGMENT|5442,5447|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|5442,5447|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|5442,5447|false|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|5467,5473|false|false|false|C1547311|Patient Condition Code - Stable|stable
Finding|Idea or Concept|SIMPLE_SEGMENT|5488,5493|false|false|false|C1552828|Table Frame - above|above
Event|Event|SIMPLE_SEGMENT|5494,5501|false|false|false|||regimen
Finding|Intellectual Product|SIMPLE_SEGMENT|5494,5501|false|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5494,5501|false|false|false|C0040808|Treatment Protocols|regimen
Event|Event|SIMPLE_SEGMENT|5510,5519|false|false|false|||scheduled
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|5525,5532|false|false|false|C1705970|Electrical Current|current
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5533,5536|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|5533,5536|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5533,5536|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5533,5536|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|SIMPLE_SEGMENT|5533,5536|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|5533,5536|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|SIMPLE_SEGMENT|5533,5536|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5533,5536|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|SIMPLE_SEGMENT|5533,5536|false|false|false|||PCP
Finding|Gene or Genome|SIMPLE_SEGMENT|5533,5536|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|SIMPLE_SEGMENT|5533,5536|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Event|SIMPLE_SEGMENT|5546,5551|false|false|false|||check
Event|Event|SIMPLE_SEGMENT|5557,5566|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|5557,5566|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|5557,5566|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|5557,5566|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|5557,5566|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|SIMPLE_SEGMENT|5578,5587|false|false|false|||scheduled
Finding|Finding|SIMPLE_SEGMENT|5592,5595|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|5592,5595|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5596,5599|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|5596,5599|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5596,5599|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5596,5599|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|SIMPLE_SEGMENT|5596,5599|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|5596,5599|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|SIMPLE_SEGMENT|5596,5599|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5596,5599|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|SIMPLE_SEGMENT|5596,5599|false|false|false|||PCP
Finding|Gene or Genome|SIMPLE_SEGMENT|5596,5599|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|SIMPLE_SEGMENT|5596,5599|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Event|SIMPLE_SEGMENT|5625,5631|false|false|false|||follow
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5638,5643|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|Liver
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5638,5643|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|Liver
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5638,5643|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|Liver
Drug|Organic Chemical|SIMPLE_SEGMENT|5638,5643|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|Liver
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5638,5643|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|Liver
Drug|Vitamin|SIMPLE_SEGMENT|5638,5643|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|Liver
Finding|Finding|SIMPLE_SEGMENT|5638,5643|false|false|false|C0577060|Liver problem|Liver
Procedure|Health Care Activity|SIMPLE_SEGMENT|5638,5643|false|false|false|C0872387|Procedures on liver|Liver
Event|Event|SIMPLE_SEGMENT|5654,5662|false|false|false|||schedule
Finding|Intellectual Product|SIMPLE_SEGMENT|5654,5662|false|false|false|C0086960|Schedule (document)|schedule
Procedure|Health Care Activity|SIMPLE_SEGMENT|5654,5662|false|false|false|C1446911|Scheduling (procedure)|schedule
Finding|Classification|SIMPLE_SEGMENT|5663,5673|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|5663,5673|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|SIMPLE_SEGMENT|5674,5683|false|false|false|||screening
Finding|Finding|SIMPLE_SEGMENT|5674,5683|false|false|false|C0220909;C1305399;C1409616|Aspects of disease screening;Screening - procedure intent;Special screening finding|screening
Finding|Functional Concept|SIMPLE_SEGMENT|5674,5683|false|false|false|C0220909;C1305399;C1409616|Aspects of disease screening;Screening - procedure intent;Special screening finding|screening
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5674,5683|false|false|false|C0199230;C0220908;C1698960;C1710031;C1710032|Disease Screening;Screening;Screening for cancer;Screening procedure;research subject screening|screening
Procedure|Health Care Activity|SIMPLE_SEGMENT|5674,5683|false|false|false|C0199230;C0220908;C1698960;C1710031;C1710032|Disease Screening;Screening;Screening for cancer;Screening procedure;research subject screening|screening
Procedure|Research Activity|SIMPLE_SEGMENT|5674,5683|false|false|false|C0199230;C0220908;C1698960;C1710031;C1710032|Disease Screening;Screening;Screening for cancer;Screening procedure;research subject screening|screening
Event|Event|SIMPLE_SEGMENT|5684,5687|false|false|false|||EGD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5684,5687|false|false|false|C0079304|Esophagogastroduodenoscopy|EGD
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5706,5717|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5706,5717|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|5706,5717|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|5706,5717|false|false|false|C4284232|Medications|Medications
Finding|Finding|SIMPLE_SEGMENT|5706,5730|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|SIMPLE_SEGMENT|5721,5730|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|5721,5730|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5749,5759|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|5749,5759|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|5749,5764|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|SIMPLE_SEGMENT|5760,5764|false|false|false|||list
Finding|Intellectual Product|SIMPLE_SEGMENT|5760,5764|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|SIMPLE_SEGMENT|5768,5776|false|false|false|||accurate
Drug|Organic Chemical|SIMPLE_SEGMENT|5781,5789|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5781,5789|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|SIMPLE_SEGMENT|5781,5789|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|SIMPLE_SEGMENT|5781,5789|false|false|false|||complete
Finding|Functional Concept|SIMPLE_SEGMENT|5781,5789|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|SIMPLE_SEGMENT|5781,5789|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Organic Chemical|SIMPLE_SEGMENT|5794,5804|false|false|false|C0016860|furosemide|Furosemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5794,5804|false|false|false|C0016860|furosemide|Furosemide
Drug|Organic Chemical|SIMPLE_SEGMENT|5824,5838|false|false|false|C0037982|spironolactone|Spironolactone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5824,5838|false|false|false|C0037982|spironolactone|Spironolactone
Drug|Organic Chemical|SIMPLE_SEGMENT|5858,5867|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5858,5867|false|false|false|C0001927|albuterol|Albuterol
Finding|Functional Concept|SIMPLE_SEGMENT|5868,5875|false|false|false|C4319647|Inhaler (unit of presentation)|Inhaler
Finding|Gene or Genome|SIMPLE_SEGMENT|5890,5893|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|SIMPLE_SEGMENT|5894,5902|false|false|false|||wheezing
Finding|Sign or Symptom|SIMPLE_SEGMENT|5894,5902|false|false|false|C0043144|Wheezing|wheezing
Event|Event|SIMPLE_SEGMENT|5904,5907|false|false|false|||SOB
Finding|Sign or Symptom|SIMPLE_SEGMENT|5904,5907|false|false|false|C0013404|Dyspnea|SOB
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|5912,5923|false|false|false|C1871526|raltegravir|Raltegravir
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5912,5923|false|false|false|C1871526|raltegravir|Raltegravir
Event|Event|SIMPLE_SEGMENT|5912,5923|false|false|false|||Raltegravir
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|5934,5937|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5934,5937|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5934,5937|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|5934,5937|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|5934,5937|false|false|false|C1332410|BID gene|BID
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|5942,5955|false|false|false|C0909839|emtricitabine|Emtricitabine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5942,5955|false|false|false|C0909839|emtricitabine|Emtricitabine
Drug|Organic Chemical|SIMPLE_SEGMENT|5942,5965|false|false|false|C1532298|Emtricitabine- and tenofovir-containing product|Emtricitabine-Tenofovir
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5942,5965|false|false|false|C1532298|Emtricitabine- and tenofovir-containing product|Emtricitabine-Tenofovir
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|5956,5965|false|false|false|C0384228|tenofovir|Tenofovir
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5956,5965|false|false|false|C0384228|tenofovir|Tenofovir
Event|Event|SIMPLE_SEGMENT|5956,5965|false|false|false|||Tenofovir
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|5967,5974|false|false|false|C1528494|Truvada|Truvada
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5967,5974|false|false|false|C1528494|Truvada|Truvada
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5978,5981|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|SIMPLE_SEGMENT|5978,5981|false|false|false|||TAB
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|5995,6003|false|false|false|C0028040|nicotine|Nicotine
Drug|Organic Chemical|SIMPLE_SEGMENT|5995,6003|false|false|false|C0028040|nicotine|Nicotine
Event|Event|SIMPLE_SEGMENT|5995,6003|false|false|false|||Nicotine
Drug|Clinical Drug|SIMPLE_SEGMENT|5995,6009|false|false|false|C0358855|Nicotine Transdermal Patch|Nicotine Patch
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6004,6009|false|false|false|C0445403;C1533128;C1707974|Body tissue patch material;Human patch material;Patch - Extended Release Film|Patch
Event|Event|SIMPLE_SEGMENT|6004,6009|false|false|false|||Patch
Finding|Finding|SIMPLE_SEGMENT|6004,6009|false|false|false|C0332461|Plaque (lesion)|Patch
Drug|Organic Chemical|SIMPLE_SEGMENT|6029,6040|false|false|false|C0027235|ipratropium|Ipratropium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6029,6040|false|false|false|C0027235|ipratropium|Ipratropium
Event|Event|SIMPLE_SEGMENT|6029,6040|false|false|false|||Ipratropium
Drug|Organic Chemical|SIMPLE_SEGMENT|6029,6048|false|false|false|C0700580|ipratropium bromide|Ipratropium Bromide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6029,6048|false|false|false|C0700580|ipratropium bromide|Ipratropium Bromide
Drug|Inorganic Chemical|SIMPLE_SEGMENT|6041,6048|false|false|false|C0006222|Bromides|Bromide
Event|Event|SIMPLE_SEGMENT|6041,6048|false|false|false|||Bromide
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6041,6048|false|false|false|C0202341|Bromides measurement|Bromide
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6049,6052|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6049,6052|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6049,6052|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Event|Event|SIMPLE_SEGMENT|6049,6052|false|false|false|||Neb
Finding|Cell Function|SIMPLE_SEGMENT|6049,6052|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Finding|Gene or Genome|SIMPLE_SEGMENT|6049,6052|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6055,6058|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6055,6058|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6055,6058|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Event|Event|SIMPLE_SEGMENT|6055,6058|false|false|false|||NEB
Finding|Cell Function|SIMPLE_SEGMENT|6055,6058|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|SIMPLE_SEGMENT|6055,6058|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Event|Event|SIMPLE_SEGMENT|6066,6069|false|false|false|||SOB
Finding|Sign or Symptom|SIMPLE_SEGMENT|6066,6069|false|false|false|C0013404|Dyspnea|SOB
Event|Event|SIMPLE_SEGMENT|6074,6083|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|6074,6083|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|6074,6083|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|6074,6083|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|6074,6083|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|6074,6095|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6084,6095|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6084,6095|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|6084,6095|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|6084,6095|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|SIMPLE_SEGMENT|6100,6109|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6100,6109|false|false|false|C0001927|albuterol|Albuterol
Finding|Functional Concept|SIMPLE_SEGMENT|6110,6117|false|false|false|C4319647|Inhaler (unit of presentation)|Inhaler
Finding|Gene or Genome|SIMPLE_SEGMENT|6132,6135|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|SIMPLE_SEGMENT|6136,6144|false|false|false|||wheezing
Finding|Sign or Symptom|SIMPLE_SEGMENT|6136,6144|false|false|false|C0043144|Wheezing|wheezing
Event|Event|SIMPLE_SEGMENT|6146,6149|false|false|false|||SOB
Finding|Sign or Symptom|SIMPLE_SEGMENT|6146,6149|false|false|false|C0013404|Dyspnea|SOB
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|6154,6167|false|false|false|C0909839|emtricitabine|Emtricitabine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6154,6167|false|false|false|C0909839|emtricitabine|Emtricitabine
Drug|Organic Chemical|SIMPLE_SEGMENT|6154,6177|false|false|false|C1532298|Emtricitabine- and tenofovir-containing product|Emtricitabine-Tenofovir
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6154,6177|false|false|false|C1532298|Emtricitabine- and tenofovir-containing product|Emtricitabine-Tenofovir
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|6168,6177|false|false|false|C0384228|tenofovir|Tenofovir
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6168,6177|false|false|false|C0384228|tenofovir|Tenofovir
Event|Event|SIMPLE_SEGMENT|6168,6177|false|false|false|||Tenofovir
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|6179,6186|false|false|false|C1528494|Truvada|Truvada
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6179,6186|false|false|false|C1528494|Truvada|Truvada
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6190,6193|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|SIMPLE_SEGMENT|6190,6193|false|false|false|||TAB
Drug|Organic Chemical|SIMPLE_SEGMENT|6207,6217|false|false|false|C0016860|furosemide|Furosemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6207,6217|false|false|false|C0016860|furosemide|Furosemide
Event|Event|SIMPLE_SEGMENT|6234,6236|false|false|false|||RX
Drug|Organic Chemical|SIMPLE_SEGMENT|6238,6248|false|false|false|C0016860|furosemide|furosemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6238,6248|false|false|false|C0016860|furosemide|furosemide
Event|Event|SIMPLE_SEGMENT|6238,6248|false|false|false|||furosemide
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6257,6263|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|SIMPLE_SEGMENT|6267,6275|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6270,6275|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|6270,6275|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6292,6298|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|6292,6298|false|false|false|||Tablet
Event|Event|SIMPLE_SEGMENT|6300,6307|false|false|false|||Refills
Finding|Idea or Concept|SIMPLE_SEGMENT|6300,6307|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|6314,6325|false|false|false|C0027235|ipratropium|Ipratropium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6314,6325|false|false|false|C0027235|ipratropium|Ipratropium
Event|Event|SIMPLE_SEGMENT|6314,6325|false|false|false|||Ipratropium
Drug|Organic Chemical|SIMPLE_SEGMENT|6314,6333|false|false|false|C0700580|ipratropium bromide|Ipratropium Bromide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6314,6333|false|false|false|C0700580|ipratropium bromide|Ipratropium Bromide
Drug|Inorganic Chemical|SIMPLE_SEGMENT|6326,6333|false|false|false|C0006222|Bromides|Bromide
Event|Event|SIMPLE_SEGMENT|6326,6333|false|false|false|||Bromide
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6326,6333|false|false|false|C0202341|Bromides measurement|Bromide
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6334,6337|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6334,6337|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6334,6337|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Event|Event|SIMPLE_SEGMENT|6334,6337|false|false|false|||Neb
Finding|Cell Function|SIMPLE_SEGMENT|6334,6337|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Finding|Gene or Genome|SIMPLE_SEGMENT|6334,6337|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6340,6343|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6340,6343|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6340,6343|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Event|Event|SIMPLE_SEGMENT|6340,6343|false|false|false|||NEB
Finding|Cell Function|SIMPLE_SEGMENT|6340,6343|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|SIMPLE_SEGMENT|6340,6343|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Event|Event|SIMPLE_SEGMENT|6351,6354|false|false|false|||SOB
Finding|Sign or Symptom|SIMPLE_SEGMENT|6351,6354|false|false|false|C0013404|Dyspnea|SOB
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|6359,6367|false|false|false|C0028040|nicotine|Nicotine
Drug|Organic Chemical|SIMPLE_SEGMENT|6359,6367|false|false|false|C0028040|nicotine|Nicotine
Drug|Clinical Drug|SIMPLE_SEGMENT|6359,6373|false|false|false|C0358855|Nicotine Transdermal Patch|Nicotine Patch
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6368,6373|false|false|false|C0445403;C1533128;C1707974|Body tissue patch material;Human patch material;Patch - Extended Release Film|Patch
Event|Event|SIMPLE_SEGMENT|6368,6373|false|false|false|||Patch
Finding|Finding|SIMPLE_SEGMENT|6368,6373|false|false|false|C0332461|Plaque (lesion)|Patch
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|6393,6404|false|false|false|C1871526|raltegravir|Raltegravir
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6393,6404|false|false|false|C1871526|raltegravir|Raltegravir
Event|Event|SIMPLE_SEGMENT|6393,6404|false|false|false|||Raltegravir
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|6415,6418|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6415,6418|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6415,6418|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|6415,6418|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|6415,6418|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|6423,6437|false|false|false|C0037982|spironolactone|Spironolactone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6423,6437|false|false|false|C0037982|spironolactone|Spironolactone
Drug|Organic Chemical|SIMPLE_SEGMENT|6457,6470|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6457,6470|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|SIMPLE_SEGMENT|6457,6470|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6457,6470|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|SIMPLE_SEGMENT|6485,6488|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6489,6493|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|6489,6493|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|6489,6493|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|6489,6493|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|6498,6507|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|6498,6507|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|6498,6507|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|6498,6507|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|6498,6507|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6498,6519|false|false|false|C4019243||Discharge Disposition
Finding|Finding|SIMPLE_SEGMENT|6498,6519|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6508,6519|false|false|false|C2926604||Disposition
Event|Event|SIMPLE_SEGMENT|6508,6519|false|false|false|||Disposition
Procedure|Health Care Activity|SIMPLE_SEGMENT|6508,6519|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|SIMPLE_SEGMENT|6521,6525|false|false|false|||Home
Finding|Idea or Concept|SIMPLE_SEGMENT|6521,6525|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|SIMPLE_SEGMENT|6521,6525|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|SIMPLE_SEGMENT|6521,6525|false|false|false|C1553498|home health encounter|Home
Event|Event|SIMPLE_SEGMENT|6528,6537|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|6528,6537|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|6528,6537|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|6528,6537|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|6528,6537|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|6528,6547|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6538,6547|false|false|false|C0945731||Diagnosis
Event|Event|SIMPLE_SEGMENT|6538,6547|false|false|false|||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|6538,6547|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|6538,6547|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6538,6547|false|false|false|C0011900|Diagnosis|Diagnosis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6549,6556|false|false|false|C0003962|Ascites|Ascites
Event|Event|SIMPLE_SEGMENT|6549,6556|false|false|false|||Ascites
Finding|Pathologic Function|SIMPLE_SEGMENT|6549,6556|false|false|false|C5441966|Peritoneal Effusion|Ascites
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6562,6568|false|false|false|C0205054|Hepatic|Portal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6569,6572|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|SIMPLE_SEGMENT|6569,6572|false|false|false|||HTN
Event|Event|SIMPLE_SEGMENT|6576,6585|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|6576,6585|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|6576,6585|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|6576,6585|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|6576,6585|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6586,6595|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6586,6595|false|false|false|C0012634|Disease|Condition
Event|Event|SIMPLE_SEGMENT|6586,6595|false|false|false|||Condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|6586,6595|false|false|false|C1705253|Logical Condition|Condition
Finding|Mental Process|SIMPLE_SEGMENT|6597,6603|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6597,6610|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|SIMPLE_SEGMENT|6597,6610|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6604,6610|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|6604,6610|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|6612,6617|false|false|false|||Clear
Finding|Idea or Concept|SIMPLE_SEGMENT|6612,6617|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|SIMPLE_SEGMENT|6622,6630|false|false|false|||coherent
Finding|Finding|SIMPLE_SEGMENT|6622,6630|false|false|false|C4068804|Coherent|coherent
Event|Event|SIMPLE_SEGMENT|6632,6637|false|false|false|||Level
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6632,6654|false|false|false|C4050479||Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|6632,6654|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|SIMPLE_SEGMENT|6641,6654|false|false|false|||Consciousness
Finding|Finding|SIMPLE_SEGMENT|6641,6654|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|SIMPLE_SEGMENT|6641,6654|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6656,6661|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|6656,6661|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6656,6661|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|SIMPLE_SEGMENT|6656,6661|false|false|false|||Alert
Finding|Finding|SIMPLE_SEGMENT|6656,6661|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|6656,6661|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|6656,6661|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|SIMPLE_SEGMENT|6666,6677|false|false|false|||interactive
Finding|Functional Concept|SIMPLE_SEGMENT|6666,6677|false|false|false|C1704675|Interaction|interactive
Event|Activity|SIMPLE_SEGMENT|6679,6687|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|6679,6687|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|SIMPLE_SEGMENT|6679,6687|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6688,6694|false|false|false|C5889824||Status
Event|Event|SIMPLE_SEGMENT|6688,6694|false|false|false|||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|6688,6694|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|6696,6706|false|false|false|||Ambulatory
Finding|Functional Concept|SIMPLE_SEGMENT|6696,6706|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|SIMPLE_SEGMENT|6696,6706|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|SIMPLE_SEGMENT|6696,6706|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|SIMPLE_SEGMENT|6696,6706|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|SIMPLE_SEGMENT|6709,6720|false|false|false|||Independent
Finding|Finding|SIMPLE_SEGMENT|6709,6720|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|SIMPLE_SEGMENT|6709,6720|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Event|Event|SIMPLE_SEGMENT|6725,6734|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|6725,6734|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|6725,6734|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|6725,6734|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|6725,6734|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6725,6747|false|false|false|C3669312||Discharge Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|6725,6747|false|false|false|C4282220|Discharge instructions|Discharge Instructions
Procedure|Health Care Activity|SIMPLE_SEGMENT|6725,6747|false|false|false|C2266673|hospital discharge instructions (treatment)|Discharge Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6735,6747|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|6735,6747|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|6735,6747|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Finding|Gene or Genome|SIMPLE_SEGMENT|6749,6753|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Event|Event|SIMPLE_SEGMENT|6772,6780|false|false|false|||pleasure
Finding|Intellectual Product|SIMPLE_SEGMENT|6772,6780|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|SIMPLE_SEGMENT|6772,6780|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|SIMPLE_SEGMENT|6788,6792|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|6788,6792|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|6788,6792|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|6788,6792|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|6788,6795|false|false|false|C1555558|care of - AddressPartType|care of
Event|Event|SIMPLE_SEGMENT|6805,6809|false|false|false|||came
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6822,6829|false|false|false|C0038351;C3714551;C4266636|Abdomen>Stomach;Stomach;Stomach structure|stomach
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6822,6829|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6822,6829|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Event|Event|SIMPLE_SEGMENT|6822,6829|false|false|false|||stomach
Finding|Finding|SIMPLE_SEGMENT|6822,6829|false|false|false|C0577027|Stomach problem|stomach
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6822,6829|false|false|false|C0872393|Procedure on stomach|stomach
Finding|Sign or Symptom|SIMPLE_SEGMENT|6822,6834|false|false|false|C0000737;C0221512|Abdominal Pain;Stomach ache|stomach pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6830,6834|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|6830,6834|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|6830,6834|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|6830,6834|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Idea or Concept|SIMPLE_SEGMENT|6839,6848|false|false|false|C1546960|Patient Outcome - Worsening|worsening
Event|Event|SIMPLE_SEGMENT|6849,6859|false|false|false|||distension
Finding|Finding|SIMPLE_SEGMENT|6849,6859|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distension
Finding|Pathologic Function|SIMPLE_SEGMENT|6849,6859|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distension
Event|Event|SIMPLE_SEGMENT|6891,6903|false|false|false|||paracentesis
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6891,6903|false|false|false|C0034115|Paracentesis|paracentesis
Event|Event|SIMPLE_SEGMENT|6907,6913|false|false|false|||remove
Drug|Substance|SIMPLE_SEGMENT|6922,6927|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|6922,6927|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|6922,6927|false|false|false|C1546638|Fluid Specimen Code|fluid
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6938,6943|false|false|false|C0224086|Belly of skeletal muscle|belly
Event|Event|SIMPLE_SEGMENT|6954,6960|false|false|false|||placed
Drug|Organic Chemical|SIMPLE_SEGMENT|6981,6986|false|false|false|C0699992|Lasix|Lasix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6981,6986|false|false|false|C0699992|Lasix|Lasix
Drug|Organic Chemical|SIMPLE_SEGMENT|7000,7009|false|false|false|C0591054|Aldactone|Aldactone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7000,7009|false|false|false|C0591054|Aldactone|Aldactone
Event|Event|SIMPLE_SEGMENT|7014,7018|false|false|false|||help
Finding|Intellectual Product|SIMPLE_SEGMENT|7014,7018|false|false|false|C1552861|Help document|help
Event|Event|SIMPLE_SEGMENT|7023,7030|false|false|false|||urinate
Finding|Pathologic Function|SIMPLE_SEGMENT|7035,7047|false|false|false|C0013604;C0546817|Edema;Hypervolemia (finding)|excess fluid
Drug|Substance|SIMPLE_SEGMENT|7042,7047|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|7042,7047|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|7042,7047|false|false|false|C1546638|Fluid Specimen Code|fluid
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7048,7053|false|false|false|C1410088|Still|still
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7062,7067|false|false|false|C0224086|Belly of skeletal muscle|belly
Event|Event|SIMPLE_SEGMENT|7076,7085|false|false|false|||discussed
Event|Event|SIMPLE_SEGMENT|7112,7116|false|false|false|||dose
Drug|Organic Chemical|SIMPLE_SEGMENT|7120,7125|false|false|true|C0699992|Lasix|lasix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7120,7125|false|false|true|C0699992|Lasix|lasix
Event|Event|SIMPLE_SEGMENT|7120,7125|false|false|false|||lasix
Event|Event|SIMPLE_SEGMENT|7126,7134|false|false|false|||required
Event|Event|SIMPLE_SEGMENT|7139,7143|false|false|false|||make
Event|Event|SIMPLE_SEGMENT|7149,7156|false|false|false|||urinate
Event|Event|SIMPLE_SEGMENT|7166,7172|false|false|false|||likely
Finding|Finding|SIMPLE_SEGMENT|7166,7172|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|7166,7172|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|SIMPLE_SEGMENT|7199,7203|false|false|false|||high
Finding|Finding|SIMPLE_SEGMENT|7199,7203|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|SIMPLE_SEGMENT|7199,7203|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|SIMPLE_SEGMENT|7199,7203|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Event|Event|SIMPLE_SEGMENT|7212,7216|false|false|false|||dose
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7236,7247|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7236,7247|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|7236,7247|false|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|7236,7247|false|false|false|C4284232|Medications|medications
Event|Event|SIMPLE_SEGMENT|7262,7268|false|false|false|||excess
Drug|Substance|SIMPLE_SEGMENT|7270,7275|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|7270,7275|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|7276,7279|false|false|false|||off
Event|Event|SIMPLE_SEGMENT|7284,7287|false|false|false|||eat
Finding|Finding|SIMPLE_SEGMENT|7290,7293|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|SIMPLE_SEGMENT|7290,7293|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7290,7303|false|false|false|C0012169|Low sodium diet|low salt diet
Drug|Chemical Viewed Structurally|SIMPLE_SEGMENT|7294,7298|false|false|false|C0036140;C0037494;C0206136|Salts;Sodium Chloride, Dietary;sodium chloride|salt
Drug|Food|SIMPLE_SEGMENT|7294,7298|false|false|false|C0036140;C0037494;C0206136|Salts;Sodium Chloride, Dietary;sodium chloride|salt
Drug|Inorganic Chemical|SIMPLE_SEGMENT|7294,7298|false|false|false|C0036140;C0037494;C0206136|Salts;Sodium Chloride, Dietary;sodium chloride|salt
Drug|Food|SIMPLE_SEGMENT|7299,7303|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|SIMPLE_SEGMENT|7299,7303|false|false|false|||diet
Finding|Functional Concept|SIMPLE_SEGMENT|7299,7303|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|SIMPLE_SEGMENT|7299,7303|false|false|false|C0012159|Diet therapy|diet
Event|Event|SIMPLE_SEGMENT|7314,7320|false|false|false|||follow
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7341,7346|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7341,7346|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7341,7346|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|SIMPLE_SEGMENT|7341,7346|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7341,7346|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|SIMPLE_SEGMENT|7341,7346|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Finding|Finding|SIMPLE_SEGMENT|7341,7346|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|SIMPLE_SEGMENT|7341,7346|false|false|false|C0872387|Procedures on liver|liver
Event|Event|SIMPLE_SEGMENT|7379,7390|false|false|false|||colonoscopy
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7379,7390|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Procedure|Health Care Activity|SIMPLE_SEGMENT|7379,7390|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Event|Event|SIMPLE_SEGMENT|7396,7399|false|false|false|||EGD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7396,7399|false|false|false|C0079304|Esophagogastroduodenoscopy|EGD
Event|Event|SIMPLE_SEGMENT|7400,7409|false|false|false|||scheduled
Finding|Finding|SIMPLE_SEGMENT|7429,7435|false|false|false|C1549493;C3812891|All of the Time;Always - AcknowledgementCondition|always
Finding|Idea or Concept|SIMPLE_SEGMENT|7429,7435|false|false|false|C1549493;C3812891|All of the Time;Always - AcknowledgementCondition|always
Event|Event|SIMPLE_SEGMENT|7448,7452|false|false|false|||need
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7478,7482|false|false|false|C0339510|Vitelliform Macular Dystrophy|best
Event|Event|SIMPLE_SEGMENT|7478,7482|false|false|false|||best
Finding|Gene or Genome|SIMPLE_SEGMENT|7478,7482|false|false|false|C1826421;C5781213|BEST1 gene;BEST1 wt Allele|best
Procedure|Health Care Activity|SIMPLE_SEGMENT|7503,7511|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7512,7524|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|7512,7524|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|7512,7524|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

