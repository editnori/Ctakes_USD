 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|25,29
No|30,32
:|32,33
_|36,37
_|37,38
_|38,39
<EOL>|39,40
<EOL>|41,42
Admission|42,51
Date|52,56
:|56,57
_|59,60
_|60,61
_|61,62
Discharge|76,85
Date|86,90
:|90,91
_|94,95
_|95,96
_|96,97
<EOL>|97,98
<EOL>|99,100
Date|100,104
of|105,107
Birth|108,113
:|113,114
_|116,117
_|117,118
_|118,119
Sex|132,135
:|135,136
F|139,140
<EOL>|140,141
<EOL>|142,143
Service|143,150
:|150,151
MEDICINE|152,160
<EOL>|160,161
<EOL>|162,163
No|175,177
Known|178,183
Allergies|184,193
/|194,195
Adverse|196,203
Drug|204,208
Reactions|209,218
<EOL>|218,219
<EOL>|220,221
Attending|221,230
:|230,231
_|232,233
_|233,234
_|234,235
.|235,236
<EOL>|236,237
<EOL>|238,239
Atypical|256,264
chest|265,270
pain|271,275
<EOL>|275,276
<EOL>|277,278
Major|278,283
Surgical|284,292
or|293,295
Invasive|296,304
Procedure|305,314
:|314,315
<EOL>|315,316
Stess|316,321
Echo|322,326
<EOL>|326,327
<EOL>|327,328
<EOL>|329,330
_|358,359
_|359,360
_|360,361
y|362,363
/|363,364
o|364,365
woman|366,371
with|372,376
intermittent|377,389
chest|390,395
pain|396,400
past|401,405
several|406,413
months|414,420
.|420,421
<EOL>|422,423
Pain|423,427
is|428,430
located|431,438
on|439,441
left|442,446
posterior|447,456
shoulder|457,465
and|466,469
radiates|470,478
down|479,483
arm|484,487
<EOL>|488,489
to|489,491
fingers|492,499
where|500,505
it|506,508
turns|509,514
into|515,519
"|520,521
pins|521,525
-|525,526
n|526,527
-|527,528
needles|528,535
"|535,536
symptom|537,544
.|544,545
No|546,548
<EOL>|549,550
SOB|550,553
/|553,554
N|554,555
/|555,556
V|556,557
.|557,558
Patient|559,566
does|567,571
endorse|572,579
some|580,584
minimal|585,592
diaphoresis|593,604
and|605,608
gerd|609,613
<EOL>|614,615
like|615,619
symptoms|620,628
accompanying|629,641
it|642,644
.|644,645
Pain|646,650
has|651,654
been|655,659
controlled|660,670
with|671,675
<EOL>|676,677
tylenol|677,684
#|685,686
3|686,687
.|687,688
<EOL>|689,690
<EOL>|691,692
HTN|714,717
<EOL>|719,720
Asthma|720,726
<EOL>|728,729
Diverticulitis|729,743
several|744,751
years|752,757
ago|758,761
<EOL>|763,764
R|764,765
hip|766,769
replacement|770,781
in|782,784
_|785,786
_|786,787
_|787,788
<EOL>|790,791
<EOL>|791,792
<EOL>|793,794
:|808,809
<EOL>|809,810
_|810,811
_|811,812
_|812,813
<EOL>|813,814
:|828,829
<EOL>|829,830
Mother|830,836
:|836,837
_|838,839
_|839,840
_|840,841
,|841,842
HTN|843,846
<EOL>|848,849
Father|849,855
:|855,856
_|857,858
_|858,859
_|859,860
CA|861,863
<EOL>|865,866
Brother|866,873
:|873,874
CA|875,877
?|877,878
<EOL>|880,881
Brother|881,888
:|888,889
_|890,891
_|891,892
_|892,893
<EOL>|895,896
<EOL>|896,897
<EOL>|898,899
Physical|899,907
_|908,909
_|909,910
_|910,911
:|911,912
<EOL>|912,913
Vtals|913,918
:|918,919
T|920,921
:|921,922
97.6|923,927
BP|928,930
:|930,931
167|932,935
/|935,936
88|936,938
P|939,940
:|940,941
83|942,944
R|945,946
:|946,947
20|948,950
O2|951,953
:|953,954
99|955,957
%|957,958
2L|959,961
<EOL>|963,964
General|964,971
:|971,972
Alert|973,978
,|978,979
oriented|980,988
,|988,989
no|990,992
acute|993,998
distress|999,1007
<EOL>|1009,1010
HEENT|1010,1015
:|1015,1016
Sclera|1017,1023
anicteric|1024,1033
,|1033,1034
MMM|1035,1038
,|1038,1039
oropharynx|1040,1050
clear|1051,1056
<EOL>|1058,1059
Neck|1059,1063
:|1063,1064
supple|1065,1071
,|1071,1072
JVP|1073,1076
not|1077,1080
elevated|1081,1089
,|1089,1090
no|1091,1093
LAD|1094,1097
<EOL>|1099,1100
Lungs|1100,1105
:|1105,1106
Clear|1107,1112
to|1113,1115
auscultation|1116,1128
bilaterally|1129,1140
,|1140,1141
no|1142,1144
wheezes|1145,1152
,|1152,1153
rales|1154,1159
,|1159,1160
<EOL>|1161,1162
ronchi|1162,1168
<EOL>|1170,1171
CV|1171,1173
:|1173,1174
Regular|1175,1182
rate|1183,1187
and|1188,1191
rhythm|1192,1198
,|1198,1199
normal|1200,1206
S1|1207,1209
+|1210,1211
S2|1212,1214
,|1214,1215
no|1216,1218
murmurs|1219,1226
,|1226,1227
rubs|1228,1232
,|1232,1233
<EOL>|1234,1235
gallops|1235,1242
<EOL>|1244,1245
Abdomen|1245,1252
:|1252,1253
soft|1254,1258
,|1258,1259
non-tender|1260,1270
,|1270,1271
non-distended|1272,1285
,|1285,1286
bowel|1287,1292
sounds|1293,1299
present|1300,1307
,|1307,1308
<EOL>|1309,1310
no|1310,1312
rebound|1313,1320
tenderness|1321,1331
or|1332,1334
guarding|1335,1343
,|1343,1344
no|1345,1347
organomegaly|1348,1360
<EOL>|1362,1363
Ext|1363,1366
:|1366,1367
Warm|1368,1372
,|1372,1373
well|1374,1378
perfused|1379,1387
,|1387,1388
2|1389,1390
+|1390,1391
pulses|1392,1398
,|1398,1399
no|1400,1402
clubbing|1403,1411
,|1411,1412
cyanosis|1413,1421
or|1422,1424
<EOL>|1425,1426
edema|1426,1431
<EOL>|1433,1434
<EOL>|1434,1435
<EOL>|1436,1437
Pertinent|1437,1446
Results|1447,1454
:|1454,1455
<EOL>|1455,1456
_|1456,1457
_|1457,1458
_|1458,1459
03|1460,1462
:|1462,1463
20PM|1463,1467
BLOOD|1468,1473
WBC|1474,1477
-|1477,1478
6.2|1478,1481
RBC|1482,1485
-|1485,1486
4|1486,1487
.|1487,1488
51|1488,1490
Hgb|1491,1494
-|1494,1495
13.1|1495,1499
Hct|1500,1503
-|1503,1504
38.6|1504,1508
MCV|1509,1512
-|1512,1513
86|1513,1515
<EOL>|1516,1517
MCH|1517,1520
-|1520,1521
29.1|1521,1525
MCHC|1526,1530
-|1530,1531
33.9|1531,1535
RDW|1536,1539
-|1539,1540
15.4|1540,1544
Plt|1545,1548
_|1549,1550
_|1550,1551
_|1551,1552
<EOL>|1552,1553
_|1553,1554
_|1554,1555
_|1555,1556
07|1557,1559
:|1559,1560
15AM|1560,1564
BLOOD|1565,1570
WBC|1571,1574
-|1574,1575
6.0|1575,1578
RBC|1579,1582
-|1582,1583
4|1583,1584
.|1584,1585
91|1585,1587
Hgb|1588,1591
-|1591,1592
13.8|1592,1596
Hct|1597,1600
-|1600,1601
41.7|1601,1605
MCV|1606,1609
-|1609,1610
85|1610,1612
<EOL>|1613,1614
MCH|1614,1617
-|1617,1618
28.1|1618,1622
MCHC|1623,1627
-|1627,1628
33.0|1628,1632
RDW|1633,1636
-|1636,1637
15.1|1637,1641
Plt|1642,1645
_|1646,1647
_|1647,1648
_|1648,1649
<EOL>|1649,1650
_|1650,1651
_|1651,1652
_|1652,1653
07|1654,1656
:|1656,1657
50AM|1657,1661
BLOOD|1662,1667
WBC|1668,1671
-|1671,1672
5.2|1672,1675
RBC|1676,1679
-|1679,1680
4|1680,1681
.|1681,1682
67|1682,1684
Hgb|1685,1688
-|1688,1689
13.4|1689,1693
Hct|1694,1697
-|1697,1698
39.4|1698,1702
MCV|1703,1706
-|1706,1707
84|1707,1709
<EOL>|1710,1711
MCH|1711,1714
-|1714,1715
28.7|1715,1719
MCHC|1720,1724
-|1724,1725
34.1|1725,1729
RDW|1730,1733
-|1733,1734
15.2|1734,1738
Plt|1739,1742
_|1743,1744
_|1744,1745
_|1745,1746
<EOL>|1746,1747
_|1747,1748
_|1748,1749
_|1749,1750
03|1751,1753
:|1753,1754
20PM|1754,1758
BLOOD|1759,1764
Glucose|1765,1772
-|1772,1773
95|1773,1775
UreaN|1776,1781
-|1781,1782
21|1782,1784
*|1784,1785
Creat|1786,1791
-|1791,1792
0.8|1792,1795
Na|1796,1798
-|1798,1799
139|1799,1802
<EOL>|1803,1804
K|1804,1805
-|1805,1806
3.5|1806,1809
Cl|1810,1812
-|1812,1813
100|1813,1816
HCO3|1817,1821
-|1821,1822
30|1822,1824
AnGap|1825,1830
-|1830,1831
13|1831,1833
<EOL>|1833,1834
_|1834,1835
_|1835,1836
_|1836,1837
09|1838,1840
:|1840,1841
10PM|1841,1845
BLOOD|1846,1851
Glucose|1852,1859
-|1859,1860
120|1860,1863
*|1863,1864
UreaN|1865,1870
-|1870,1871
17|1871,1873
Creat|1874,1879
-|1879,1880
0.9|1880,1883
Na|1884,1886
-|1886,1887
137|1887,1890
<EOL>|1891,1892
K|1892,1893
-|1893,1894
3.3|1894,1897
Cl|1898,1900
-|1900,1901
99|1901,1903
HCO3|1904,1908
-|1908,1909
31|1909,1911
AnGap|1912,1917
-|1917,1918
10|1918,1920
<EOL>|1920,1921
_|1921,1922
_|1922,1923
_|1923,1924
07|1925,1927
:|1927,1928
15AM|1928,1932
BLOOD|1933,1938
Glucose|1939,1946
-|1946,1947
100|1947,1950
UreaN|1951,1956
-|1956,1957
15|1957,1959
Creat|1960,1965
-|1965,1966
0.8|1966,1969
Na|1970,1972
-|1972,1973
138|1973,1976
<EOL>|1977,1978
K|1978,1979
-|1979,1980
4.4|1980,1983
Cl|1984,1986
-|1986,1987
98|1987,1989
HCO3|1990,1994
-|1994,1995
35|1995,1997
*|1997,1998
AnGap|1999,2004
-|2004,2005
9|2005,2006
<EOL>|2006,2007
_|2007,2008
_|2008,2009
_|2009,2010
03|2011,2013
:|2013,2014
20PM|2014,2018
BLOOD|2019,2024
cTropnT|2025,2032
-|2032,2033
<|2033,2034
0|2034,2035
.|2035,2036
01|2036,2038
<EOL>|2038,2039
_|2039,2040
_|2040,2041
_|2041,2042
09|2043,2045
:|2045,2046
10PM|2046,2050
BLOOD|2051,2056
CK|2057,2059
-|2059,2060
MB|2060,2062
-|2062,2063
3|2063,2064
cTropnT|2065,2072
-|2072,2073
<|2073,2074
0|2074,2075
.|2075,2076
01|2076,2078
<EOL>|2078,2079
_|2079,2080
_|2080,2081
_|2081,2082
07|2083,2085
:|2085,2086
15AM|2086,2090
BLOOD|2091,2096
CK|2097,2099
-|2099,2100
MB|2100,2102
-|2102,2103
4|2103,2104
cTropnT|2105,2112
-|2112,2113
<|2113,2114
0.01|2114,2118
<EOL>|2118,2119
.|2119,2120
<EOL>|2120,2121
_|2121,2122
_|2122,2123
_|2123,2124
_|2125,2126
_|2126,2127
_|2127,2128
F|2129,2130
_|2132,2133
_|2133,2134
_|2134,2135
_|2137,2138
_|2138,2139
_|2139,2140
<EOL>|2141,2142
<EOL>|2143,2144
Cardiology|2144,2154
Report|2155,2161
Stress|2162,2168
Study|2169,2174
Date|2175,2179
of|2180,2182
_|2183,2184
_|2184,2185
_|2185,2186
<EOL>|2189,2190
<EOL>|2191,2192
<EOL>|2194,2195
EXERCISE|2195,2203
RESULTS|2204,2211
<EOL>|2212,2213
<EOL>|2213,2214
<EOL>|2215,2216
<EOL>|2218,2219
RESTING|2219,2226
DATA|2227,2231
<EOL>|2232,2233
EKG|2233,2236
:|2236,2237
SINUS|2239,2244
WITH|2245,2249
AEA|2250,2253
,|2253,2254
LBBB|2255,2259
<EOL>|2262,2263
HEART|2263,2268
RATE|2269,2273
:|2273,2274
68|2276,2278
BLOOD|2279,2284
PRESSURE|2285,2293
:|2293,2294
146|2296,2299
/|2299,2300
86|2300,2302
<EOL>|2303,2304
<EOL>|2306,2307
PROTOCOL|2307,2315
MODIFIED|2316,2324
_|2325,2326
_|2326,2327
_|2327,2328
-|2329,2330
TREAD|2331,2336
_|2336,2337
_|2337,2338
_|2338,2339
<EOL>|2340,2341
STAGE|2341,2346
TIME|2347,2351
SPEED|2352,2357
ELEVATION|2358,2367
HEART|2368,2373
BLOOD|2374,2379
RPP|2380,2383
<EOL>|2384,2385
(|2387,2388
MIN|2388,2391
)|2391,2392
(|2393,2394
MPH|2394,2397
)|2397,2398
(|2399,2400
%|2400,2401
)|2401,2402
RATE|2403,2407
PRESSURE|2408,2416
<EOL>|2419,2420
0|2420,2421
_|2422,2423
_|2423,2424
_|2424,2425
1.0|2426,2429
8|2430,2431
100|2432,2435
176|2436,2439
/|2439,2440
88|2440,2442
_|2443,2444
_|2444,2445
_|2445,2446
<EOL>|2447,2448
1|2448,2449
_|2450,2451
_|2451,2452
_|2452,2453
1.7|2454,2457
10|2458,2460
114|2461,2464
178|2465,2468
/|2468,2469
92|2469,2471
_|2472,2473
_|2473,2474
_|2474,2475
2.5|2476,2479
12|2480,2482
126|2483,2486
184|2487,2490
/|2490,2491
98|2491,2493
_|2494,2495
_|2495,2496
_|2496,2497
<EOL>|2498,2499
<EOL>|2501,2502
TOTAL|2502,2507
EXERCISE|2508,2516
TIME|2517,2521
:|2521,2522
9|2524,2525
%|2526,2527
MAX|2528,2531
HRT|2532,2535
RATE|2536,2540
ACHIEVED|2541,2549
:|2549,2550
83|2552,2554
<EOL>|2555,2556
<EOL>|2557,2558
SYMPTOMS|2558,2566
:|2566,2567
ATYPICAL|2568,2576
PEAK|2577,2581
INTENSITY|2582,2591
:|2591,2592
_|2593,2594
_|2594,2595
_|2595,2596
<EOL>|2597,2598
<EOL>|2599,2600
<EOL>|2602,2603
INTERPRETATION|2603,2617
:|2617,2618
_|2619,2620
_|2620,2621
_|2621,2622
yo|2623,2625
woman|2626,2631
was|2632,2635
referred|2636,2644
to|2645,2647
evaluate|2648,2656
an|2657,2659
atypical|2660,2668
<EOL>|2669,2670
<EOL>|2670,2671
chest|2671,2676
discomfort|2677,2687
.|2687,2688
The|2689,2692
patient|2693,2700
completed|2701,2710
9|2711,2712
minutes|2713,2720
of|2721,2723
a|2724,2725
Gervino|2726,2733
<EOL>|2734,2735
protocol|2735,2743
<EOL>|2744,2745
representing|2745,2757
a|2758,2759
fair|2760,2764
exercise|2765,2773
tolerance|2774,2783
for|2784,2787
her|2788,2791
age|2792,2795
;|2795,2796
~|2797,2798
_|2799,2800
_|2800,2801
_|2801,2802
METS|2803,2807
.|2807,2808
<EOL>|2809,2810
The|2810,2813
<EOL>|2814,2815
exercise|2815,2823
test|2824,2828
was|2829,2832
stopped|2833,2840
at|2841,2843
the|2844,2847
patient|2848,2855
's|2855,2857
request|2858,2865
secondary|2866,2875
to|2876,2878
<EOL>|2879,2880
fatigue|2880,2887
.|2887,2888
<EOL>|2889,2890
During|2890,2896
exercise|2897,2905
,|2905,2906
the|2907,2910
patient|2911,2918
reported|2919,2927
a|2928,2929
non-progressive|2930,2945
,|2945,2946
<EOL>|2947,2948
isolated|2948,2956
upper|2957,2962
<EOL>|2963,2964
left|2964,2968
-|2968,2969
sided|2969,2974
chest|2975,2980
discomfort|2981,2991
;|2991,2992
_|2993,2994
_|2994,2995
_|2995,2996
.|2996,2997
The|2998,3001
area|3002,3006
of|3007,3009
discomfort|3010,3020
was|3021,3024
<EOL>|3025,3026
reportedly|3026,3036
<EOL>|3037,3038
tender|3038,3044
to|3045,3047
palpation|3048,3057
.|3057,3058
This|3059,3063
discomfort|3064,3074
resolved|3075,3083
with|3084,3088
rest|3089,3093
and|3094,3097
was|3098,3101
<EOL>|3102,3103
absent|3103,3109
<EOL>|3110,3111
2.5|3111,3114
minutes|3115,3122
post-exercise|3123,3136
.|3136,3137
In|3138,3140
the|3141,3144
presence|3145,3153
of|3154,3156
the|3157,3160
LBBB|3161,3165
,|3165,3166
the|3167,3170
ST|3171,3173
<EOL>|3174,3175
segments|3175,3183
<EOL>|3184,3185
are|3185,3188
uninterpretable|3189,3204
for|3205,3208
ischemia|3209,3217
.|3217,3218
The|3219,3222
rhythm|3223,3229
was|3230,3233
sinus|3234,3239
with|3240,3244
<EOL>|3245,3246
frequent|3246,3254
<EOL>|3255,3256
isolated|3256,3264
APDs|3265,3269
and|3270,3273
occasional|3274,3284
atrial|3285,3291
couplets|3292,3300
and|3301,3304
atrial|3305,3311
<EOL>|3312,3313
triplets|3313,3321
.|3321,3322
<EOL>|3323,3324
Resting|3324,3331
mild|3332,3336
systolic|3337,3345
hypertension|3346,3358
with|3359,3363
normal|3364,3370
blood|3371,3376
pressure|3377,3385
<EOL>|3386,3387
response|3387,3395
<EOL>|3396,3397
to|3397,3399
exercise|3400,3408
.|3408,3409
The|3410,3413
heart|3414,3419
rate|3420,3424
response|3425,3433
to|3434,3436
exercise|3437,3445
was|3446,3449
mildly|3450,3456
<EOL>|3457,3458
blunted|3458,3465
.|3465,3466
<EOL>|3467,3468
<EOL>|3470,3471
IMPRESSION|3471,3481
:|3481,3482
Fair|3483,3487
exercise|3488,3496
tolerance|3497,3506
.|3506,3507
No|3508,3510
anginal|3511,3518
symptoms|3519,3527
with|3528,3532
<EOL>|3533,3534
uninterpretable|3534,3549
ECG|3550,3553
to|3554,3556
achieved|3557,3565
workload|3566,3574
.|3574,3575
Resting|3576,3583
mild|3584,3588
systolic|3589,3597
<EOL>|3598,3599
hypertension|3599,3611
with|3612,3616
appropriate|3617,3628
blood|3629,3634
pressure|3635,3643
response|3644,3652
to|3653,3655
<EOL>|3656,3657
exercise|3657,3665
.|3665,3666
<EOL>|3667,3668
Suboptimal|3668,3678
study|3679,3684
-|3685,3686
target|3687,3693
heart|3694,3699
rate|3700,3704
not|3705,3708
achieved|3709,3717
.|3717,3718
<EOL>|3719,3720
<EOL>|3721,3722
SIGNED|3722,3728
:|3728,3729
_|3731,3732
_|3732,3733
_|3733,3734
<EOL>|3735,3736
<EOL>|3737,3738
<EOL>|3738,3739
<EOL>|3740,3741
_|3764,3765
_|3765,3766
_|3766,3767
_|3768,3769
_|3769,3770
_|3770,3771
with|3772,3776
several|3777,3784
month|3785,3790
history|3791,3798
of|3799,3801
left|3802,3806
sided|3807,3812
arm|3813,3816
and|3817,3820
chest|3821,3826
<EOL>|3827,3828
wall|3828,3832
pain|3833,3837
in|3838,3840
the|3841,3844
setting|3845,3852
of|3853,3855
LBBB|3856,3860
presenting|3861,3871
for|3872,3875
_|3876,3877
_|3877,3878
_|3878,3879
.|3879,3880
<EOL>|3882,3883
.|3883,3884
<EOL>|3886,3887
.|3887,3888
<EOL>|3890,3891
#|3891,3892
Chest|3893,3898
Pain|3899,3903
:|3903,3904
The|3904,3907
patient|3908,3915
's|3915,3917
symptoms|3918,3926
were|3927,3931
not|3932,3935
typically|3936,3945
anginal|3946,3953
<EOL>|3954,3955
in|3955,3957
nature|3958,3964
to|3965,3967
suggest|3968,3975
ACS|3976,3979
.|3979,3980
However|3981,3988
she|3989,3992
does|3993,3997
have|3998,4002
several|4003,4010
cardiac|4011,4018
<EOL>|4019,4020
risk|4020,4024
factors|4025,4032
and|4033,4036
a|4037,4038
LBBB|4039,4043
,|4043,4044
so|4045,4047
physicians|4049,4059
could|4060,4065
not|4067,4070
r|4071,4072
/|4072,4073
oMI|4073,4076
with|4077,4081
<EOL>|4082,4083
EKG|4083,4086
alone|4087,4092
.|4092,4093
Trop|4094,4098
.|4098,4099
results|4100,4107
were|4108,4112
negative|4113,4121
x3|4122,4124
.|4124,4125
Stress|4126,4132
Echo|4133,4137
revealed|4138,4146
<EOL>|4147,4148
new|4148,4151
regional|4152,4160
dysfunction|4161,4172
with|4173,4177
hypokinesis|4178,4189
of|4190,4192
the|4193,4196
inferior|4197,4205
and|4206,4209
<EOL>|4210,4211
inferolateral|4211,4224
walls|4225,4230
consistent|4231,4241
with|4242,4246
single|4247,4253
vessel|4254,4260
disease|4261,4268
in|4269,4271
the|4272,4275
<EOL>|4276,4277
PDA|4277,4280
distribution|4281,4293
.|4293,4294
A|4295,4296
cardiology|4297,4307
consult|4308,4315
was|4316,4319
obtained|4320,4328
and|4329,4332
they|4333,4337
<EOL>|4338,4339
felt|4339,4343
she|4344,4347
could|4348,4353
be|4354,4356
managed|4357,4364
medically|4365,4374
.|4374,4375
Patient|4376,4383
was|4384,4387
already|4388,4395
on|4396,4398
an|4399,4401
<EOL>|4402,4403
aspirin|4403,4410
,|4410,4411
and|4412,4415
a|4416,4417
statin|4418,4424
.|4424,4425
Given|4426,4431
history|4432,4439
to|4440,4442
suggest|4443,4450
asthma|4451,4457
B|4458,4459
-|4459,4460
blocker|4460,4467
<EOL>|4468,4469
was|4469,4472
contraindicated|4473,4488
.|4488,4489
She|4490,4493
was|4494,4497
discharged|4498,4508
on|4509,4511
120|4512,4515
mg|4516,4518
extended|4519,4527
<EOL>|4528,4529
release|4529,4536
diltiazem|4537,4546
with|4547,4551
instructions|4552,4564
to|4565,4567
follow|4568,4574
up|4575,4577
in|4578,4580
cardiology|4581,4591
<EOL>|4592,4593
and|4593,4596
with|4597,4601
her|4602,4605
PCP|4606,4609
.|4609,4610
<EOL>|4611,4612
.|4612,4613
<EOL>|4613,4614
#|4614,4615
Supraventricular|4616,4632
tachycardia|4633,4644
:|4644,4645
The|4646,4649
patient|4650,4657
had|4658,4661
multiple|4662,4670
runs|4671,4675
of|4676,4678
<EOL>|4679,4680
SVT|4680,4683
that|4684,4688
was|4689,4692
likley|4693,4699
MAT|4700,4703
in|4704,4706
the|4707,4710
setting|4711,4718
of|4719,4721
severe|4722,4728
obstructive|4729,4740
<EOL>|4741,4742
lung|4742,4746
disease|4747,4754
and|4755,4758
chronic|4759,4766
theophylline|4767,4779
use|4780,4783
.|4783,4784
Cardiology|4785,4795
<EOL>|4796,4797
reccomended|4797,4808
that|4809,4813
we|4814,4816
discontinue|4817,4828
her|4829,4832
theophylline|4833,4845
.|4845,4846
We|4847,4849
spoke|4850,4855
with|4856,4860
<EOL>|4861,4862
her|4862,4865
pulmonologist|4866,4879
who|4880,4883
agreed|4884,4890
this|4891,4895
would|4896,4901
be|4902,4904
the|4905,4908
best|4909,4913
course|4914,4920
of|4921,4923
<EOL>|4924,4925
action|4925,4931
for|4932,4935
her|4936,4939
.|4939,4940
She|4941,4944
was|4945,4948
discharged|4949,4959
with|4960,4964
instructions|4965,4977
to|4978,4980
<EOL>|4981,4982
discontinue|4982,4993
use|4994,4997
of|4998,5000
theophylline|5001,5013
and|5014,5017
follow|5018,5024
up|5025,5027
with|5028,5032
her|5033,5036
<EOL>|5037,5038
pulmonologist|5038,5051
and|5052,5055
cardiology|5056,5066
.|5066,5067
<EOL>|5067,5068
<EOL>|5068,5069
<EOL>|5070,5071
Medications|5071,5082
on|5083,5085
Admission|5086,5095
:|5095,5096
<EOL>|5096,5097
Tylenol|5097,5104
_|5105,5106
_|5106,5107
_|5107,5108
Q4h|5109,5112
PRN|5113,5116
pain|5117,5121
<EOL>|5123,5124
Albuterol|5124,5133
Sulfate|5134,5141
2|5142,5143
puffs|5144,5149
q4|5150,5152
-|5152,5153
6h|5153,5155
PRN|5156,5159
SOB|5160,5163
<EOL>|5165,5166
Fluticasone|5166,5177
50|5178,5180
mcg|5181,5184
spray|5185,5190
/|5190,5191
suspension|5191,5201
2|5202,5203
whiffs|5204,5210
PRN|5211,5214
allergies|5215,5224
<EOL>|5226,5227
Adviar|5227,5233
500|5234,5237
/|5237,5238
50|5238,5240
1|5241,5242
INH|5243,5246
BID|5247,5250
<EOL>|5252,5253
HCTZ|5253,5257
50mg|5258,5262
One|5263,5266
PO|5267,5269
daily|5270,5275
<EOL>|5277,5278
Singulari|5278,5287
10mg|5288,5292
tablet|5293,5299
One|5300,5303
PO|5304,5306
QD|5307,5309
<EOL>|5311,5312
omeprazole|5312,5322
20mg|5323,5327
1|5328,5329
PO|5330,5332
QD|5333,5335
<EOL>|5337,5338
simvastatin|5338,5349
20mg|5350,5354
1|5355,5356
PO|5357,5359
QD|5360,5362
<EOL>|5364,5365
theophylline|5365,5377
200mg|5378,5383
sustained|5384,5393
release|5394,5401
one|5402,5405
PO|5406,5408
TID|5409,5412
<EOL>|5414,5415
spiriva|5415,5422
18|5423,5425
mcg|5426,5429
w|5430,5431
/|5431,5432
inhalation|5433,5443
<EOL>|5445,5446
ASA|5446,5449
81mg|5450,5454
<EOL>|5456,5457
Calcium|5457,5464
sig|5465,5468
unknown|5469,5476
<EOL>|5478,5479
Cod|5479,5482
liver|5483,5488
oil|5489,5492
Sig|5493,5496
unk|5497,5500
<EOL>|5502,5503
Multivitamin|5503,5515
<EOL>|5517,5518
<EOL>|5518,5519
<EOL>|5520,5521
Discharge|5521,5530
Medications|5531,5542
:|5542,5543
<EOL>|5543,5544
1.|5544,5546
acetaminophen|5547,5560
325|5561,5564
mg|5565,5567
Tablet|5568,5574
Sig|5575,5578
:|5578,5579
One|5580,5583
(|5584,5585
1|5585,5586
)|5586,5587
Tablet|5588,5594
PO|5595,5597
Q4H|5598,5601
(|5602,5603
every|5603,5608
<EOL>|5609,5610
4|5610,5611
hours|5612,5617
)|5617,5618
as|5619,5621
needed|5622,5628
for|5629,5632
pain|5633,5637
.|5637,5638
<EOL>|5640,5641
2.|5641,5643
albuterol|5644,5653
sulfate|5654,5661
90|5662,5664
mcg|5665,5668
/|5668,5669
Actuation|5669,5678
HFA|5679,5682
Aerosol|5683,5690
Inhaler|5691,5698
Sig|5699,5702
:|5702,5703
<EOL>|5704,5705
Two|5705,5708
(|5709,5710
2|5710,5711
)|5711,5712
Puff|5713,5717
Inhalation|5718,5728
Q6H|5729,5732
(|5733,5734
every|5734,5739
6|5740,5741
hours|5742,5747
)|5747,5748
as|5749,5751
needed|5752,5758
for|5759,5762
SOB|5763,5766
<EOL>|5767,5768
wheeze|5768,5774
.|5774,5775
<EOL>|5777,5778
3.|5778,5780
fluticasone|5781,5792
-|5792,5793
salmeterol|5793,5803
500|5804,5807
-|5807,5808
50|5808,5810
mcg|5811,5814
/|5814,5815
dose|5815,5819
Disk|5820,5824
with|5825,5829
Device|5830,5836
Sig|5837,5840
:|5840,5841
<EOL>|5842,5843
One|5843,5846
(|5847,5848
1|5848,5849
)|5849,5850
Disk|5851,5855
with|5856,5860
Device|5861,5867
Inhalation|5868,5878
BID|5879,5882
(|5883,5884
2|5884,5885
times|5886,5891
a|5892,5893
day|5894,5897
)|5897,5898
.|5898,5899
<EOL>|5901,5902
4.|5902,5904
fluticasone|5905,5916
50|5917,5919
mcg|5920,5923
/|5923,5924
Actuation|5924,5933
Spray|5934,5939
,|5939,5940
Suspension|5941,5951
Sig|5952,5955
:|5955,5956
_|5957,5958
_|5958,5959
_|5959,5960
<EOL>|5962,5963
Nasal|5963,5968
once|5969,5973
a|5974,5975
day|5976,5979
as|5980,5982
needed|5983,5989
for|5990,5993
allergy|5994,6001
symptoms|6002,6010
.|6010,6011
<EOL>|6013,6014
5.|6014,6016
hydrochlorothiazide|6017,6036
50|6037,6039
mg|6040,6042
Tablet|6043,6049
Sig|6050,6053
:|6053,6054
One|6055,6058
(|6059,6060
1|6060,6061
)|6061,6062
Tablet|6063,6069
PO|6070,6072
once|6073,6077
<EOL>|6078,6079
a|6079,6080
day|6081,6084
.|6084,6085
<EOL>|6087,6088
6.|6088,6090
omeprazole|6091,6101
20|6102,6104
mg|6105,6107
Capsule|6108,6115
,|6115,6116
Delayed|6117,6124
Release|6125,6132
(|6132,6133
E.C|6133,6136
.|6136,6137
)|6137,6138
Sig|6139,6142
:|6142,6143
One|6144,6147
(|6148,6149
1|6149,6150
)|6150,6151
<EOL>|6152,6153
Capsule|6153,6160
,|6160,6161
Delayed|6162,6169
Release|6170,6177
(|6177,6178
E.C|6178,6181
.|6181,6182
)|6182,6183
PO|6184,6186
DAILY|6187,6192
(|6193,6194
Daily|6194,6199
)|6199,6200
.|6200,6201
<EOL>|6203,6204
7.|6204,6206
simvastatin|6207,6218
20|6219,6221
mg|6222,6224
Tablet|6225,6231
Sig|6232,6235
:|6235,6236
One|6237,6240
(|6241,6242
1|6242,6243
)|6243,6244
Tablet|6245,6251
PO|6252,6254
once|6255,6259
a|6260,6261
day|6262,6265
.|6265,6266
<EOL>|6268,6269
8.|6269,6271
tiotropium|6272,6282
bromide|6283,6290
18|6291,6293
mcg|6294,6297
Capsule|6298,6305
,|6305,6306
w|6307,6308
/|6308,6309
Inhalation|6309,6319
Device|6320,6326
Sig|6327,6330
:|6330,6331
<EOL>|6332,6333
One|6333,6336
(|6337,6338
1|6338,6339
)|6339,6340
Cap|6341,6344
Inhalation|6345,6355
DAILY|6356,6361
(|6362,6363
Daily|6363,6368
)|6368,6369
.|6369,6370
<EOL>|6372,6373
9.|6373,6375
aspirin|6376,6383
81|6384,6386
mg|6387,6389
Tablet|6390,6396
Sig|6397,6400
:|6400,6401
One|6402,6405
(|6406,6407
1|6407,6408
)|6408,6409
Tablet|6410,6416
PO|6417,6419
once|6420,6424
a|6425,6426
day|6427,6430
.|6430,6431
<EOL>|6433,6434
10.|6434,6437
multivitamin|6438,6450
Tablet|6455,6461
Sig|6462,6465
:|6465,6466
One|6467,6470
(|6471,6472
1|6472,6473
)|6473,6474
Tablet|6475,6481
PO|6482,6484
DAILY|6485,6490
<EOL>|6491,6492
(|6492,6493
Daily|6493,6498
)|6498,6499
.|6499,6500
<EOL>|6502,6503
11.|6503,6506
diltiazem|6507,6516
HCl|6517,6520
120|6521,6524
mg|6525,6527
Tablet|6528,6534
Sustained|6535,6544
Release|6545,6552
24|6553,6555
hr|6556,6558
Sig|6559,6562
:|6562,6563
One|6564,6567
<EOL>|6568,6569
(|6569,6570
1|6570,6571
)|6571,6572
Tablet|6573,6579
Sustained|6580,6589
Release|6590,6597
24|6598,6600
hr|6601,6603
PO|6604,6606
once|6607,6611
a|6612,6613
day|6614,6617
.|6617,6618
<EOL>|6618,6619
Disp|6619,6623
:|6623,6624
*|6624,6625
30|6625,6627
Tablet|6628,6634
Sustained|6635,6644
Release|6645,6652
24|6653,6655
hr|6656,6658
(|6658,6659
s|6659,6660
)|6660,6661
*|6661,6662
Refills|6663,6670
:|6670,6671
*|6671,6672
2|6672,6673
*|6673,6674
<EOL>|6674,6675
12.|6675,6678
nitroglycerin|6679,6692
0.3|6693,6696
mg|6697,6699
Tablet|6700,6706
,|6706,6707
Sublingual|6708,6718
Sig|6719,6722
:|6722,6723
One|6724,6727
(|6728,6729
1|6729,6730
)|6730,6731
<EOL>|6733,6734
Sublingual|6734,6744
every|6745,6750
5|6751,6752
min|6753,6756
as|6757,6759
needed|6760,6766
for|6767,6770
chest|6771,6776
pain|6777,6781
:|6781,6782
take|6783,6787
one|6788,6791
at|6792,6794
<EOL>|6795,6796
onset|6796,6801
of|6802,6804
chest|6805,6810
pain|6811,6815
.|6815,6816
_|6817,6818
_|6818,6819
_|6819,6820
repeat|6821,6827
every|6828,6833
5|6834,6835
min|6836,6839
x3|6840,6842
with|6843,6847
continued|6848,6857
<EOL>|6858,6859
chest|6859,6864
pain|6865,6869
.|6869,6870
Call|6871,6875
PCP|6876,6879
if|6880,6882
chest|6883,6888
pain|6889,6893
persists|6894,6902
.|6902,6903
<EOL>|6903,6904
Disp|6904,6908
:|6908,6909
*|6909,6910
30|6910,6912
tabs|6913,6917
*|6917,6918
Refills|6919,6926
:|6926,6927
*|6927,6928
0|6928,6929
*|6929,6930
<EOL>|6930,6931
<EOL>|6931,6932
<EOL>|6933,6934
Discharge|6934,6943
Disposition|6944,6955
:|6955,6956
<EOL>|6956,6957
Home|6957,6961
<EOL>|6961,6962
<EOL>|6963,6964
Discharge|6964,6973
Diagnosis|6974,6983
:|6983,6984
<EOL>|6984,6985
Coronary|6985,6993
Artery|6994,7000
Disease|7001,7008
<EOL>|7008,7009
<EOL>|7009,7010
<EOL>|7011,7012
Mental|7033,7039
Status|7040,7046
:|7046,7047
Clear|7048,7053
and|7054,7057
coherent|7058,7066
.|7066,7067
<EOL>|7067,7068
Level|7068,7073
of|7074,7076
Consciousness|7077,7090
:|7090,7091
Alert|7092,7097
and|7098,7101
interactive|7102,7113
.|7113,7114
<EOL>|7114,7115
Activity|7115,7123
Status|7124,7130
:|7130,7131
Ambulatory|7132,7142
-|7143,7144
Independent|7145,7156
.|7156,7157
<EOL>|7157,7158
<EOL>|7158,7159
<EOL>|7160,7161
You|7185,7188
were|7189,7193
admitted|7194,7202
to|7203,7205
_|7206,7207
_|7207,7208
_|7208,7209
because|7210,7217
you|7218,7221
had|7222,7225
back|7226,7230
and|7231,7234
arm|7235,7238
pain|7239,7243
<EOL>|7244,7245
that|7245,7249
was|7250,7253
worrisome|7254,7263
for|7264,7267
heart|7268,7273
disease|7274,7281
.|7281,7282
A|7283,7284
strees|7285,7291
test|7292,7296
found|7297,7302
that|7303,7307
<EOL>|7308,7309
you|7309,7312
have|7313,7317
coronary|7318,7326
artery|7327,7333
disease|7334,7341
.|7341,7342
You|7343,7346
were|7347,7351
started|7352,7359
on|7360,7362
a|7363,7364
new|7365,7368
<EOL>|7369,7370
blood|7370,7375
pressure|7376,7384
medication|7385,7395
and|7396,7399
tolerated|7400,7409
this|7410,7414
well|7415,7419
.|7419,7420
You|7421,7424
should|7425,7431
<EOL>|7432,7433
keep|7433,7437
all|7438,7441
of|7442,7444
you|7445,7448
follow|7449,7455
up|7456,7458
appointments|7459,7471
as|7472,7474
listed|7475,7481
below|7482,7487
.|7487,7488
<EOL>|7489,7490
.|7490,7491
<EOL>|7491,7492
While|7492,7497
you|7498,7501
were|7502,7506
here|7507,7511
we|7512,7514
made|7515,7519
the|7520,7523
following|7524,7533
changes|7534,7541
to|7542,7544
your|7545,7549
<EOL>|7550,7551
.|7564,7565
<EOL>|7565,7566
We|7566,7568
STARTED|7569,7576
you|7577,7580
on|7581,7583
Diltiazem|7584,7593
120mg|7594,7599
once|7600,7604
a|7605,7606
day|7607,7610
<EOL>|7610,7611
.|7611,7612
<EOL>|7612,7613
We|7613,7615
STOPPED|7616,7623
_|7624,7625
_|7625,7626
_|7626,7627
theophylline|7628,7640
<EOL>|7640,7641
.|7641,7642
<EOL>|7642,7643
We|7643,7645
STARTED|7646,7653
nitroglycerine|7654,7668
to|7669,7671
take|7672,7676
when|7677,7681
you|7682,7685
have|7686,7690
chest|7691,7696
pain|7697,7701
<EOL>|7701,7702
.|7702,7703
<EOL>|7703,7704
YOU|7704,7707
NEED|7708,7712
TO|7713,7715
STOP|7716,7720
SMOKING|7721,7728
.|7728,7729
IT|7730,7732
WILL|7733,7737
KILL|7738,7742
YOU|7743,7746
.|7746,7747
<EOL>|7747,7748
<EOL>|7749,7750
Followup|7750,7758
Instructions|7759,7771
:|7771,7772
<EOL>|7772,7773
_|7773,7774
_|7774,7775
_|7775,7776
<EOL>|7776,7777

