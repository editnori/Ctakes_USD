CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Pharmaceutical Preparations|Drug|false|false||MEDICINEnull|Medicine|Title|false|false||MEDICINEnull|Dyes|Drug|false|false||Dyenull|Iodine, Homeopathic preparation|Drug|false|false||Iodine
null|iodine|Drug|false|false||Iodine
null|iodine|Drug|false|false||Iodine
null|iodine|Drug|false|false||Iodinenull|Containing (qualifier value)|Finding|false|false||Containingnull|Contain (action)|Event|false|false||Containingnull|Contrast Media|Drug|false|false|C1254021;C0162867|Contrast Medianull|Contrast Media|Drug|false|false||Contrastnull|Contrast|Modifier|false|false||Contrastnull|Communications Media|Finding|false|false|C1254021;C0162867|Media
null|PAMS Media|Finding|false|false|C1254021;C0162867|Medianull|Tunica Media|Anatomy|false|false|C0009924;C0524222;C0677540;C0009458|Media
null|Media layer|Anatomy|false|false|C0009924;C0524222;C0677540;C0009458|Medianull|oxycodone|Drug|false|false||Oxycodone
null|oxycodone|Drug|false|false||Oxycodonenull|Oxycodone measurement|Procedure|false|false|C1254021;C0162867|Oxycodonenull|cilostazol|Drug|false|false||cilostazol
null|cilostazol|Drug|false|false||cilostazolnull|varenicline|Drug|false|false||Varenicline
null|varenicline|Drug|false|false||Vareniclinenull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|null|Finding|false|false||Dyspnea
null|Dyspnea|Finding|false|false||Dyspneanull|Atrial Fibrillation|Disorder|false|false|C0018792|Atrial Fibrillationnull|null|Attribute|false|false|C0018792|Atrial Fibrillationnull|Atrial Fibrillation by ECG Finding|Lab|false|false|C0018792|Atrial Fibrillationnull|Heart Atrium|Anatomy|false|false|C0344434;C0004238;C2926591;C0232197|Atrialnull|Fibrillation|Disorder|false|false|C0018792|Fibrillationnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|Hypertensive disease|Disorder|false|false||htnnull|Atrial Fibrillation|Disorder|false|false||afibnull|Atrial Fibrillation by ECG Finding|Lab|false|false||afibnull|null|Finding|false|false||dyspnea
null|Dyspnea|Finding|false|false||dyspneanull|Current (present time)|Time|false|false||currentlynull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|Atrial Fibrillation|Disorder|false|false||Afibnull|Atrial Fibrillation by ECG Finding|Lab|false|false||Afibnull|Rapid Virologic Response|Finding|false|false||RVR
null|NR1D2 wt Allele|Finding|false|false||RVR
null|NR1D2 gene|Finding|false|false||RVRnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|Flare|Finding|false|false||flare
null|Exacerbation of cGVHD|Finding|false|false||flarenull|prednisone|Drug|false|false||prednisone
null|prednisone|Drug|false|false||prednisone
null|prednisone|Drug|false|false||prednisonenull|null|Procedure|false|false||tapernull|Current (present time)|Time|false|false||currentlynull|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED|Drug|false|false||azithromycin
null|azithromycin|Drug|false|false||azithromycin
null|azithromycin|Drug|false|false||azithromycinnull|Initially|Time|false|false||initiallynull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|Rest Dyspnea|Finding|false|false||dyspnea at restnull|null|Finding|false|false||dyspnea
null|Dyspnea|Finding|false|false||dyspneanull|At rest (qualifier value)|Finding|false|false||at restnull|REST protein, human|Drug|false|false||rest
null|REST protein, human|Drug|false|false||restnull|REST gene|Finding|false|false||rest
null|site-specific telomere resolvase activity|Finding|false|false||rest
null|Rest|Finding|false|false||restnull|Exertion|Finding|false|false||exertionnull|Inhaler|Device|false|false||inhalersnull|Dyspnea|Finding|false|false||SOBnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Consistent with|Finding|false|false||consistent withnull|Compatible|Modifier|false|false||consistent withnull|Consistent with|Finding|false|false||consistentnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|Clinic|Device|false|false||clinic
null|Ambulatory Care Facilities|Device|false|false||clinicnull|Clinic|Entity|false|false||clinic
null|Ambulatory Care Facilities|Entity|false|false||clinicnull|Patient location type - Clinic|Modifier|false|false||clinic
null|Person location type - Clinic|Modifier|false|false||clinicnull|Atrial Fibrillation|Disorder|false|false||Afibnull|Atrial Fibrillation by ECG Finding|Lab|false|false||Afibnull|Rapid Virologic Response|Finding|false|false||RVR
null|NR1D2 wt Allele|Finding|false|false||RVR
null|NR1D2 gene|Finding|false|false||RVRnull|Amount type - Rate|Finding|false|false||ratenull|Rating (action)|Event|false|false||ratenull|Rate|LabModifier|false|false||ratenull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Atrial Fibrillation|Disorder|false|false||afibnull|Atrial Fibrillation by ECG Finding|Lab|false|false||afibnull|Persistent|Time|false|false||persistentnull|Dyspnea|Finding|false|false||SOBnull|Atrial Fibrillation|Disorder|false|false||afibnull|Atrial Fibrillation by ECG Finding|Lab|false|false||afibnull|Rapid Virologic Response|Finding|false|false||RVR
null|NR1D2 wt Allele|Finding|false|false||RVR
null|NR1D2 gene|Finding|false|false||RVRnull|Compliance behavior|Finding|false|false||compliantnull|Compliant (qualifier value)|Modifier|false|false||compliantnull|Nebulizer solution|Drug|false|false||nebsnull|Steroid [EPC]|Drug|false|false||steroid
null|Steroids|Drug|false|false||steroid
null|Steroids|Drug|false|false||steroidnull|GDC Regimen Terminology|Finding|false|false||regimennull|Treatment Protocols|Procedure|false|false||regimennull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|sleeping upright or using specific number of extra pillows (orthopnea)|Finding|false|false||orthopnea
null|Orthopnea|Finding|false|false||orthopneanull|Recent|Time|false|false||recentnull|travel|Finding|true|false||travelnull|travel charge|Procedure|true|false||travelnull|Operative Surgical Procedures|Procedure|false|false||surgeriesnull|Episode of|Time|false|false||episode ofnull|Episode of|Time|false|false||episodenull|Chest tightness|Finding|false|false|C1527391;C0817096|chest tightnessnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0232292;C0741025|chest
null|Anterior thoracic region|Anatomy|false|false|C0232292;C0741025|chestnull|Tightness sensation quality|Modifier|false|false||tightnessnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|Fever|Finding|true|false||feversnull|Coughing|Finding|true|false||coughingnull|Production Processing ID|Finding|false|false||productionnull|production|Event|false|false||productionnull|Specimen Type - Sputum|Finding|false|false||sputum
null|null|Finding|false|false||sputum
null|Sputum|Finding|false|false||sputumnull|Asthma|Disorder|false|false||ASTHMAnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|Atypical chest pain|Finding|false|false|C1527391;C0817096|ATYPICAL CHEST PAINnull|atypia morphology|Finding|false|false|C1527391;C0817096|ATYPICALnull|Atypical|Modifier|false|false||ATYPICALnull|Chest Pain|Finding|false|false|C1527391;C0817096|CHEST PAINnull|null|Attribute|false|false|C1527391;C0817096|CHEST PAINnull|Chest problem|Finding|false|false|C1527391;C0817096|CHESTnull|Chest|Anatomy|false|false|C0741025;C0008031;C1549543;C0030193;C0741302;C2598155;C0262384;C2926613|CHEST
null|Anterior thoracic region|Anatomy|false|false|C0741025;C0008031;C1549543;C0030193;C0741302;C2598155;C0262384;C2926613|CHESTnull|Administration Method - Pain|Finding|false|false|C1527391;C0817096|PAIN
null|Pain|Finding|false|false|C1527391;C0817096|PAINnull|null|Attribute|false|false|C1527391;C0817096|PAINnull|Cervical radiculitis|Disorder|false|false|C0027530|CERVICAL RADICULITISnull|Neck|Anatomy|false|false|C0034544;C0263884|CERVICALnull|Cervical|Modifier|false|false||CERVICALnull|Radiculitis|Disorder|false|false|C0027530|RADICULITISnull|Cervical spondylosis without myelopathy|Disorder|false|false|C0027530|CERVICAL SPONDYLOSIS
null|Cervical spondylosis|Disorder|false|false|C0027530|CERVICAL SPONDYLOSISnull|Neck|Anatomy|false|false|C0038019;C0158241;C1384641|CERVICALnull|Cervical|Modifier|false|false||CERVICALnull|Spondylosis|Disorder|false|false|C0027530|SPONDYLOSISnull|Coronary Artery Disease|Disorder|false|false|C0226004;C0003842;C0205042;C0018787|CORONARY ARTERY DISEASE
null|Coronary Arteriosclerosis|Disorder|false|false|C0226004;C0003842;C0205042;C0018787|CORONARY ARTERY DISEASEnull|Coronary artery|Anatomy|false|false|C1956346;C0010054;C0012634;C0852949|CORONARY ARTERYnull|Heart|Anatomy|false|false|C0852949;C0012634;C1956346;C0010054|CORONARYnull|Coronary|Modifier|false|false||CORONARYnull|Arteriopathic disease|Disorder|false|false|C0018787;C0205042;C0226004;C0003842|ARTERY DISEASEnull|Arterial system|Anatomy|false|false|C1956346;C0010054;C0012634;C0852949|ARTERY
null|Arteries|Anatomy|false|false|C1956346;C0010054;C0012634;C0852949|ARTERYnull|Disease|Disorder|false|false|C0018787;C0205042;C0226004;C0003842|DISEASEnull|Headache|Finding|false|false||HEADACHEnull|Prosthetic arthroplasty of hip (procedure)|Procedure|false|false|C0022122;C0228391;C0019552;C4299095|HIP REPLACEMENTnull|heme iron polypeptide|Drug|false|false|C0022122;C0228391;C0019552;C4299095|HIP
null|ST13 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|HIP
null|ST13 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|HIP
null|RPL29 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|HIP
null|RPL29 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|HIP
null|HHIP protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|HIP
null|HHIP protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|HIP
null|heme iron polypeptide|Drug|false|false|C0022122;C0228391;C0019552;C4299095|HIPnull|RPL29 wt Allele|Finding|false|false|C0022122;C0228391;C0019552;C4299095|HIP
null|REG3A gene|Finding|false|false|C0022122;C0228391;C0019552;C4299095|HIP
null|RPL29 gene|Finding|false|false|C0022122;C0228391;C0019552;C4299095|HIP
null|ST13 wt Allele|Finding|false|false|C0022122;C0228391;C0019552;C4299095|HIP
null|ST13 gene|Finding|false|false|C0022122;C0228391;C0019552;C4299095|HIP
null|HHIP gene|Finding|false|false|C0022122;C0228391;C0019552;C4299095|HIP
null|HHIP wt Allele|Finding|false|false|C0022122;C0228391;C0019552;C4299095|HIP
null|REG3A wt Allele|Finding|false|false|C0022122;C0228391;C0019552;C4299095|HIPnull|Procedure on hip|Procedure|false|false|C0022122;C0228391;C0019552;C4299095|HIPnull|Lower extremity>Hip|Anatomy|false|false|C1292890;C0559956;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C1555302;C0035139;C0392806;C1430701;C0529134;C1505163;C1654726|HIP
null|Hip structure|Anatomy|false|false|C1292890;C0559956;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C1555302;C0035139;C0392806;C1430701;C0529134;C1505163;C1654726|HIP
null|Structure of habenulopeduncular tract|Anatomy|false|false|C1292890;C0559956;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C1555302;C0035139;C0392806;C1430701;C0529134;C1505163;C1654726|HIP
null|Bone structure of ischium|Anatomy|false|false|C1292890;C0559956;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C1555302;C0035139;C0392806;C1430701;C0529134;C1505163;C1654726|HIPnull|Replacement|Finding|false|false|C0022122;C0228391;C0019552;C4299095|REPLACEMENTnull|Replacement - supply|Procedure|false|false|C0022122;C0228391;C0019552;C4299095|REPLACEMENT
null|Surgical Replantation|Procedure|false|false|C0022122;C0228391;C0019552;C4299095|REPLACEMENTnull|Hyperlipidemia|Disorder|false|false||HYPERLIPIDEMIA
null|Hyperlipoproteinemias|Disorder|false|false||HYPERLIPIDEMIAnull|Serum lipids high (finding)|Finding|false|false||HYPERLIPIDEMIAnull|Hypertensive disease|Disorder|false|false||HYPERTENSIONnull|Degenerative polyarthritis|Disorder|false|false||OSTEOARTHRITISnull|Herpes zoster (disorder)|Disorder|false|false||HERPES ZOSTER
null|herpesvirus 3, human|Disorder|false|false||HERPES ZOSTERnull|Herpes simplex dermatitis|Disorder|false|false||HERPES
null|null|Disorder|false|false||HERPESnull|Herpes <Hyperinae>|Entity|false|false||HERPESnull|Herpes zoster (disorder)|Disorder|false|false||ZOSTERnull|Atrial Fibrillation|Disorder|false|false|C0018792|ATRIAL FIBRILLATIONnull|null|Attribute|false|false|C0018792|ATRIAL FIBRILLATIONnull|Atrial Fibrillation by ECG Finding|Lab|false|false|C0018792|ATRIAL FIBRILLATIONnull|Heart Atrium|Anatomy|false|false|C0344434;C2926591;C0004238;C0232197|ATRIALnull|Fibrillation|Disorder|false|false|C0018792|FIBRILLATIONnull|Anxiety Disorders|Disorder|false|false||ANXIETY
null|Anxiety|Disorder|false|false||ANXIETYnull|Anxiety symptoms|Finding|false|false||ANXIETYnull|Gastrointestinal Hemorrhage|Finding|false|false||GASTROINTESTINAL BLEEDINGnull|Gastrointestinal attachment|Finding|false|false||GASTROINTESTINALnull|gastrointestinal|Modifier|false|false||GASTROINTESTINALnull|Hemorrhage|Finding|false|false||BLEEDINGnull|Degenerative polyarthritis|Disorder|false|false||OSTEOARTHRITISnull|Atherosclerosis|Disorder|false|false|C0007226;C3887460|ATHEROSCLEROTIC CARDIOVASCULAR DISEASEnull|atherosclerotic|Finding|false|false|C0007226;C3887460|ATHEROSCLEROTICnull|Cardiovascular Diseases|Disorder|false|false|C0007226;C3887460|CARDIOVASCULAR DISEASEnull|Cardiovascular system|Anatomy|false|false|C0012634;C0007222;C0004153;C0333482|CARDIOVASCULAR
null|Cardiovascular|Anatomy|false|false|C0012634;C0007222;C0004153;C0333482|CARDIOVASCULARnull|Disease|Disorder|false|false|C0007226;C3887460|DISEASEnull|Peripheral Vascular Diseases|Disorder|false|false|C0005847|PERIPHERAL VASCULAR DISEASEnull|Peripheral|Modifier|false|false||PERIPHERALnull|Vascular Diseases|Disorder|false|false|C0005847|VASCULAR DISEASEnull|Blood Vessel|Anatomy|false|false|C0042373;C0085096;C0012634|VASCULARnull|Vascular|Modifier|false|false||VASCULARnull|Disease|Disorder|false|false|C0005847|DISEASEnull|Relationship - Mother|Finding|false|false||Mothernull|Mother (person)|Subject|false|false||Mothernull|Hypertensive disease|Disorder|false|false||HTNnull|Indirect exposure mechanism - Father|Finding|false|false||Father
null|Relationship - Father|Finding|false|false||Father
null|Father - courtesy title|Finding|false|false||Fathernull|Father (person)|Subject|false|false||Fathernull|Brother - courtesy title|Finding|false|false||Brother
null|Relationship - Brother|Finding|false|false||Brothernull|Brothers|Subject|false|false||Brothernull|Brother - courtesy title|Finding|false|false||Brother
null|Relationship - Brother|Finding|false|false||Brothernull|Brothers|Subject|false|false||Brothernull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|physical examination (physical finding)|Finding|false|false||PHYSICAL EXAMnull|Physical Examination|Procedure|false|false||PHYSICAL EXAMnull|physical examination (physical finding)|Finding|false|false||PHYSICAL
null|Physical|Finding|false|false||PHYSICALnull|Physical Examination|Procedure|false|false||PHYSICALnull|Exam|Finding|false|false||EXAMnull|Medical Examination|Procedure|false|false||EXAMnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||GENERALnull|General medical service|Procedure|false|false||GENERALnull|Generalized|Modifier|false|false||GENERALnull|Well (answer to question)|Finding|false|false||Wellnull|Well (container)|Device|false|false||Wellnull|Microplate Well|Modifier|false|false||Well
null|Good|Modifier|false|false||Well
null|Healthy|Modifier|false|false||Wellnull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|Use of accessory muscles|Finding|true|false|C4083049;C0026845|accessory muscle usenull|Accessory skeletal muscle|Disorder|true|false|C4083049;C0026845|accessory musclenull|Accessory|Device|true|false||accessorynull|Muscle (organ)|Anatomy|false|false|C0158784;C1947944;C0042153;C0457083;C1821466|muscle
null|Muscle Tissue|Anatomy|false|false|C0158784;C1947944;C0042153;C0457083;C1821466|musclenull|Use - dosing instruction imperative|Finding|true|false|C4083049;C0026845|use
null|utilization qualifier|Finding|true|false|C4083049;C0026845|use
null|Usage|Finding|true|false|C4083049;C0026845|usenull|HEENT|Anatomy|false|false||HEENTnull|Scleral Diseases|Disorder|false|false|C0036410|Scleranull|examination of sclera|Procedure|false|false|C0036410|Scleranull|Sclera|Anatomy|false|false|C0205180;C2228481;C0036412|Scleranull|Anicteric|Finding|false|false|C0036410|anictericnull|Pupil equal round and reacting to light|Finding|false|false||PERRLnull|Passive joint movement of neck (finding)|Finding|false|false|C0027530;C3159206|NECK
null|Neck problem|Finding|false|false|C0027530;C3159206|NECKnull|dendritic spine neck|Anatomy|false|false|C0812434;C0684335|NECK
null|Neck|Anatomy|false|false|C0812434;C0684335|NECKnull|Jugular venous engorgement|Finding|true|false||JVDnull|Cardiac attachment|Finding|false|false|C0018787|CARDIACnull|Heart|Anatomy|false|false|C1314974|CARDIACnull|Cardiac - anatomy qualifier|Modifier|false|false||CARDIACnull|Irregular|Modifier|false|false||Irregularnull|Rhythm|Finding|false|false||rhythm
null|rhythmic process (biological)|Finding|false|false||rhythmnull|Amount type - Rate|Finding|false|false||ratenull|Rating (action)|Event|false|false||ratenull|Rate|LabModifier|false|false||ratenull|Heart murmur|Finding|false|false||murmursnull|Pericardial friction rub|Finding|false|false||rubsnull|Lung|Anatomy|false|false||LUNGSnull|Air (substance)|Drug|false|false||air
null|air|Drug|false|false||air
null|air|Drug|false|false||airnull|ACUTE INSULIN RESPONSE|Finding|false|false||air
null|AIRN gene|Finding|false|false||air
null|AI/RHEUM|Finding|false|false||airnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Sequence Chromatogram|Finding|false|false||Tracenull|Trace Dosing Unit|LabModifier|false|false||Trace
null|trace amount|LabModifier|false|false||Trace
null|unknown - trace|LabModifier|false|false||Tracenull|Inspiratory wheezing|Finding|false|false||inspiratory wheezingnull|Inspiration (function)|Finding|false|false||inspiratorynull|Wheezing|Finding|false|false||wheezingnull|Expiratory wheezing|Finding|false|false||expiratory wheezingnull|Expiration, Respiratory|Finding|false|false||expiratorynull|Wheezing|Finding|false|false||wheezingnull|Lung diseases|Disorder|false|false|C4037972;C0024109|lungnull|Lung Problem|Finding|false|false|C4037972;C0024109|lungnull|Chest>Lung|Anatomy|false|false|C0740941;C0024115|lung
null|Lung|Anatomy|false|false|C0740941;C0024115|lungnull|Basilar Rales|Finding|false|false||crackles
null|Rales|Finding|false|false||cracklesnull|Rhonchi|Finding|false|false||rhonchinull|Malignant neoplasm of abdomen|Disorder|false|false|C0230168;C0000726|ABDOMENnull|Abdomen problem|Finding|false|false|C0230168;C0000726|ABDOMENnull|Abdomen|Anatomy|false|false|C0941288;C0153662|ABDOMEN
null|Abdominal Cavity|Anatomy|false|false|C0941288;C0153662|ABDOMENnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||Softnull|Soft|Modifier|false|false||Softnull|LRRC4B gene|Finding|true|false||HSMnull|Emotional tenderness|Finding|true|false||tenderness
null|Sore to touch|Finding|true|false||tendernessnull|All extremities|Anatomy|false|false||EXTREMITIES
null|Limb structure|Anatomy|false|false||EXTREMITIESnull|Femur|Anatomy|false|false|C0006318|femoralnull|Bruit|Finding|true|false|C0015811|bruitsnull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|physical examination (physical finding)|Finding|false|false||PHYSICAL EXAMnull|Physical Examination|Procedure|false|false||PHYSICAL EXAMnull|physical examination (physical finding)|Finding|false|false||PHYSICAL
null|Physical|Finding|false|false||PHYSICALnull|Physical Examination|Procedure|false|false||PHYSICALnull|Exam|Finding|false|false||EXAMnull|Medical Examination|Procedure|false|false||EXAMnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||GENERALnull|General medical service|Procedure|false|false||GENERALnull|Generalized|Modifier|false|false||GENERALnull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|HEENT|Anatomy|false|false||HEENTnull|Scleral Diseases|Disorder|false|false|C0036410|Scleranull|examination of sclera|Procedure|false|false|C0036410|Scleranull|Sclera|Anatomy|false|false|C0205180;C2228481;C0036412|Scleranull|Anicteric|Finding|false|false|C0036410|anictericnull|Remote control command - Clear|Finding|false|false||clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|Passive joint movement of neck (finding)|Finding|false|false|C0027530;C3159206|NECK
null|Neck problem|Finding|false|false|C0027530;C3159206|NECKnull|dendritic spine neck|Anatomy|false|false|C0812434;C0684335|NECK
null|Neck|Anatomy|false|false|C0812434;C0684335|NECKnull|Jugular venous engorgement|Finding|true|false||JVDnull|Cardiac attachment|Finding|false|false|C0018787|CARDIACnull|Heart|Anatomy|false|false|C1314974|CARDIACnull|Cardiac - anatomy qualifier|Modifier|false|false||CARDIACnull|Heart murmur|Finding|true|false||murmursnull|Pericardial friction rub|Finding|true|false||rubsnull|Lung|Anatomy|false|false||LUNGSnull|MILDLY|Modifier|false|false||Mildly
null|Mild (qualifier value)|Modifier|false|false||Mildlynull|Air Movements|Phenomenon|false|false||air movementnull|Air (substance)|Drug|false|false||air
null|air|Drug|false|false||air
null|air|Drug|false|false||airnull|ACUTE INSULIN RESPONSE|Finding|false|false||air
null|AIRN gene|Finding|false|false||air
null|AI/RHEUM|Finding|false|false||airnull|Movement|Finding|false|false||movementnull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|Wheezing|Finding|false|false||wheezingnull|Rhonchi|Finding|false|false||rhonchinull|Basilar Rales|Finding|true|false||crackles
null|Rales|Finding|true|false||cracklesnull|Malignant neoplasm of abdomen|Disorder|false|false|C0230168;C0000726|ABDOMENnull|Abdomen problem|Finding|false|false|C0230168;C0000726|ABDOMENnull|Abdomen|Anatomy|false|false|C0941288;C0153662|ABDOMEN
null|Abdominal Cavity|Anatomy|false|false|C0941288;C0153662|ABDOMENnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||Softnull|Soft|Modifier|false|false||Softnull|LRRC4B gene|Finding|true|false||HSMnull|Emotional tenderness|Finding|true|false||tenderness
null|Sore to touch|Finding|true|false||tendernessnull|All extremities|Anatomy|false|false||EXTREMITIES
null|Limb structure|Anatomy|false|false||EXTREMITIESnull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|Laboratory test finding|Lab|false|false||LABSnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0005768;C0229664;C0005767;C0851353|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C1114281;C0014792|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Lymph|Finding|false|false||Lymphsnull|Monos|Drug|false|false||Monos
null|Mono-S|Drug|false|false||Monos
null|Monos|Drug|false|false||Monosnull|SARCOIDOSIS, EARLY-ONSET|Disorder|false|false||Eos
null|Familial eosinophilia|Disorder|false|false||Eosnull|PRSS33 gene|Finding|false|false||Eos
null|IKZF4 gene|Finding|false|false||Eosnull|Eos <Loriini>|Entity|false|false||Eosnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood calcium measurement|Procedure|false|false||BLOOD Calciumnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Laboratory test finding|Lab|false|false||LABSnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MB
null|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MBnull|creatine kinase activity|Finding|false|false||CK-MBnull|Serum creatine phosphokinase MB isoenzyme measurement|Procedure|false|false||CK-MB
null|Creatine kinase MB measurement|Procedure|false|false||CK-MBnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Thyrotropin-Releasing Hormone, human|Drug|false|false||TRF
null|IL5 protein, human|Drug|false|false||TRF
null|IL5 protein, human|Drug|false|false||TRF
null|thyrotropin-releasing hormone|Drug|false|false||TRF
null|thyrotropin-releasing hormone|Drug|false|false||TRF
null|thyrotropin-releasing hormone|Drug|false|false||TRF
null|Tocotrienol-rich Fraction|Drug|false|false||TRF
null|Thyrotropin-Releasing Hormone, human|Drug|false|false||TRFnull|TERF1 wt Allele|Finding|false|false||TRF
null|TERF1 gene|Finding|false|false||TRF
null|IL5 gene|Finding|false|false||TRFnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|thyrotropin|Drug|false|false||TSH
null|thyrotropin|Drug|false|false||TSH
null|thyrotropin|Drug|false|false||TSHnull|Thyroid stimulating hormone measurement|Procedure|false|false||TSHnull|null|Attribute|false|false||TSHnull|Mandibular right second molar abutment mesial hemisection|Device|false|false||31AMnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Partial pressure of Oxygen|Finding|false|false||pO2
null|US Military enlisted E5|Finding|false|false||pO2null|PO2 measurement|Procedure|false|false||pO2null|Carbon dioxide measurement, partial pressure|Procedure|false|false||pCO2null|Carbon dioxide, partial pressure|Lab|false|false||pCO2null|nitrogenous base|Drug|false|false|C2987514|Base
null|Base|Drug|false|false|C2987514|Base
null|Dental Base|Drug|false|false|C2987514|Base
null|base - RoleClass|Drug|false|false|C2987514|Basenull|Base - General Qualifier|Finding|false|false|C2987514|Base
null|BPIFA4P gene|Finding|false|false|C2987514|Base
null|Base - RX Component Type|Finding|false|false|C2987514|Basenull|Anatomical base|Anatomy|false|false|C1549548;C1705938;C1843354;C1704464;C0178499;C1550601;C1880279|Basenull|Base - unit of product usage|LabModifier|false|false||Basenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Free of (attribute)|Finding|false|false||FREEnull|Empty (qualifier)|Modifier|false|false||FREEnull|Direct - PostalAddressUse|Finding|false|false||DIRECT
null|direct address|Finding|false|false||DIRECTnull|Direct type of relationship|Modifier|false|false||DIRECT
null|Direct (qualifier)|Modifier|false|false||DIRECTnull|Dialysis Method of Administration|Finding|false|false|C4318744|DIALYSISnull|Dialysis procedure|Procedure|false|false|C4318744|DIALYSIS
null|Renal Dialysis|Procedure|false|false|C4318744|DIALYSISnull|dialysis device|Device|false|false||DIALYSISnull|Physical Dialysis|Phenomenon|false|false||DIALYSISnull|Dialysis <Coenomyiinae>|Entity|false|false||DIALYSISnull|Tests (qualifier value)|Finding|false|false|C4318744|Test
null|Testing|Finding|false|false|C4318744|Testnull|Laboratory Procedures|Procedure|false|false|C4318744|Testnull|Test - temporal region|Anatomy|false|false|C0456984;C0039593;C0392366;C0022885;C4723631;C0011946;C4551529|Testnull|Test Result|Lab|false|false|C4318744|Testnull|Test Dosing Unit|LabModifier|false|false||Testnull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|Laboratory test finding|Lab|false|false||LABSnull|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0005768;C0229664;C0005767;C0851353|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C1114281;C0014792|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood calcium measurement|Procedure|false|false||BLOOD Calciumnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Imaging problem|Finding|false|false||IMAGINGnull|Diagnostic Imaging|Procedure|false|false||IMAGING
null|Imaging Techniques|Procedure|false|false||IMAGINGnull|Imaging Technology|Title|false|false||IMAGINGnull|Plain chest X-ray|Procedure|false|false|C1527391;C0817096|Chest X raynull|Chest problem|Finding|false|false|C1527391;C0817096|Chestnull|Chest|Anatomy|false|false|C1428870;C5444437;C0043309;C1962945;C1306645;C0851346;C0741025;C0039985|Chest
null|Anterior thoracic region|Anatomy|false|false|C1428870;C5444437;C0043309;C1962945;C1306645;C0851346;C0741025;C0039985|Chestnull|Plain x-ray|Procedure|false|false|C1527391;C0817096|X ray
null|Radiographic imaging procedure|Procedure|false|false|C1527391;C0817096|X raynull|Roentgen Rays|Phenomenon|false|false|C1527391;C0817096|X raynull|RAB35 wt Allele|Finding|false|false|C1527391;C0817096|ray
null|SH3YL1 gene|Finding|false|false|C1527391;C0817096|raynull|Radiation|Phenomenon|false|false|C1527391;C0817096|raynull|Dipturus trachyderma|Entity|false|false||ray
null|Rajiformes|Entity|false|false||raynull|Living Arrangement - Relative|Finding|false|false|C4037972;C0024109|Relativenull|null|Attribute|false|false||Relativenull|Relative (related person)|Subject|false|false||Relativenull|Relative|Modifier|false|false||Relativenull|Increase|Finding|false|false|C4037972;C0024109|increasenull|Abnormally opaque structure (morphologic abnormality)|Finding|false|false||opacity
null|Decreased translucency|Finding|false|false||opacitynull|Lung diseases|Disorder|false|false|C4037972;C0024109|lungnull|Lung Problem|Finding|false|false|C4037972;C0024109|lungnull|Chest>Lung|Anatomy|false|false|C1546849;C0740941;C0024115;C0442805|lung
null|Lung|Anatomy|false|false|C1546849;C0740941;C0024115;C0442805|lungnull|Base|Drug|false|false||basesnull|Base - unit of product usage|LabModifier|false|false||basesnull|Neck+Chest>Soft tissue|Anatomy|false|false|C1547928;C3542022|soft tissue
null|soft tissue|Anatomy|false|false|C1547928;C3542022|soft tissuenull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false|C0040300;C0225317;C4532079|softnull|Soft|Modifier|false|false||softnull|Tissue Specimen Code|Finding|false|false|C0225317;C4532079;C0040300|tissuenull|Body tissue|Anatomy|false|false|C3542022;C1547928|tissuenull|Lung consolidation|Disorder|false|false||consolidationnull|Consolidation|Modifier|false|false||consolidationnull|Lateral|Modifier|false|false||Lateralnull|View|Modifier|false|false||viewnull|Helpful|Modifier|false|false||helpfulnull|confirmation - ResponseLevel|Finding|false|false||confirmation
null|Confirmation|Finding|false|false||confirmationnull|Confirmation of|Modifier|false|false||confirmationnull|Plain chest X-ray|Procedure|false|false|C1527391;C0817096|Chest X raynull|Chest problem|Finding|false|false|C1527391;C0817096|Chestnull|Chest|Anatomy|false|false|C1962945;C1306645;C0043309;C1428870;C5444437;C0741025;C0039985;C0851346|Chest
null|Anterior thoracic region|Anatomy|false|false|C1962945;C1306645;C0043309;C1428870;C5444437;C0741025;C0039985;C0851346|Chestnull|Plain x-ray|Procedure|false|false|C1527391;C0817096|X ray
null|Radiographic imaging procedure|Procedure|false|false|C1527391;C0817096|X raynull|Roentgen Rays|Phenomenon|false|false|C1527391;C0817096|X raynull|RAB35 wt Allele|Finding|false|false|C1527391;C0817096|ray
null|SH3YL1 gene|Finding|false|false|C1527391;C0817096|raynull|Radiation|Phenomenon|false|false|C1527391;C0817096|raynull|Dipturus trachyderma|Entity|false|false||ray
null|Rajiformes|Entity|false|false||raynull|Hyperdistention|Disorder|false|false||hyperinflationnull|Pneumothorax|Disorder|false|false||pneumothoraxnull|Effusion (substance)|Finding|false|false||effusion
null|null|Finding|false|false||effusion
null|effusion|Finding|false|false||effusionnull|Lung consolidation|Disorder|false|false||consolidationnull|Consolidation|Modifier|false|false||consolidationnull|Congestive heart failure|Disorder|false|false|C0262212|CHFnull|Choroidal fissure|Anatomy|false|false|C0018802|CHFnull|Probable diagnosis|Finding|false|false||probablenull|Probability|LabModifier|false|false||probablenull|Osteopenia|Disorder|false|false||osteopenianull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Peripheral Vascular Diseases|Disorder|false|false||PVDnull|Pomalidomide/Bortezomib/Dexamethasone Regimen|Procedure|false|false||PVDnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false|C1527391;C0817096|history
null|History of previous events|Finding|false|false|C1527391;C0817096|history
null|Historical aspects qualifier|Finding|false|false|C1527391;C0817096|history
null|Medical History|Finding|false|false|C1527391;C0817096|history
null|Concept History|Finding|false|false|C1527391;C0817096|historynull|History|Subject|false|false||historynull|Recurrent|Time|false|false||recurrent
null|Episodic|Time|false|false||recurrentnull|Chest Pain|Finding|false|false|C1527391;C0817096|chest painnull|null|Attribute|false|false|C1527391;C0817096|chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0262926;C1705255;C0019665;C0262512;C2004062;C0741025;C1549543;C0030193;C0008031;C2926613|chest
null|Anterior thoracic region|Anatomy|false|false|C0262926;C1705255;C0019665;C0262512;C2004062;C0741025;C1549543;C0030193;C0008031;C2926613|chestnull|Administration Method - Pain|Finding|false|false|C1527391;C0817096|pain
null|Pain|Finding|false|false|C1527391;C0817096|painnull|null|Attribute|false|false||painnull|Atrial Fibrillation|Disorder|false|false||afibnull|Atrial Fibrillation by ECG Finding|Lab|false|false||afibnull|Rapid Virologic Response|Finding|false|false||RVR
null|NR1D2 wt Allele|Finding|false|false||RVR
null|NR1D2 gene|Finding|false|false||RVRnull|COPD exacerbation|Disorder|false|false||COPD exacerbationnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|Exacerbation|Finding|false|false||exacerbationnull|Admission Level of Care Code - Acute|Finding|false|false||ACUTE
null|Acute - Triage Code|Finding|false|false||ACUTEnull|acute|Time|false|false||ACUTEnull|Problems - What subject filter|Finding|false|false||PROBLEMSnull|COPD exacerbation|Disorder|false|false||COPD exacerbationnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|Exacerbation|Finding|false|false||exacerbationnull|Recent|Time|false|false||recentnull|Visit|Finding|false|false||visitsnull|Patient Visit|Procedure|false|false||visitsnull|COPD exacerbation|Disorder|false|false||COPD exacerbationnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|Exacerbation|Finding|false|false||exacerbationnull|Recent|Time|false|false||recentlynull|prednisone|Drug|false|false||prednisone
null|prednisone|Drug|false|false||prednisone
null|prednisone|Drug|false|false||prednisonenull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|Address type - Office|Finding|false|false||officenull|Office|Device|false|false||officenull|Organization unit type - Office|Entity|false|false||officenull|null|Finding|false|false||dyspnea
null|Dyspnea|Finding|false|false||dyspneanull|Therapy Object (animal model)|Finding|false|false||therapy
null|therapeutic aspects|Finding|false|false||therapynull|Therapeutic procedure|Procedure|false|false||therapynull|Nasal congestion (finding)|Finding|false|false|C0028429|nasal congestionnull|Nasal brand of oxymetazoline|Drug|false|false|C0028429|nasal
null|Nasal brand of oxymetazoline|Drug|false|false|C0028429|nasal
null|Nasal dosage form|Drug|false|false|C0028429|nasalnull|Nasal Route of Administration|Finding|false|false|C0028429|nasal
null|Nasal (intended site)|Finding|false|false|C0028429|nasalnull|null|Anatomy|false|false|C0027424;C0700148;C4520890;C1522019;C1272939;C0721966|nasalnull|Congestion|Finding|false|false|C0028429|congestionnull|Viral|Finding|false|false||viralnull|Upper Respiratory Infections|Disorder|false|false||URInull|Uniform Resource Identifier|Finding|false|false||URI
null|URI1 gene|Finding|false|false||URI
null|URI1 wt Allele|Finding|false|false||URInull|Precipitating Factors|Attribute|false|false||triggernull|Triggered by|Modifier|false|false||triggernull|Clinic|Device|false|false||clinic
null|Ambulatory Care Facilities|Device|false|false||clinicnull|Clinic|Entity|false|false||clinic
null|Ambulatory Care Facilities|Entity|false|false||clinicnull|Patient location type - Clinic|Modifier|false|false||clinic
null|Person location type - Clinic|Modifier|false|false||clinicnull|Atrial Fibrillation|Disorder|false|false||afibnull|Atrial Fibrillation by ECG Finding|Lab|false|false||afibnull|Rapid Virologic Response|Finding|false|false||RVR
null|NR1D2 wt Allele|Finding|false|false||RVR
null|NR1D2 gene|Finding|false|false||RVRnull|Control brand of phenylpropanolamine|Drug|false|false||control
null|CONTROL veterinary product|Drug|false|false||control
null|control substance|Drug|false|false||control
null|Control brand of phenylpropanolamine|Drug|false|false||controlnull|Control - Relationship modifier|Finding|false|false||control
null|Control function|Finding|false|false||control
null|Scientific Control|Finding|false|false||controlnull|Control Groups|Subject|false|false||controlnull|True Control Status|Modifier|false|false||control
null|control aspects|Modifier|false|false||controlnull|null|Finding|false|false|C4037974;C0018787|heart ratenull|examination of heart rate|Procedure|false|false|C4037974;C0018787|heart ratenull|heart rate|Attribute|false|false|C4037974;C0018787|heart rate
null|null|Attribute|false|false|C4037974;C0018787|heart ratenull|Mean Heart Rate|LabModifier|false|false||heart ratenull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787|heart
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787|heartnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|heartnull|Chest>Heart|Anatomy|false|false|C1549480;C2041121;C0795691;C2197023;C0153957;C0153500;C0018810;C0488794|heart
null|Heart|Anatomy|false|false|C1549480;C2041121;C0795691;C2197023;C0153957;C0153500;C0018810;C0488794|heartnull|Amount type - Rate|Finding|false|false|C4037974;C0018787|ratenull|Rating (action)|Event|false|false||ratenull|Rate|LabModifier|false|false||ratenull|On admission|Time|false|false||On admissionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Floor (anatomic)|Anatomy|false|false||floornull|floor (object)|Device|false|false||floornull|Floor - story of building|Entity|false|false||floornull|Wheezing|Finding|false|false||wheezingnull|Increased work of breathing|Finding|false|false||increased work of breathingnull|Increased (finding)|Finding|false|false||increased
null|Increase|Finding|false|false||increasednull|Increased|LabModifier|false|false||increasednull|Work of Breathing|Finding|false|false||work of breathingnull|Work|Event|false|false||worknull|outcomes otolaryngology breathing|Finding|false|false||breathing
null|Inspiration (function)|Finding|false|false||breathing
null|Respiration|Finding|false|false||breathingnull|null|Attribute|false|false||breathingnull|respiratory system process|Phenomenon|false|false||breathingnull|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group|Finding|false|false||poor
null|Patient Condition Code - Poor|Finding|false|false||poornull|Poverty|Subject|false|false||poornull|Language Proficiency - Poor|Modifier|false|false||poor
null|Specimen Quality - Poor|Modifier|false|false||poor
null|Poor - grade|Modifier|false|false||poor
null|Poor - qualifier|Modifier|false|false||poornull|Air Movements|Phenomenon|false|false||air movementnull|Air (substance)|Drug|false|false||air
null|air|Drug|false|false||air
null|air|Drug|false|false||airnull|ACUTE INSULIN RESPONSE|Finding|false|false||air
null|AIRN gene|Finding|false|false||air
null|AI/RHEUM|Finding|false|false||airnull|Movement|Finding|false|false||movementnull|Solu-Medrol|Drug|false|false||solumedrol
null|Solu-Medrol|Drug|false|false||solumedrolnull|prednisone|Drug|false|false||prednisone
null|prednisone|Drug|false|false||prednisone
null|prednisone|Drug|false|false||prednisonenull|Daily|Time|false|false||dailynull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|theophylline|Drug|false|false||theophylline
null|theophylline|Drug|false|false||theophyllinenull|Assay of theophylline|Procedure|false|false||theophyllinenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Tachyarrhythmia|Finding|false|false||tachyarrhythmianull|ipratropium|Drug|false|false||ipratropium
null|ipratropium|Drug|false|false||ipratropiumnull|Nebulizer solution|Drug|false|false||nebsnull|Every six hours|Time|false|false||q6hnull|albuterol|Drug|false|false||albuterol
null|albuterol|Drug|false|false||albuterolnull|Nebulizer solution|Drug|false|false||nebsnull|Every two hours|Time|false|false||q2hnull|fluticasone / salmeterol|Drug|false|false||fluticasone-salmeterolnull|fluticasone|Drug|false|false||fluticasone
null|fluticasone|Drug|false|false||fluticasonenull|salmeterol|Drug|false|false||salmeterol
null|salmeterol|Drug|false|false||salmeterolnull|Pulmonary (intended site)|Finding|false|false|C0024109|Pulmonarynull|Lung|Anatomy|false|false|C4522268;C2707265|Pulmonarynull|null|Attribute|false|false|C0024109|Pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||Pulmonarynull|Clinical Trials|Procedure|false|false||trialnull|Diuresis|Finding|false|false||diuresisnull|Lasix|Drug|false|false||Lasix
null|Lasix|Drug|false|false||Lasixnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED|Drug|false|false||Azithromycin
null|azithromycin|Drug|false|false||Azithromycin
null|azithromycin|Drug|false|false||Azithromycinnull|theophylline|Drug|false|false||theophylline
null|theophylline|Drug|false|false||theophyllinenull|Assay of theophylline|Procedure|false|false||theophyllinenull|amiodarone|Drug|false|false||amiodarone
null|amiodarone|Drug|false|false||amiodaronenull|Drug assay amiodarone|Procedure|false|false||amiodaronenull|Corrected QT Interval|LabModifier|false|false||QTcnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Course|Time|false|false||coursenull|ceftriaxone|Drug|false|false||ceftriaxone
null|ceftriaxone|Drug|false|false||ceftriaxonenull|Course|Time|false|false||coursenull|cefpodoxime|Drug|false|false||cefpodoxime
null|cefpodoxime|Drug|false|false||cefpodoximenull|prednisone|Drug|false|false||prednisone
null|prednisone|Drug|false|false||prednisone
null|prednisone|Drug|false|false||prednisonenull|null|Procedure|false|false||tapernull|Every three days|Time|false|false||q3dnull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|Pulmonary ventilator management|Procedure|false|false||pulmnull|Follow-up status|Finding|false|false||follow upnull|follow-up|Procedure|false|false||follow upnull|Follow - dosing instruction imperative|Finding|false|false||follow
null|Follow|Finding|false|false||follownull|Followed by|Time|false|false||follownull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Pulmonary (intended site)|Finding|false|false|C0024109|pulmonarynull|Lung|Anatomy|false|false|C4522268|pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Rehabilitation therapy|Procedure|false|false||rehabnull|Pulmonologists|Subject|false|false||pulmonologistnull|Supplement|Finding|false|false||supplementalnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Atrial Fibrillation|Disorder|false|false|C0018792|Atrial fibrillationnull|null|Attribute|false|false|C0018792|Atrial fibrillationnull|Atrial Fibrillation by ECG Finding|Lab|false|false|C0018792|Atrial fibrillationnull|Heart Atrium|Anatomy|false|false|C0344434;C0004238;C0232197;C2926591|Atrialnull|Fibrillation|Disorder|false|false|C0018792|fibrillationnull|Heart Atrium|Anatomy|false|false||atrialnull|Fibrillation|Disorder|false|false||fibrillationnull|amiodarone|Drug|false|false||amiodarone
null|amiodarone|Drug|false|false||amiodaronenull|Drug assay amiodarone|Procedure|false|false||amiodaronenull|apixaban|Drug|false|false||apixaban
null|apixaban|Drug|false|false||apixabannull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|Address type - Office|Finding|false|false||officenull|Office|Device|false|false||officenull|Organization unit type - Office|Entity|false|false||officenull|Prompting|Finding|false|false||promptingnull|Referral to|Procedure|false|false||referral tonull|Patient referral|Procedure|false|false||referralnull|COPD exacerbation|Disorder|false|false||COPD exacerbationnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|Exacerbation|Finding|false|false||exacerbationnull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Possible|Finding|false|false||possiblynull|Possible diagnosis|Modifier|false|false||possiblynull|theophylline|Drug|false|false||theophylline
null|theophylline|Drug|false|false||theophyllinenull|Assay of theophylline|Procedure|false|false||theophyllinenull|diltiazem|Drug|false|false||diltiazem
null|diltiazem|Drug|false|false||diltiazemnull|Drops - Drug Form|Drug|false|false||gttnull|Gestational Trophoblastic Neoplasms|Disorder|false|false||gttnull|Glucose tolerance test|Procedure|false|false||gttnull|Drop Dosing Unit|LabModifier|false|false||gtt
null|Medical Drop|LabModifier|false|false||gttnull|diltiazem|Drug|false|false||diltiazem
null|diltiazem|Drug|false|false||diltiazemnull|Every six hours|Time|false|false||q6hnull|arrival - ActRelationshipType|Finding|false|false|C3714591|arrivalnull|null|Event|false|false||arrivalnull|Floor (anatomic)|Anatomy|false|false|C1555577|floornull|floor (object)|Device|false|false||floornull|Floor - story of building|Entity|false|false||floornull|amiodarone|Drug|false|false||amiodarone
null|amiodarone|Drug|false|false||amiodaronenull|Drug assay amiodarone|Procedure|false|false||amiodaronenull|apixaban|Drug|false|false||apixaban
null|apixaban|Drug|false|false||apixabannull|theophylline|Drug|false|false||theophylline
null|theophylline|Drug|false|false||theophyllinenull|Assay of theophylline|Procedure|false|false||theophyllinenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Iron deficiency anemia|Disorder|false|false||Iron deficiency anemianull|Iron deficiency anemia|Disorder|false|false||Iron deficiency
null|Iron deficiency|Disorder|false|false||Iron deficiencynull|Iron Drug Class|Drug|false|false||Iron
null|iron|Drug|false|false||Iron
null|iron|Drug|false|false||Iron
null|iron|Drug|false|false||Iron
null|Ferrum metallicum, Homeopathic preparation|Drug|false|false||Ironnull|Iron measurement|Procedure|false|false||Ironnull|Deficiency anemias|Disorder|false|false||deficiency anemianull|Malnutrition|Disorder|false|false||deficiencynull|Deficiency|Finding|false|false||deficiencynull|deficiency aspects|Modifier|false|false||deficiencynull|Anemia|Disorder|false|false||anemianull|Anemia <Anemiaceae>|Entity|false|false||anemianull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|microcytic|Finding|false|false||microcyticnull|Anemia|Disorder|false|false||anemianull|Anemia <Anemiaceae>|Entity|false|false||anemianull|Iron low|Finding|false|false||low ironnull|IPSS-R Risk Category Low|Finding|false|false||low
null|IPSS Risk Category Low|Finding|false|false||low
null|low confidentiality|Finding|false|false||lownull|Low - MessageWaitingPriority|Modifier|false|false||low
null|low|Modifier|false|false||low
null|low exposure|Modifier|false|false||lownull|null|LabModifier|false|false||lownull|Iron Drug Class|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|Ferrum metallicum, Homeopathic preparation|Drug|false|false||ironnull|Iron measurement|Procedure|false|false||ironnull|Ferritin|Drug|false|false||ferritin
null|Ferritin|Drug|false|false||ferritin
null|Ferritin|Drug|false|false||ferritinnull|Ferritin measurement|Procedure|false|false||ferritinnull|On IV|Finding|false|false||on IVnull|ferryl iron|Drug|false|false||IV ironnull|Iron Drug Class|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|Ferrum metallicum, Homeopathic preparation|Drug|false|false||ironnull|Iron measurement|Procedure|false|false||ironnull|ferric gluconate|Drug|false|false||ferric gluconate
null|ferric gluconate|Drug|false|false||ferric gluconatenull|ferric cation|Drug|false|false||ferric
null|ferric cation|Drug|false|false||ferricnull|gluconate|Drug|false|false||gluconate
null|Gluconates|Drug|false|false||gluconate
null|Gluconates|Drug|false|false||gluconate
null|gluconate|Drug|false|false||gluconate
null|gluconate|Drug|false|false||gluconatenull|Dosage|LabModifier|false|false||dosesnull|Iron Drug Class|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|Ferrum metallicum, Homeopathic preparation|Drug|false|false||ironnull|Iron measurement|Procedure|false|false||ironnull|Bowel Regimen|Procedure|false|false|C0021853|bowel regimennull|Intestines|Anatomy|false|false|C0040808;C5979615|bowelnull|GDC Regimen Terminology|Finding|false|false||regimennull|Treatment Protocols|Procedure|false|false|C0021853|regimennull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Hemorrhage|Finding|true|false||bleedingnull|Marketing basis - Transitional|Finding|false|false||Transitionalnull|Transitional cell morphology|Modifier|false|false||Transitionalnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|prednisone|Drug|false|false||prednisone
null|prednisone|Drug|false|false||prednisone
null|prednisone|Drug|false|false||prednisonenull|null|Procedure|false|false||tapernull|Reduced|Finding|false|false||decreasenull|Decrease|LabModifier|false|false||decreasenull|3 Days|Time|false|false||3 daysnull|day|Time|false|false||daysnull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|Pulmonary Medicine|Title|false|false||pulmonologynull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Infantile Neuroaxonal Dystrophy|Disorder|false|false||plannull|Treatment Plan|Finding|false|false||plan
null|Planned|Finding|false|false||plan
null|null|Finding|false|false||plannull|Pulmonary Medicine|Title|false|false||pulmonologynull|Pulmonary (intended site)|Finding|false|false|C0024109|pulmonarynull|Lung|Anatomy|false|false|C4522268;C2707265;C0034991|pulmonarynull|null|Attribute|false|false|C0024109|pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Rehabilitation therapy|Procedure|false|false|C0024109|rehabnull|Appointments|Event|false|false||appointmentnull|Pulmonary (intended site)|Finding|false|false|C0024109|pulmonarynull|Lung|Anatomy|false|false|C0034991;C2707265;C4522268|pulmonarynull|null|Attribute|false|false|C0024109|pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Rehabilitation therapy|Procedure|false|false|C0024109|rehabnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|2 Days|Time|false|false||2 daysnull|day|Time|false|false||daysnull|cefpodoxime|Drug|false|false||cefpodoxime
null|cefpodoxime|Drug|false|false||cefpodoximenull|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||completenull|Completion Status for valid values - Complete|Finding|false|false||complete
null|Data operation - complete|Finding|false|false||complete
null|Finish - dosing instruction imperative|Finding|false|false||completenull|Complete|Modifier|false|false||completenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Course|Time|false|false||coursenull|Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE|Drug|false|false||antibiotics
null|Antibiotics|Drug|false|false||antibiotics
null|Antibiotics, ophthalmologic|Drug|false|false||antibiotics
null|Antibiotics, Gynecological|Drug|false|false||antibiotics
null|antibiotics, intestinal|Drug|false|false||antibiotics
null|Antibiotic throat preparations|Drug|false|false||antibiotics
null|Antibiotics, Antitubercular|Drug|false|false||antibiotics
null|Antibiotics for systemic use|Drug|false|false||antibiotics
null|Antifungal Antibiotics, Topical|Drug|false|false||antibioticsnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|COPD exacerbation|Disorder|false|false||COPD exacerbationnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|Exacerbation|Finding|false|false||exacerbationnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Concentrator Device|Device|false|false||concentratornull|Continuous|Finding|false|false||continuousnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|theophylline|Drug|false|false||theophylline
null|theophylline|Drug|false|false||theophyllinenull|Assay of theophylline|Procedure|false|false||theophyllinenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Atrial Fibrillation|Disorder|false|false||afibnull|Atrial Fibrillation by ECG Finding|Lab|false|false||afibnull|Rapid Virologic Response|Finding|false|false||RVR
null|NR1D2 wt Allele|Finding|false|false||RVR
null|NR1D2 gene|Finding|false|false||RVRnull|Further|Modifier|false|false||furthernull|theophylline|Drug|false|false||theophylline
null|theophylline|Drug|false|false||theophyllinenull|Assay of theophylline|Procedure|false|false||theophyllinenull|Weaning|Finding|false|false||weannull|In addition to|Finding|false|false||addition
null|Add - instruction imperative|Finding|false|false||additionnull|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED|Drug|false|false||azithromycin
null|azithromycin|Drug|false|false||azithromycin
null|azithromycin|Drug|false|false||azithromycinnull|Corrected QT Interval|LabModifier|false|false||QTcnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|amiodarone|Drug|false|false||amiodarone
null|amiodarone|Drug|false|false||amiodaronenull|Drug assay amiodarone|Procedure|false|false||amiodaronenull|roflumilast|Drug|false|false||roflumilast
null|roflumilast|Drug|false|false||roflumilastnull|Therapy Object (animal model)|Finding|false|false||therapy
null|therapeutic aspects|Finding|false|false||therapynull|Therapeutic procedure|Procedure|false|false||therapynull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Iron Drug Class|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|Ferrum metallicum, Homeopathic preparation|Drug|false|false||ironnull|Iron measurement|Procedure|false|false||ironnull|Deficiency|Finding|false|false||deficientnull|On IV|Finding|false|false||on IVnull|ferryl iron|Drug|false|false||IV ironnull|Iron Drug Class|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|Ferrum metallicum, Homeopathic preparation|Drug|false|false||ironnull|Iron measurement|Procedure|false|false||ironnull|Iron Drug Class|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|Ferrum metallicum, Homeopathic preparation|Drug|false|false||ironnull|Iron measurement|Procedure|false|false||ironnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Raised TSH level|Finding|false|false||elevated TSHnull|Elevated|Modifier|false|false||elevated
null|High|Modifier|false|false||elevatednull|thyrotropin|Drug|false|false||TSH
null|thyrotropin|Drug|false|false||TSH
null|thyrotropin|Drug|false|false||TSHnull|Thyroid stimulating hormone measurement|Procedure|false|false||TSHnull|null|Attribute|false|false||TSHnull|T4 free measurement|Procedure|false|false||free T4null|Free of (attribute)|Finding|false|false||freenull|Empty (qualifier)|Modifier|false|false||freenull|Pending - Allergy Clinical Status|Finding|false|false||pending
null|Pending - referral status|Finding|false|false||pendingnull|Pending - status|Time|false|false||pendingnull|pending - ManagedParticipationStatus|Modifier|false|false||pending
null|pending - RoleStatus|Modifier|false|false||pending
null|Pending - Day type|Modifier|false|false||pendingnull|On discharge|Time|false|false||on dischargenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|MDF Attribute Type - Code|Finding|false|false||Code
null|A Codes|Finding|false|false||Code
null|Code|Finding|false|false||Codenull|Coding|Event|false|false||Codenull|Full|Modifier|false|false||fullnull|emergency contact|Finding|false|false||Emergency Contactnull|Consent Non-Disclosure Reason - Emergency|Finding|false|false||Emergency
null|Admission Type - Emergency|Finding|false|false||Emergency
null|Referral category - Emergency|Finding|false|false||Emergency
null|Emergencies [Disease/Finding]|Finding|false|false||Emergency
null|Consent Bypass Reason - Emergency|Finding|false|false||Emergency
null|Level of Care - Emergency|Finding|false|false||Emergency
null|Certification patient type - Emergency|Finding|false|false||Emergency
null|Encounter Admission Source - emergency|Finding|false|false||Emergency
null|Patient Class - Emergency|Finding|false|false||Emergency
null|Visit Priority Code - Emergency|Finding|false|false||Emergencynull|emergency encounter|Procedure|false|false||Emergencynull|Emergency Situation|Phenomenon|false|false||Emergencynull|Specialty Type - Emergency|Title|false|false||Emergencynull|Bale out|Time|false|false||Emergencynull|Contact - HL7 Attribution|Finding|false|false||Contact
null|Contact with|Finding|false|false||Contact
null|Communication Contact|Finding|false|false||Contactnull|contact person|Subject|false|false||Contactnull|Physical contact|Phenomenon|false|false||Contactnull|Personal Contact|Event|false|false||Contactnull|husband|Subject|false|false||Husbandnull|Daughter|Subject|false|false||Daughternull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|MEDICATION LIST|Finding|false|false||Medication listnull|Pharmaceutical Preparations|Drug|false|false||Medicationnull|medication - HL7 publishing domain|Finding|false|false||Medication
null|Medications|Finding|false|false||Medicationnull|List|Finding|false|false||list
null|Sequence Data Type|Finding|false|false||listnull|Accurate (qualifier value)|Modifier|false|false||accuratenull|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||completenull|Completion Status for valid values - Complete|Finding|false|false||complete
null|Data operation - complete|Finding|false|false||complete
null|Finish - dosing instruction imperative|Finding|false|false||completenull|Complete|Modifier|false|false||completenull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|apixaban|Drug|false|false||Apixaban
null|apixaban|Drug|false|false||Apixabannull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|albuterol|Drug|false|false||Albuterol
null|albuterol|Drug|false|false||Albuterolnull|NEB protein, human|Drug|false|false||Neb
null|NEB protein, human|Drug|false|false||Neb
null|Nebulizer solution|Drug|false|false||Nebnull|NEB gene|Finding|false|false||Neb
null|mitotic nuclear membrane disassembly|Finding|false|false||Nebnull|NEB protein, human|Drug|false|false||NEB
null|NEB protein, human|Drug|false|false||NEB
null|Nebulizer solution|Drug|false|false||NEBnull|NEB gene|Finding|false|false||NEB
null|mitotic nuclear membrane disassembly|Finding|false|false||NEBnull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Breath|Finding|false|false||breathnull|amiodarone|Drug|false|false||Amiodarone
null|amiodarone|Drug|false|false||Amiodaronenull|Drug assay amiodarone|Procedure|false|false||Amiodaronenull|Daily|Time|false|false||DAILYnull|atorvastatin|Drug|false|false||Atorvastatin
null|atorvastatin|Drug|false|false||Atorvastatinnull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|artificial tears (medication)|Drug|false|false||Artificial Tears
null|Lubricant Eye Drops|Drug|false|false||Artificial Tears
null|Artificial Tears|Drug|false|false||Artificial Tearsnull|Artificial (qualifier value)|Modifier|false|false||Artificialnull|Tears (substance)|Finding|false|false||Tears
null|null|Finding|false|false||Tears
null|Tears specimen|Finding|false|false||Tearsnull|Drops - Drug Form|Drug|false|false||DROPnull|Dropping|Event|false|false||DROPnull|Drop (unit of presentation)|LabModifier|false|false||DROP
null|Drop British|LabModifier|false|false||DROP
null|Drop Dosing Unit|LabModifier|false|false||DROP
null|Medical Drop|LabModifier|false|false||DROP
null|Drop Unit of Volume|LabModifier|false|false||DROPnull|Structure of both eyes|Anatomy|false|false||BOTH EYESnull|Eye|Anatomy|false|false|C5848506|EYESnull|null|Attribute|false|false|C0015392|EYESnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Have Vulvar Irritation question|Finding|false|false||irritation
null|Irritability - emotion|Finding|false|false||irritation
null|Irritation (finding)|Finding|false|false||irritationnull|Irritation|Phenomenon|false|false||irritationnull|latanoprost|Drug|false|false||Latanoprost
null|latanoprost|Drug|false|false||Latanoprostnull|Ophthalmic Route of Administration|Finding|false|false||Ophthnull|Drops - Drug Form|Drug|false|false|C0229090|DROPnull|Dropping|Event|false|false|C0229090|DROPnull|Drop (unit of presentation)|LabModifier|false|false||DROP
null|Drop British|LabModifier|false|false||DROP
null|Drop Dosing Unit|LabModifier|false|false||DROP
null|Medical Drop|LabModifier|false|false||DROP
null|Drop Unit of Volume|LabModifier|false|false||DROPnull|examination of left eye|Procedure|false|false|C0229090;C4266572;C0015392;C0700042|LEFT EYEnull|Left eye structure|Anatomy|false|false|C2141124;C0154094;C0015397;C1552822;C1705648;C1550636;C1546630;C0262477;C0991568|LEFT EYEnull|Table Cell Horizontal Align - left|Finding|false|false|C0229090;C4266572;C0015392;C0700042|LEFTnull|Left sided|Modifier|false|false||LEFT
null|Left|Modifier|false|false||LEFTnull|Carcinoma in situ of eye|Disorder|false|false|C4266572;C0015392;C0700042;C0229090|EYE
null|Disorder of eye|Disorder|false|false|C4266572;C0015392;C0700042;C0229090|EYEnull|Eye - Specimen Source Code|Finding|false|false|C4266572;C0015392;C0700042;C0229090|EYE
null|Eye problem|Finding|false|false|C4266572;C0015392;C0700042;C0229090|EYE
null|Eye Specimen|Finding|false|false|C4266572;C0015392;C0700042;C0229090|EYEnull|Head>Eye|Anatomy|false|false|C0154094;C0015397;C1550636;C1546630;C0262477;C2141124;C1552822|EYE
null|Eye|Anatomy|false|false|C0154094;C0015397;C1550636;C1546630;C0262477;C2141124;C1552822|EYE
null|Orbital region|Anatomy|false|false|C0154094;C0015397;C1550636;C1546630;C0262477;C2141124;C1552822|EYEnull|Once a day, at bedtime|Time|false|false||QHSnull|diltiazem|Drug|false|false||Diltiazem
null|diltiazem|Drug|false|false||Diltiazemnull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|fluticasone propionate|Drug|false|false||Fluticasone Propionate
null|fluticasone propionate|Drug|false|false||Fluticasone Propionatenull|fluticasone|Drug|false|false||Fluticasone
null|fluticasone|Drug|false|false||Fluticasonenull|propionate|Drug|false|false||Propionate
null|Propionates|Drug|false|false||Propionatenull|Nasal brand of oxymetazoline|Drug|false|false|C0028429|NASAL
null|Nasal brand of oxymetazoline|Drug|false|false|C0028429|NASAL
null|Nasal dosage form|Drug|false|false|C0028429|NASALnull|Nasal Route of Administration|Finding|false|false|C0028429|NASAL
null|Nasal (intended site)|Finding|false|false|C0028429|NASALnull|null|Anatomy|false|false|C4520890;C1522019;C1332410;C1272939;C0721966;C4546282|NASALnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false|C0028429|BIDnull|BID gene|Finding|false|false|C0028429|BIDnull|Twice a day|Time|false|false||BIDnull|Fluticasone-Salmeterol Diskus|Drug|false|false||Fluticasone-Salmeterol Diskus
null|Fluticasone-Salmeterol Diskus|Drug|false|false||Fluticasone-Salmeterol Diskusnull|fluticasone / salmeterol|Drug|false|false||Fluticasone-Salmeterolnull|fluticasone|Drug|false|false||Fluticasone
null|fluticasone|Drug|false|false||Fluticasonenull|salmeterol|Drug|false|false||Salmeterol
null|salmeterol|Drug|false|false||Salmeterolnull|Diskus|Device|false|false||Diskusnull|Inhalant dose form|Drug|false|false||INH
null|isoniazid|Drug|false|false||INH
null|isoniazid|Drug|false|false||INHnull|Inhalation Route of Administration|Finding|false|false||INHnull|Ingush language|Entity|false|false||INHnull|Inhalation Dosing Unit|LabModifier|false|false||INHnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|hydrochlorothiazide|Drug|false|false||Hydrochlorothiazide
null|hydrochlorothiazide|Drug|false|false||Hydrochlorothiazidenull|Daily|Time|false|false||DAILYnull|isosorbide mononitrate|Drug|false|false||Isosorbide Mononitrate
null|isosorbide mononitrate|Drug|false|false||Isosorbide Mononitratenull|isosorbide|Drug|false|false||Isosorbide
null|isosorbide|Drug|false|false||Isosorbidenull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Daily|Time|false|false||DAILYnull|lorazepam|Drug|false|false||Lorazepam
null|lorazepam|Drug|false|false||Lorazepamnull|Once a day, at bedtime|Time|false|false||QHSnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Insomnia homeopathic medication|Drug|false|false||insomnianull|Sleeplessness|Finding|false|false||insomnianull|Theophylline ER|Drug|false|false||Theophylline ER
null|Theophylline ER|Drug|false|false||Theophylline ERnull|theophylline|Drug|false|false||Theophylline
null|theophylline|Drug|false|false||Theophyllinenull|Assay of theophylline|Procedure|false|false||Theophyllinenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|ranitidine|Drug|false|false||Ranitidine
null|ranitidine|Drug|false|false||Ranitidinenull|Daily|Time|false|false||DAILYnull|tiotropium bromide|Drug|false|false||Tiotropium Bromide
null|tiotropium bromide|Drug|false|false||Tiotropium Bromidenull|tiotropium|Drug|false|false||Tiotropium
null|tiotropium|Drug|false|false||Tiotropiumnull|Bromides|Drug|false|false||Bromidenull|Bromides measurement|Procedure|false|false||Bromidenull|capsule (pharmacologic)|Drug|false|false||CAPnull|CATARACT, ANTERIOR POLAR|Disorder|false|false||CAPnull|BRD4 wt Allele|Finding|false|false||CAP
null|HACD1 gene|Finding|false|false||CAP
null|SERPINB6 gene|Finding|false|false||CAP
null|BRD4 gene|Finding|false|false||CAP
null|CAP1 gene|Finding|false|false||CAP
null|SORBS1 gene|Finding|false|false||CAP
null|LNPEP gene|Finding|false|false||CAPnull|CAP Regimen|Procedure|false|false||CAP
null|cisplatin/cyclophosphamide/doxorubicin protocol|Procedure|false|false||CAP
null|cyclophosphamide/doxorubicin/prednisone protocol|Procedure|false|false||CAPnull|Cap (physical object)|Device|false|false||CAP
null|Syringe Caps|Device|false|false||CAP
null|Cap device|Device|false|false||CAPnull|College of American Pathologists|Subject|false|false||CAPnull|Controlled Attenuation Parameter|Modifier|false|false||CAPnull|Capsule Dosing Unit|LabModifier|false|false||CAPnull|Daily|Time|false|false||DAILYnull|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin Drug Class|Drug|false|false||Multivitamins
null|Multivitamin Drug Class|Drug|false|false||Multivitaminsnull|Minerals|Drug|false|false||mineralsnull|Tablet Dosage Form|Drug|false|false||TABnull|Tablet Dosing Unit|LabModifier|false|false||TABnull|Daily|Time|false|false||DAILYnull|aspirin|Drug|false|false||Aspirin
null|aspirin|Drug|false|false||Aspirinnull|Daily|Time|false|false||DAILYnull|dorzolamide|Drug|false|false||Dorzolamide
null|dorzolamide|Drug|false|false||Dorzolamidenull|Ophthalmic Route of Administration|Finding|false|false||Ophthnull|Drops - Drug Form|Drug|false|false||DROPnull|Dropping|Event|false|false|C0229118|DROPnull|Drop (unit of presentation)|LabModifier|false|false||DROP
null|Drop British|LabModifier|false|false||DROP
null|Drop Dosing Unit|LabModifier|false|false||DROP
null|Medical Drop|LabModifier|false|false||DROP
null|Drop Unit of Volume|LabModifier|false|false||DROPnull|Structure of both eyes|Anatomy|false|false|C1705648|BOTH EYESnull|Eye|Anatomy|false|false|C5848506;C4546282|EYESnull|null|Attribute|false|false|C0015392|EYESnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false|C0015392|BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|Continuous|Finding|false|false|C0028429|continuousnull|Oxygen nasal cannula|Device|false|false||nasal cannula
null|Nasal Cannula|Device|false|false||nasal cannulanull|Nasal brand of oxymetazoline|Drug|false|false|C0028429|nasal
null|Nasal brand of oxymetazoline|Drug|false|false|C0028429|nasal
null|Nasal dosage form|Drug|false|false|C0028429|nasalnull|Nasal Route of Administration|Finding|false|false|C0028429|nasal
null|Nasal (intended site)|Finding|false|false|C0028429|nasalnull|null|Anatomy|false|false|C1272939;C0721966;C0549178;C4520890;C1522019;C1550622;C1546577|nasalnull|Specimen Type - Cannula|Finding|false|false|C1550232;C0028429|cannula
null|null|Finding|false|false|C1550232;C0028429|cannulanull|Body Parts - Cannula|Anatomy|false|false|C1550622;C1546577|cannulanull|Cannula device|Device|false|false||cannulanull|Calamus <grasshoppers>|Entity|false|false||cannulanull|Exertion|Finding|false|false||exertionnull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Chronic Obstructive Airway Disease|Disorder|false|false|C0024109|chronic obstructive pulmonary diseasenull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Lung Diseases, Obstructive|Disorder|false|false|C0024109|obstructive pulmonary diseasenull|Obstructed|Finding|false|false||obstructivenull|Lung diseases|Disorder|false|false|C0024109|pulmonary diseasenull|History of - respiratory disease|Finding|false|false|C0024109|pulmonary diseasenull|Pulmonary (intended site)|Finding|false|false|C0024109|pulmonarynull|Lung|Anatomy|false|false|C0024117;C0024115;C4522268;C2707265;C0600260;C0455540;C0012634|pulmonarynull|null|Attribute|false|false|C0024109|pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Disease|Disorder|false|false|C0024109|diseasenull|Length|LabModifier|false|false||Lengthnull|Patient need for (contextual qualifier)|Finding|false|false||Needsnull|Needs|Modifier|false|false||Needsnull|Continuous|Finding|false|false||ongoingnull|year|Time|false|false||yearsnull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|amiodarone|Drug|false|false||Amiodarone
null|amiodarone|Drug|false|false||Amiodaronenull|Drug assay amiodarone|Procedure|false|false||Amiodaronenull|Daily|Time|false|false||DAILYnull|apixaban|Drug|false|false||Apixaban
null|apixaban|Drug|false|false||Apixabannull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|albuterol|Drug|false|false||Albuterol
null|albuterol|Drug|false|false||Albuterolnull|NEB protein, human|Drug|false|false||Neb
null|NEB protein, human|Drug|false|false||Neb
null|Nebulizer solution|Drug|false|false||Nebnull|NEB gene|Finding|false|false||Neb
null|mitotic nuclear membrane disassembly|Finding|false|false||Nebnull|NEB protein, human|Drug|false|false||NEB
null|NEB protein, human|Drug|false|false||NEB
null|Nebulizer solution|Drug|false|false||NEBnull|NEB gene|Finding|false|false||NEB
null|mitotic nuclear membrane disassembly|Finding|false|false||NEBnull|Every two hours|Time|false|false||Q2Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Breath|Finding|false|false||breathnull|artificial tears (medication)|Drug|false|false||Artificial Tears
null|Lubricant Eye Drops|Drug|false|false||Artificial Tears
null|Artificial Tears|Drug|false|false||Artificial Tearsnull|Artificial (qualifier value)|Modifier|false|false||Artificialnull|Tears (substance)|Finding|false|false||Tears
null|null|Finding|false|false||Tears
null|Tears specimen|Finding|false|false||Tearsnull|Drops - Drug Form|Drug|false|false||DROPnull|Dropping|Event|false|false||DROPnull|Drop (unit of presentation)|LabModifier|false|false||DROP
null|Drop British|LabModifier|false|false||DROP
null|Drop Dosing Unit|LabModifier|false|false||DROP
null|Medical Drop|LabModifier|false|false||DROP
null|Drop Unit of Volume|LabModifier|false|false||DROPnull|Structure of both eyes|Anatomy|false|false||BOTH EYESnull|Eye|Anatomy|false|false|C5848506|EYESnull|null|Attribute|false|false|C0015392|EYESnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Have Vulvar Irritation question|Finding|false|false||irritation
null|Irritability - emotion|Finding|false|false||irritation
null|Irritation (finding)|Finding|false|false||irritationnull|Irritation|Phenomenon|false|false||irritationnull|aspirin|Drug|false|false||Aspirin
null|aspirin|Drug|false|false||Aspirinnull|Daily|Time|false|false||DAILYnull|atorvastatin|Drug|false|false||Atorvastatin
null|atorvastatin|Drug|false|false||Atorvastatinnull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|diltiazem|Drug|false|false||Diltiazem
null|diltiazem|Drug|false|false||Diltiazemnull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|dorzolamide|Drug|false|false||Dorzolamide
null|dorzolamide|Drug|false|false||Dorzolamidenull|Ophthalmic Route of Administration|Finding|false|false||Ophthnull|Drops - Drug Form|Drug|false|false||DROPnull|Dropping|Event|false|false|C0229118|DROPnull|Drop (unit of presentation)|LabModifier|false|false||DROP
null|Drop British|LabModifier|false|false||DROP
null|Drop Dosing Unit|LabModifier|false|false||DROP
null|Medical Drop|LabModifier|false|false||DROP
null|Drop Unit of Volume|LabModifier|false|false||DROPnull|Structure of both eyes|Anatomy|false|false|C1705648;C4546282;C1332410|BOTH EYESnull|Eye|Anatomy|false|false|C5848506;C1332410;C4546282|EYESnull|null|Attribute|false|false|C0015392|EYESnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false|C0229118;C0015392|BIDnull|BID gene|Finding|false|false|C0015392;C0229118|BIDnull|Twice a day|Time|false|false||BIDnull|fluticasone propionate|Drug|false|false||Fluticasone Propionate
null|fluticasone propionate|Drug|false|false||Fluticasone Propionatenull|fluticasone|Drug|false|false||Fluticasone
null|fluticasone|Drug|false|false||Fluticasonenull|propionate|Drug|false|false||Propionate
null|Propionates|Drug|false|false||Propionatenull|Nasal brand of oxymetazoline|Drug|false|false|C0028429|NASAL
null|Nasal brand of oxymetazoline|Drug|false|false|C0028429|NASAL
null|Nasal dosage form|Drug|false|false|C0028429|NASALnull|Nasal Route of Administration|Finding|false|false|C0028429|NASAL
null|Nasal (intended site)|Finding|false|false|C0028429|NASALnull|null|Anatomy|false|false|C4546282;C1332410;C4520890;C1522019;C1272939;C0721966|NASALnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false|C0028429|BIDnull|BID gene|Finding|false|false|C0028429|BIDnull|Twice a day|Time|false|false||BIDnull|Fluticasone-Salmeterol Diskus|Drug|false|false||Fluticasone-Salmeterol Diskus
null|Fluticasone-Salmeterol Diskus|Drug|false|false||Fluticasone-Salmeterol Diskusnull|fluticasone / salmeterol|Drug|false|false||Fluticasone-Salmeterolnull|fluticasone|Drug|false|false||Fluticasone
null|fluticasone|Drug|false|false||Fluticasonenull|salmeterol|Drug|false|false||Salmeterol
null|salmeterol|Drug|false|false||Salmeterolnull|Diskus|Device|false|false||Diskusnull|Inhalant dose form|Drug|false|false||INH
null|isoniazid|Drug|false|false||INH
null|isoniazid|Drug|false|false||INHnull|Inhalation Route of Administration|Finding|false|false||INHnull|Ingush language|Entity|false|false||INHnull|Inhalation Dosing Unit|LabModifier|false|false||INHnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|hydrochlorothiazide|Drug|false|false||Hydrochlorothiazide
null|hydrochlorothiazide|Drug|false|false||Hydrochlorothiazidenull|Daily|Time|false|false||DAILYnull|isosorbide mononitrate|Drug|false|false||Isosorbide Mononitrate
null|isosorbide mononitrate|Drug|false|false||Isosorbide Mononitratenull|isosorbide|Drug|false|false||Isosorbide
null|isosorbide|Drug|false|false||Isosorbidenull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Daily|Time|false|false||DAILYnull|latanoprost|Drug|false|false||Latanoprost
null|latanoprost|Drug|false|false||Latanoprostnull|Ophthalmic Route of Administration|Finding|false|false||Ophthnull|Drops - Drug Form|Drug|false|false|C0229090|DROPnull|Dropping|Event|false|false|C0229090|DROPnull|Drop (unit of presentation)|LabModifier|false|false||DROP
null|Drop British|LabModifier|false|false||DROP
null|Drop Dosing Unit|LabModifier|false|false||DROP
null|Medical Drop|LabModifier|false|false||DROP
null|Drop Unit of Volume|LabModifier|false|false||DROPnull|examination of left eye|Procedure|false|false|C0229090;C4266572;C0015392;C0700042|LEFT EYEnull|Left eye structure|Anatomy|false|false|C2141124;C0154094;C0015397;C0991568;C1552822;C1705648;C1550636;C1546630;C0262477|LEFT EYEnull|Table Cell Horizontal Align - left|Finding|false|false|C0229090;C4266572;C0015392;C0700042|LEFTnull|Left sided|Modifier|false|false||LEFT
null|Left|Modifier|false|false||LEFTnull|Carcinoma in situ of eye|Disorder|false|false|C0229090;C4266572;C0015392;C0700042|EYE
null|Disorder of eye|Disorder|false|false|C0229090;C4266572;C0015392;C0700042|EYEnull|Eye - Specimen Source Code|Finding|false|false|C0229090;C4266572;C0015392;C0700042|EYE
null|Eye problem|Finding|false|false|C0229090;C4266572;C0015392;C0700042|EYE
null|Eye Specimen|Finding|false|false|C0229090;C4266572;C0015392;C0700042|EYEnull|Head>Eye|Anatomy|false|false|C1552822;C0154094;C0015397;C1550636;C1546630;C0262477;C2141124|EYE
null|Eye|Anatomy|false|false|C1552822;C0154094;C0015397;C1550636;C1546630;C0262477;C2141124|EYE
null|Orbital region|Anatomy|false|false|C1552822;C0154094;C0015397;C1550636;C1546630;C0262477;C2141124|EYEnull|Once a day, at bedtime|Time|false|false||QHSnull|lorazepam|Drug|false|false||Lorazepam
null|lorazepam|Drug|false|false||Lorazepamnull|Once a day, at bedtime|Time|false|false||QHSnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Insomnia homeopathic medication|Drug|false|false||insomnianull|Sleeplessness|Finding|false|false||insomnianull|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin Drug Class|Drug|false|false||Multivitamins
null|Multivitamin Drug Class|Drug|false|false||Multivitaminsnull|Minerals|Drug|false|false||mineralsnull|Tablet Dosage Form|Drug|false|false||TABnull|Tablet Dosing Unit|LabModifier|false|false||TABnull|Daily|Time|false|false||DAILYnull|ranitidine|Drug|false|false||Ranitidine
null|ranitidine|Drug|false|false||Ranitidinenull|Daily|Time|false|false||DAILYnull|tiotropium bromide|Drug|false|false||Tiotropium Bromide
null|tiotropium bromide|Drug|false|false||Tiotropium Bromidenull|tiotropium|Drug|false|false||Tiotropium
null|tiotropium|Drug|false|false||Tiotropiumnull|Bromides|Drug|false|false||Bromidenull|Bromides measurement|Procedure|false|false||Bromidenull|capsule (pharmacologic)|Drug|false|false||CAPnull|CATARACT, ANTERIOR POLAR|Disorder|false|false||CAPnull|BRD4 wt Allele|Finding|false|false||CAP
null|HACD1 gene|Finding|false|false||CAP
null|SERPINB6 gene|Finding|false|false||CAP
null|BRD4 gene|Finding|false|false||CAP
null|CAP1 gene|Finding|false|false||CAP
null|SORBS1 gene|Finding|false|false||CAP
null|LNPEP gene|Finding|false|false||CAPnull|CAP Regimen|Procedure|false|false||CAP
null|cisplatin/cyclophosphamide/doxorubicin protocol|Procedure|false|false||CAP
null|cyclophosphamide/doxorubicin/prednisone protocol|Procedure|false|false||CAPnull|Cap (physical object)|Device|false|false||CAP
null|Syringe Caps|Device|false|false||CAP
null|Cap device|Device|false|false||CAPnull|College of American Pathologists|Subject|false|false||CAPnull|Controlled Attenuation Parameter|Modifier|false|false||CAPnull|Capsule Dosing Unit|LabModifier|false|false||CAPnull|Daily|Time|false|false||DAILYnull|Theophylline SR|Drug|false|false||Theophylline SR
null|Theophylline SR|Drug|false|false||Theophylline SRnull|theophylline|Drug|false|false||Theophylline
null|theophylline|Drug|false|false||Theophyllinenull|Assay of theophylline|Procedure|false|false||Theophyllinenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|theophylline|Drug|false|false||theophylline
null|theophylline|Drug|false|false||theophyllinenull|Assay of theophylline|Procedure|false|false||theophyllinenull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false|C0230028;C0226896|by mouthnull|Oral cavity|Anatomy|false|false|C1527415|mouth
null|Oral region|Anatomy|false|false|C1527415|mouthnull|Twice a day|Time|false|false||twice a daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|PRSS30P gene|Finding|false|false||Dispnull|Dispense (activity)|Event|false|false||Dispnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|cefpodoxime proxetil|Drug|false|false||Cefpodoxime Proxetil
null|cefpodoxime proxetil|Drug|false|false||Cefpodoxime Proxetilnull|cefpodoxime|Drug|false|false||Cefpodoxime
null|cefpodoxime|Drug|false|false||Cefpodoximenull|Every twelve hours|Time|false|false||Q12Hnull|Duration brand of oxymetazoline|Drug|false|false||Durationnull|Duration (temporal concept)|Time|false|false||Durationnull|2 Days|Time|false|false||2 Daysnull|day|Time|false|false||Daysnull|cefpodoxime|Drug|false|false||cefpodoxime
null|cefpodoxime|Drug|false|false||cefpodoximenull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false|C0230028;C0226896|by mouthnull|Oral cavity|Anatomy|false|false|C1561538;C1561539;C1527415|mouth
null|Oral region|Anatomy|false|false|C1561538;C1561539;C1527415|mouthnull|Twice a day|Time|false|false||twice a daynull|Transaction counts and value totals - day|Finding|false|false|C0230028;C0226896|day
null|Precision - day|Finding|false|false|C0230028;C0226896|daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|ferrous sulfate|Drug|false|false||Ferrous Sulfate
null|ferrous sulfate|Drug|false|false||Ferrous Sulfatenull|Ferrous|Drug|false|false||Ferrousnull|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||Sulfate
null|Sulfates, Inorganic|Drug|false|false||Sulfate
null|sulfate ion|Drug|false|false||Sulfate
null|sulfate ion|Drug|false|false||Sulfate
null|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||Sulfatenull|Daily|Time|false|false||DAILYnull|ferrous sulfate|Drug|false|false||ferrous sulfate
null|ferrous sulfate|Drug|false|false||ferrous sulfatenull|Ferrous|Drug|false|false||ferrousnull|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||sulfate
null|Sulfates, Inorganic|Drug|false|false||sulfate
null|sulfate ion|Drug|false|false||sulfate
null|sulfate ion|Drug|false|false||sulfate
null|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||sulfatenull|Iron Drug Class|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|Ferrum metallicum, Homeopathic preparation|Drug|false|false||ironnull|Iron measurement|Procedure|false|false||ironnull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false|C0230028;C0226896|by mouthnull|Oral cavity|Anatomy|false|false|C1527415|mouth
null|Oral region|Anatomy|false|false|C1527415|mouthnull|Daily|Time|false|false||dailynull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|docusate sodium|Drug|false|false||Docusate Sodium
null|docusate sodium|Drug|false|false||Docusate Sodiumnull|docusate|Drug|false|false||Docusate
null|docusate|Drug|false|false||Docusatenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|docusate sodium|Drug|false|false||docusate sodium
null|docusate sodium|Drug|false|false||docusate sodiumnull|docusate|Drug|false|false||docusate
null|docusate|Drug|false|false||docusatenull|Sodium supplements|Drug|false|false||sodium
null|sodium|Drug|false|false||sodium
null|sodium|Drug|false|false||sodium
null|Sodium Drug Class|Drug|false|false||sodiumnull|Sodium metabolic function|Finding|false|false||sodiumnull|Sodium measurement|Procedure|false|false||sodiumnull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0006935|capsule
null|Structure of organ capsule|Anatomy|false|false|C0006935|capsulenull|Capsule Shape|Modifier|false|false||capsulenull|Capsule (unit of presentation)|LabModifier|false|false||capsule
null|Capsule Dosing Unit|LabModifier|false|false||capsulenull|Oral Route of Administration|Finding|false|false|C0230028;C0226896|by mouthnull|Oral cavity|Anatomy|false|false|C1527415|mouth
null|Oral region|Anatomy|false|false|C1527415|mouthnull|Twice a day|Time|false|false||twice a daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0006935|Capsule
null|Structure of organ capsule|Anatomy|false|false|C0006935|Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|refill|Finding|false|false||Refillsnull|polyethylene glycols|Drug|false|false||Polyethylene Glycol
null|polyethylene glycols|Drug|false|false||Polyethylene Glycolnull|high-density polyethylene|Drug|false|false||Polyethylene
null|high-density polyethylene|Drug|false|false||Polyethylene
null|polyethylenes|Drug|false|false||Polyethylene
null|polyethylenes|Drug|false|false||Polyethylene
null|Polyethylene|Drug|false|false||Polyethylene
null|Polyethylene|Drug|false|false||Polyethylenenull|ethylene glycol|Drug|false|false||Glycol
null|Glycol|Drug|false|false||Glycol
null|ethylene glycol|Drug|false|false||Glycol
null|Glycols|Drug|false|false||Glycolnull|Daily|Time|false|false||DAILYnull|polyethylene glycol 3350|Drug|false|false||polyethylene glycol 3350
null|polyethylene glycol 3350|Drug|false|false||polyethylene glycol 3350null|polyethylene glycols|Drug|false|false||polyethylene glycol
null|polyethylene glycols|Drug|false|false||polyethylene glycolnull|high-density polyethylene|Drug|false|false||polyethylene
null|high-density polyethylene|Drug|false|false||polyethylene
null|polyethylenes|Drug|false|false||polyethylene
null|polyethylenes|Drug|false|false||polyethylene
null|Polyethylene|Drug|false|false||polyethylene
null|Polyethylene|Drug|false|false||polyethylenenull|ethylene glycol|Drug|false|false||glycol
null|Glycol|Drug|false|false||glycol
null|ethylene glycol|Drug|false|false||glycol
null|Glycols|Drug|false|false||glycolnull|gram|LabModifier|false|false||gramnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Powder dose form|Drug|false|false||powder
null|powder physical state|Drug|false|false||powdernull|Oral Route of Administration|Finding|false|false|C0230028;C0226896|by mouthnull|Oral cavity|Anatomy|false|false|C1527415|mouth
null|Oral region|Anatomy|false|false|C1527415|mouthnull|Daily|Time|false|false||dailynull|refill|Finding|false|false||Refillsnull|ipratropium bromide|Drug|false|false||Ipratropium Bromide
null|ipratropium bromide|Drug|false|false||Ipratropium Bromidenull|ipratropium|Drug|false|false||Ipratropium
null|ipratropium|Drug|false|false||Ipratropiumnull|Bromides|Drug|false|false||Bromidenull|Bromides measurement|Procedure|false|false||Bromidenull|NEB protein, human|Drug|false|false||Neb
null|NEB protein, human|Drug|false|false||Neb
null|Nebulizer solution|Drug|false|false||Nebnull|NEB gene|Finding|false|false||Neb
null|mitotic nuclear membrane disassembly|Finding|false|false||Nebnull|NEB protein, human|Drug|false|false||NEB
null|NEB protein, human|Drug|false|false||NEB
null|Nebulizer solution|Drug|false|false||NEBnull|NEB gene|Finding|false|false||NEB
null|mitotic nuclear membrane disassembly|Finding|false|false||NEBnull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|null|Finding|false|false||dyspnea
null|Dyspnea|Finding|false|false||dyspneanull|Wheezing|Finding|false|false||wheezingnull|ipratropium bromide|Drug|false|false||ipratropium bromide
null|ipratropium bromide|Drug|false|false||ipratropium bromidenull|ipratropium|Drug|false|false||ipratropium
null|ipratropium|Drug|false|false||ipratropiumnull|Bromides|Drug|false|false||bromidenull|Bromides measurement|Procedure|false|false||bromidenull|Kilogram per Cubic Meter|LabModifier|false|false||mg/mLnull|per milliliter|LabModifier|false|false||/mLnull|NEB protein, human|Drug|false|false||neb
null|NEB protein, human|Drug|false|false||neb
null|Nebulizer solution|Drug|false|false||nebnull|NEB gene|Finding|false|false||neb
null|mitotic nuclear membrane disassembly|Finding|false|false||nebnull|Inhalant dose form|Drug|false|false||INH
null|isoniazid|Drug|false|false||INH
null|isoniazid|Drug|false|false||INHnull|Inhalation Route of Administration|Finding|false|false||INHnull|Ingush language|Entity|false|false||INHnull|Inhalation Dosing Unit|LabModifier|false|false||INHnull|Every - dosing instruction fragment|Finding|false|false||Everynull|Every (qualifier)|Modifier|false|false||Everynull|Hour|Time|false|false||hoursnull|Nebule Dosing Unit|LabModifier|false|false||Nebulenull|refill|Finding|false|false||Refillsnull|prednisone|Drug|false|false||PredniSONE
null|prednisone|Drug|false|false||PredniSONE
null|prednisone|Drug|false|false||PredniSONEnull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|Continuous|Finding|false|false||ongoingnull|null|Procedure|false|false||Taperednull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|prednisone|Drug|false|false||prednisone
null|prednisone|Drug|false|false||prednisone
null|prednisone|Drug|false|false||prednisonenull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false|C0230028;C0226896|by mouthnull|Oral cavity|Anatomy|false|false|C1527415|mouth
null|Oral region|Anatomy|false|false|C1527415|mouthnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|ADMIN.FACILITY|Finding|false|false||Facilitynull|Facility (object)|Device|false|false||Facilitynull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Chronic Obstructive Airway Disease|Disorder|false|false|C0024109|Chronic obstructive pulmonary diseasenull|Chronic - Admission Level of Care Code|Finding|false|false||Chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||Chronicnull|chronic|Time|false|false||Chronicnull|Lung Diseases, Obstructive|Disorder|false|false|C0024109|obstructive pulmonary diseasenull|Obstructed|Finding|false|false||obstructivenull|Lung diseases|Disorder|false|false|C0024109|pulmonary diseasenull|History of - respiratory disease|Finding|false|false|C0024109|pulmonary diseasenull|Pulmonary (intended site)|Finding|false|false|C0024109|pulmonarynull|Lung|Anatomy|false|false|C2707265;C0455540;C0024117;C0012634;C0600260;C4522268;C0024115|pulmonarynull|null|Attribute|false|false|C0024109|pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Disease|Disorder|false|false|C0024109|diseasenull|Atrial fibrillation with rapid ventricular response|Disorder|false|false|C0018827;C0018792|Atrial fibrillation with rapid ventricular responsenull|continuous electrocardiogram monitoring atrial fibrillation with rapid ventricular response|Procedure|false|false|C0018827;C0018792|Atrial fibrillation with rapid ventricular responsenull|Atrial Fibrillation|Disorder|false|false|C0018792|Atrial fibrillationnull|null|Attribute|false|false|C0018792|Atrial fibrillationnull|Atrial Fibrillation by ECG Finding|Lab|false|false|C0018792|Atrial fibrillationnull|Heart Atrium|Anatomy|false|false|C2926591;C3853730;C0232197;C1142306;C0004238;C0344434|Atrialnull|Fibrillation|Disorder|false|false|C0018792|fibrillationnull|rapid ventricular response|Disorder|false|false|C0018827|rapid ventricular responsenull|Rapid|Modifier|false|false||rapidnull|Heart Ventricle|Anatomy|false|false|C0748243;C3853730;C1142306|ventricularnull|Ventricular|Modifier|false|false||ventricularnull|Communication Response|Finding|false|false||response
null|Disease Response|Finding|false|false||response
null|Answer (statement)|Finding|false|false||responsenull|Response process|Subject|false|false||responsenull|Neoplasm Metastasis|Disorder|false|false||Secondarynull|metastatic qualifier|Finding|false|false||Secondarynull|Secondary to|Modifier|false|false||Secondarynull|second (number)|LabModifier|false|false||Secondarynull|Diagnosis|Procedure|false|false||diagnosesnull|Hypertensive disease|Disorder|false|false||Hypertensionnull|Coronary Artery Disease|Disorder|false|false|C0018787;C0226004;C0003842;C0205042|Coronary artery disease
null|Coronary Arteriosclerosis|Disorder|false|false|C0018787;C0226004;C0003842;C0205042|Coronary artery diseasenull|Coronary artery|Anatomy|false|false|C0012634;C0852949;C1956346;C0010054|Coronary arterynull|Heart|Anatomy|false|false|C1956346;C0010054|Coronarynull|Coronary|Modifier|false|false||Coronarynull|Arteriopathic disease|Disorder|false|false|C0226004;C0003842;C0205042|artery diseasenull|Arterial system|Anatomy|false|false|C0012634;C1956346;C0010054;C0852949|artery
null|Arteries|Anatomy|false|false|C0012634;C1956346;C0010054;C0852949|arterynull|Disease|Disorder|false|false|C0226004;C0003842;C0205042|diseasenull|Peripheral Vascular Diseases|Disorder|false|false|C0005847|Peripheral vascular diseasenull|Peripheral|Modifier|false|false||Peripheralnull|Vascular Diseases|Disorder|false|false|C0005847|vascular diseasenull|Blood Vessel|Anatomy|false|false|C0012634;C0042373;C0085096|vascularnull|Vascular|Modifier|false|false||vascularnull|Disease|Disorder|false|false|C0005847|diseasenull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Coordination of Benefits - Independent|Finding|false|false||Independent
null|Religious Affiliation - Independent|Finding|false|false||Independent
null|Independence|Finding|false|false||Independent
null|Independently able|Finding|false|false||Independentnull|FBXW7-AS1 gene|Finding|false|false||Dearnull|Respiratory distress|Finding|false|false||difficulty breathing
null|Dyspnea|Finding|false|false||difficulty breathingnull|Has difficulty doing (qualifier value)|Finding|false|false||difficultynull|outcomes otolaryngology breathing|Finding|false|false||breathing
null|Inspiration (function)|Finding|false|false||breathing
null|Respiration|Finding|false|false||breathingnull|null|Attribute|false|false||breathingnull|respiratory system process|Phenomenon|false|false||breathingnull|Clinic|Device|false|false||clinic
null|Ambulatory Care Facilities|Device|false|false||clinicnull|Clinic|Entity|false|false||clinic
null|Ambulatory Care Facilities|Entity|false|false||clinicnull|Patient location type - Clinic|Modifier|false|false||clinic
null|Person location type - Clinic|Modifier|false|false||clinicnull|Tachycardia|Finding|false|false|C4037974;C0018787|fast heart ratenull|Fas-activated serine/threonine kinase activity|Finding|false|false||fast
null|FASTK Gene|Finding|false|false||fast
null|FOXD3-AS1 gene|Finding|false|false||fast
null|FASTK wt Allele|Finding|false|false||fast
null|Fasting|Finding|false|false||fastnull|Rapid|Modifier|false|false||fastnull|null|Finding|false|false|C4037974;C0018787|heart ratenull|examination of heart rate|Procedure|false|false|C4037974;C0018787|heart ratenull|heart rate|Attribute|false|false|C4037974;C0018787|heart rate
null|null|Attribute|false|false|C4037974;C0018787|heart ratenull|Mean Heart Rate|LabModifier|false|false||heart ratenull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787|heart
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787|heartnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|heartnull|Chest>Heart|Anatomy|false|false|C0018810;C0488794;C0153957;C0153500;C0039231;C2041121;C1549480;C2197023;C0795691|heart
null|Heart|Anatomy|false|false|C0018810;C0488794;C0153957;C0153500;C0039231;C2041121;C1549480;C2197023;C0795691|heartnull|Amount type - Rate|Finding|false|false|C4037974;C0018787|ratenull|Rating (action)|Event|false|false||ratenull|Rate|LabModifier|false|false||ratenull|Respiratory distress|Finding|false|false||difficulty breathing
null|Dyspnea|Finding|false|false||difficulty breathingnull|Has difficulty doing (qualifier value)|Finding|false|false||difficultynull|outcomes otolaryngology breathing|Finding|false|false||breathing
null|Inspiration (function)|Finding|false|false||breathing
null|Respiration|Finding|false|false||breathingnull|null|Attribute|false|false||breathingnull|respiratory system process|Phenomenon|false|false||breathingnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|Tachycardia|Finding|false|false|C4037974;C0018787|fast heart ratenull|Fas-activated serine/threonine kinase activity|Finding|false|false||fast
null|FASTK Gene|Finding|false|false||fast
null|FOXD3-AS1 gene|Finding|false|false||fast
null|FASTK wt Allele|Finding|false|false||fast
null|Fasting|Finding|false|false||fastnull|Rapid|Modifier|false|false||fastnull|null|Finding|false|false|C4037974;C0018787|heart ratenull|examination of heart rate|Procedure|false|false|C4037974;C0018787|heart ratenull|heart rate|Attribute|false|false|C4037974;C0018787|heart rate
null|null|Attribute|false|false|C4037974;C0018787|heart ratenull|Mean Heart Rate|LabModifier|false|false||heart ratenull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787|heart
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787|heartnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|heartnull|Chest>Heart|Anatomy|false|false|C0153957;C0153500;C0039231;C2197023;C0018810;C0488794;C0795691;C2041121|heart
null|Heart|Anatomy|false|false|C0153957;C0153500;C0039231;C2197023;C0018810;C0488794;C0795691;C2041121|heartnull|Amount type - Rate|Finding|false|false||ratenull|Rating (action)|Event|false|false||ratenull|Rate|LabModifier|false|false||ratenull|Atrial Fibrillation|Disorder|false|false|C0018792|atrial fibrillationnull|null|Attribute|false|false|C0018792|atrial fibrillationnull|Atrial Fibrillation by ECG Finding|Lab|false|false|C0018792|atrial fibrillationnull|Heart Atrium|Anatomy|false|false|C0232197;C0344434;C2926591;C0004238|atrialnull|Fibrillation|Disorder|false|false|C0018792|fibrillationnull|Irregular heart beat|Finding|false|false|C4037974;C0018787|irregular heart ratenull|Irregular|Modifier|false|false||irregularnull|null|Finding|false|false|C4037974;C0018787|heart ratenull|examination of heart rate|Procedure|false|false|C4037974;C0018787|heart ratenull|heart rate|Attribute|false|false|C4037974;C0018787|heart rate
null|null|Attribute|false|false|C4037974;C0018787|heart ratenull|Mean Heart Rate|LabModifier|false|false||heart ratenull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787|heart
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787|heartnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|heartnull|Chest>Heart|Anatomy|false|false|C0237314;C0795691;C2197023;C0153957;C0153500;C0018810;C0488794;C2041121;C1549480|heart
null|Heart|Anatomy|false|false|C0237314;C0795691;C2197023;C0153957;C0153500;C0018810;C0488794;C2041121;C1549480|heartnull|Amount type - Rate|Finding|false|false|C4037974;C0018787|ratenull|Rating (action)|Event|false|false||ratenull|Rate|LabModifier|false|false||ratenull|Sometimes|Time|false|false||sometimesnull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787|heart
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787|heartnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|heartnull|Chest>Heart|Anatomy|false|false|C0795691;C0153957;C0153500|heart
null|Heart|Anatomy|false|false|C0795691;C0153957;C0153500|heartnull|Very|Modifier|false|false||verynull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|theophylline|Drug|false|false||theophylline
null|theophylline|Drug|false|false||theophyllinenull|Assay of theophylline|Procedure|false|false||theophyllinenull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|null|Finding|false|false|C4037974;C0018787|heart ratenull|examination of heart rate|Procedure|false|false|C4037974;C0018787|heart ratenull|heart rate|Attribute|false|false|C4037974;C0018787|heart rate
null|null|Attribute|false|false|C4037974;C0018787|heart ratenull|Mean Heart Rate|LabModifier|false|false||heart ratenull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787|heart
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787|heartnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|heartnull|Chest>Heart|Anatomy|false|false|C0795691;C0153957;C0153500;C1549480;C2041121;C2197023;C0018810;C0488794|heart
null|Heart|Anatomy|false|false|C0795691;C0153957;C0153500;C1549480;C2041121;C2197023;C0018810;C0488794|heartnull|Amount type - Rate|Finding|false|false|C4037974;C0018787|ratenull|Rating (action)|Event|false|false||ratenull|Rate|LabModifier|false|false||ratenull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|At home|Finding|false|false||at homenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|diltiazem|Drug|false|false||diltiazem
null|diltiazem|Drug|false|false||diltiazemnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Cold brand of chlorpheniramine-phenylpropanolamine|Drug|false|false||cold
null|Cold brand of chlorpheniramine-phenylpropanolamine|Drug|false|false||coldnull|Common Cold|Disorder|false|false||cold
null|Chronic Obstructive Airway Disease|Disorder|false|false||coldnull|Cold Sensation|Finding|false|false||coldnull|Cold Therapy|Procedure|false|false||coldnull|Cold Temperature|Phenomenon|false|false||coldnull|Flare|Finding|false|false||flare
null|Exacerbation of cGVHD|Finding|false|false||flarenull|Very|Modifier|false|false||verynull|Equipment Alert Level - Serious|Finding|false|false||serious
null|Device Alert Level - Serious|Finding|false|false||serious
null|Alert level - Serious|Finding|false|false||seriousnull|Serious|Modifier|false|false||seriousnull|Steroids|Drug|false|false||steroids
null|Steroids|Drug|false|false||steroidsnull|Inspiration (function)|Finding|false|false||inhalednull|Therapeutic procedure|Procedure|false|false||treatmentsnull|Lung diseases|Disorder|false|false|C4037972;C0024109|lungnull|Lung Problem|Finding|false|false|C4037972;C0024109|lungnull|Chest>Lung|Anatomy|false|false|C0024115;C0740941|lung
null|Lung|Anatomy|false|false|C0024115;C0740941|lungnull|Physicians|Subject|false|false||doctorsnull|Pulmonary (intended site)|Finding|false|false|C0024109|pulmonarynull|Lung|Anatomy|false|false|C2707265;C4522268|pulmonarynull|null|Attribute|false|false|C0024109|pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Rehabilitation therapy|Procedure|false|false||rehabnull|SURE Test|Finding|false|false||surenull|Certain (qualifier value)|Modifier|false|false||surenull|Lung diseases|Disorder|false|false|C4037972;C0024109|lung diseasenull|Lung diseases|Disorder|false|false|C4037972;C0024109|lungnull|Lung Problem|Finding|false|false|C4037972;C0024109|lungnull|Chest>Lung|Anatomy|false|false|C0024115;C0024115;C0740941|lung
null|Lung|Anatomy|false|false|C0024115;C0024115;C0740941|lungnull|Disease|Disorder|false|false||diseasenull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Possible|Finding|false|false||possiblenull|Possibly Related to Intervention|Modifier|false|false||possible
null|Possible diagnosis|Modifier|false|false||possiblenull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Often - answer to question|Finding|false|false||oftennull|Frequently|Time|false|false||oftennull|Appointments|Event|false|false||appointmentnull|Production Class Code - Pleasure|Finding|false|false||pleasure
null|pleasurable emotion|Finding|false|false||pleasurenull|Pleasure - Animals raised for recreation|Entity|false|false||pleasurenull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Vitelliform Macular Dystrophy|Disorder|false|false||bestnull|BEST1 wt Allele|Finding|false|false||best
null|BEST1 gene|Finding|false|false||bestnull|best (quality)|Modifier|false|false||bestnull|Future|Time|false|false||futurenull|Team|Subject|false|false||teamnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions