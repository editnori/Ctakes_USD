 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|22,26
No|27,29
:|29,30
_|33,34
_|34,35
_|35,36
<EOL>|36,37
<EOL>|38,39
Admission|39,48
Date|49,53
:|53,54
_|56,57
_|57,58
_|58,59
Discharge|73,82
Date|83,87
:|87,88
_|91,92
_|92,93
_|93,94
<EOL>|94,95
<EOL>|96,97
Date|97,101
of|102,104
Birth|105,110
:|110,111
_|113,114
_|114,115
_|115,116
Sex|129,132
:|132,133
F|136,137
<EOL>|137,138
<EOL>|139,140
Service|140,147
:|147,148
MEDICINE|149,157
<EOL>|157,158
<EOL>|159,160
No|172,174
Known|175,180
Allergies|181,190
/|191,192
Adverse|193,200
Drug|201,205
Reactions|206,215
<EOL>|215,216
<EOL>|217,218
Attending|218,227
:|227,228
_|229,230
_|230,231
_|231,232
.|232,233
<EOL>|233,234
<EOL>|235,236
Dyspnea|253,260
and|261,264
chest|265,270
tightness|271,280
<EOL>|280,281
<EOL>|282,283
Major|283,288
Surgical|289,297
or|298,300
Invasive|301,309
Procedure|310,319
:|319,320
<EOL>|320,321
_|321,322
_|322,323
_|323,324
Pharmacologic|325,338
nuclear|339,346
stress|347,353
test|354,358
<EOL>|358,359
<EOL>|360,361
_|389,390
_|390,391
_|391,392
year|393,397
old|398,401
female|402,408
with|409,413
history|414,421
of|422,424
HTN|425,428
,|428,429
HLD|430,433
,|433,434
hx|435,437
of|438,440
CVA|441,444
,|444,445
CAD|446,449
s|450,451
/|451,452
p|452,453
<EOL>|454,455
BMS|455,458
to|459,461
circumflex|462,472
and|473,476
POBA|477,481
(|482,483
_|483,484
_|484,485
_|485,486
)|486,487
,|487,488
on|489,491
Aspirin|492,499
and|500,503
Plavix|504,510
,|510,511
CHF|512,515
<EOL>|516,517
(|517,518
EF|518,520
45|521,523
%|523,524
in|525,527
_|528,529
_|529,530
_|530,531
,|531,532
diabetes|533,541
,|541,542
presenting|543,553
with|554,558
acute|559,564
onset|565,570
<EOL>|571,572
shortness|572,581
of|582,584
breath|585,591
and|592,595
substernal|596,606
chest|607,612
tightness|613,622
since|623,628
_|629,630
_|630,631
_|631,632
<EOL>|633,634
evening|634,641
.|641,642
<EOL>|643,644
<EOL>|644,645
Patient|645,652
notes|653,658
that|659,663
_|664,665
_|665,666
_|666,667
evening|668,675
had|676,679
a|680,681
large|682,687
seafood|688,695
dinner|696,702
<EOL>|703,704
which|704,709
is|710,712
not|713,716
usual|717,722
for|723,726
her|727,730
,|730,731
and|732,735
then|736,740
later|741,746
around|747,753
10pm|754,758
had|759,762
acute|763,768
<EOL>|769,770
onset|770,775
of|776,778
SOB|779,782
feeling|783,790
like|791,795
she|796,799
could|800,805
not|806,809
take|810,814
deep|815,819
breaths|820,827
with|828,832
<EOL>|833,834
chest|834,839
tightness|840,849
(|850,851
patient|851,858
notes|859,864
this|865,869
is|870,872
her|873,876
"|877,878
angina|878,884
"|884,885
)|885,886
.|886,887
Denies|888,894
<EOL>|895,896
pleuritic|896,905
component|906,915
to|916,918
CP|919,921
,|921,922
described|923,932
as|933,935
central|936,943
and|944,947
across|948,954
lower|955,960
<EOL>|961,962
rib|962,965
cage|966,970
,|970,971
persistent|972,982
since|983,988
onset|989,994
,|994,995
no|996,998
radiation|999,1008
to|1009,1011
the|1012,1015
<EOL>|1016,1017
shoulders|1017,1026
/|1026,1027
jaw|1027,1030
/|1030,1031
back|1031,1035
,|1035,1036
no|1037,1039
diaphoreses|1040,1051
.|1051,1052
Worsens|1053,1060
with|1061,1065
activity|1066,1074
,|1074,1075
<EOL>|1076,1077
improves|1077,1085
somewhat|1086,1094
with|1095,1099
rest|1100,1104
.|1104,1105
Patient|1106,1113
does|1114,1118
not|1119,1122
it|1123,1125
feels|1126,1131
like|1132,1136
<EOL>|1137,1138
other|1138,1143
episodes|1144,1152
when|1153,1157
she|1158,1161
then|1162,1166
required|1167,1175
her|1176,1179
stent|1180,1185
placement|1186,1195
.|1195,1196
Took|1197,1201
<EOL>|1202,1203
a|1203,1204
SLNx1|1205,1210
,|1210,1211
which|1212,1217
improved|1218,1226
her|1227,1230
symptoms|1231,1239
though|1240,1246
these|1247,1252
persisted|1253,1262
,|1262,1263
but|1264,1267
<EOL>|1268,1269
almost|1269,1275
immediately|1276,1287
led|1288,1291
to|1292,1294
abdominal|1295,1304
discomfort|1305,1315
with|1316,1320
vomiting|1321,1329
x1|1330,1332
,|1332,1333
<EOL>|1334,1335
nonbloody|1335,1344
with|1345,1349
dinner|1350,1356
pieces|1357,1363
.|1363,1364
_|1365,1366
_|1366,1367
_|1367,1368
,|1368,1369
1|1370,1371
day|1372,1375
prior|1376,1381
to|1382,1384
admission|1385,1394
,|1394,1395
<EOL>|1396,1397
decided|1397,1404
to|1405,1407
see|1408,1411
if|1412,1414
her|1415,1418
pain|1419,1423
improved|1424,1432
on|1433,1435
its|1436,1439
own|1440,1443
,|1443,1444
then|1445,1449
when|1450,1454
it|1455,1457
<EOL>|1458,1459
persisted|1459,1468
on|1469,1471
_|1472,1473
_|1473,1474
_|1474,1475
,|1475,1476
husband|1477,1484
arranged|1485,1493
for|1494,1497
UC|1498,1500
appt|1501,1505
at|1506,1508
_|1509,1510
_|1510,1511
_|1511,1512
<EOL>|1513,1514
_|1514,1515
_|1515,1516
_|1516,1517
.|1517,1518
At|1519,1521
PCP|1522,1525
,|1525,1526
_|1527,1528
_|1528,1529
_|1529,1530
,|1530,1531
SBP|1532,1535
up|1536,1538
to|1539,1541
200s|1542,1546
,|1546,1547
EKG|1548,1551
with|1552,1556
ST|1557,1559
<EOL>|1560,1561
depressions|1561,1572
in|1573,1575
the|1576,1579
precordial|1580,1590
leads|1591,1596
,|1596,1597
specifically|1598,1610
V3|1611,1613
,|1613,1614
V4|1615,1617
and|1618,1621
V5|1622,1624
,|1624,1625
<EOL>|1626,1627
given|1627,1632
full|1633,1637
dose|1638,1642
ASA|1643,1646
and|1647,1650
SLNx1|1651,1656
,|1656,1657
and|1658,1661
sent|1662,1666
to|1667,1669
the|1670,1673
ED|1674,1676
given|1677,1682
concern|1683,1690
<EOL>|1691,1692
for|1692,1695
ACS|1696,1699
versus|1700,1706
HTN|1707,1710
emergency|1711,1720
.|1720,1721
<EOL>|1722,1723
<EOL>|1723,1724
Patient|1724,1731
reporting|1732,1741
baseline|1742,1750
sleeps|1751,1757
with|1758,1762
2|1763,1764
pillows|1765,1772
,|1772,1773
unchanged|1774,1783
<EOL>|1784,1785
recently|1785,1793
,|1793,1794
no|1795,1797
cough|1798,1803
,|1803,1804
PND|1805,1808
,|1808,1809
orthopnea|1810,1819
with|1820,1824
2|1825,1826
pillows|1827,1834
.|1834,1835
Worsening|1836,1845
DOE|1846,1849
<EOL>|1850,1851
since|1851,1856
onset|1857,1862
of|1863,1865
symptoms|1866,1874
,|1874,1875
now|1876,1879
unable|1880,1886
to|1887,1889
complete|1890,1898
a|1899,1900
block|1901,1906
where|1907,1912
<EOL>|1913,1914
she|1914,1917
used|1918,1922
to|1923,1925
be|1926,1928
able|1929,1933
to|1934,1936
walk|1937,1941
a|1942,1943
few|1944,1947
blocks|1948,1954
at|1955,1957
a|1958,1959
time|1960,1964
without|1965,1972
<EOL>|1973,1974
stopping|1974,1982
_|1983,1984
_|1984,1985
_|1985,1986
SOB|1987,1990
/|1990,1991
CP|1991,1993
.|1993,1994
Denies|1995,2001
new|2002,2005
_|2006,2007
_|2007,2008
_|2008,2009
edema|2010,2015
(|2016,2017
baseline|2017,2025
says|2026,2030
L|2031,2032
leg|2033,2036
>|2037,2038
<EOL>|2039,2040
R|2040,2041
)|2041,2042
.|2042,2043
<EOL>|2043,2044
<EOL>|2044,2045
Also|2045,2049
had|2050,2053
emesis|2054,2060
last|2061,2065
night|2066,2071
x|2072,2073
1|2074,2075
;|2075,2076
no|2077,2079
diaphoresis|2080,2091
,|2091,2092
no|2093,2095
chest|2096,2101
pain|2102,2106
,|2106,2107
<EOL>|2108,2109
no|2109,2111
radiation|2112,2121
of|2122,2124
symptoms|2125,2133
anywhere|2134,2142
.|2142,2143
No|2144,2146
diarrhea|2147,2155
or|2156,2158
constipation|2159,2171
,|2171,2172
<EOL>|2173,2174
no|2174,2176
dysuria|2177,2184
,|2184,2185
no|2186,2188
focal|2189,2194
weakness|2195,2203
/|2203,2204
numbness|2204,2212
.|2212,2213
On|2214,2216
ROS|2217,2220
,|2220,2221
also|2222,2226
with|2227,2231
some|2232,2236
L|2237,2238
<EOL>|2239,2240
leg|2240,2243
tingling|2244,2252
intermittently|2253,2267
,|2267,2268
stable|2269,2275
and|2276,2279
chronic|2280,2287
.|2287,2288
Had|2289,2292
diarrhea|2293,2301
x1|2302,2304
<EOL>|2305,2306
on|2306,2308
_|2309,2310
_|2310,2311
_|2311,2312
following|2313,2322
_|2323,2324
_|2324,2325
_|2325,2326
seafood|2327,2334
dinner|2335,2341
,|2341,2342
normal|2343,2349
BMs|2350,2353
since|2354,2359
<EOL>|2360,2361
then|2361,2365
.|2365,2366
<EOL>|2367,2368
<EOL>|2369,2370
In|2370,2372
the|2373,2376
ED|2377,2379
initial|2380,2387
vital|2388,2393
signs|2394,2399
;|2399,2400
T|2401,2402
98|2403,2405
P|2406,2407
88|2408,2410
BP|2411,2413
190|2414,2417
/|2417,2418
120|2418,2421
R|2422,2423
18|2424,2426
O2|2427,2429
Sat|2430,2433
<EOL>|2434,2435
98|2435,2437
%|2437,2438
3L|2439,2441
nasal|2442,2447
cannula|2448,2455
.|2455,2456
Labs|2457,2461
notable|2462,2469
for|2470,2473
Cr|2474,2476
2.1|2477,2480
(|2481,2482
baseline|2482,2490
<EOL>|2491,2492
2.1|2492,2495
-|2495,2496
2.7|2496,2499
)|2499,2500
,|2500,2501
BUN|2502,2505
29|2506,2508
.|2508,2509
wbc|2510,2513
4.3|2514,2517
,|2517,2518
H|2519,2520
/|2520,2521
H|2521,2522
8.6|2523,2526
/|2526,2527
26|2527,2529
.|2529,2530
0|2530,2531
,|2531,2532
Plt|2533,2536
147|2537,2540
.|2540,2541
Initial|2542,2549
and|2550,2553
<EOL>|2554,2555
rpt|2555,2558
Tn|2559,2561
<|2562,2563
0.01|2563,2567
.|2567,2568
BNP|2569,2572
4279|2573,2577
.|2577,2578
CXR|2579,2582
showed|2583,2589
no|2590,2592
pulmonary|2593,2602
edema|2603,2608
,|2608,2609
pleural|2610,2617
<EOL>|2618,2619
effusions|2619,2628
,|2628,2629
or|2630,2632
consolidation|2633,2646
,|2646,2647
borderline|2648,2658
cardiomegaly|2659,2671
.|2671,2672
The|2673,2676
<EOL>|2677,2678
patient|2678,2685
received|2686,2694
carvedilol|2695,2705
,|2705,2706
nebulizers|2707,2717
,|2717,2718
and|2719,2722
IV|2723,2725
lasix|2726,2731
.|2731,2732
It|2733,2735
is|2736,2738
<EOL>|2739,2740
unclear|2740,2747
how|2748,2751
much|2752,2756
UOP|2757,2760
the|2761,2764
patient|2765,2772
has|2773,2776
as|2777,2779
it|2780,2782
was|2783,2786
not|2787,2790
documented|2791,2801
in|2802,2804
<EOL>|2805,2806
the|2806,2809
ED|2810,2812
.|2812,2813
<EOL>|2814,2815
<EOL>|2815,2816
The|2816,2819
patient|2820,2827
was|2828,2831
seen|2832,2836
by|2837,2839
cardiology|2840,2850
in|2851,2853
the|2854,2857
ED|2858,2860
who|2861,2864
felt|2865,2869
that|2870,2874
in|2875,2877
<EOL>|2878,2879
the|2879,2882
setting|2883,2890
of|2891,2893
systolic|2894,2902
heart|2903,2908
failure|2909,2916
,|2916,2917
her|2918,2921
dyspnea|2922,2929
was|2930,2933
likely|2934,2940
<EOL>|2941,2942
due|2942,2945
to|2946,2948
a|2949,2950
CHF|2951,2954
exacerbation|2955,2967
in|2968,2970
the|2971,2974
setting|2975,2982
of|2983,2985
dietary|2986,2993
<EOL>|2994,2995
indiscretion|2995,3007
.|3007,3008
Diuresis|3009,3017
was|3018,3021
recommended|3022,3033
in|3034,3036
addition|3037,3045
to|3046,3048
increasing|3049,3059
<EOL>|3060,3061
carvedilol|3061,3071
to|3072,3074
12.5|3075,3079
mg|3079,3081
BID|3082,3085
,|3085,3086
as|3087,3089
well|3090,3094
as|3095,3097
a|3098,3099
nuclear|3100,3107
stress|3108,3114
test|3115,3119
this|3120,3124
<EOL>|3125,3126
morning|3126,3133
.|3133,3134
<EOL>|3134,3135
<EOL>|3135,3136
On|3136,3138
the|3139,3142
floor|3143,3148
,|3148,3149
the|3150,3153
patient|3154,3161
c|3162,3163
/|3163,3164
o|3164,3165
of|3166,3168
some|3169,3173
improved|3174,3182
dyspnea|3183,3190
/|3190,3191
chest|3191,3196
<EOL>|3197,3198
tightness|3198,3207
as|3208,3210
well|3211,3215
as|3216,3218
wheezing|3219,3227
(|3228,3229
no|3229,3231
COPD|3232,3236
/|3236,3237
asthma|3237,3243
history|3244,3251
,|3251,3252
no|3253,3255
<EOL>|3256,3257
significant|3257,3268
smoking|3269,3276
history|3277,3284
)|3284,3285
,|3285,3286
but|3287,3290
otherwise|3291,3300
has|3301,3304
no|3305,3307
acute|3308,3313
<EOL>|3314,3315
complaints|3315,3325
.|3325,3326
Given|3327,3332
her|3333,3336
continued|3337,3346
SOB|3347,3350
and|3351,3354
wheezing|3355,3363
,|3363,3364
she|3365,3368
was|3369,3372
<EOL>|3373,3374
written|3374,3381
for|3382,3385
nebulizers|3386,3396
and|3397,3400
steroids|3401,3409
for|3410,3413
reactive|3414,3422
airway|3423,3429
disease|3430,3437
<EOL>|3438,3439
overnight|3439,3448
.|3448,3449
<EOL>|3449,3450
<EOL>|3451,3452
-|3474,3475
hypertension|3476,3488
<EOL>|3490,3491
-|3491,3492
diabetes|3493,3501
<EOL>|3503,3504
-|3504,3505
hx|3506,3508
CVA|3509,3512
(|3513,3514
cerebellar|3514,3524
-|3524,3525
medullary|3525,3534
stroke|3535,3541
in|3542,3544
_|3545,3546
_|3546,3547
_|3547,3548
<EOL>|3550,3551
-|3551,3552
CAD|3553,3556
(|3557,3558
hx|3558,3560
of|3561,3563
MI|3564,3566
in|3567,3569
_|3570,3571
_|3571,3572
_|3572,3573
BMS|3574,3577
to|3578,3580
circumflex|3581,3591
and|3592,3595
POBA|3596,3600
_|3601,3602
_|3602,3603
_|3603,3604
<EOL>|3606,3607
-|3607,3608
peripheral|3609,3619
arterial|3620,3628
disease|3629,3636
-|3636,3637
claudication|3638,3650
,|3650,3651
followed|3652,3660
by|3661,3663
<EOL>|3664,3665
vascular|3665,3673
,|3673,3674
managed|3675,3682
conservatively|3683,3697
<EOL>|3697,3698
-|3698,3699
stage|3700,3705
IV|3706,3708
CKD|3709,3712
(|3713,3714
baseline|3714,3722
2.1|3723,3726
-|3726,3727
2.6|3727,3730
)|3730,3731
<EOL>|3733,3734
-|3734,3735
GERD|3736,3740
/|3740,3741
esophageal|3741,3751
rings|3752,3757
<EOL>|3757,3758
<EOL>|3759,3760
:|3774,3775
<EOL>|3775,3776
_|3776,3777
_|3777,3778
_|3778,3779
<EOL>|3779,3780
:|3794,3795
<EOL>|3795,3796
Niece|3796,3801
had|3802,3805
some|3806,3810
sort|3811,3815
of|3816,3818
cancer|3819,3825
.|3825,3826
Father|3827,3833
died|3834,3838
in|3839,3841
his|3842,3845
_|3846,3847
_|3847,3848
_|3848,3849
due|3850,3853
to|3854,3856
<EOL>|3857,3858
lung|3858,3862
disease|3863,3870
.|3870,3871
Mother|3873,3879
died|3880,3884
in|3885,3887
her|3888,3891
_|3892,3893
_|3893,3894
_|3894,3895
due|3896,3899
to|3900,3902
an|3903,3905
unknown|3906,3913
cause|3914,3919
.|3919,3920
<EOL>|3922,3923
No|3923,3925
early|3926,3931
CAD|3932,3935
or|3936,3938
sudden|3939,3945
cardiac|3946,3953
death|3954,3959
.|3959,3960
No|3961,3963
other|3964,3969
known|3970,3975
history|3976,3983
of|3984,3986
<EOL>|3987,3988
cancer|3988,3994
.|3994,3995
<EOL>|3995,3996
<EOL>|3997,3998
ADMISSION|4013,4022
PHYSICAL|4023,4031
EXAM|4032,4036
:|4036,4037
<EOL>|4037,4038
=|4038,4039
=|4039,4040
=|4040,4041
=|4041,4042
=|4042,4043
=|4043,4044
=|4044,4045
=|4045,4046
=|4046,4047
=|4047,4048
=|4048,4049
=|4049,4050
=|4050,4051
=|4051,4052
=|4052,4053
=|4053,4054
=|4054,4055
=|4055,4056
=|4056,4057
=|4057,4058
=|4058,4059
=|4059,4060
=|4060,4061
=|4061,4062
=|4062,4063
=|4063,4064
=|4064,4065
<EOL>|4065,4066
Vitals|4066,4072
:|4072,4073
Tm|4074,4076
98|4077,4079
,|4079,4080
Tc|4081,4083
98|4084,4086
,|4086,4087
HR|4088,4090
68|4091,4093
(|4094,4095
68|4095,4097
-|4097,4098
78|4098,4100
)|4100,4101
,|4101,4102
BP|4103,4105
191|4106,4109
/|4109,4110
103|4110,4113
<EOL>|4114,4115
(|4115,4116
163|4116,4119
-|4119,4120
191|4120,4123
/|4123,4124
86|4124,4126
-|4126,4127
103|4127,4130
)|4130,4131
,|4131,4132
RR|4133,4135
18|4136,4138
(|4139,4140
24|4140,4142
on|4143,4145
my|4146,4148
check|4149,4154
)|4154,4155
,|4155,4156
O2|4157,4159
Sat|4160,4163
94|4164,4166
-|4166,4167
100|4167,4170
%|4170,4171
RA|4171,4173
<EOL>|4173,4174
FSBS|4174,4178
250s|4179,4183
<EOL>|4183,4184
General|4184,4191
:|4191,4192
Obese|4193,4198
woman|4199,4204
lying|4205,4210
in|4211,4213
bed|4214,4217
in|4218,4220
NAD|4221,4224
,|4224,4225
audible|4226,4233
wheezing|4234,4242
with|4243,4247
<EOL>|4248,4249
some|4249,4253
tachypnea|4254,4263
.|4263,4264
Speaking|4265,4273
in|4274,4276
_|4277,4278
_|4278,4279
_|4279,4280
word|4281,4285
sentences|4286,4295
with|4296,4300
slow|4301,4305
speech|4306,4312
.|4312,4313
<EOL>|4313,4314
HEENT|4314,4319
:|4319,4320
PERRL|4321,4326
,|4326,4327
EOMI|4328,4332
with|4333,4337
_|4338,4339
_|4339,4340
_|4340,4341
beats|4342,4347
of|4348,4350
nystagmus|4351,4360
on|4361,4363
rightward|4364,4373
gaze|4374,4378
<EOL>|4379,4380
in|4380,4382
both|4383,4387
eyes|4388,4392
,|4392,4393
no|4394,4396
other|4397,4402
nystagmus|4403,4412
,|4412,4413
sclera|4414,4420
anicteris|4421,4430
,|4430,4431
some|4432,4436
<EOL>|4437,4438
conjunctibal|4438,4450
pallor|4451,4457
,|4457,4458
MMM|4459,4462
,|4462,4463
clear|4464,4469
posterior|4470,4479
OP|4480,4482
,|4482,4483
no|4484,4486
lesions|4487,4494
,|4494,4495
<EOL>|4496,4497
symmetric|4497,4506
palate|4507,4513
elevation|4514,4523
,|4523,4524
tongue|4525,4531
midline|4532,4539
.|4539,4540
<EOL>|4540,4541
Neck|4541,4545
:|4545,4546
No|4547,4549
cervical|4550,4558
/|4558,4559
supraclavicular|4559,4574
LAD|4575,4578
,|4578,4579
no|4580,4582
notable|4583,4590
JVD|4591,4594
(|4595,4596
difficult|4596,4605
<EOL>|4606,4607
to|4607,4609
assess|4610,4616
_|4617,4618
_|4618,4619
_|4619,4620
body|4621,4625
habitus|4626,4633
)|4633,4634
<EOL>|4634,4635
CV|4635,4637
:|4637,4638
RRR|4639,4642
,|4642,4643
soft|4644,4648
S1|4649,4651
,|4651,4652
normal|4653,4659
S2|4660,4662
,|4662,4663
no|4664,4666
murmurs|4667,4674
noted|4675,4680
.|4680,4681
<EOL>|4681,4682
Lungs|4682,4687
:|4687,4688
Diffuse|4689,4696
expiratory|4697,4707
rhonchi|4708,4715
this|4716,4720
morning|4721,4728
,|4728,4729
no|4730,4732
wheezing|4733,4741
on|4742,4744
<EOL>|4745,4746
lung|4746,4750
exam|4751,4755
,|4755,4756
with|4757,4761
crackles|4762,4770
in|4771,4773
bilateral|4774,4783
bases|4784,4789
up|4790,4792
_|4793,4794
_|4794,4795
_|4795,4796
of|4797,4799
back|4800,4804
.|4804,4805
Poor|4806,4810
<EOL>|4811,4812
air|4812,4815
movement|4816,4824
overall|4825,4832
.|4832,4833
<EOL>|4833,4834
Abdomen|4834,4841
:|4841,4842
soft|4843,4847
,|4847,4848
obese|4849,4854
,|4854,4855
nontender|4856,4865
,|4865,4866
nondistended|4867,4879
,|4879,4880
+|4881,4882
BS|4882,4884
.|4884,4885
Unable|4886,4892
to|4893,4895
<EOL>|4896,4897
adequately|4897,4907
assess|4908,4914
organomegaly|4915,4927
.|4927,4928
<EOL>|4928,4929
GU|4929,4931
:|4931,4932
No|4933,4935
foley|4936,4941
<EOL>|4941,4942
Ext|4942,4945
:|4945,4946
wwp|4947,4950
,|4950,4951
2|4952,4953
+|4953,4954
peripheral|4955,4965
pulses|4966,4972
,|4972,4973
3|4974,4975
+|4975,4976
pitting|4977,4984
edema|4985,4990
to|4991,4993
knee|4994,4998
on|4999,5001
L|5002,5003
,|5003,5004
<EOL>|5005,5006
2|5006,5007
+|5007,5008
pitting|5009,5016
edema|5017,5022
in|5023,5025
R|5026,5027
leg|5028,5031
.|5031,5032
<EOL>|5032,5033
Neuro|5033,5038
:|5038,5039
CN2|5040,5043
-|5043,5044
12|5044,5046
notable|5047,5054
for|5055,5058
rightward|5059,5068
gaze|5069,5073
nystagmus|5074,5083
_|5084,5085
_|5085,5086
_|5086,5087
beats|5088,5093
)|5093,5094
,|5094,5095
<EOL>|5096,5097
otheriwse|5097,5106
intact|5107,5113
.|5113,5114
A|5115,5116
+|5116,5117
O|5117,5118
to|5119,5121
person|5122,5128
,|5128,5129
hospital|5130,5138
,|5138,5139
month|5140,5145
,|5145,5146
year|5147,5151
(|5152,5153
date|5153,5157
was|5158,5161
<EOL>|5162,5163
wrong|5163,5168
on|5169,5171
calendar|5172,5180
so|5181,5183
did|5184,5187
not|5188,5191
know|5192,5196
date|5197,5201
)|5201,5202
.|5202,5203
No|5204,5206
pronator|5207,5215
drift|5216,5221
,|5221,5222
some|5223,5227
<EOL>|5228,5229
positional|5229,5239
tremor|5240,5246
in|5247,5249
bilateral|5250,5259
hands|5260,5265
.|5265,5266
FNF|5267,5270
with|5271,5275
hesitancy|5276,5285
at|5286,5288
<EOL>|5289,5290
end|5290,5293
-|5293,5294
action|5294,5300
.|5300,5301
No|5302,5304
asterixis|5305,5314
.|5314,5315
Sensation|5316,5325
to|5326,5328
light|5329,5334
touch|5335,5340
grossly|5341,5348
<EOL>|5349,5350
intact|5350,5356
in|5357,5359
all|5360,5363
extremities|5364,5375
.|5375,5376
No|5377,5379
truncal|5380,5387
ataxia|5388,5394
sitting|5395,5402
upright|5403,5410
in|5411,5413
<EOL>|5414,5415
bed|5415,5418
during|5419,5425
exam|5426,5430
.|5430,5431
Gait|5432,5436
testing|5437,5444
deferred|5445,5453
.|5453,5454
Noted|5455,5460
to|5461,5463
have|5464,5468
repetitive|5469,5479
<EOL>|5480,5481
movements|5481,5490
at|5491,5493
rest|5494,5498
with|5499,5503
L|5504,5505
hand|5506,5510
(|5511,5512
wringing|5512,5520
sheets|5521,5527
,|5527,5528
tapping|5529,5536
,|5536,5537
etc|5538,5541
.|5541,5542
<EOL>|5543,5544
seemingly|5544,5553
patient|5554,5561
unaware|5562,5569
)|5569,5570
.|5570,5571
<EOL>|5571,5572
Skin|5572,5576
:|5576,5577
No|5578,5580
obvious|5581,5588
rashes|5589,5595
/|5595,5596
excoriations|5596,5608
on|5609,5611
extremities|5612,5623
and|5624,5627
<EOL>|5628,5629
abdomen|5629,5636
/|5636,5637
back|5637,5641
.|5641,5642
<EOL>|5642,5643
<EOL>|5643,5644
DISCHARGE|5644,5653
PHYSICAL|5654,5662
EXAM|5663,5667
:|5667,5668
<EOL>|5668,5669
=|5669,5670
=|5670,5671
=|5671,5672
=|5672,5673
=|5673,5674
=|5674,5675
=|5675,5676
=|5676,5677
=|5677,5678
=|5678,5679
=|5679,5680
=|5680,5681
=|5681,5682
=|5682,5683
=|5683,5684
=|5684,5685
=|5685,5686
=|5686,5687
=|5687,5688
=|5688,5689
=|5689,5690
=|5690,5691
=|5691,5692
=|5692,5693
=|5693,5694
=|5694,5695
=|5695,5696
<EOL>|5696,5697
Vitals|5697,5703
:|5703,5704
Tm|5705,5707
98.1|5708,5712
,|5712,5713
146|5714,5717
/|5717,5718
64|5718,5720
(|5721,5722
SBP|5722,5725
110|5726,5729
-|5729,5730
146|5730,5733
)|5733,5734
,|5734,5735
70|5736,5738
-|5738,5739
76|5739,5741
,|5741,5742
18|5743,5745
,|5745,5746
98|5747,5749
%|5749,5750
RA|5750,5752
<EOL>|5752,5753
Weight|5753,5759
:|5759,5760
75.9|5761,5765
kg|5766,5768
<EOL>|5768,5769
General|5769,5776
:|5776,5777
Obese|5778,5783
woman|5784,5789
in|5790,5792
NAD|5793,5796
.|5796,5797
<EOL>|5798,5799
HEENT|5799,5804
:|5804,5805
PERRL|5806,5811
,|5811,5812
EOMI|5813,5817
with|5818,5822
_|5823,5824
_|5824,5825
_|5825,5826
beats|5827,5832
of|5833,5835
nystagmus|5836,5845
on|5846,5848
rightward|5849,5858
gaze|5859,5863
<EOL>|5864,5865
in|5865,5867
both|5868,5872
eyes|5873,5877
,|5877,5878
no|5879,5881
other|5882,5887
nystagmus|5888,5897
,|5897,5898
sclera|5899,5905
anicteris|5906,5915
,|5915,5916
some|5917,5921
<EOL>|5922,5923
conjunctibal|5923,5935
pallor|5936,5942
,|5942,5943
MMM|5944,5947
,|5947,5948
clear|5949,5954
posterior|5955,5964
OP|5965,5967
,|5967,5968
no|5969,5971
lesions|5972,5979
,|5979,5980
<EOL>|5981,5982
symmetric|5982,5991
palate|5992,5998
elevation|5999,6008
,|6008,6009
tongue|6010,6016
midline|6017,6024
.|6024,6025
<EOL>|6027,6028
Neck|6028,6032
:|6032,6033
No|6034,6036
notable|6037,6044
JVD|6045,6048
(|6049,6050
difficult|6050,6059
to|6060,6062
assess|6063,6069
_|6070,6071
_|6071,6072
_|6072,6073
body|6074,6078
habitus|6079,6086
)|6086,6087
<EOL>|6087,6088
CV|6088,6090
:|6090,6091
RRR|6092,6095
,|6095,6096
soft|6097,6101
S1|6102,6104
,|6104,6105
normal|6106,6112
S2|6113,6115
,|6115,6116
no|6117,6119
murmurs|6120,6127
noted|6128,6133
.|6133,6134
<EOL>|6134,6135
Lungs|6135,6140
:|6140,6141
CTAB|6142,6146
<EOL>|6147,6148
Abdomen|6148,6155
:|6155,6156
soft|6157,6161
,|6161,6162
obese|6163,6168
,|6168,6169
nontender|6170,6179
,|6179,6180
nondistended|6181,6193
,|6193,6194
+|6195,6196
BS|6196,6198
.|6198,6199
Unable|6200,6206
to|6207,6209
<EOL>|6210,6211
adequately|6211,6221
assess|6222,6228
organomegaly|6229,6241
.|6241,6242
<EOL>|6242,6243
Ext|6243,6246
:|6246,6247
wwp|6248,6251
,|6251,6252
2|6253,6254
+|6254,6255
peripheral|6256,6266
pulses|6267,6273
,|6273,6274
no|6275,6277
pitting|6278,6285
edema|6286,6291
<EOL>|6291,6292
<EOL>|6293,6294
Pertinent|6294,6303
Results|6304,6311
:|6311,6312
<EOL>|6312,6313
=|6313,6314
=|6314,6315
=|6315,6316
=|6316,6317
ADMISSION|6318,6327
LABS|6328,6332
=|6333,6334
=|6334,6335
=|6335,6336
=|6336,6337
<EOL>|6337,6338
_|6338,6339
_|6339,6340
_|6340,6341
04|6342,6344
:|6344,6345
00PM|6345,6349
BLOOD|6350,6355
WBC|6356,6359
-|6359,6360
4.3|6360,6363
RBC|6364,6367
-|6367,6368
2|6368,6369
.|6369,6370
84|6370,6372
*|6372,6373
Hgb|6374,6377
-|6377,6378
8|6378,6379
.|6379,6380
6|6380,6381
*|6381,6382
Hct|6383,6386
-|6386,6387
26|6387,6389
.|6389,6390
0|6390,6391
*|6391,6392
<EOL>|6393,6394
MCV|6394,6397
-|6397,6398
92|6398,6400
MCH|6401,6404
-|6404,6405
30.4|6405,6409
MCHC|6410,6414
-|6414,6415
33.2|6415,6419
RDW|6420,6423
-|6423,6424
14.2|6424,6428
Plt|6429,6432
_|6433,6434
_|6434,6435
_|6435,6436
<EOL>|6436,6437
_|6437,6438
_|6438,6439
_|6439,6440
04|6441,6443
:|6443,6444
00PM|6444,6448
BLOOD|6449,6454
Neuts|6455,6460
-|6460,6461
71|6461,6463
.|6463,6464
5|6464,6465
*|6465,6466
_|6467,6468
_|6468,6469
_|6469,6470
Monos|6471,6476
-|6476,6477
4.5|6477,6480
Eos|6481,6484
-|6484,6485
2.6|6485,6488
<EOL>|6489,6490
Baso|6490,6494
-|6494,6495
0.1|6495,6498
<EOL>|6498,6499
_|6499,6500
_|6500,6501
_|6501,6502
04|6503,6505
:|6505,6506
00PM|6506,6510
BLOOD|6511,6516
_|6517,6518
_|6518,6519
_|6519,6520
PTT|6521,6524
-|6524,6525
24|6525,6527
.|6527,6528
5|6528,6529
*|6529,6530
_|6531,6532
_|6532,6533
_|6533,6534
<EOL>|6534,6535
_|6535,6536
_|6536,6537
_|6537,6538
04|6539,6541
:|6541,6542
00PM|6542,6546
BLOOD|6547,6552
Glucose|6553,6560
-|6560,6561
325|6561,6564
*|6564,6565
UreaN|6566,6571
-|6571,6572
29|6572,6574
*|6574,6575
Creat|6576,6581
-|6581,6582
2|6582,6583
.|6583,6584
1|6584,6585
*|6585,6586
Na|6587,6589
-|6589,6590
141|6590,6593
<EOL>|6594,6595
K|6595,6596
-|6596,6597
4.0|6597,6600
Cl|6601,6603
-|6603,6604
106|6604,6607
HCO3|6608,6612
-|6612,6613
24|6613,6615
AnGap|6616,6621
-|6621,6622
15|6622,6624
<EOL>|6624,6625
_|6625,6626
_|6626,6627
_|6627,6628
07|6629,6631
:|6631,6632
55AM|6632,6636
BLOOD|6637,6642
Calcium|6643,6650
-|6650,6651
9.5|6651,6654
Phos|6655,6659
-|6659,6660
3|6660,6661
.|6661,6662
5|6662,6663
#|6663,6664
Mg|6665,6667
-|6667,6668
1.5|6668,6671
*|6671,6672
<EOL>|6672,6673
<EOL>|6673,6674
_|6674,6675
_|6675,6676
_|6676,6677
07|6678,6680
:|6680,6681
00PM|6681,6685
URINE|6686,6691
Color|6692,6697
-|6697,6698
Yellow|6698,6704
Appear|6705,6711
-|6711,6712
Clear|6712,6717
Sp|6718,6720
_|6721,6722
_|6722,6723
_|6723,6724
<EOL>|6724,6725
_|6725,6726
_|6726,6727
_|6727,6728
07|6729,6731
:|6731,6732
00PM|6732,6736
URINE|6737,6742
Blood|6743,6748
-|6748,6749
NEG|6749,6752
Nitrite|6753,6760
-|6760,6761
NEG|6761,6764
Protein|6765,6772
-|6772,6773
100|6773,6776
<EOL>|6777,6778
Glucose|6778,6785
-|6785,6786
300|6786,6789
Ketone|6790,6796
-|6796,6797
NEG|6797,6800
Bilirub|6801,6808
-|6808,6809
NEG|6809,6812
Urobiln|6813,6820
-|6820,6821
NEG|6821,6824
pH|6825,6827
-|6827,6828
6.0|6828,6831
Leuks|6832,6837
-|6837,6838
SM|6838,6840
<EOL>|6841,6842
_|6842,6843
_|6843,6844
_|6844,6845
07|6846,6848
:|6848,6849
00PM|6849,6853
URINE|6854,6859
RBC|6860,6863
-|6863,6864
2|6864,6865
WBC|6866,6869
-|6869,6870
4|6870,6871
Bacteri|6872,6879
-|6879,6880
FEW|6880,6883
Yeast|6884,6889
-|6889,6890
NONE|6890,6894
Epi|6895,6898
-|6898,6899
1|6899,6900
<EOL>|6900,6901
_|6901,6902
_|6902,6903
_|6903,6904
07|6905,6907
:|6907,6908
00PM|6908,6912
URINE|6913,6918
CastHy|6919,6925
-|6925,6926
6|6926,6927
*|6927,6928
<EOL>|6928,6929
<EOL>|6929,6930
_|6930,6931
_|6931,6932
_|6932,6933
04|6934,6936
:|6936,6937
00PM|6937,6941
BLOOD|6942,6947
cTropnT|6948,6955
-|6955,6956
<|6956,6957
0|6957,6958
.|6958,6959
01|6959,6961
proBNP|6962,6968
-|6968,6969
4279|6969,6973
*|6973,6974
<EOL>|6974,6975
_|6975,6976
_|6976,6977
_|6977,6978
09|6979,6981
:|6981,6982
30PM|6982,6986
BLOOD|6987,6992
cTropnT|6993,7000
-|7000,7001
<|7001,7002
0|7002,7003
.|7003,7004
01|7004,7006
<EOL>|7006,7007
<EOL>|7007,7008
=|7008,7009
=|7009,7010
=|7010,7011
=|7011,7012
IMAGING|7013,7020
=|7021,7022
=|7022,7023
=|7023,7024
=|7024,7025
<EOL>|7025,7026
<EOL>|7026,7027
_|7027,7028
_|7028,7029
_|7029,7030
CHEST|7031,7036
(|7037,7038
PA|7038,7040
AND|7041,7044
LAT|7045,7048
)|7048,7049
:|7049,7050
<EOL>|7050,7051
The|7051,7054
lungs|7055,7060
are|7061,7064
clear|7065,7070
of|7071,7073
consolidation|7074,7087
,|7087,7088
effusion|7089,7097
,|7097,7098
or|7099,7101
edema|7102,7107
.|7107,7108
<EOL>|7109,7110
Cardiac|7110,7117
silhouette|7118,7128
is|7129,7131
top|7132,7135
normal|7136,7142
.|7142,7143
Descending|7144,7154
thoracic|7155,7163
aorta|7164,7169
is|7170,7172
<EOL>|7173,7174
tortuous|7174,7182
with|7183,7187
atherosclerotic|7188,7203
calcification|7204,7217
seen|7218,7222
at|7223,7225
the|7226,7229
arch|7230,7234
.|7234,7235
No|7236,7238
<EOL>|7239,7240
acute|7240,7245
osseous|7246,7253
abnormalities|7254,7267
identified|7268,7278
.|7278,7279
<EOL>|7280,7281
No|7295,7297
acute|7298,7303
cardiopulmonary|7304,7319
process|7320,7327
.|7327,7328
<EOL>|7328,7329
<EOL>|7329,7330
_|7330,7331
_|7331,7332
_|7332,7333
P|7334,7335
-|7335,7336
MIBI|7336,7340
:|7340,7341
<EOL>|7341,7342
Clinical|7342,7350
Indication|7351,7361
:|7361,7362
SS|7363,7365
CHEST|7366,7371
TIGHTNESS|7372,7381
ASSESS|7382,7388
FOR|7389,7392
EVIDENCE|7393,7401
OF|7402,7404
<EOL>|7405,7406
ISCHEMIA|7406,7414
<EOL>|7416,7417
HISTORY|7417,7424
:|7424,7425
_|7426,7427
_|7427,7428
_|7428,7429
yo|7430,7432
woman|7433,7438
with|7439,7443
a|7444,7445
history|7446,7453
of|7454,7456
CAD|7457,7460
and|7461,7464
CHF|7465,7468
referred|7469,7477
for|7478,7481
<EOL>|7482,7483
evaluation|7483,7493
of|7494,7496
chest|7497,7502
pain|7503,7507
and|7508,7511
dyspnea|7512,7519
.|7519,7520
<EOL>|7520,7521
<EOL>|7521,7522
SUMMARY|7522,7529
FROM|7530,7534
THE|7535,7538
EXERCISE|7539,7547
LAB|7548,7551
:|7551,7552
<EOL>|7553,7554
For|7554,7557
pharmacologic|7558,7571
coronary|7572,7580
vasodilatation|7581,7595
dipyridamole|7596,7608
was|7609,7612
<EOL>|7613,7614
infused|7614,7621
intravenously|7622,7635
for|7636,7639
4|7640,7641
minutes|7642,7649
at|7650,7652
a|7653,7654
dose|7655,7659
of|7660,7662
0.142|7663,7668
<EOL>|7669,7670
milligram|7670,7679
/|7679,7680
kilogram|7680,7688
/|7688,7689
min|7689,7692
.|7692,7693
She|7694,7697
had|7698,7701
no|7702,7704
anginal|7705,7712
symptoms|7713,7721
or|7722,7724
ischemic|7725,7733
<EOL>|7734,7735
ECG|7735,7738
changes|7739,7746
.|7746,7747
<EOL>|7747,7748
<EOL>|7748,7749
ISOTOPE|7761,7768
DATA|7769,7773
:|7773,7774
(|7775,7776
_|7776,7777
_|7777,7778
_|7778,7779
)|7779,7780
11.0|7781,7785
mCi|7786,7789
Tc|7790,7792
-|7792,7793
99m|7793,7796
Sestamibi|7797,7806
Rest|7807,7811
;|7811,7812
<EOL>|7813,7814
(|7814,7815
_|7815,7816
_|7816,7817
_|7817,7818
)|7818,7819
29.6|7820,7824
mCi|7825,7828
Tc|7829,7831
-|7831,7832
99m|7832,7835
Sestamibi|7836,7845
Stress|7846,7852
;|7852,7853
DRUG|7854,7858
DATA|7859,7863
:|7863,7864
(|7865,7866
Non-NM|7866,7872
<EOL>|7873,7874
admin|7874,7879
)|7879,7880
Dipyridamole|7881,7893
;|7893,7894
<EOL>|7894,7895
<EOL>|7895,7896
IMAGING|7896,7903
METHOD|7904,7910
:|7910,7911
<EOL>|7911,7912
Resting|7912,7919
perfusion|7920,7929
images|7930,7936
were|7937,7941
obtained|7942,7950
with|7951,7955
Tc|7956,7958
-|7958,7959
99m|7959,7962
sestamibi|7963,7972
.|7972,7973
<EOL>|7974,7975
Tracer|7975,7981
was|7982,7985
injected|7986,7994
approximately|7995,8008
45|8009,8011
minutes|8012,8019
prior|8020,8025
to|8026,8028
obtaining|8029,8038
<EOL>|8039,8040
the|8040,8043
resting|8044,8051
images|8052,8058
.|8058,8059
<EOL>|8060,8061
Following|8061,8070
resting|8071,8078
images|8079,8085
and|8086,8089
following|8090,8099
intravenous|8100,8111
infusion|8112,8120
,|8120,8121
<EOL>|8122,8123
approximately|8123,8136
three|8137,8142
times|8143,8148
the|8149,8152
resting|8153,8160
dose|8161,8165
of|8166,8168
Tc|8169,8171
-|8171,8172
99m|8172,8175
sestamibi|8176,8185
<EOL>|8186,8187
was|8187,8190
administered|8191,8203
intravenously|8204,8217
.|8217,8218
Stress|8219,8225
images|8226,8232
were|8233,8237
obtained|8238,8246
<EOL>|8247,8248
approximately|8248,8261
30|8262,8264
minutes|8265,8272
following|8273,8282
tracer|8283,8289
injection|8290,8299
.|8299,8300
<EOL>|8301,8302
Imaging|8302,8309
protocol|8310,8318
:|8318,8319
Gated|8320,8325
SPECT|8326,8331
.|8331,8332
<EOL>|8333,8334
This|8334,8338
study|8339,8344
was|8345,8348
interpreted|8349,8360
using|8361,8366
the|8367,8370
17|8371,8373
-|8373,8374
segment|8374,8381
myocardial|8382,8392
<EOL>|8393,8394
perfusion|8394,8403
model|8404,8409
.|8409,8410
<EOL>|8411,8412
<EOL>|8412,8413
:|8421,8422
<EOL>|8423,8424
The|8424,8427
image|8428,8433
quality|8434,8441
is|8442,8444
adequate|8445,8453
but|8454,8457
limited|8458,8465
due|8466,8469
to|8470,8472
soft|8473,8477
tissue|8478,8484
and|8485,8488
<EOL>|8489,8490
breast|8490,8496
attenuation|8497,8508
.|8508,8509
<EOL>|8509,8510
Left|8510,8514
ventricular|8515,8526
cavity|8527,8533
size|8534,8538
is|8539,8541
increased|8542,8551
.|8551,8552
<EOL>|8552,8553
Rest|8553,8557
and|8558,8561
stress|8562,8568
perfusion|8569,8578
images|8579,8585
reveal|8586,8592
uniform|8593,8600
tracer|8601,8607
uptake|8608,8614
<EOL>|8615,8616
throughout|8616,8626
the|8627,8630
left|8631,8635
ventricular|8636,8647
myocardium|8648,8658
.|8658,8659
<EOL>|8660,8661
Gated|8661,8666
images|8667,8673
reveal|8674,8680
normal|8681,8687
wall|8688,8692
motion|8693,8699
.|8699,8700
<EOL>|8701,8702
The|8702,8705
calculated|8706,8716
left|8717,8721
ventricular|8722,8733
ejection|8734,8742
fraction|8743,8751
is|8752,8754
59|8755,8757
%|8757,8758
with|8759,8763
an|8764,8766
<EOL>|8767,8768
EDV|8768,8771
of|8772,8774
117|8775,8778
ml|8779,8781
.|8781,8782
<EOL>|8782,8783
<EOL>|8783,8784
1.|8796,8798
Normal|8799,8805
myocardial|8806,8816
perfusion|8817,8826
.|8826,8827
<EOL>|8828,8829
2.|8829,8831
Increased|8832,8841
left|8842,8846
ventricular|8847,8858
cavity|8859,8865
size|8866,8870
with|8871,8875
normal|8876,8882
systolic|8883,8891
<EOL>|8892,8893
function|8893,8901
.|8901,8902
<EOL>|8902,8903
Compared|8903,8911
with|8912,8916
prior|8917,8922
study|8923,8928
of|8929,8931
_|8932,8933
_|8933,8934
_|8934,8935
,|8935,8936
the|8937,8940
cavity|8941,8947
size|8948,8952
is|8953,8955
<EOL>|8956,8957
larger|8957,8963
.|8963,8964
<EOL>|8964,8965
<EOL>|8966,8967
<EOL>|8968,8969
_|8992,8993
_|8993,8994
_|8994,8995
year|8996,9000
old|9001,9004
female|9005,9011
with|9012,9016
history|9017,9024
of|9025,9027
HTN|9028,9031
,|9031,9032
CVA|9033,9036
,|9036,9037
CAD|9038,9041
(|9042,9043
s|9043,9044
/|9044,9045
p|9045,9046
BMS|9047,9050
to|9051,9053
<EOL>|9054,9055
circumflex|9055,9065
in|9066,9068
_|9069,9070
_|9070,9071
_|9071,9072
,|9072,9073
CHF|9074,9077
(|9078,9079
EF|9079,9081
45|9082,9084
%|9084,9085
in|9086,9088
_|9089,9090
_|9090,9091
_|9091,9092
who|9093,9096
presented|9097,9106
<EOL>|9107,9108
with|9108,9112
acute|9113,9118
onset|9119,9124
shortness|9125,9134
of|9135,9137
breath|9138,9144
and|9145,9148
substernal|9149,9159
chest|9160,9165
<EOL>|9166,9167
tightness|9167,9176
.|9176,9177
<EOL>|9177,9178
<EOL>|9178,9179
#|9179,9180
Shortness|9181,9190
of|9191,9193
breath|9194,9200
:|9200,9201
<EOL>|9201,9202
Patient|9202,9209
with|9210,9214
acute|9215,9220
onset|9221,9226
SOB|9227,9230
following|9231,9240
seafood|9241,9248
meal|9249,9253
with|9254,9258
<EOL>|9259,9260
associated|9260,9270
chest|9271,9276
tightness|9277,9286
(|9287,9288
see|9288,9291
below|9292,9297
)|9297,9298
.|9298,9299
Patient|9300,9307
with|9308,9312
crackles|9313,9321
<EOL>|9322,9323
and|9323,9326
expiratory|9327,9337
rhonchi|9338,9345
on|9346,9348
lung|9349,9353
exam|9354,9358
.|9358,9359
CXR|9360,9363
did|9364,9367
not|9368,9371
show|9372,9376
<EOL>|9377,9378
significant|9378,9389
pulmonary|9390,9399
edema|9400,9405
,|9405,9406
pleural|9407,9414
effusions|9415,9424
,|9424,9425
or|9426,9428
consolidation|9429,9442
<EOL>|9443,9444
although|9444,9452
her|9453,9456
BNP|9457,9460
was|9461,9464
elevated|9465,9473
.|9473,9474
Per|9475,9478
pharmacy|9479,9487
records|9488,9495
,|9495,9496
patient|9497,9504
had|9505,9508
<EOL>|9509,9510
not|9510,9513
refilled|9514,9522
lasix|9523,9528
prescription|9529,9541
since|9542,9547
_|9548,9549
_|9549,9550
_|9550,9551
.|9551,9552
Overall|9553,9560
,|9560,9561
<EOL>|9562,9563
presentation|9563,9575
was|9576,9579
most|9580,9584
consistent|9585,9595
with|9596,9600
a|9601,9602
mild|9603,9607
CHF|9608,9611
exacerbation|9612,9624
.|9624,9625
<EOL>|9626,9627
She|9627,9630
received|9631,9639
treatment|9640,9649
with|9650,9654
IV|9655,9657
lasix|9658,9663
and|9664,9667
her|9668,9671
shortness|9672,9681
of|9682,9684
breath|9685,9691
<EOL>|9692,9693
subsequently|9693,9705
improved|9706,9714
quickly|9715,9722
.|9722,9723
She|9724,9727
was|9728,9731
able|9732,9736
to|9737,9739
be|9740,9742
transitioned|9743,9755
<EOL>|9756,9757
to|9757,9759
a|9760,9761
PO|9762,9764
regimen|9765,9772
of|9773,9775
lasix|9776,9781
40mg|9782,9786
qday|9787,9791
on|9792,9794
_|9795,9796
_|9796,9797
_|9797,9798
(|9799,9800
day|9800,9803
of|9804,9806
discharge|9807,9816
)|9816,9817
.|9817,9818
<EOL>|9819,9820
Dry|9820,9823
weight|9824,9830
on|9831,9833
day|9834,9837
of|9838,9840
discharge|9841,9850
was|9851,9854
75.9|9855,9859
kg|9859,9861
.|9861,9862
<EOL>|9862,9863
<EOL>|9863,9864
#|9864,9865
Chest|9866,9871
Tightness|9872,9881
:|9881,9882
<EOL>|9882,9883
Patient|9883,9890
reported|9891,9899
chest|9900,9905
tightness|9906,9915
associated|9916,9926
with|9927,9931
her|9932,9935
shortness|9936,9945
<EOL>|9946,9947
of|9947,9949
breath|9950,9956
.|9956,9957
Was|9958,9961
given|9962,9967
aspirin|9968,9975
and|9976,9979
SL|9980,9982
nitroglycerin|9983,9996
in|9997,9999
her|10000,10003
PCP|10004,10007
's|10007,10009
<EOL>|10010,10011
office|10011,10017
prior|10018,10023
to|10024,10026
being|10027,10032
directed|10033,10041
to|10042,10044
the|10045,10048
ED|10049,10051
.|10051,10052
Troponin|10053,10061
was|10062,10065
negative|10066,10074
<EOL>|10075,10076
x2|10076,10078
.|10078,10079
EKG|10080,10083
without|10084,10091
evidence|10092,10100
of|10101,10103
acute|10104,10109
ischemia|10110,10118
.|10118,10119
Due|10120,10123
to|10124,10126
her|10127,10130
<EOL>|10131,10132
significant|10132,10143
CAD|10144,10147
history|10148,10155
,|10155,10156
she|10157,10160
underwent|10161,10170
a|10171,10172
P|10173,10174
-|10174,10175
MIBI|10175,10179
on|10180,10182
_|10183,10184
_|10184,10185
_|10185,10186
which|10187,10192
<EOL>|10193,10194
was|10194,10197
unremarkable|10198,10210
.|10210,10211
Her|10212,10215
chest|10216,10221
tightness|10222,10231
was|10232,10235
thought|10236,10243
to|10244,10246
be|10247,10249
of|10250,10252
<EOL>|10253,10254
non-cardiac|10254,10265
etiology|10266,10274
.|10274,10275
<EOL>|10275,10276
<EOL>|10276,10277
#|10277,10278
HTN|10279,10282
:|10282,10283
<EOL>|10283,10284
Patient|10284,10291
presented|10292,10301
with|10302,10306
SBP|10307,10310
of|10311,10313
190|10314,10317
-|10317,10318
200|10318,10321
.|10321,10322
Cardiology|10323,10333
was|10334,10337
consulted|10338,10347
<EOL>|10348,10349
and|10349,10352
recommended|10353,10364
increasing|10365,10375
her|10376,10379
carvedilol|10380,10390
from|10391,10395
6.25|10396,10400
mg|10400,10402
BID|10403,10406
to|10407,10409
<EOL>|10410,10411
12.5|10411,10415
mg|10415,10417
BID|10418,10421
.|10421,10422
With|10423,10427
this|10428,10432
change|10433,10439
,|10439,10440
and|10441,10444
continuation|10445,10457
of|10458,10460
her|10461,10464
other|10465,10470
home|10471,10475
<EOL>|10476,10477
medications|10477,10488
,|10488,10489
her|10490,10493
blood|10494,10499
pressure|10500,10508
decreased|10509,10518
to|10519,10521
systolics|10522,10531
in|10532,10534
range|10535,10540
<EOL>|10541,10542
of|10542,10544
110|10545,10548
-|10548,10549
146|10549,10552
on|10553,10555
day|10556,10559
of|10560,10562
discharge|10563,10572
.|10572,10573
It|10574,10576
is|10577,10579
unclear|10580,10587
whether|10588,10595
her|10596,10599
very|10600,10604
<EOL>|10605,10606
elevated|10606,10614
BP|10615,10617
on|10618,10620
admission|10621,10630
was|10631,10634
occurring|10635,10644
in|10645,10647
the|10648,10651
setting|10652,10659
of|10660,10662
<EOL>|10663,10664
medication|10664,10674
non-compliance|10675,10689
.|10689,10690
Nifedipine|10691,10701
was|10702,10705
decreased|10706,10715
from|10716,10720
BID|10721,10724
to|10725,10727
<EOL>|10728,10729
daily|10729,10734
given|10735,10740
increased|10741,10750
carvedilol|10751,10761
and|10762,10765
addition|10766,10774
of|10775,10777
Lasix|10778,10783
(|10784,10785
which|10785,10790
<EOL>|10791,10792
patient|10792,10799
was|10800,10803
believed|10804,10812
to|10813,10815
have|10816,10820
been|10821,10825
non-compliant|10826,10839
with|10840,10844
prior|10845,10850
to|10851,10853
<EOL>|10854,10855
this|10855,10859
admission|10860,10869
)|10869,10870
.|10870,10871
<EOL>|10871,10872
<EOL>|10872,10873
=|10873,10874
=|10874,10875
=|10875,10876
=|10876,10877
TRANSITIONAL|10878,10890
ISSUES|10891,10897
=|10898,10899
=|10899,10900
=|10900,10901
=|10901,10902
<EOL>|10902,10903
<EOL>|10903,10904
#|10904,10905
CHF|10906,10909
:|10909,10910
<EOL>|10910,10911
-|10911,10912
_|10913,10914
_|10914,10915
_|10915,10916
services|10917,10925
for|10926,10929
medication|10930,10940
teaching|10941,10949
and|10950,10953
pill|10954,10958
-|10958,10959
box|10959,10962
,|10962,10963
as|10964,10966
well|10967,10971
as|10972,10974
<EOL>|10975,10976
weights|10976,10983
<EOL>|10983,10984
-|10984,10985
Follow|10986,10992
up|10993,10995
with|10996,11000
her|11001,11004
cardiologist|11005,11017
Dr.|11018,11021
_|11022,11023
_|11023,11024
_|11024,11025
on|11026,11028
_|11029,11030
_|11030,11031
_|11031,11032
<EOL>|11032,11033
-|11033,11034
Please|11035,11041
check|11042,11047
repeat|11048,11054
Chem|11055,11059
-|11059,11060
10|11060,11062
and|11063,11066
CBC|11067,11070
on|11071,11073
_|11074,11075
_|11075,11076
_|11076,11077
<EOL>|11077,11078
-|11078,11079
Continue|11080,11088
furosemide|11089,11099
40mg|11100,11104
qday|11105,11109
<EOL>|11109,11110
<EOL>|11110,11111
#|11111,11112
Hct|11113,11116
Drop|11117,11121
:|11121,11122
Patient|11123,11130
with|11131,11135
chronic|11136,11143
anemia|11144,11150
and|11151,11154
Hgb|11155,11158
drop|11159,11163
on|11164,11166
day|11167,11170
of|11171,11173
<EOL>|11174,11175
discharge|11175,11184
from|11185,11189
9.3|11190,11193
to|11194,11196
8.5|11197,11200
.|11200,11201
<EOL>|11201,11202
-|11202,11203
Repeat|11204,11210
CBC|11211,11214
check|11215,11220
on|11221,11223
_|11224,11225
_|11225,11226
_|11226,11227
<EOL>|11227,11228
<EOL>|11228,11229
#|11229,11230
HTN|11231,11234
:|11234,11235
<EOL>|11235,11236
-|11236,11237
Increased|11238,11247
carvedilol|11248,11258
to|11259,11261
12.5|11262,11266
mg|11266,11268
BID|11269,11272
<EOL>|11272,11273
-|11273,11274
Nifedipine|11275,11285
was|11286,11289
decreased|11290,11299
from|11300,11304
BID|11305,11308
to|11309,11311
daily|11312,11317
given|11318,11323
increased|11324,11333
<EOL>|11334,11335
carvedilol|11335,11345
and|11346,11349
addition|11350,11358
of|11359,11361
lasix|11362,11367
(|11368,11369
with|11369,11373
which|11374,11379
patient|11380,11387
was|11388,11391
likely|11392,11398
<EOL>|11399,11400
non-compliant|11400,11413
prior|11414,11419
to|11420,11422
this|11423,11427
admission|11428,11437
)|11437,11438
.|11438,11439
<EOL>|11439,11440
<EOL>|11440,11441
#|11441,11442
Health|11443,11449
Screening|11450,11459
<EOL>|11459,11460
-|11460,11461
Patient|11462,11469
is|11470,11472
due|11473,11476
for|11477,11480
colonoscopy|11481,11492
this|11493,11497
year|11498,11502
.|11502,11503
<EOL>|11503,11504
-|11504,11505
PCP|11506,11509
follow|11510,11516
up|11517,11519
with|11520,11524
Dr.|11525,11528
_|11529,11530
_|11530,11531
_|11531,11532
on|11533,11535
_|11536,11537
_|11537,11538
_|11538,11539
<EOL>|11539,11540
<EOL>|11540,11541
#|11541,11542
Weight|11543,11549
at|11550,11552
discharge|11553,11562
:|11562,11563
75.9|11564,11568
kg|11569,11571
<EOL>|11571,11572
<EOL>|11572,11573
#|11573,11574
Code|11575,11579
:|11579,11580
Full|11581,11585
(|11586,11587
confirmed|11587,11596
with|11597,11601
patient|11602,11609
)|11609,11610
<EOL>|11610,11611
#|11611,11612
Emergency|11613,11622
Contacts|11623,11631
:|11631,11632
<EOL>|11632,11633
-|11633,11634
_|11635,11636
_|11636,11637
_|11637,11638
,|11638,11639
_|11640,11641
_|11641,11642
_|11642,11643
(|11644,11645
_|11645,11646
_|11646,11647
_|11647,11648
)|11648,11649
<EOL>|11649,11650
-|11650,11651
Alternate|11652,11661
HCP|11662,11665
_|11666,11667
_|11667,11668
_|11668,11669
_|11669,11670
_|11670,11671
_|11671,11672
)|11672,11673
<EOL>|11673,11674
<EOL>|11675,11676
Medications|11676,11687
on|11688,11690
Admission|11691,11700
:|11700,11701
<EOL>|11701,11702
The|11702,11705
Preadmission|11706,11718
Medication|11719,11729
list|11730,11734
is|11735,11737
accurate|11738,11746
and|11747,11750
complete|11751,11759
.|11759,11760
<EOL>|11760,11761
1.|11761,11763
Aspirin|11764,11771
81|11772,11774
mg|11775,11777
PO|11778,11780
DAILY|11781,11786
<EOL>|11787,11788
2.|11788,11790
Clopidogrel|11791,11802
75|11803,11805
mg|11806,11808
PO|11809,11811
DAILY|11812,11817
<EOL>|11818,11819
3.|11819,11821
Furosemide|11822,11832
40|11833,11835
mg|11836,11838
PO|11839,11841
DAILY|11842,11847
<EOL>|11848,11849
4.|11849,11851
Multivitamins|11852,11865
1|11866,11867
TAB|11868,11871
PO|11872,11874
DAILY|11875,11880
<EOL>|11881,11882
5.|11882,11884
Ranitidine|11885,11895
300|11896,11899
mg|11900,11902
PO|11903,11905
DAILY|11906,11911
<EOL>|11912,11913
6.|11913,11915
Atorvastatin|11916,11928
80|11929,11931
mg|11932,11934
PO|11935,11937
DAILY|11938,11943
<EOL>|11944,11945
7.|11945,11947
HumuLIN|11948,11955
70|11956,11958
/|11958,11959
30|11959,11961
(|11962,11963
insulin|11963,11970
NPH|11971,11974
and|11975,11978
regular|11979,11986
human|11987,11992
)|11992,11993
30|11994,11996
units|11997,12002
<EOL>|12003,12004
subcutaneous|12004,12016
daily|12017,12022
<EOL>|12023,12024
8.|12024,12026
Nitroglycerin|12027,12040
SL|12041,12043
0.3|12044,12047
mg|12048,12050
SL|12051,12053
PRN|12054,12057
chest|12058,12063
pain|12064,12068
<EOL>|12069,12070
9.|12070,12072
Vitamin|12073,12080
D|12081,12082
_|12083,12084
_|12084,12085
_|12085,12086
UNIT|12087,12091
PO|12092,12094
DAILY|12095,12100
<EOL>|12101,12102
10.|12102,12105
NIFEdipine|12106,12116
CR|12117,12119
60|12120,12122
mg|12123,12125
PO|12126,12128
BID|12129,12132
<EOL>|12133,12134
11.|12134,12137
Lisinopril|12138,12148
40|12149,12151
mg|12152,12154
PO|12155,12157
DAILY|12158,12163
<EOL>|12164,12165
12.|12165,12168
Allopurinol|12169,12180
_|12181,12182
_|12182,12183
_|12183,12184
mg|12185,12187
PO|12188,12190
DAILY|12191,12196
<EOL>|12197,12198
13.|12198,12201
Ferrous|12202,12209
Sulfate|12210,12217
325|12218,12221
mg|12222,12224
PO|12225,12227
DAILY|12228,12233
<EOL>|12234,12235
14.|12235,12238
Carvedilol|12239,12249
6.25|12250,12254
mg|12255,12257
PO|12258,12260
BID|12261,12264
<EOL>|12265,12266
<EOL>|12266,12267
<EOL>|12268,12269
Discharge|12269,12278
Medications|12279,12290
:|12290,12291
<EOL>|12291,12292
1.|12292,12294
Outpatient|12295,12305
Lab|12306,12309
Work|12310,12314
<EOL>|12314,12315
Please|12315,12321
draw|12322,12326
Chem|12327,12331
-|12331,12332
10|12332,12334
and|12335,12338
CBC|12339,12342
on|12343,12345
_|12346,12347
_|12347,12348
_|12348,12349
.|12349,12350
<EOL>|12350,12351
Indication|12351,12361
:|12361,12362
428.0|12363,12368
(|12369,12370
CHF|12370,12373
)|12373,12374
and|12375,12378
anemia|12379,12385
(|12386,12387
280.1|12387,12392
)|12392,12393
<EOL>|12393,12394
Send|12394,12398
results|12399,12406
to|12407,12409
Dr.|12410,12413
_|12414,12415
_|12415,12416
_|12416,12417
(|12418,12419
fax|12419,12422
:|12422,12423
_|12424,12425
_|12425,12426
_|12426,12427
<EOL>|12427,12428
2.|12428,12430
Nitroglycerin|12431,12444
SL|12445,12447
0.3|12448,12451
mg|12452,12454
SL|12455,12457
PRN|12458,12461
chest|12462,12467
pain|12468,12472
<EOL>|12473,12474
3.|12474,12476
Vitamin|12477,12484
D|12485,12486
_|12487,12488
_|12488,12489
_|12489,12490
UNIT|12491,12495
PO|12496,12498
DAILY|12499,12504
<EOL>|12505,12506
4.|12506,12508
Ranitidine|12509,12519
300|12520,12523
mg|12524,12526
PO|12527,12529
DAILY|12530,12535
<EOL>|12536,12537
5.|12537,12539
NIFEdipine|12540,12550
CR|12551,12553
60|12554,12556
mg|12557,12559
PO|12560,12562
DAILY|12563,12568
<EOL>|12569,12570
6.|12570,12572
Multivitamins|12573,12586
1|12587,12588
TAB|12589,12592
PO|12593,12595
DAILY|12596,12601
<EOL>|12602,12603
7.|12603,12605
Allopurinol|12606,12617
_|12618,12619
_|12619,12620
_|12620,12621
mg|12622,12624
PO|12625,12627
DAILY|12628,12633
<EOL>|12634,12635
8.|12635,12637
Aspirin|12638,12645
81|12646,12648
mg|12649,12651
PO|12652,12654
DAILY|12655,12660
<EOL>|12661,12662
9.|12662,12664
Atorvastatin|12665,12677
80|12678,12680
mg|12681,12683
PO|12684,12686
DAILY|12687,12692
<EOL>|12693,12694
10.|12694,12697
Clopidogrel|12698,12709
75|12710,12712
mg|12713,12715
PO|12716,12718
DAILY|12719,12724
<EOL>|12725,12726
11.|12726,12729
Ferrous|12730,12737
Sulfate|12738,12745
325|12746,12749
mg|12750,12752
PO|12753,12755
DAILY|12756,12761
<EOL>|12762,12763
12.|12763,12766
Furosemide|12767,12777
40|12778,12780
mg|12781,12783
PO|12784,12786
DAILY|12787,12792
<EOL>|12793,12794
RX|12794,12796
*|12797,12798
furosemide|12798,12808
40|12809,12811
mg|12812,12814
1|12815,12816
tablet|12817,12823
(|12823,12824
s|12824,12825
)|12825,12826
by|12827,12829
mouth|12830,12835
qday|12836,12840
Disp|12841,12845
#|12846,12847
*|12847,12848
30|12848,12850
Tablet|12851,12857
<EOL>|12858,12859
Refills|12859,12866
:|12866,12867
*|12867,12868
0|12868,12869
<EOL>|12869,12870
13.|12870,12873
HumuLIN|12874,12881
70|12882,12884
/|12884,12885
30|12885,12887
(|12888,12889
insulin|12889,12896
NPH|12897,12900
and|12901,12904
regular|12905,12912
human|12913,12918
)|12918,12919
30|12920,12922
units|12923,12928
<EOL>|12929,12930
subcutaneous|12930,12942
daily|12943,12948
<EOL>|12949,12950
14.|12950,12953
Lisinopril|12954,12964
40|12965,12967
mg|12968,12970
PO|12971,12973
DAILY|12974,12979
<EOL>|12980,12981
15.|12981,12984
Carvedilol|12985,12995
12.5|12996,13000
mg|13001,13003
PO|13004,13006
BID|13007,13010
<EOL>|13011,13012
RX|13012,13014
*|13015,13016
carvedilol|13016,13026
12.5|13027,13031
mg|13032,13034
1|13035,13036
tablet|13037,13043
(|13043,13044
s|13044,13045
)|13045,13046
by|13047,13049
mouth|13050,13055
twice|13056,13061
a|13062,13063
day|13064,13067
Disp|13068,13072
<EOL>|13073,13074
#|13074,13075
*|13075,13076
60|13076,13078
Tablet|13079,13085
Refills|13086,13093
:|13093,13094
*|13094,13095
0|13095,13096
<EOL>|13096,13097
<EOL>|13097,13098
<EOL>|13099,13100
Discharge|13100,13109
Disposition|13110,13121
:|13121,13122
<EOL>|13122,13123
Home|13123,13127
With|13128,13132
Service|13133,13140
<EOL>|13140,13141
<EOL>|13142,13143
Facility|13143,13151
:|13151,13152
<EOL>|13152,13153
_|13153,13154
_|13154,13155
_|13155,13156
<EOL>|13156,13157
<EOL>|13158,13159
Discharge|13159,13168
Diagnosis|13169,13178
:|13178,13179
<EOL>|13179,13180
-|13199,13200
Acute|13201,13206
on|13207,13209
chronic|13210,13217
decompensated|13218,13231
systolic|13232,13240
heart|13241,13246
failure|13247,13254
<EOL>|13254,13255
<EOL>|13255,13256
<EOL>|13257,13258
Mental|13279,13285
Status|13286,13292
:|13292,13293
Clear|13294,13299
and|13300,13303
coherent|13304,13312
.|13312,13313
<EOL>|13313,13314
Level|13314,13319
of|13320,13322
Consciousness|13323,13336
:|13336,13337
Alert|13338,13343
and|13344,13347
interactive|13348,13359
.|13359,13360
<EOL>|13360,13361
Activity|13361,13369
Status|13370,13376
:|13376,13377
Ambulatory|13378,13388
-|13389,13390
Independent|13391,13402
.|13402,13403
<EOL>|13403,13404
<EOL>|13404,13405
<EOL>|13406,13407
Dear|13431,13435
_|13436,13437
_|13437,13438
_|13438,13439
,|13439,13440
<EOL>|13440,13441
<EOL>|13441,13442
_|13442,13443
_|13443,13444
_|13444,13445
were|13446,13450
admitted|13451,13459
to|13460,13462
_|13463,13464
_|13464,13465
_|13465,13466
on|13467,13469
_|13470,13471
_|13471,13472
_|13472,13473
with|13474,13478
shortness|13479,13488
of|13489,13491
breath|13492,13498
.|13498,13499
<EOL>|13500,13501
_|13501,13502
_|13502,13503
_|13503,13504
were|13505,13509
diagnosed|13510,13519
with|13520,13524
an|13525,13527
exacerbation|13528,13540
of|13541,13543
your|13544,13548
heart|13549,13554
failure|13555,13562
,|13562,13563
a|13564,13565
<EOL>|13566,13567
result|13567,13573
of|13574,13576
retaining|13577,13586
too|13587,13590
much|13591,13595
fluid|13596,13601
.|13601,13602
_|13603,13604
_|13604,13605
_|13605,13606
were|13607,13611
treated|13612,13619
with|13620,13624
<EOL>|13625,13626
diuretics|13626,13635
and|13636,13639
removal|13640,13647
of|13648,13650
this|13651,13655
fluid|13656,13661
with|13662,13666
subsequent|13667,13677
improvement|13678,13689
<EOL>|13690,13691
in|13691,13693
your|13694,13698
symptoms|13699,13707
.|13707,13708
We|13709,13711
also|13712,13716
increased|13717,13726
your|13727,13731
carvedilol|13732,13742
dose|13743,13747
for|13748,13751
<EOL>|13752,13753
better|13753,13759
blood|13760,13765
pressure|13766,13774
control|13775,13782
.|13782,13783
<EOL>|13783,13784
<EOL>|13784,13785
It|13785,13787
is|13788,13790
very|13791,13795
important|13796,13805
that|13806,13810
_|13811,13812
_|13812,13813
_|13813,13814
weigh|13815,13820
yourself|13821,13829
every|13830,13835
morning|13836,13843
,|13843,13844
call|13845,13849
<EOL>|13850,13851
MD|13851,13853
if|13854,13856
weight|13857,13863
goes|13864,13868
up|13869,13871
more|13872,13876
than|13877,13881
3|13882,13883
lbs|13884,13887
.|13887,13888
Taking|13889,13895
your|13896,13900
furosemide|13901,13911
<EOL>|13912,13913
will|13913,13917
keep|13918,13922
_|13923,13924
_|13924,13925
_|13925,13926
from|13927,13931
retaining|13932,13941
fluid|13942,13947
.|13947,13948
<EOL>|13948,13949
<EOL>|13949,13950
Sincerely|13950,13959
,|13959,13960
<EOL>|13960,13961
Your|13961,13965
_|13966,13967
_|13967,13968
_|13968,13969
Team|13970,13974
<EOL>|13974,13975
<EOL>|13976,13977
Followup|13977,13985
Instructions|13986,13998
:|13998,13999
<EOL>|13999,14000
_|14000,14001
_|14001,14002
_|14002,14003
<EOL>|14003,14004

