 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|26,30
No|31,33
:|33,34
_|37,38
_|38,39
_|39,40
<EOL>|40,41
<EOL>|42,43
Admission|43,52
Date|53,57
:|57,58
_|60,61
_|61,62
_|62,63
Discharge|77,86
Date|87,91
:|91,92
_|95,96
_|96,97
_|97,98
<EOL>|98,99
<EOL>|100,101
Date|101,105
of|106,108
Birth|109,114
:|114,115
_|117,118
_|118,119
_|119,120
Sex|133,136
:|136,137
F|140,141
<EOL>|141,142
<EOL>|143,144
Service|144,151
:|151,152
MEDICINE|153,161
<EOL>|161,162
<EOL>|163,164
Allergies|164,173
:|173,174
<EOL>|175,176
No|176,178
Known|179,184
Allergies|185,194
/|195,196
Adverse|197,204
Drug|205,209
Reactions|210,219
<EOL>|219,220
<EOL>|221,222
Attending|222,231
:|231,232
_|233,234
_|234,235
_|235,236
.|236,237
<EOL>|237,238
<EOL>|239,240
Chief|240,245
Complaint|246,255
:|255,256
<EOL>|256,257
Hematuria|257,266
,|266,267
weakness|268,276
<EOL>|276,277
<EOL>|278,279
Major|279,284
Surgical|285,293
or|294,296
Invasive|297,305
Procedure|306,315
:|315,316
<EOL>|316,317
None|317,321
<EOL>|321,322
<EOL>|322,323
<EOL>|324,325
History|325,332
of|333,335
Present|336,343
Illness|344,351
:|351,352
<EOL>|352,353
_|353,354
_|354,355
_|355,356
y|357,358
/|358,359
o|359,360
female|361,367
with|368,372
h|373,374
/|374,375
o|375,376
PE|377,379
(|380,381
on|381,383
lovenox|384,391
)|391,392
,|392,393
bladder|394,401
cancer|402,408
s|409,410
/|410,411
p|411,412
<EOL>|414,415
Robotic|415,422
TAH|423,426
-|426,427
BSO|427,430
,|430,431
lap|432,435
radical|436,443
cystectomy|444,454
with|455,459
ileal|460,465
loop|466,470
<EOL>|471,472
diversion|472,481
and|482,485
anterior|486,494
vaginectomy|495,506
in|507,509
_|510,511
_|511,512
_|512,513
c|514,515
/|515,516
b|516,517
abdominal|518,527
<EOL>|528,529
fluid|529,534
requiring|535,544
placement|545,554
of|555,557
drainage|558,566
catheters|567,576
.|576,577
Recent|578,584
<EOL>|585,586
abdominal|586,595
imaging|596,603
noted|604,609
worsening|610,619
of|620,622
her|623,626
bilateral|627,636
severe|637,643
<EOL>|644,645
hydronephrosis|645,659
and|660,663
her|664,667
Cr|668,670
was|671,674
noted|675,680
to|681,683
have|684,688
risen|689,694
from|695,699
0.8|700,703
to|704,706
<EOL>|707,708
1.3|708,711
(|711,712
outside|712,719
lab|720,723
value|724,729
)|729,730
.|730,731
Patient|732,739
recently|740,748
underwent|749,758
bilateral|759,768
<EOL>|769,770
nephrostomy|770,781
tube|782,786
placement|787,796
by|797,799
_|800,801
_|801,802
_|802,803
on|804,806
_|807,808
_|808,809
_|809,810
.|810,811
<EOL>|811,812
<EOL>|812,813
She|813,816
first|817,822
started|823,830
feeling|831,838
weak|839,843
during|844,850
_|851,852
_|852,853
_|853,854
yesterday|855,864
doing|865,870
the|871,874
<EOL>|875,876
exercises|876,885
.|885,886
Had|887,890
palpitations|891,903
with|904,908
ambulation|909,919
.|919,920
Has|921,924
tightness|925,934
in|935,937
<EOL>|938,939
chest|939,944
with|945,949
ambulating|950,960
since|961,966
yesterday|967,976
.|976,977
Felt|978,982
light|983,988
headed|989,995
with|996,1000
<EOL>|1001,1002
ambulation|1002,1012
.|1012,1013
SNF|1014,1017
noticed|1018,1025
increased|1026,1035
hematuria|1036,1045
with|1046,1050
R|1051,1052
bag|1053,1056
darker|1057,1063
<EOL>|1064,1065
than|1065,1069
L|1070,1071
bag|1072,1075
since|1076,1081
yesterday|1082,1091
.|1091,1092
Her|1093,1096
Urostomy|1097,1105
(|1106,1107
placed|1107,1113
in|1114,1116
_|1117,1118
_|1118,1119
_|1119,1120
<EOL>|1121,1122
also|1122,1126
positive|1127,1135
for|1136,1139
hematuria|1140,1149
.|1149,1150
She|1151,1154
was|1155,1158
transferred|1159,1170
to|1171,1173
_|1174,1175
_|1175,1176
_|1176,1177
ED|1178,1180
for|1181,1184
<EOL>|1185,1186
further|1186,1193
management|1194,1204
.|1204,1205
<EOL>|1205,1206
<EOL>|1206,1207
In|1207,1209
the|1210,1213
ED|1214,1216
,|1216,1217
initial|1218,1225
vitals|1226,1232
were|1233,1237
:|1237,1238
<EOL>|1240,1241
<EOL>|1241,1242
Temp|1242,1246
.|1246,1247
98.1|1248,1252
,|1252,1253
HR|1254,1256
72|1257,1259
,|1259,1260
BP|1261,1263
139|1264,1267
/|1267,1268
56|1268,1270
,|1270,1271
RR|1272,1274
16|1275,1277
,|1277,1278
99|1279,1281
%|1281,1282
RA|1283,1285
<EOL>|1285,1286
<EOL>|1288,1289
-|1289,1290
Labs|1291,1295
notable|1296,1303
for|1304,1307
:|1307,1308
<EOL>|1310,1311
WBC|1311,1314
5.9|1315,1318
,|1318,1319
Hg|1320,1322
8.1|1323,1326
,|1326,1327
platelets|1328,1337
374|1338,1341
.|1341,1342
Na|1343,1345
140|1346,1349
,|1349,1350
K|1351,1352
4.3|1353,1356
,|1356,1357
Cl|1358,1360
103|1361,1364
,|1364,1365
biacrb|1366,1372
<EOL>|1373,1374
22|1374,1376
,|1376,1377
BUN|1378,1381
29|1382,1384
,|1384,1385
Cr|1386,1388
1.0|1389,1392
<EOL>|1392,1393
<EOL>|1393,1394
UA|1394,1396
from|1397,1401
bilateral|1402,1411
nephrostomy|1412,1423
tubes|1424,1429
with|1430,1434
>|1435,1436
100|1437,1440
WBC|1441,1444
,|1444,1445
moderate|1446,1454
<EOL>|1455,1456
leukocytes|1456,1466
,|1466,1467
and|1468,1471
large|1472,1477
blood|1478,1483
.|1483,1484
<EOL>|1484,1485
<EOL>|1485,1486
-|1486,1487
Imaging|1488,1495
was|1496,1499
notable|1500,1507
for|1508,1511
:|1511,1512
<EOL>|1513,1514
CT|1514,1516
abd|1517,1520
/|1520,1521
pelvis|1521,1527
w|1528,1529
/|1529,1530
o|1530,1531
contrast|1532,1540
:|1540,1541
<EOL>|1541,1542
Interval|1542,1550
placement|1551,1560
of|1561,1563
bilateral|1564,1573
percutaneous|1574,1586
nephroureterostomy|1587,1605
<EOL>|1606,1607
tubes|1607,1612
with|1613,1617
resolved|1618,1626
hydroureteronephrosis|1627,1648
.|1648,1649
No|1650,1652
RP|1653,1655
hematoma|1656,1664
.|1664,1665
<EOL>|1665,1666
<EOL>|1667,1668
-|1668,1669
Patient|1670,1677
was|1678,1681
given|1682,1687
:|1687,1688
<EOL>|1690,1691
LR|1691,1693
<EOL>|1693,1694
<EOL>|1694,1695
Upon|1695,1699
arrival|1700,1707
to|1708,1710
the|1711,1714
floor|1715,1720
,|1720,1721
patient|1722,1729
reports|1730,1737
that|1738,1742
she|1743,1746
noticed|1747,1754
<EOL>|1755,1756
shortness|1756,1765
of|1766,1768
breath|1769,1775
today|1776,1781
with|1782,1786
walking|1787,1794
in|1795,1797
conjunction|1798,1809
with|1810,1814
<EOL>|1815,1816
bloody|1816,1822
output|1823,1829
from|1830,1834
her|1835,1838
ostomy|1839,1845
tubes|1846,1851
.|1851,1852
She|1853,1856
notes|1857,1862
that|1863,1867
the|1868,1871
output|1872,1878
<EOL>|1879,1880
from|1880,1884
her|1885,1888
nephrostomy|1889,1900
tubes|1901,1906
was|1907,1910
pink|1911,1915
tinged|1916,1922
when|1923,1927
she|1928,1931
left|1932,1936
the|1937,1940
<EOL>|1941,1942
hospital|1942,1950
2|1951,1952
days|1953,1957
ago|1958,1961
.|1961,1962
She|1963,1966
also|1967,1971
endorses|1972,1980
associated|1981,1991
chest|1992,1997
<EOL>|1998,1999
tightness|1999,2008
but|2009,2012
no|2013,2015
pain|2016,2020
or|2021,2023
pressure|2024,2032
.|2032,2033
She|2034,2037
denies|2038,2044
cough|2045,2050
,|2050,2051
fever|2052,2057
,|2057,2058
<EOL>|2059,2060
chills|2060,2066
,|2066,2067
abdominal|2068,2077
pain|2078,2082
,|2082,2083
or|2084,2086
diarrhea|2087,2095
.|2095,2096
She|2097,2100
notes|2101,2106
that|2107,2111
she|2112,2115
has|2116,2119
an|2120,2122
<EOL>|2123,2124
ostomy|2124,2130
and|2131,2134
nephroureterostomy|2135,2153
without|2154,2161
sensation|2162,2171
of|2172,2174
dysuria|2175,2182
.|2182,2183
<EOL>|2184,2185
Patient|2185,2192
notes|2193,2198
feeling|2199,2206
dizzy|2207,2212
and|2213,2216
lightheaded|2217,2228
previously|2229,2239
though|2240,2246
is|2247,2249
<EOL>|2250,2251
currently|2251,2260
asymptomatic|2261,2273
.|2273,2274
<EOL>|2275,2276
<EOL>|2276,2277
<EOL>|2278,2279
Past|2279,2283
Medical|2284,2291
History|2292,2299
:|2299,2300
<EOL>|2300,2301
-|2301,2302
Hypertension|2303,2315
<EOL>|2317,2318
-|2319,2320
s|2321,2322
/|2322,2323
p|2323,2324
lap|2325,2328
chole|2329,2334
<EOL>|2336,2337
-|2338,2339
s|2340,2341
/|2341,2342
p|2342,2343
left|2344,2348
knee|2349,2353
replacement|2354,2365
<EOL>|2367,2368
-|2369,2370
s|2371,2372
/|2372,2373
p|2373,2374
laminectomy|2375,2386
of|2387,2389
L5|2390,2392
-|2392,2393
S1|2393,2395
at|2396,2398
age|2399,2402
_|2403,2404
_|2404,2405
_|2405,2406
<EOL>|2408,2409
-|2410,2411
Bladder|2412,2419
Cancer|2420,2426
high|2427,2431
grade|2432,2437
TCC|2438,2441
,|2441,2442
T1|2443,2445
diagnosed|2446,2455
in|2456,2458
_|2459,2460
_|2460,2461
_|2461,2462
,|2462,2463
then|2464,2468
<EOL>|2469,2470
_|2470,2471
_|2471,2472
_|2472,2473
pelvic|2474,2480
MRI|2481,2484
w|2485,2486
/|2486,2487
invasion|2487,2495
into|2496,2500
bladder|2501,2508
wall|2509,2513
,|2513,2514
perivesical|2515,2526
<EOL>|2527,2528
soft|2528,2532
tissue|2533,2539
and|2540,2543
anterior|2544,2552
vaginal|2553,2560
wall|2561,2565
c|2566,2567
/|2567,2568
w|2568,2569
T4|2570,2572
staging|2573,2580
<EOL>|2582,2583
-|2584,2585
s|2586,2587
/|2587,2588
p|2588,2589
hysterectomy|2590,2602
and|2603,2606
bilateral|2607,2616
oophorectomy|2617,2629
for|2630,2633
large|2634,2639
uterus|2640,2646
<EOL>|2647,2648
w|2648,2649
/|2649,2650
fibroid|2650,2657
,|2657,2658
s|2659,2660
/|2660,2661
p|2661,2662
laparascopic|2663,2675
b|2676,2677
/|2677,2678
l|2678,2679
pelvic|2680,2686
lymph|2687,2692
node|2693,2697
resection|2698,2707
,|2707,2708
s|2709,2710
/|2710,2711
p|2711,2712
<EOL>|2713,2714
radical|2714,2721
cystectomy|2722,2732
and|2733,2736
anterior|2737,2745
vaginectomy|2746,2757
with|2758,2762
vaginal|2763,2770
<EOL>|2771,2772
reconstruction|2772,2786
with|2787,2791
ileal|2792,2797
conduit|2798,2805
creation|2806,2814
_|2815,2816
_|2816,2817
_|2817,2818
,|2818,2819
course|2820,2826
<EOL>|2827,2828
complicated|2828,2839
by|2840,2842
bacteremia|2843,2853
and|2854,2857
development|2858,2869
of|2870,2872
intra-abdominal|2873,2888
<EOL>|2889,2890
fluid|2890,2895
collection|2896,2906
,|2906,2907
no|2908,2910
s|2911,2912
/|2912,2913
p|2913,2914
drain|2915,2920
placement|2921,2930
by|2931,2933
_|2934,2935
_|2935,2936
_|2936,2937
_|2938,2939
_|2939,2940
_|2940,2941
<EOL>|2943,2944
-|2945,2946
h|2947,2948
/|2948,2949
o|2949,2950
LLE|2951,2954
DVT|2955,2958
and|2959,2962
PE|2963,2965
on|2966,2968
lovenox|2969,2976
<EOL>|2978,2979
<EOL>|2979,2980
<EOL>|2981,2982
Social|2982,2988
History|2989,2996
:|2996,2997
<EOL>|2997,2998
_|2998,2999
_|2999,3000
_|3000,3001
<EOL>|3001,3002
Family|3002,3008
History|3009,3016
:|3016,3017
<EOL>|3017,3018
Negative|3018,3026
for|3027,3030
bladder|3031,3038
CA|3039,3041
.|3041,3042
<EOL>|3042,3043
<EOL>|3043,3044
<EOL>|3045,3046
Physical|3046,3054
Exam|3055,3059
:|3059,3060
<EOL>|3060,3061
=|3061,3062
=|3062,3063
=|3063,3064
=|3064,3065
=|3065,3066
=|3066,3067
=|3067,3068
=|3068,3069
=|3069,3070
=|3070,3071
=|3071,3072
=|3072,3073
=|3073,3074
=|3074,3075
=|3075,3076
=|3076,3077
=|3077,3078
=|3078,3079
=|3079,3080
=|3080,3081
=|3081,3082
=|3082,3083
=|3083,3084
=|3084,3085
=|3085,3086
<EOL>|3086,3087
ADMISSION|3087,3096
PHYSICAL|3097,3105
EXAM|3106,3110
:|3110,3111
<EOL>|3112,3113
=|3113,3114
=|3114,3115
=|3115,3116
=|3116,3117
=|3117,3118
=|3118,3119
=|3119,3120
=|3120,3121
=|3121,3122
=|3122,3123
=|3123,3124
=|3124,3125
=|3125,3126
=|3126,3127
=|3127,3128
=|3128,3129
=|3129,3130
=|3130,3131
=|3131,3132
=|3132,3133
=|3133,3134
=|3134,3135
=|3135,3136
=|3136,3137
=|3137,3138
<EOL>|3139,3140
VITAL|3140,3145
SIGNS|3146,3151
:|3151,3152
Temp|3153,3157
.|3157,3158
98.1|3159,3163
PO|3164,3166
BP|3167,3169
158|3170,3173
/|3174,3175
66|3176,3178
HR|3179,3181
72|3182,3184
RR|3185,3187
18|3188,3190
Spo2|3191,3195
95|3196,3198
RA|3199,3201
<EOL>|3202,3203
GENERAL|3203,3210
:|3210,3211
well|3212,3216
-|3216,3217
appearing|3217,3226
elderly|3227,3234
woman|3235,3240
in|3241,3243
no|3244,3246
acute|3247,3252
distress|3253,3261
<EOL>|3262,3263
CARDIAC|3263,3270
:|3270,3271
RRR|3272,3275
,|3275,3276
no|3277,3279
murmurs|3280,3287
<EOL>|3287,3288
LUNGS|3288,3293
:|3293,3294
clear|3295,3300
to|3301,3303
auscultation|3304,3316
bilaterally|3317,3328
<EOL>|3329,3330
ABDOMEN|3330,3337
:|3337,3338
soft|3339,3343
,|3343,3344
non-tender|3345,3355
to|3356,3358
palpation|3359,3368
,|3368,3369
normal|3370,3376
bowel|3377,3382
sounds|3383,3389
.|3389,3390
<EOL>|3391,3392
Ostomy|3392,3398
draining|3399,3407
brown|3408,3413
stool|3414,3419
.|3419,3420
Nephroureterostomy|3421,3439
draining|3440,3448
dark|3449,3453
<EOL>|3454,3455
red|3455,3458
bloody|3459,3465
urine|3466,3471
.|3471,3472
Bilateral|3473,3482
nephrostomy|3483,3494
tubes|3495,3500
draining|3501,3509
blood|3510,3515
<EOL>|3516,3517
urine|3517,3522
.|3522,3523
<EOL>|3524,3525
EXTREMITIES|3525,3536
:|3536,3537
No|3538,3540
edema|3541,3546
,|3546,3547
warm|3548,3552
and|3553,3556
well|3557,3561
-|3561,3562
perfused|3562,3570
.|3570,3571
<EOL>|3571,3572
<EOL>|3572,3573
=|3573,3574
=|3574,3575
=|3575,3576
=|3576,3577
=|3577,3578
=|3578,3579
=|3579,3580
=|3580,3581
=|3581,3582
=|3582,3583
=|3583,3584
=|3584,3585
=|3585,3586
=|3586,3587
=|3587,3588
=|3588,3589
=|3589,3590
=|3590,3591
=|3591,3592
=|3592,3593
=|3593,3594
=|3594,3595
=|3595,3596
=|3596,3597
=|3597,3598
<EOL>|3598,3599
DISCHARGE|3599,3608
PHYSICAL|3609,3617
EXAM|3618,3622
:|3622,3623
<EOL>|3624,3625
=|3625,3626
=|3626,3627
=|3627,3628
=|3628,3629
=|3629,3630
=|3630,3631
=|3631,3632
=|3632,3633
=|3633,3634
=|3634,3635
=|3635,3636
=|3636,3637
=|3637,3638
=|3638,3639
=|3639,3640
=|3640,3641
=|3641,3642
=|3642,3643
=|3643,3644
=|3644,3645
=|3645,3646
=|3646,3647
=|3647,3648
=|3648,3649
=|3649,3650
<EOL>|3651,3652
VS|3652,3654
-|3655,3656
98.3|3658,3662
PO|3663,3665
139|3666,3669
/|3669,3670
67|3670,3672
71|3673,3675
18|3676,3678
94|3679,3681
RA|3682,3684
<EOL>|3685,3686
GENERAL|3686,3693
:|3693,3694
well|3695,3699
-|3699,3700
appearing|3700,3709
elderly|3710,3717
woman|3718,3723
in|3724,3726
no|3727,3729
acute|3730,3735
distress|3736,3744
<EOL>|3745,3746
CARDIAC|3746,3753
:|3753,3754
RRR|3755,3758
,|3758,3759
no|3760,3762
murmurs|3763,3770
<EOL>|3770,3771
LUNGS|3771,3776
:|3776,3777
clear|3778,3783
to|3784,3786
auscultation|3787,3799
bilaterally|3800,3811
<EOL>|3812,3813
ABDOMEN|3813,3820
:|3820,3821
soft|3822,3826
,|3826,3827
non-tender|3828,3838
to|3839,3841
palpation|3842,3851
,|3851,3852
normal|3853,3859
bowel|3860,3865
sounds|3866,3872
.|3872,3873
<EOL>|3875,3876
Nephroureterostomy|3876,3894
draining|3895,3903
dark|3904,3908
red|3909,3912
bloody|3913,3919
urine|3920,3925
.|3925,3926
Bilateral|3927,3936
<EOL>|3937,3938
nephrostomy|3938,3949
tubes|3950,3955
capped|3956,3962
.|3962,3963
<EOL>|3964,3965
EXTREMITIES|3965,3976
:|3976,3977
No|3978,3980
edema|3981,3986
,|3986,3987
warm|3988,3992
and|3993,3996
well|3997,4001
-|4001,4002
perfused|4002,4010
<EOL>|4010,4011
<EOL>|4011,4012
<EOL>|4013,4014
Pertinent|4014,4023
Results|4024,4031
:|4031,4032
<EOL>|4032,4033
=|4033,4034
=|4034,4035
=|4035,4036
=|4036,4037
=|4037,4038
=|4038,4039
=|4039,4040
=|4040,4041
=|4041,4042
=|4042,4043
=|4043,4044
=|4044,4045
=|4045,4046
=|4046,4047
=|4047,4048
=|4048,4049
<EOL>|4049,4050
ADMISSION|4050,4059
LABS|4060,4064
<EOL>|4064,4065
=|4065,4066
=|4066,4067
=|4067,4068
=|4068,4069
=|4069,4070
=|4070,4071
=|4071,4072
=|4072,4073
=|4073,4074
=|4074,4075
=|4075,4076
=|4076,4077
=|4077,4078
=|4078,4079
=|4079,4080
=|4080,4081
<EOL>|4081,4082
_|4082,4083
_|4083,4084
_|4084,4085
05|4086,4088
:|4088,4089
20PM|4089,4093
BLOOD|4094,4099
WBC|4100,4103
-|4103,4104
5.9|4104,4107
RBC|4108,4111
-|4111,4112
2|4112,4113
.|4113,4114
90|4114,4116
*|4116,4117
Hgb|4118,4121
-|4121,4122
8|4122,4123
.|4123,4124
1|4124,4125
*|4125,4126
Hct|4127,4130
-|4130,4131
26|4131,4133
.|4133,4134
6|4134,4135
*|4135,4136
<EOL>|4137,4138
MCV|4138,4141
-|4141,4142
92|4142,4144
MCH|4145,4148
-|4148,4149
27.9|4149,4153
MCHC|4154,4158
-|4158,4159
30|4159,4161
.|4161,4162
5|4162,4163
*|4163,4164
RDW|4165,4168
-|4168,4169
15.4|4169,4173
RDWSD|4174,4179
-|4179,4180
51|4180,4182
.|4182,4183
2|4183,4184
*|4184,4185
Plt|4186,4189
_|4190,4191
_|4191,4192
_|4192,4193
<EOL>|4193,4194
_|4194,4195
_|4195,4196
_|4196,4197
05|4198,4200
:|4200,4201
48AM|4201,4205
BLOOD|4206,4211
WBC|4212,4215
-|4215,4216
4.6|4216,4219
RBC|4220,4223
-|4223,4224
2|4224,4225
.|4225,4226
46|4226,4228
*|4228,4229
Hgb|4230,4233
-|4233,4234
7|4234,4235
.|4235,4236
0|4236,4237
*|4237,4238
Hct|4239,4242
-|4242,4243
22|4243,4245
.|4245,4246
6|4246,4247
*|4247,4248
<EOL>|4249,4250
MCV|4250,4253
-|4253,4254
92|4254,4256
MCH|4257,4260
-|4260,4261
28.5|4261,4265
MCHC|4266,4270
-|4270,4271
31|4271,4273
.|4273,4274
0|4274,4275
*|4275,4276
RDW|4277,4280
-|4280,4281
15.3|4281,4285
RDWSD|4286,4291
-|4291,4292
51|4292,4294
.|4294,4295
7|4295,4296
*|4296,4297
Plt|4298,4301
_|4302,4303
_|4303,4304
_|4304,4305
<EOL>|4305,4306
_|4306,4307
_|4307,4308
_|4308,4309
05|4310,4312
:|4312,4313
20PM|4313,4317
BLOOD|4318,4323
Neuts|4324,4329
-|4329,4330
56.3|4330,4334
_|4335,4336
_|4336,4337
_|4337,4338
Monos|4339,4344
-|4344,4345
12.6|4345,4349
Eos|4350,4353
-|4353,4354
1.5|4354,4357
<EOL>|4358,4359
Baso|4359,4363
-|4363,4364
0.3|4364,4367
Im|4368,4370
_|4371,4372
_|4372,4373
_|4373,4374
AbsNeut|4375,4382
-|4382,4383
3|4383,4384
.|4384,4385
29|4385,4387
#|4387,4388
AbsLymp|4389,4396
-|4396,4397
1|4397,4398
.|4398,4399
69|4399,4401
AbsMono|4402,4409
-|4409,4410
0|4410,4411
.|4411,4412
74|4412,4414
<EOL>|4415,4416
AbsEos|4416,4422
-|4422,4423
0|4423,4424
.|4424,4425
09|4425,4427
AbsBaso|4428,4435
-|4435,4436
0|4436,4437
.|4437,4438
02|4438,4440
<EOL>|4440,4441
_|4441,4442
_|4442,4443
_|4443,4444
05|4445,4447
:|4447,4448
20PM|4448,4452
BLOOD|4453,4458
Glucose|4459,4466
-|4466,4467
101|4467,4470
*|4470,4471
UreaN|4472,4477
-|4477,4478
29|4478,4480
*|4480,4481
Creat|4482,4487
-|4487,4488
1.0|4488,4491
Na|4492,4494
-|4494,4495
140|4495,4498
<EOL>|4499,4500
K|4500,4501
-|4501,4502
4.3|4502,4505
Cl|4506,4508
-|4508,4509
103|4509,4512
HCO3|4513,4517
-|4517,4518
22|4518,4520
AnGap|4521,4526
-|4526,4527
19|4527,4529
<EOL>|4529,4530
<EOL>|4530,4531
=|4531,4532
=|4532,4533
=|4533,4534
=|4534,4535
=|4535,4536
=|4536,4537
=|4537,4538
=|4538,4539
=|4539,4540
=|4540,4541
=|4541,4542
=|4542,4543
=|4543,4544
=|4544,4545
=|4545,4546
=|4546,4547
=|4547,4548
<EOL>|4548,4549
IMAGING|4549,4556
/|4556,4557
STUDIES|4557,4564
<EOL>|4564,4565
=|4565,4566
=|4566,4567
=|4567,4568
=|4568,4569
=|4569,4570
=|4570,4571
=|4571,4572
=|4572,4573
=|4573,4574
=|4574,4575
=|4575,4576
=|4576,4577
=|4577,4578
=|4578,4579
=|4579,4580
=|4580,4581
=|4581,4582
<EOL>|4582,4583
<EOL>|4583,4584
_|4584,4585
_|4585,4586
_|4586,4587
CT|4588,4590
Abd|4591,4594
/|4594,4595
Pel|4595,4598
w|4599,4600
/|4600,4601
o|4601,4602
Contrast|4603,4611
:|4611,4612
<EOL>|4613,4614
IMPRESSION|4614,4624
:|4624,4625
<EOL>|4628,4629
1.|4629,4631
Interval|4632,4640
placement|4641,4650
of|4651,4653
bilateral|4654,4663
percutaneous|4664,4676
<EOL>|4677,4678
nephroureterostomy|4678,4696
tubes|4697,4702
with|4703,4707
resolved|4708,4716
hydroureteronephrosis|4717,4738
.|4738,4739
<EOL>|4741,4742
No|4742,4744
RP|4745,4747
hematoma|4748,4756
.|4756,4757
<EOL>|4758,4759
2.|4759,4761
Partially|4762,4771
imaged|4772,4778
nodular|4779,4786
opacity|4787,4794
in|4795,4797
the|4798,4801
right|4802,4807
middle|4808,4814
lobe|4815,4819
<EOL>|4820,4821
which|4821,4826
can|4827,4830
be|4831,4833
<EOL>|4834,4835
further|4835,4842
assessed|4843,4851
on|4852,4854
a|4855,4856
nonemergent|4857,4868
dedicated|4869,4878
CT|4879,4881
chest|4882,4887
.|4887,4888
<EOL>|4889,4890
<EOL>|4890,4891
_|4891,4892
_|4892,4893
_|4893,4894
CXR|4895,4898
<EOL>|4898,4899
AP|4899,4901
portable|4902,4910
upright|4911,4918
view|4919,4923
of|4924,4926
the|4927,4930
chest|4931,4936
.|4936,4937
Right|4940,4945
upper|4946,4951
extremity|4952,4961
<EOL>|4962,4963
access|4963,4969
PICC|4970,4974
<EOL>|4975,4976
line|4976,4980
is|4981,4983
seen|4984,4988
with|4989,4993
its|4994,4997
tip|4998,5001
in|5002,5004
the|5005,5008
upper|5009,5014
SVC|5015,5018
.|5018,5019
Overlying|5021,5030
EKG|5031,5034
leads|5035,5040
<EOL>|5041,5042
are|5042,5045
present|5046,5053
.|5053,5054
Lungs|5056,5061
are|5062,5065
clear|5066,5071
.|5071,5072
Cardiomediastinal|5074,5091
silhouette|5092,5102
is|5103,5105
<EOL>|5106,5107
stable|5107,5113
.|5113,5114
Bony|5116,5120
structures|5121,5131
are|5132,5135
intact|5136,5142
.|5142,5143
<EOL>|5144,5145
<EOL>|5145,5146
=|5146,5147
=|5147,5148
=|5148,5149
=|5149,5150
=|5150,5151
=|5151,5152
=|5152,5153
=|5153,5154
=|5154,5155
=|5155,5156
=|5156,5157
=|5157,5158
=|5158,5159
=|5159,5160
<EOL>|5160,5161
MICROBIOLOGY|5161,5173
<EOL>|5173,5174
=|5174,5175
=|5175,5176
=|5176,5177
=|5177,5178
=|5178,5179
=|5179,5180
=|5180,5181
=|5181,5182
=|5182,5183
=|5183,5184
=|5184,5185
=|5185,5186
=|5186,5187
=|5187,5188
<EOL>|5188,5189
_|5189,5190
_|5190,5191
_|5191,5192
6|5193,5194
:|5194,5195
35|5195,5197
pm|5198,5200
URINE|5201,5206
LEFT|5212,5216
NEPHROSTOMY|5217,5228
TUBE|5229,5233
.|5233,5234
<EOL>|5235,5236
*|5264,5265
*|5265,5266
FINAL|5266,5271
REPORT|5272,5278
_|5279,5280
_|5280,5281
_|5281,5282
<EOL>|5282,5283
URINE|5286,5291
CULTURE|5292,5299
(|5300,5301
Final|5301,5306
_|5307,5308
_|5308,5309
_|5309,5310
:|5310,5311
NO|5315,5317
GROWTH|5318,5324
.|5324,5325
<EOL>|5326,5327
<EOL>|5327,5328
=|5328,5329
=|5329,5330
=|5330,5331
=|5331,5332
=|5332,5333
=|5333,5334
=|5334,5335
=|5335,5336
=|5336,5337
=|5337,5338
=|5338,5339
=|5339,5340
=|5340,5341
=|5341,5342
=|5342,5343
=|5343,5344
<EOL>|5344,5345
DISCHARGE|5345,5354
LABS|5355,5359
<EOL>|5359,5360
=|5360,5361
=|5361,5362
=|5362,5363
=|5363,5364
=|5364,5365
=|5365,5366
=|5366,5367
=|5367,5368
=|5368,5369
=|5369,5370
=|5370,5371
=|5371,5372
=|5372,5373
=|5373,5374
=|5374,5375
=|5375,5376
<EOL>|5376,5377
_|5377,5378
_|5378,5379
_|5379,5380
05|5381,5383
:|5383,5384
08AM|5384,5388
BLOOD|5389,5394
WBC|5395,5398
-|5398,5399
5.4|5399,5402
RBC|5403,5406
-|5406,5407
2|5407,5408
.|5408,5409
86|5409,5411
*|5411,5412
Hgb|5413,5416
-|5416,5417
8|5417,5418
.|5418,5419
2|5419,5420
*|5420,5421
Hct|5422,5425
-|5425,5426
26|5426,5428
.|5428,5429
5|5429,5430
*|5430,5431
<EOL>|5432,5433
MCV|5433,5436
-|5436,5437
93|5437,5439
MCH|5440,5443
-|5443,5444
28.7|5444,5448
MCHC|5449,5453
-|5453,5454
30|5454,5456
.|5456,5457
9|5457,5458
*|5458,5459
RDW|5460,5463
-|5463,5464
15.3|5464,5468
RDWSD|5469,5474
-|5474,5475
51|5475,5477
.|5477,5478
8|5478,5479
*|5479,5480
Plt|5481,5484
_|5485,5486
_|5486,5487
_|5487,5488
<EOL>|5488,5489
_|5489,5490
_|5490,5491
_|5491,5492
05|5493,5495
:|5495,5496
08AM|5496,5500
BLOOD|5501,5506
Glucose|5507,5514
-|5514,5515
94|5515,5517
UreaN|5518,5523
-|5523,5524
29|5524,5526
*|5526,5527
Creat|5528,5533
-|5533,5534
0.9|5534,5537
Na|5538,5540
-|5540,5541
143|5541,5544
<EOL>|5545,5546
K|5546,5547
-|5547,5548
4.0|5548,5551
Cl|5552,5554
-|5554,5555
106|5555,5558
HCO3|5559,5563
-|5563,5564
26|5564,5566
AnGap|5567,5572
-|5572,5573
15|5573,5575
<EOL>|5575,5576
_|5576,5577
_|5577,5578
_|5578,5579
05|5580,5582
:|5582,5583
08AM|5583,5587
BLOOD|5588,5593
Calcium|5594,5601
-|5601,5602
8.8|5602,5605
Phos|5606,5610
-|5610,5611
5|5611,5612
.|5612,5613
2|5613,5614
*|5614,5615
Mg|5616,5618
-|5618,5619
2.1|5619,5622
<EOL>|5622,5623
<EOL>|5624,5625
Brief|5625,5630
Hospital|5631,5639
Course|5640,5646
:|5646,5647
<EOL>|5647,5648
Ms.|5648,5651
_|5652,5653
_|5653,5654
_|5654,5655
is|5656,5658
an|5659,5661
_|5662,5663
_|5663,5664
_|5664,5665
year|5666,5670
old|5671,5674
woman|5675,5680
with|5681,5685
history|5686,5693
of|5694,5696
provoked|5697,5705
<EOL>|5706,5707
DVT|5707,5710
/|5710,5711
PE|5711,5713
(|5714,5715
on|5715,5717
lovenox|5718,5725
)|5725,5726
,|5726,5727
bladder|5728,5735
cancer|5736,5742
s|5743,5744
/|5744,5745
p|5745,5746
Robotic|5747,5754
TAH|5755,5758
-|5758,5759
BSO|5759,5762
,|5762,5763
lap|5764,5767
<EOL>|5768,5769
radical|5769,5776
cystectomy|5777,5787
with|5788,5792
ileal|5793,5798
loop|5799,5803
diversion|5804,5813
and|5814,5817
anterior|5818,5826
<EOL>|5827,5828
vaginectomy|5828,5839
in|5840,5842
_|5843,5844
_|5844,5845
_|5845,5846
c|5847,5848
/|5848,5849
b|5849,5850
abdominal|5851,5860
fluid|5861,5866
requiring|5867,5876
<EOL>|5877,5878
placement|5878,5887
of|5888,5890
drainage|5891,5899
catheters|5900,5909
,|5909,5910
and|5911,5914
recent|5915,5921
hydronephrosis|5922,5936
<EOL>|5937,5938
requiring|5938,5947
placement|5948,5957
of|5958,5960
bilateral|5961,5970
PCN|5971,5974
tubes|5975,5980
on|5981,5983
_|5984,5985
_|5985,5986
_|5986,5987
,|5987,5988
presenting|5989,5999
<EOL>|6000,6001
from|6001,6005
rehab|6006,6011
with|6012,6016
hematuria|6017,6026
and|6027,6030
weakness|6031,6039
.|6039,6040
<EOL>|6040,6041
<EOL>|6041,6042
On|6042,6044
arrival|6045,6052
,|6052,6053
pt|6054,6056
had|6057,6060
evidence|6061,6069
of|6070,6072
frank|6073,6078
hematuria|6079,6088
in|6089,6091
her|6092,6095
urostomy|6096,6104
<EOL>|6105,6106
bag|6106,6109
and|6110,6113
PCN|6114,6117
tubes|6118,6123
.|6123,6124
Her|6125,6128
hemoglobin|6129,6139
was|6140,6143
initially|6144,6153
8.1|6154,6157
,|6157,6158
which|6159,6164
<EOL>|6165,6166
subsequently|6166,6178
dropped|6179,6186
to|6187,6189
7.0|6190,6193
Her|6194,6197
lovenox|6198,6205
was|6206,6209
held|6210,6214
,|6214,6215
and|6216,6219
she|6220,6223
was|6224,6227
<EOL>|6228,6229
transfused|6229,6239
with|6240,6244
1|6245,6246
U|6247,6248
PRBC|6249,6253
with|6254,6258
an|6259,6261
appropriate|6262,6273
hemoglobin|6274,6284
bump|6285,6289
to|6290,6292
<EOL>|6293,6294
8.2|6294,6297
.|6297,6298
Hematuria|6299,6308
was|6309,6312
likely|6313,6319
caused|6320,6326
by|6327,6329
recent|6330,6336
instrumentation|6337,6352
in|6353,6355
<EOL>|6356,6357
the|6357,6360
setting|6361,6368
of|6369,6371
anticoagulation|6372,6387
.|6387,6388
Her|6389,6392
hematuria|6393,6402
improved|6403,6411
,|6411,6412
as|6413,6415
did|6416,6419
<EOL>|6420,6421
her|6421,6424
dizziness|6425,6434
/|6434,6435
weakness|6435,6443
.|6443,6444
_|6445,6446
_|6446,6447
_|6447,6448
was|6449,6452
consulted|6453,6462
and|6463,6466
recommending|6467,6479
<EOL>|6480,6481
capping|6481,6488
her|6489,6492
PCN|6493,6496
tubes|6497,6502
.|6502,6503
After|6504,6509
discussion|6510,6520
with|6521,6525
the|6526,6529
patient|6530,6537
's|6537,6539
<EOL>|6540,6541
hematologist|6541,6553
,|6553,6554
it|6555,6557
was|6558,6561
decided|6562,6569
to|6570,6572
stop|6573,6577
her|6578,6581
lovenox|6582,6589
treatment|6590,6599
given|6600,6605
<EOL>|6606,6607
that|6607,6611
her|6612,6615
DVT|6616,6619
/|6619,6620
PE|6620,6622
were|6623,6627
provoked|6628,6636
in|6637,6639
the|6640,6643
setting|6644,6651
of|6652,6654
her|6655,6658
recovery|6659,6667
<EOL>|6668,6669
from|6669,6673
surgery|6674,6681
,|6681,6682
and|6683,6686
that|6687,6691
she|6692,6695
had|6696,6699
received|6700,6708
almost|6709,6715
6|6716,6717
months|6718,6724
of|6725,6727
<EOL>|6728,6729
treatment|6729,6738
.|6738,6739
<EOL>|6739,6740
<EOL>|6740,6741
Secondary|6741,6750
Issues|6751,6757
:|6757,6758
<EOL>|6758,6759
<EOL>|6759,6760
#|6760,6761
Asymptomatic|6762,6774
bacteruria|6775,6785
:|6785,6786
Patient|6787,6794
with|6795,6799
asymptomatic|6800,6812
bacteruria|6813,6823
<EOL>|6824,6825
in|6825,6827
setting|6828,6835
of|6836,6838
recent|6839,6845
procedural|6846,6856
manipulation|6857,6869
.|6869,6870
She|6871,6874
was|6875,6878
afebrile|6879,6887
<EOL>|6888,6889
and|6889,6892
without|6893,6900
leukocytosis|6901,6913
,|6913,6914
so|6915,6917
treatment|6918,6927
with|6928,6932
antibiotics|6933,6944
was|6945,6948
<EOL>|6949,6950
deferred|6950,6958
.|6958,6959
<EOL>|6959,6960
<EOL>|6960,6961
#|6961,6962
Hyperlipidemia|6963,6977
:|6977,6978
continued|6979,6988
atorvastatin|6989,7001
10|7002,7004
mg|7005,7007
daily|7008,7013
<EOL>|7013,7014
<EOL>|7014,7015
#|7015,7016
Hypothyroidism|7017,7031
:|7031,7032
continue|7033,7041
levothyroxine|7042,7055
175|7056,7059
mcg|7060,7063
daily|7064,7069
<EOL>|7069,7070
<EOL>|7070,7071
=|7071,7072
=|7072,7073
=|7073,7074
=|7074,7075
=|7075,7076
=|7076,7077
=|7077,7078
=|7078,7079
=|7079,7080
=|7080,7081
=|7081,7082
=|7082,7083
=|7083,7084
=|7084,7085
=|7085,7086
=|7086,7087
=|7087,7088
=|7088,7089
=|7089,7090
<EOL>|7090,7091
TRANSITIONAL|7091,7103
ISSUES|7104,7110
<EOL>|7110,7111
=|7111,7112
=|7112,7113
=|7113,7114
=|7114,7115
=|7115,7116
=|7116,7117
=|7117,7118
=|7118,7119
=|7119,7120
=|7120,7121
=|7121,7122
=|7122,7123
=|7123,7124
=|7124,7125
=|7125,7126
=|7126,7127
=|7127,7128
=|7128,7129
=|7129,7130
<EOL>|7130,7131
Medication|7131,7141
Changes|7142,7149
:|7149,7150
Lovenox|7151,7158
stopped|7159,7166
<EOL>|7167,7168
[|7168,7169
]|7170,7171
CT|7172,7174
Abdomen|7175,7182
/|7182,7183
Pelvis|7183,7189
showed|7190,7196
partially|7197,7206
imaged|7207,7213
nodular|7214,7221
opacity|7222,7229
in|7230,7232
<EOL>|7233,7234
the|7234,7237
right|7238,7243
middle|7244,7250
lobe|7251,7255
which|7256,7261
can|7262,7265
be|7266,7268
further|7269,7276
assessed|7277,7285
on|7286,7288
a|7289,7290
<EOL>|7291,7292
nonemergent|7292,7303
dedicated|7304,7313
CT|7314,7316
chest|7317,7322
.|7322,7323
<EOL>|7324,7325
[|7325,7326
]|7327,7328
Pt|7329,7331
's|7331,7333
PCN|7334,7337
tubes|7338,7343
were|7344,7348
capped|7349,7355
per|7356,7359
_|7360,7361
_|7361,7362
_|7362,7363
recommendation|7364,7378
during|7379,7385
her|7386,7389
<EOL>|7390,7391
hospitalization|7391,7406
;|7406,7407
she|7408,7411
was|7412,7415
discharged|7416,7426
with|7427,7431
scheduled|7432,7441
followup|7442,7450
to|7451,7453
<EOL>|7454,7455
decide|7455,7461
on|7462,7464
long|7465,7469
term|7470,7474
management|7475,7485
<EOL>|7485,7486
[|7486,7487
]|7488,7489
If|7490,7492
pt|7493,7495
develops|7496,7504
hematuria|7505,7514
and|7515,7518
/|7518,7519
or|7519,7521
lightheadedness|7522,7537
or|7538,7540
other|7541,7546
<EOL>|7547,7548
symptoms|7548,7556
of|7557,7559
anemia|7560,7566
,|7566,7567
a|7568,7569
CBC|7570,7573
should|7574,7580
be|7581,7583
rechecked|7584,7593
to|7594,7596
assess|7597,7603
for|7604,7607
<EOL>|7608,7609
bleeding|7609,7617
<EOL>|7617,7618
[|7618,7619
]|7620,7621
Hemoglobin|7622,7632
/|7632,7633
Hematocrit|7633,7643
on|7644,7646
discharge|7647,7656
:|7656,7657
8.2|7658,7661
/|7661,7662
26.5|7662,7666
<EOL>|7666,7667
<EOL>|7667,7668
#|7668,7669
CODE|7670,7674
:|7674,7675
presumed|7676,7684
full|7685,7689
<EOL>|7689,7690
#|7690,7691
CONTACT|7692,7699
:|7699,7700
_|7701,7702
_|7702,7703
_|7703,7704
(|7705,7706
MD|7706,7708
)|7708,7709
_|7710,7711
_|7711,7712
_|7712,7713
(|7714,7715
cell|7715,7719
)|7719,7720
<EOL>|7721,7722
_|7722,7723
_|7723,7724
_|7724,7725
(|7726,7727
home|7727,7731
)|7731,7732
<EOL>|7733,7734
<EOL>|7734,7735
<EOL>|7736,7737
Medications|7737,7748
on|7749,7751
Admission|7752,7761
:|7761,7762
<EOL>|7762,7763
The|7763,7766
Preadmission|7767,7779
Medication|7780,7790
list|7791,7795
is|7796,7798
accurate|7799,7807
and|7808,7811
complete|7812,7820
.|7820,7821
<EOL>|7821,7822
1.|7822,7824
Atorvastatin|7825,7837
10|7838,7840
mg|7841,7843
PO|7844,7846
QPM|7847,7850
<EOL>|7851,7852
2.|7852,7854
Enoxaparin|7855,7865
Sodium|7866,7872
70|7873,7875
mg|7876,7878
SC|7879,7881
Q12H|7882,7886
<EOL>|7887,7888
Start|7888,7893
:|7893,7894
_|7895,7896
_|7896,7897
_|7897,7898
,|7898,7899
First|7900,7905
Dose|7906,7910
:|7910,7911
Next|7912,7916
Routine|7917,7924
Administration|7925,7939
Time|7940,7944
<EOL>|7945,7946
3.|7946,7948
Levothyroxine|7949,7962
Sodium|7963,7969
175|7970,7973
mcg|7974,7977
PO|7978,7980
DAILY|7981,7986
<EOL>|7987,7988
4.|7988,7990
Multivitamins|7991,8004
1|8005,8006
TAB|8007,8010
PO|8011,8013
DAILY|8014,8019
<EOL>|8020,8021
5.|8021,8023
Probiotic|8024,8033
-|8033,8034
Digestive|8034,8043
Enzymes|8044,8051
(|8052,8053
L.|8053,8055
acidophilus|8056,8067
-|8067,8068
dig|8068,8071
_|8072,8073
_|8073,8074
_|8074,8075
5|8076,8077
)|8077,8078
<EOL>|8079,8080
_|8080,8081
_|8081,8082
_|8082,8083
mg|8084,8086
oral|8087,8091
daily|8092,8097
<EOL>|8098,8099
<EOL>|8099,8100
<EOL>|8101,8102
Discharge|8102,8111
Medications|8112,8123
:|8123,8124
<EOL>|8124,8125
1.|8125,8127
Atorvastatin|8129,8141
10|8142,8144
mg|8145,8147
PO|8148,8150
QPM|8151,8154
<EOL>|8156,8157
2.|8157,8159
Levothyroxine|8161,8174
Sodium|8175,8181
175|8182,8185
mcg|8186,8189
PO|8190,8192
DAILY|8193,8198
<EOL>|8200,8201
3.|8201,8203
Multivitamins|8205,8218
1|8219,8220
TAB|8221,8224
PO|8225,8227
DAILY|8228,8233
<EOL>|8235,8236
4.|8236,8238
Probiotic|8240,8249
-|8249,8250
Digestive|8250,8259
Enzymes|8260,8267
(|8268,8269
L.|8269,8271
acidophilus|8272,8283
-|8283,8284
dig|8284,8287
_|8288,8289
_|8289,8290
_|8290,8291
5|8292,8293
)|8293,8294
<EOL>|8295,8296
_|8296,8297
_|8297,8298
_|8298,8299
mg|8300,8302
oral|8303,8307
daily|8308,8313
<EOL>|8315,8316
<EOL>|8316,8317
<EOL>|8318,8319
Discharge|8319,8328
Disposition|8329,8340
:|8340,8341
<EOL>|8341,8342
Extended|8342,8350
Care|8351,8355
<EOL>|8355,8356
<EOL>|8357,8358
Facility|8358,8366
:|8366,8367
<EOL>|8367,8368
_|8368,8369
_|8369,8370
_|8370,8371
<EOL>|8371,8372
<EOL>|8373,8374
Discharge|8374,8383
Diagnosis|8384,8393
:|8393,8394
<EOL>|8394,8395
Primary|8395,8402
Diagnoses|8403,8412
:|8412,8413
Hematuria|8414,8423
,|8423,8424
anemia|8425,8431
<EOL>|8431,8432
<EOL>|8432,8433
Secondary|8433,8442
Diagnoses|8443,8452
:|8452,8453
Bladder|8454,8461
cancer|8462,8468
,|8468,8469
hydronephrosis|8470,8484
,|8484,8485
<EOL>|8486,8487
hypothyroidism|8487,8501
,|8501,8502
DVT|8503,8506
/|8506,8507
PE|8507,8509
<EOL>|8509,8510
<EOL>|8510,8511
<EOL>|8512,8513
Discharge|8513,8522
Condition|8523,8532
:|8532,8533
<EOL>|8533,8534
Mental|8534,8540
Status|8541,8547
:|8547,8548
Clear|8549,8554
and|8555,8558
coherent|8559,8567
.|8567,8568
<EOL>|8568,8569
Level|8569,8574
of|8575,8577
Consciousness|8578,8591
:|8591,8592
Alert|8593,8598
and|8599,8602
interactive|8603,8614
.|8614,8615
<EOL>|8615,8616
Activity|8616,8624
Status|8625,8631
:|8631,8632
Ambulatory|8633,8643
-|8644,8645
Independent|8646,8657
.|8657,8658
<EOL>|8658,8659
<EOL>|8659,8660
<EOL>|8661,8662
Discharge|8662,8671
Instructions|8672,8684
:|8684,8685
<EOL>|8685,8686
Dear|8686,8690
Ms.|8691,8694
_|8695,8696
_|8696,8697
_|8697,8698
,|8698,8699
<EOL>|8700,8701
<EOL>|8701,8702
It|8702,8704
was|8705,8708
a|8709,8710
pleasure|8711,8719
taking|8720,8726
care|8727,8731
of|8732,8734
you|8735,8738
at|8739,8741
_|8742,8743
_|8743,8744
_|8744,8745
.|8745,8746
<EOL>|8747,8748
<EOL>|8748,8749
WHY|8749,8752
DID|8753,8756
YOU|8757,8760
COME|8761,8765
TO|8766,8768
THE|8769,8772
HOSPITAL|8773,8781
?|8781,8782
<EOL>|8782,8783
You|8783,8786
noticed|8787,8794
blood|8795,8800
in|8801,8803
your|8804,8808
urine|8809,8814
,|8814,8815
and|8816,8819
you|8820,8823
were|8824,8828
feeling|8829,8836
<EOL>|8837,8838
weak|8838,8842
/|8842,8843
lightheaded|8843,8854
.|8854,8855
<EOL>|8855,8856
<EOL>|8856,8857
WHAT|8857,8861
HAPPENED|8862,8870
WHILE|8871,8876
YOU|8877,8880
WERE|8881,8885
HERE|8886,8890
?|8890,8891
<EOL>|8891,8892
We|8892,8894
did|8895,8898
not|8899,8902
give|8903,8907
you|8908,8911
your|8912,8916
blood|8917,8922
thinner|8923,8930
medication|8931,8941
(|8942,8943
Lovenox|8943,8950
)|8950,8951
,|8951,8952
and|8953,8956
<EOL>|8957,8958
we|8958,8960
gave|8961,8965
you|8966,8969
a|8970,8971
unit|8972,8976
of|8977,8979
blood|8980,8985
.|8985,8986
The|8987,8990
blood|8991,8996
in|8997,8999
your|9000,9004
urine|9005,9010
cleared|9011,9018
up|9019,9021
.|9021,9022
<EOL>|9023,9024
<EOL>|9024,9025
<EOL>|9025,9026
WHAT|9026,9030
SHOULD|9031,9037
YOU|9038,9041
DO|9042,9044
WHEN|9045,9049
YOU|9050,9053
LEAVE|9054,9059
THE|9060,9063
HOSPITAL|9064,9072
?|9072,9073
<EOL>|9073,9074
Along|9074,9079
with|9080,9084
your|9085,9089
oncologist|9090,9100
Dr.|9101,9104
_|9105,9106
_|9106,9107
_|9107,9108
have|9109,9113
decided|9114,9121
that|9122,9126
you|9127,9130
<EOL>|9131,9132
no|9132,9134
longer|9135,9141
need|9142,9146
to|9147,9149
take|9150,9154
any|9155,9158
Lovenox|9159,9166
.|9166,9167
You|9168,9171
should|9172,9178
continue|9179,9187
to|9188,9190
<EOL>|9191,9192
follow|9192,9198
up|9199,9201
with|9202,9206
your|9207,9211
doctors|9212,9219
,|9219,9220
and|9221,9224
take|9225,9229
all|9230,9233
of|9234,9236
your|9237,9241
medications|9242,9253
as|9254,9256
<EOL>|9257,9258
prescribed|9258,9268
.|9268,9269
Your|9270,9274
followup|9275,9283
appointments|9284,9296
are|9297,9300
listed|9301,9307
below|9308,9313
.|9313,9314
<EOL>|9314,9315
<EOL>|9315,9316
Again|9316,9321
,|9321,9322
it|9323,9325
was|9326,9329
a|9330,9331
pleasure|9332,9340
taking|9341,9347
care|9348,9352
of|9353,9355
you|9356,9359
!|9359,9360
<EOL>|9360,9361
<EOL>|9361,9362
Sincerely|9362,9371
,|9371,9372
<EOL>|9373,9374
<EOL>|9374,9375
Your|9375,9379
_|9380,9381
_|9381,9382
_|9382,9383
Team|9384,9388
<EOL>|9388,9389
<EOL>|9390,9391
Followup|9391,9399
Instructions|9400,9412
:|9412,9413
<EOL>|9413,9414
_|9414,9415
_|9415,9416
_|9416,9417
<EOL>|9417,9418

