 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|49,58|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|49,58|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|49,63|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|83,92|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|83,92|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|83,92|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|83,92|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|83,92|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|83,97|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|115,120|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|115,120|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|115,120|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|139,142|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|139,142|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|139,142|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|139,142|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|139,142|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|150,157|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|150,157|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|159,167|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Event|Event|Allergies|188,197|false|false|false|||Attending
Finding|Functional Concept|Allergies|188,197|false|false|false|C1999232|Attending (action)|Attending
Anatomy|Body Location or Region|Chief Complaint|223,232|false|false|false|C0000726|Abdomen|Abdominal
Finding|Sign or Symptom|Chief Complaint|223,237|false|false|false|C0000737|Abdominal Pain|Abdominal pain
Attribute|Clinical Attribute|Chief Complaint|233,237|false|false|false|C2598155||pain
Event|Event|Chief Complaint|233,237|false|false|false|||pain
Finding|Functional Concept|Chief Complaint|233,237|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Chief Complaint|233,237|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Classification|Chief Complaint|241,246|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|247,255|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|247,255|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|259,277|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|268,277|false|false|false|C0945766||Procedure
Event|Event|Chief Complaint|268,277|false|false|false|||Procedure
Event|Occupational Activity|Chief Complaint|268,277|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|268,277|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|268,277|false|false|false|C0184661|Interventional procedure|Procedure
Event|Event|Chief Complaint|279,290|false|false|false|||Colonoscopy
Procedure|Diagnostic Procedure|Chief Complaint|279,290|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|Colonoscopy
Procedure|Health Care Activity|Chief Complaint|279,290|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|Colonoscopy
Procedure|Diagnostic Procedure|Chief Complaint|279,302|false|false|false|C0372088;C0810150|Colonoscopy and Biopsy;Colonoscopy through stoma; with biopsy, single or multiple|Colonoscopy with biopsy
Event|Event|Chief Complaint|296,302|false|false|false|||biopsy
Finding|Finding|Chief Complaint|296,302|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Finding|Intellectual Product|Chief Complaint|296,302|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Procedure|Diagnostic Procedure|Chief Complaint|296,302|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Procedure|Health Care Activity|Chief Complaint|296,302|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Finding|Body Substance|History of Present Illness|343,350|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|343,350|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|343,350|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|360,364|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|History of Present Illness|360,364|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Event|Event|History of Present Illness|365,368|false|false|false|||old
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|387,394|false|false|false|C0227391|Sigmoid colon|sigmoid
Disorder|Disease or Syndrome|History of Present Illness|396,410|false|false|false|C0012813|Diverticulitis|diverticulitis
Event|Event|History of Present Illness|396,410|false|false|false|||diverticulitis
Event|Event|History of Present Illness|415,424|false|false|false|||resection
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|415,424|false|false|false|C0015252;C0728940|Excision;removal technique|resection
Event|Event|History of Present Illness|437,446|false|false|false|||complains
Anatomy|Body Location or Region|History of Present Illness|450,453|false|false|false|C0230178|Structure of right lower quadrant of abdomen|RLQ
Anatomy|Body Location or Region|History of Present Illness|455,464|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|History of Present Illness|455,469|false|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|History of Present Illness|465,469|false|false|false|C2598155||pain
Event|Event|History of Present Illness|465,469|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|465,469|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|465,469|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Body Substance|History of Present Illness|475,482|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|475,482|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|475,482|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|483,489|false|false|false|||states
Attribute|Clinical Attribute|History of Present Illness|499,503|false|false|false|C2598155||pain
Event|Event|History of Present Illness|499,503|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|499,503|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|499,503|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|History of Present Illness|504,509|false|false|false|||began
Event|Event|History of Present Illness|521,530|false|false|false|||afternoon
Event|Event|History of Present Illness|532,540|false|false|false|||worsened
Event|Event|History of Present Illness|555,562|false|false|false|||causing
Event|Event|History of Present Illness|570,577|false|false|false|||present
Finding|Finding|History of Present Illness|570,577|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|History of Present Illness|570,577|false|false|false|C0150312;C0449450|Present;Presentation|present
Event|Event|History of Present Illness|586,588|false|false|false|||ED
Event|Event|History of Present Illness|596,599|false|false|false|||3AM
Event|Event|History of Present Illness|605,614|false|false|false|||describes
Event|Event|History of Present Illness|624,631|false|false|false|||gnawing
Finding|Finding|History of Present Illness|624,631|false|false|false|C1444776|Gnawing sensation quality|gnawing
Attribute|Clinical Attribute|History of Present Illness|633,637|false|false|false|C2598155||pain
Event|Event|History of Present Illness|633,637|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|633,637|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|633,637|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|History of Present Illness|640,652|false|false|false|||nonradiating
Event|Event|History of Present Illness|654,662|false|false|false|||constant
Finding|Intellectual Product|History of Present Illness|654,662|false|false|false|C1720529|Constant - dosing instruction fragment|constant
Event|Event|History of Present Illness|671,680|false|false|false|||intensity
Event|Event|History of Present Illness|686,692|false|false|false|||states
Event|Event|History of Present Illness|699,704|false|false|false|||feels
Event|Event|History of Present Illness|705,712|false|false|false|||similar
Event|Event|History of Present Illness|720,727|false|false|false|||episode
Disorder|Disease or Syndrome|History of Present Illness|731,745|false|false|false|C0012813|Diverticulitis|diverticulitis
Event|Event|History of Present Illness|731,745|false|false|false|||diverticulitis
Finding|Gene or Genome|History of Present Illness|761,764|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Event|Event|History of Present Illness|774,781|false|false|false|||present
Finding|Finding|History of Present Illness|774,781|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|History of Present Illness|774,781|false|false|false|C0150312;C0449450|Present;Presentation|present
Anatomy|Body Location or Region|History of Present Illness|807,814|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|abdomen
Disorder|Neoplastic Process|History of Present Illness|807,814|false|false|false|C0153662|Malignant neoplasm of abdomen|abdomen
Event|Event|History of Present Illness|807,814|false|false|false|||abdomen
Finding|Finding|History of Present Illness|807,814|false|false|false|C0941288|Abdomen problem|abdomen
Event|Event|History of Present Illness|821,827|true|false|false|||denies
Event|Event|History of Present Illness|832,837|true|false|false|||fever
Finding|Finding|History of Present Illness|832,837|true|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|History of Present Illness|832,837|true|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Attribute|Clinical Attribute|History of Present Illness|839,845|true|false|false|C4255480||nausea
Event|Event|History of Present Illness|839,845|true|false|false|||nausea
Finding|Sign or Symptom|History of Present Illness|839,845|true|false|false|C0027497|Nausea|nausea
Event|Event|History of Present Illness|847,855|true|false|false|||vomiting
Finding|Sign or Symptom|History of Present Illness|847,855|true|false|false|C0042963|Vomiting|vomiting
Event|Event|History of Present Illness|857,860|true|false|false|||SOB
Finding|Sign or Symptom|History of Present Illness|857,860|true|false|false|C0013404|Dyspnea|SOB
Anatomy|Body Location or Region|History of Present Illness|862,867|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|History of Present Illness|862,867|false|false|false|C0741025|Chest problem|Chest
Attribute|Clinical Attribute|History of Present Illness|862,872|true|false|false|C2926613||Chest pain
Finding|Sign or Symptom|History of Present Illness|862,872|true|false|false|C0008031|Chest Pain|Chest pain
Attribute|Clinical Attribute|History of Present Illness|868,872|true|false|false|C2598155||pain
Event|Event|History of Present Illness|868,872|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|868,872|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|868,872|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Disorder|Disease or Syndrome|History of Present Illness|874,879|true|false|false|C0018932|Hematochezia|BRBPR
Event|Event|History of Present Illness|874,879|false|false|false|||BRBPR
Attribute|Clinical Attribute|History of Present Illness|899,909|false|false|false|C2979880||subjective
Finding|Finding|History of Present Illness|899,909|false|false|false|C2266644|subjective (symptom)|subjective
Event|Event|History of Present Illness|910,917|false|false|false|||feeling
Finding|Mental Process|History of Present Illness|910,917|false|false|false|C1527305|Feelings|feeling
Event|Event|History of Present Illness|921,927|false|false|false|||chills
Finding|Sign or Symptom|History of Present Illness|921,927|false|false|false|C0085593|Chills|chills
Phenomenon|Natural Phenomenon or Process|History of Present Illness|948,955|false|false|false|C1705970|Electrical Current|current
Finding|Body Substance|History of Present Illness|969,976|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|969,976|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|969,976|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|977,984|false|false|false|||reports
Anatomy|Body Space or Junction|History of Present Illness|996,1001|false|false|false|C0030471;C1305231|Nasal sinus;Sinus - general anatomical term|sinus
Disorder|Anatomical Abnormality|History of Present Illness|996,1001|false|false|false|C0016169|pathologic fistula|sinus
Drug|Organic Chemical|History of Present Illness|996,1001|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Drug|Pharmacologic Substance|History of Present Illness|996,1001|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Disorder|Disease or Syndrome|History of Present Illness|996,1011|false|false|false|C0037199|Sinusitis|sinus infection
Disorder|Disease or Syndrome|History of Present Illness|1002,1011|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|History of Present Illness|1002,1011|false|false|false|||infection
Finding|Pathologic Function|History of Present Illness|1002,1011|false|false|false|C3714514|Infection|infection
Finding|Gene or Genome|History of Present Illness|1027,1030|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Event|Event|History of Present Illness|1036,1044|false|false|false|||resolved
Finding|Intellectual Product|History of Present Illness|1054,1058|false|false|false|C1561540|Transaction counts and value totals - week|week
Finding|Gene or Genome|History of Present Illness|1060,1063|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Finding|Gene or Genome|History of Present Illness|1079,1082|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Event|Event|History of Present Illness|1092,1097|false|false|false|||began
Event|Event|History of Present Illness|1098,1104|false|false|false|||taking
Finding|Finding|History of Present Illness|1107,1110|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|History of Present Illness|1107,1110|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1116,1119|false|false|false|C0228217|Structure of occipital pole|OCP
Disorder|Disease or Syndrome|History of Present Illness|1116,1119|false|false|false|C1282359|Ocular Cicatricial Pemphigoid|OCP
Event|Event|History of Present Illness|1116,1119|false|false|false|||OCP
Event|Activity|History of Present Illness|1124,1129|false|false|false|C1705178|Order (action)|order
Finding|Classification|History of Present Illness|1124,1129|false|false|false|C1546465;C1705175;C1705177;C4284072;C5444833|Medical Order;Order (document);Order (record artifact);Order (taxonomic);What subject filter - Order|order
Finding|Idea or Concept|History of Present Illness|1124,1129|false|false|false|C1546465;C1705175;C1705177;C4284072;C5444833|Medical Order;Order (document);Order (record artifact);Order (taxonomic);What subject filter - Order|order
Finding|Intellectual Product|History of Present Illness|1124,1129|false|false|false|C1546465;C1705175;C1705177;C4284072;C5444833|Medical Order;Order (document);Order (record artifact);Order (taxonomic);What subject filter - Order|order
Phenomenon|Natural Phenomenon or Process|History of Present Illness|1124,1129|false|false|false|C1373200|Order [PK]|order
Event|Event|History of Present Illness|1133,1139|false|false|false|||treate
Finding|Finding|History of Present Illness|1140,1154|false|false|false|C3839366|Perimenopausal state|perimenopausal
Event|Event|History of Present Illness|1155,1163|false|false|false|||cramping
Finding|Sign or Symptom|History of Present Illness|1155,1163|false|false|false|C0026821|Muscle Cramp|cramping
Finding|Functional Concept|History of Present Illness|1172,1178|false|false|false|C1522484;C1561503;C1705190|Precision - second;Second Suffix;metastatic qualifier|second
Finding|Idea or Concept|History of Present Illness|1172,1178|false|false|false|C1522484;C1561503;C1705190|Precision - second;Second Suffix;metastatic qualifier|second
Finding|Intellectual Product|History of Present Illness|1172,1178|false|false|false|C1522484;C1561503;C1705190|Precision - second;Second Suffix;metastatic qualifier|second
Finding|Intellectual Product|History of Present Illness|1179,1183|false|false|false|C1561540|Transaction counts and value totals - week|week
Event|Event|History of Present Illness|1189,1196|false|false|false|||started
Event|Event|History of Present Illness|1205,1213|false|false|false|||spotting
Finding|Functional Concept|History of Present Illness|1205,1213|false|false|false|C0025874;C0312414;C1704255|Menstrual spotting;Metrorrhagia;Spotting|spotting
Finding|Pathologic Function|History of Present Illness|1205,1213|false|false|false|C0025874;C0312414;C1704255|Menstrual spotting;Metrorrhagia;Spotting|spotting
Finding|Sign or Symptom|History of Present Illness|1205,1213|false|false|false|C0025874;C0312414;C1704255|Menstrual spotting;Metrorrhagia;Spotting|spotting
Event|Event|History of Present Illness|1233,1241|false|false|false|||bleeding
Finding|Pathologic Function|History of Present Illness|1233,1241|false|false|false|C0019080|Hemorrhage|bleeding
Finding|Intellectual Product|History of Present Illness|1260,1264|false|false|false|C1561540|Transaction counts and value totals - week|week
Event|Event|History of Present Illness|1277,1284|false|false|false|||episode
Event|Event|History of Present Illness|1288,1296|false|false|false|||diarrhea
Finding|Finding|History of Present Illness|1288,1296|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|History of Present Illness|1288,1296|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Intellectual Product|History of Present Illness|1301,1305|false|false|false|C1561540|Transaction counts and value totals - week|week
Finding|Gene or Genome|History of Present Illness|1306,1309|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Event|Event|History of Present Illness|1334,1343|false|false|false|||nonbloody
Event|Event|History of Present Illness|1348,1356|false|false|false|||resolved
Finding|Finding|History of Present Illness|1364,1367|false|false|false|C5939094|Own|own
Event|Event|History of Present Illness|1400,1407|false|false|false|||feeling
Finding|Mental Process|History of Present Illness|1400,1407|false|false|false|C1527305|Feelings|feeling
Event|Event|History of Present Illness|1412,1427|false|false|false|||lightheadedness
Finding|Sign or Symptom|History of Present Illness|1412,1427|false|false|false|C0220870|Lightheadedness|lightheadedness
Event|Event|History of Present Illness|1430,1440|false|false|false|||associated
Event|Event|History of Present Illness|1446,1457|false|false|false|||diaphoresis
Finding|Finding|History of Present Illness|1446,1457|false|false|false|C0700590|Increased sweating|diaphoresis
Attribute|Clinical Attribute|History of Present Illness|1462,1468|false|false|false|C4255480||nausea
Event|Event|History of Present Illness|1462,1468|false|false|false|||nausea
Finding|Sign or Symptom|History of Present Illness|1462,1468|false|false|false|C0027497|Nausea|nausea
Finding|Idea or Concept|History of Present Illness|1487,1494|false|false|false|C1555582|Initial (abbreviation)|initial
Finding|Body Substance|History of Present Illness|1530,1537|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|1530,1537|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|1530,1537|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|History of Present Illness|1543,1548|false|false|false|||given
Drug|Organic Chemical|History of Present Illness|1549,1557|false|false|false|C0026549|morphine|morphine
Drug|Pharmacologic Substance|History of Present Illness|1549,1557|false|false|false|C0026549|morphine|morphine
Event|Event|History of Present Illness|1549,1557|false|false|false|||morphine
Drug|Organic Chemical|History of Present Illness|1567,1575|false|false|false|C0728755|Dilaudid|dilaudid
Drug|Pharmacologic Substance|History of Present Illness|1567,1575|false|false|false|C0728755|Dilaudid|dilaudid
Event|Event|History of Present Illness|1567,1575|false|false|false|||dilaudid
Drug|Organic Chemical|History of Present Illness|1591,1597|false|false|false|C0206046|Zofran|zofran
Drug|Pharmacologic Substance|History of Present Illness|1591,1597|false|false|false|C0206046|Zofran|zofran
Event|Event|History of Present Illness|1591,1597|false|false|false|||zofran
Finding|Functional Concept|History of Present Illness|1634,1642|true|false|false|C1511117|Bimanual|bimanual
Event|Event|History of Present Illness|1643,1647|true|false|false|||exam
Finding|Functional Concept|History of Present Illness|1643,1647|true|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|History of Present Illness|1643,1647|true|false|false|C0582103|Medical Examination|exam
Event|Event|History of Present Illness|1677,1682|true|false|false|||signs
Finding|Finding|History of Present Illness|1677,1682|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|History of Present Illness|1677,1682|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Event|Event|History of Present Illness|1686,1690|true|false|false|||mass
Finding|Finding|History of Present Illness|1686,1690|true|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|History of Present Illness|1686,1690|true|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|History of Present Illness|1686,1690|true|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Drug|Organic Chemical|History of Present Illness|1692,1695|true|false|false|C1154262|CMT brand of Choline Magnesium Trisalicylate|CMT
Drug|Pharmacologic Substance|History of Present Illness|1692,1695|true|false|false|C1154262|CMT brand of Choline Magnesium Trisalicylate|CMT
Event|Event|History of Present Illness|1692,1695|true|false|false|||CMT
Finding|Sign or Symptom|History of Present Illness|1692,1695|true|false|false|C0238953|CERVICAL MOTION TENDERNESS|CMT
Finding|Finding|History of Present Illness|1700,1718|false|false|false|C0238594|Adnexal tenderness|adnexal tenderness
Event|Event|History of Present Illness|1708,1718|false|false|false|||tenderness
Finding|Mental Process|History of Present Illness|1708,1718|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|History of Present Illness|1708,1718|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Lab|Laboratory or Test Result|History of Present Illness|1720,1724|false|false|false|C0587081|Laboratory test finding|Labs
Event|Event|History of Present Illness|1731,1738|false|false|false|||notable
Disorder|Disease or Syndrome|History of Present Illness|1745,1757|false|false|false|C0023518|Leukocytosis|leukocytosis
Event|Event|History of Present Illness|1745,1757|false|false|false|||leukocytosis
Finding|Finding|History of Present Illness|1745,1757|false|false|false|C0750426|Blood leukocyte number above reference range|leukocytosis
Event|Event|History of Present Illness|1785,1797|false|false|false|||unremarkable
Attribute|Clinical Attribute|History of Present Illness|1799,1809|false|false|false|C1644645||CT abdomen
Procedure|Diagnostic Procedure|History of Present Illness|1799,1809|false|false|false|C0412620|CT of abdomen|CT abdomen
Anatomy|Body Location or Region|History of Present Illness|1802,1809|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|abdomen
Disorder|Neoplastic Process|History of Present Illness|1802,1809|false|false|false|C0153662|Malignant neoplasm of abdomen|abdomen
Event|Event|History of Present Illness|1802,1809|false|false|false|||abdomen
Finding|Finding|History of Present Illness|1802,1809|false|false|false|C0941288|Abdomen problem|abdomen
Event|Event|History of Present Illness|1810,1816|false|false|false|||showed
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1824,1832|false|false|false|C0003617;C4037994|Abdomen+Pelvis>Appendix;Appendix|appendix
Disorder|Neoplastic Process|History of Present Illness|1824,1832|false|false|false|C0348899;C0496779;C0496860|Benign neoplasm of appendix;Malignant neoplasm of appendix;Neoplasm of uncertain or unknown behavior of appendix|appendix
Event|Event|History of Present Illness|1824,1832|false|false|false|||appendix
Finding|Intellectual Product|History of Present Illness|1824,1832|false|false|false|C1552860|appendix - HTML link|appendix
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1824,1832|false|false|false|C0869813|Procedure on appendix|appendix
Finding|Finding|History of Present Illness|1837,1849|false|false|false|C4697736|Thick-walled|thick-walled
Event|Event|History of Present Illness|1843,1849|false|false|false|||walled
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1851,1856|false|false|false|C0007531|Cecum|cecum
Disorder|Neoplastic Process|History of Present Illness|1851,1856|false|false|false|C0153437;C0496859|Benign neoplasm of cecum;Malignant neoplasm of cecum|cecum
Event|Event|History of Present Illness|1851,1856|false|false|false|||cecum
Attribute|Clinical Attribute|History of Present Illness|1862,1872|false|false|false|C0550215||appearance
Event|Event|History of Present Illness|1862,1872|false|false|false|||appearance
Procedure|Health Care Activity|History of Present Illness|1862,1872|false|false|false|C2051406|patient appearance regarding mental status exam|appearance
Finding|Finding|History of Present Illness|1876,1884|false|false|false|C0332149|Possible|possible
Event|Event|History of Present Illness|1885,1889|false|false|false|||mass
Finding|Finding|History of Present Illness|1885,1889|false|true|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|History of Present Illness|1885,1889|false|true|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|History of Present Illness|1885,1889|false|true|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1891,1897|true|false|false|C0030797|Pelvis|Pelvic
Procedure|Diagnostic Procedure|History of Present Illness|1891,1908|true|false|false|C0948766|Ultrasound pelvis|Pelvic ultrasound
Event|Event|History of Present Illness|1898,1908|true|false|false|||ultrasound
Finding|Functional Concept|History of Present Illness|1898,1908|true|false|false|C0220934|Ultrasonic|ultrasound
Phenomenon|Natural Phenomenon or Process|History of Present Illness|1898,1908|true|false|false|C0041621;C1456803|Ultrasonic Shockwave;Ultrasonics (sound)|ultrasound
Procedure|Diagnostic Procedure|History of Present Illness|1898,1908|true|false|false|C0041618;C1315081|Ultrasonography;Urological ultrasound|ultrasound
Event|Event|History of Present Illness|1918,1922|true|false|false|||show
Event|Event|History of Present Illness|1927,1933|true|false|false|||source
Finding|Finding|History of Present Illness|1927,1933|true|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Finding|Functional Concept|History of Present Illness|1927,1933|true|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Finding|Intellectual Product|History of Present Illness|1927,1933|true|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Attribute|Clinical Attribute|History of Present Illness|1941,1945|true|false|false|C2598155||pain
Event|Event|History of Present Illness|1941,1945|true|false|false|||pain
Finding|Functional Concept|History of Present Illness|1941,1945|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1941,1945|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|History of Present Illness|1977,1983|true|false|false|C0723011|Relief brand of phenylephrine|relief
Drug|Pharmacologic Substance|History of Present Illness|1977,1983|true|false|false|C0723011|Relief brand of phenylephrine|relief
Event|Event|History of Present Illness|1977,1983|true|false|false|||relief
Finding|Finding|History of Present Illness|1977,1983|true|false|false|C0564405|Feeling relief|relief
Attribute|Clinical Attribute|History of Present Illness|1989,1993|true|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|1989,1993|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1989,1993|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|History of Present Illness|1994,2005|true|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|History of Present Illness|1994,2005|true|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|History of Present Illness|1994,2005|true|false|false|||medications
Finding|Intellectual Product|History of Present Illness|1994,2005|true|false|false|C4284232|Medications|medications
Event|Event|History of Present Illness|2015,2023|false|false|false|||admitted
Event|Event|History of Present Illness|2031,2038|false|false|false|||medical
Finding|Functional Concept|History of Present Illness|2031,2038|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Idea or Concept|History of Present Illness|2031,2038|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Intellectual Product|History of Present Illness|2031,2038|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Procedure|Health Care Activity|History of Present Illness|2031,2038|false|false|false|C0199168|Medical service|medical
Event|Event|History of Present Illness|2040,2047|false|false|false|||service
Event|Occupational Activity|History of Present Illness|2040,2047|false|false|false|C0557854|Services|service
Finding|Idea or Concept|History of Present Illness|2040,2047|false|false|false|C3245478|ActInformationPrivacyReason - service|service
Attribute|Clinical Attribute|History of Present Illness|2052,2056|false|false|false|C2598155||pain
Event|Event|History of Present Illness|2052,2056|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|2052,2056|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|2052,2056|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|History of Present Illness|2052,2064|false|false|false|C5548091|Demonstrates adequate pain control|pain control
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|2052,2064|false|false|false|C0002766;C1304888|Pain control;Pain management (procedure)|pain control
Drug|Organic Chemical|History of Present Illness|2057,2064|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Pharmacologic Substance|History of Present Illness|2057,2064|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Substance|History of Present Illness|2057,2064|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Event|Event|History of Present Illness|2057,2064|false|false|false|||control
Finding|Conceptual Entity|History of Present Illness|2057,2064|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Functional Concept|History of Present Illness|2057,2064|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Idea or Concept|History of Present Illness|2057,2064|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Event|Event|History of Present Illness|2072,2078|false|false|false|||Vitals
Event|Event|History of Present Illness|2082,2090|false|false|false|||transfer
Finding|Functional Concept|History of Present Illness|2082,2090|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|History of Present Illness|2082,2090|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|History of Present Illness|2082,2090|false|false|false|C4706767|Transfer (immobility management)|transfer
Anatomy|Anatomical Structure|History of Present Illness|2133,2138|false|false|false|C3714591|Floor (anatomic)|floor
Finding|Body Substance|History of Present Illness|2140,2147|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|2140,2147|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|2140,2147|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|2148,2156|false|false|false|||reported
Event|Event|History of Present Illness|2157,2166|false|false|false|||continued
Attribute|Clinical Attribute|History of Present Illness|2171,2175|false|false|false|C2598155||pain
Event|Event|History of Present Illness|2171,2175|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|2171,2175|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|2171,2175|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Anatomy|Body Location or Region|History of Present Illness|2183,2186|false|false|false|C0230178|Structure of right lower quadrant of abdomen|RLQ
Finding|Intellectual Product|History of Present Illness|2205,2209|false|false|false|C1547225|Mild Severity of Illness Code|mild
Attribute|Clinical Attribute|History of Present Illness|2210,2216|false|false|false|C4255480||nausea
Event|Event|History of Present Illness|2210,2216|false|false|false|||nausea
Finding|Sign or Symptom|History of Present Illness|2210,2216|false|false|false|C0027497|Nausea|nausea
Event|Event|History of Present Illness|2224,2230|false|false|false|||Review
Finding|Idea or Concept|History of Present Illness|2224,2230|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|Review
Finding|Intellectual Product|History of Present Illness|2224,2230|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|Review
Finding|Functional Concept|History of Present Illness|2224,2233|false|false|false|C0699752|Review of|Review of
Attribute|Clinical Attribute|History of Present Illness|2224,2241|false|false|false|C0488564;C0488565||Review of systems
Procedure|Health Care Activity|History of Present Illness|2224,2241|false|false|false|C0489633|Review of systems (procedure)|Review of systems
Event|Event|History of Present Illness|2234,2241|false|false|false|||systems
Finding|Functional Concept|History of Present Illness|2234,2241|false|false|false|C0449913|System|systems
Disorder|Disease or Syndrome|History of Present Illness|2253,2256|false|false|false|C0268529|Proline dehydrogenase deficiency|HPI
Event|Event|History of Present Illness|2253,2256|false|false|false|||HPI
Finding|Finding|History of Present Illness|2253,2256|false|false|false|C0262512;C1323983|History of present illness (finding);allene oxide synthase activity|HPI
Finding|Molecular Function|History of Present Illness|2253,2256|false|false|false|C0262512;C1323983|History of present illness (finding);allene oxide synthase activity|HPI
Event|Event|History of Present Illness|2263,2269|false|false|false|||Denies
Event|Event|History of Present Illness|2270,2275|true|false|false|||fever
Finding|Finding|History of Present Illness|2270,2275|true|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|History of Present Illness|2270,2275|true|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Event|Event|History of Present Illness|2277,2283|true|false|false|||chills
Finding|Sign or Symptom|History of Present Illness|2277,2283|true|false|false|C0085593|Chills|chills
Finding|Sign or Symptom|History of Present Illness|2285,2297|true|false|false|C0028081|Night sweats|night sweats
Event|Event|History of Present Illness|2291,2297|true|false|false|||sweats
Finding|Body Substance|History of Present Illness|2291,2297|true|false|false|C0038984;C0038990|Sweat;Sweating|sweats
Finding|Finding|History of Present Illness|2291,2297|true|false|false|C0038984;C0038990|Sweat;Sweating|sweats
Attribute|Clinical Attribute|History of Present Illness|2306,2312|false|false|false|C0944911||weight
Event|Event|History of Present Illness|2306,2312|false|false|false|||weight
Finding|Finding|History of Present Illness|2306,2312|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|History of Present Illness|2306,2312|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|History of Present Illness|2306,2312|false|false|false|C1305866|Weighing patient|weight
Finding|Finding|History of Present Illness|2306,2317|true|false|false|C1262477;C3540682|Losing Weight (question);Weight Loss|weight loss
Finding|Intellectual Product|History of Present Illness|2306,2317|true|false|false|C1262477;C3540682|Losing Weight (question);Weight Loss|weight loss
Event|Event|History of Present Illness|2313,2317|false|false|false|||loss
Finding|Finding|History of Present Illness|2313,2317|true|false|false|C5890125|Loss (adaptation)|loss
Event|Event|History of Present Illness|2322,2326|false|false|false|||gain
Event|Event|History of Present Illness|2328,2334|false|false|false|||Denies
Event|Event|History of Present Illness|2335,2343|true|false|false|||headache
Finding|Sign or Symptom|History of Present Illness|2335,2343|true|false|false|C0018681|Headache|headache
Anatomy|Body Space or Junction|History of Present Illness|2345,2350|true|false|false|C0030471;C1305231|Nasal sinus;Sinus - general anatomical term|sinus
Disorder|Anatomical Abnormality|History of Present Illness|2345,2350|true|false|false|C0016169|pathologic fistula|sinus
Drug|Organic Chemical|History of Present Illness|2345,2350|true|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Drug|Pharmacologic Substance|History of Present Illness|2345,2350|true|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Event|Event|History of Present Illness|2351,2361|true|false|false|||tenderness
Finding|Mental Process|History of Present Illness|2351,2361|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|History of Present Illness|2351,2361|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Event|Event|History of Present Illness|2363,2373|true|false|false|||rhinorrhea
Finding|Sign or Symptom|History of Present Illness|2363,2373|true|false|false|C1260880|Rhinorrhea|rhinorrhea
Event|Event|History of Present Illness|2378,2388|false|false|false|||congestion
Finding|Pathologic Function|History of Present Illness|2378,2388|false|false|false|C0700148|Congestion|congestion
Drug|Organic Chemical|History of Present Illness|2397,2402|true|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|History of Present Illness|2397,2402|true|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|History of Present Illness|2397,2402|true|false|false|||cough
Finding|Sign or Symptom|History of Present Illness|2397,2402|true|false|false|C0010200|Coughing|cough
Event|Event|History of Present Illness|2404,2413|true|false|false|||shortness
Attribute|Clinical Attribute|History of Present Illness|2404,2423|true|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|History of Present Illness|2404,2423|true|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|History of Present Illness|2417,2423|true|false|false|C0225386|Breath|breath
Event|Event|History of Present Illness|2425,2431|false|false|false|||Denied
Anatomy|Body Location or Region|History of Present Illness|2432,2437|true|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|2432,2437|true|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|History of Present Illness|2432,2442|true|false|false|C2926613||chest pain
Finding|Sign or Symptom|History of Present Illness|2432,2442|true|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|History of Present Illness|2438,2442|true|true|false|C2598155||pain
Event|Event|History of Present Illness|2438,2442|true|false|false|||pain
Finding|Functional Concept|History of Present Illness|2438,2442|true|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|2438,2442|true|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|History of Present Illness|2447,2456|true|false|false|||tightness
Event|Event|History of Present Illness|2458,2470|true|false|false|||palpitations
Finding|Finding|History of Present Illness|2458,2470|true|false|false|C0030252|Palpitations|palpitations
Event|Event|History of Present Illness|2479,2487|true|false|false|||vomiting
Finding|Sign or Symptom|History of Present Illness|2479,2487|true|false|false|C0042963|Vomiting|vomiting
Event|Event|History of Present Illness|2489,2497|true|false|false|||diarrhea
Finding|Finding|History of Present Illness|2489,2497|true|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|History of Present Illness|2489,2497|true|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Event|Event|History of Present Illness|2500,2512|true|false|false|||constipation
Finding|Sign or Symptom|History of Present Illness|2500,2512|true|false|false|C0009806|Constipation|constipation
Disorder|Disease or Syndrome|History of Present Illness|2516,2521|false|false|false|C0018932|Hematochezia|BRBPR
Event|Event|History of Present Illness|2516,2521|false|false|false|||BRBPR
Event|Event|History of Present Illness|2526,2533|true|false|false|||dysuria
Finding|Sign or Symptom|History of Present Illness|2526,2533|true|false|false|C0013428|Dysuria|dysuria
Event|Event|History of Present Illness|2542,2553|true|false|false|||arthralgias
Finding|Sign or Symptom|History of Present Illness|2542,2553|true|false|false|C0003862|Arthralgia|arthralgias
Event|Event|History of Present Illness|2558,2566|true|false|false|||myalgias
Finding|Sign or Symptom|History of Present Illness|2558,2566|true|false|false|C0231528|Myalgia|myalgias
Disorder|Disease or Syndrome|Past Medical History|2598,2612|false|false|false|C0012813|Diverticulitis|diverticulitis
Event|Event|Past Medical History|2598,2612|false|false|false|||diverticulitis
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2617,2624|false|false|false|C0227391|Sigmoid colon|sigmoid
Event|Event|Past Medical History|2625,2634|false|false|false|||resection
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2625,2634|false|false|false|C0015252;C0728940|Excision;removal technique|resection
Disorder|Mental or Behavioral Dysfunction|Past Medical History|2641,2648|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|Anxiety
Event|Event|Past Medical History|2641,2648|false|false|false|||Anxiety
Finding|Sign or Symptom|Past Medical History|2641,2648|false|false|false|C0860603|Anxiety symptoms|Anxiety
Finding|Functional Concept|Past Medical History|2651,2659|false|false|false|C0700624|Allergic|Allergic
Disorder|Disease or Syndrome|Past Medical History|2651,2668|false|false|false|C2607914|Allergic rhinitis (disorder)|Allergic rhinitis
Finding|Gene or Genome|Past Medical History|2651,2668|false|false|false|C1334103|IL13 gene|Allergic rhinitis
Disorder|Disease or Syndrome|Past Medical History|2660,2668|false|false|false|C0035455|Rhinitis|rhinitis
Event|Event|Past Medical History|2660,2668|false|false|false|||rhinitis
Disorder|Disease or Syndrome|Past Medical History|2671,2675|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Event|Event|Past Medical History|2671,2675|false|false|false|||GERD
Disorder|Disease or Syndrome|Past Medical History|2678,2684|false|false|false|C0013595|Eczema|Eczema
Event|Event|Past Medical History|2678,2684|false|false|false|||Eczema
Disorder|Disease or Syndrome|Past Medical History|2687,2695|false|false|false|C0149931|Migraine Disorders|Migraine
Disorder|Disease or Syndrome|Past Medical History|2687,2705|false|false|false|C0149931|Migraine Disorders|Migraine headaches
Event|Event|Past Medical History|2696,2705|false|false|false|||headaches
Finding|Sign or Symptom|Past Medical History|2696,2705|false|false|false|C0018681|Headache|headaches
Finding|Functional Concept|Past Medical History|2718,2722|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|tube
Finding|Gene or Genome|Past Medical History|2718,2722|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|tube
Disorder|Disease or Syndrome|Past Medical History|2723,2734|false|false|false|C3887505|DYSFUNCTION - SKIN DISORDERS|dysfunction
Event|Event|Past Medical History|2723,2734|false|false|false|||dysfunction
Finding|Conceptual Entity|Past Medical History|2723,2734|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Functional Concept|Past Medical History|2723,2734|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Pathologic Function|Past Medical History|2723,2734|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Event|Event|Family Medical History|2776,2782|false|false|false|||Father
Finding|Conceptual Entity|Family Medical History|2776,2782|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Idea or Concept|Family Medical History|2776,2782|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Disorder|Disease or Syndrome|Family Medical History|2794,2801|false|false|false|C0009319|Colitis|colitis
Event|Event|Family Medical History|2794,2801|false|false|false|||colitis
Anatomy|Body Location or Region|Family Medical History|2810,2814|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2810,2814|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Family Medical History|2810,2814|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Family Medical History|2810,2814|false|false|false|C0740941|Lung Problem|lung
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2829,2835|false|false|false|C0006141|Breast|breast
Disorder|Neoplastic Process|Family Medical History|2829,2835|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|breast
Event|Event|Family Medical History|2829,2835|false|false|false|||breast
Finding|Finding|Family Medical History|2829,2835|false|false|false|C0567499|Breast problem|breast
Procedure|Therapeutic or Preventive Procedure|Family Medical History|2829,2835|false|false|false|C0191838|Procedures on breast|breast
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2859,2866|false|false|false|C0038351;C3714551;C4266636|Abdomen>Stomach;Stomach;Stomach structure|stomach
Disorder|Disease or Syndrome|Family Medical History|2859,2866|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Disorder|Neoplastic Process|Family Medical History|2859,2866|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Finding|Finding|Family Medical History|2859,2866|false|false|false|C0577027|Stomach problem|stomach
Procedure|Therapeutic or Preventive Procedure|Family Medical History|2859,2866|false|false|false|C0872393|Procedure on stomach|stomach
Disorder|Neoplastic Process|Family Medical History|2859,2869|false|false|false|C0024623|Malignant neoplasm of stomach|stomach Ca
Event|Event|Family Medical History|2867,2869|false|false|false|||Ca
Event|Event|Family Medical History|2871,2877|false|false|false|||Mother
Finding|Idea or Concept|Family Medical History|2871,2877|false|false|false|C1546508|Relationship - Mother|Mother
Anatomy|Body Space or Junction|Family Medical History|2883,2886|false|false|false|C0262212|Choroidal fissure|CHF
Disorder|Disease or Syndrome|Family Medical History|2883,2886|false|false|false|C0018802|Congestive heart failure|CHF
Disorder|Disease or Syndrome|Family Medical History|2891,2894|false|false|false|C2931689|Dystrophia myotonica 2|DM2
Event|Event|Family Medical History|2891,2894|false|false|false|||DM2
Finding|Gene or Genome|Family Medical History|2891,2894|false|false|false|C1415938;C1824763;C3273677|CNBP gene;CNBP wt Allele;IGHD1-14 gene|DM2
Event|Event|General Exam|2966,2973|false|false|false|||General
Finding|Classification|General Exam|2966,2973|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|General Exam|2966,2973|false|false|false|C3812897|General medical service|General
Attribute|Clinical Attribute|General Exam|2975,2980|true|false|false|C5890168||Alert
Drug|Organic Chemical|General Exam|2975,2980|true|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|General Exam|2975,2980|true|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|General Exam|2975,2980|true|false|false|||Alert
Finding|Finding|General Exam|2975,2980|true|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|General Exam|2975,2980|true|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|General Exam|2975,2980|true|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|General Exam|2982,2990|true|false|false|||oriented
Finding|Intellectual Product|General Exam|2995,3000|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|General Exam|3001,3009|true|false|false|||distress
Finding|Finding|General Exam|3001,3009|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|General Exam|3001,3009|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Anatomy|Body Location or Region|General Exam|3012,3017|true|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|General Exam|3019,3025|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|General Exam|3019,3025|false|false|false|C0036412|Scleral Diseases|Sclera
Event|Event|General Exam|3019,3025|false|false|false|||Sclera
Procedure|Health Care Activity|General Exam|3019,3025|false|false|false|C2228481|examination of sclera|Sclera
Event|Event|General Exam|3026,3035|false|false|false|||anicteric
Finding|Finding|General Exam|3026,3035|false|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Part, Organ, or Organ Component|General Exam|3037,3040|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|General Exam|3037,3040|false|false|false|C0026987|Myelofibrosis|MMM
Anatomy|Body Location or Region|General Exam|3042,3052|false|false|false|C0521367|Oropharyngeal|oropharynx
Event|Event|General Exam|3053,3058|false|false|false|||clear
Finding|Idea or Concept|General Exam|3053,3058|false|false|false|C1550016|Remote control command - Clear|clear
Anatomy|Body Location or Region|General Exam|3061,3065|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Anatomy|Cell Component|General Exam|3061,3065|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Finding|Finding|General Exam|3061,3065|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|Neck
Event|Event|General Exam|3067,3073|true|false|false|||supple
Finding|Functional Concept|General Exam|3067,3073|true|false|false|C0332254|Supple|supple
Event|Event|General Exam|3075,3078|true|false|false|||JVP
Finding|Finding|General Exam|3075,3078|true|false|false|C0428897|Jugular venous pressure|JVP
Event|Event|General Exam|3083,3091|true|false|false|||elevated
Anatomy|Body Part, Organ, or Organ Component|General Exam|3096,3099|true|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|General Exam|3096,3099|true|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|General Exam|3096,3099|true|false|false|||LAD
Finding|Gene or Genome|General Exam|3096,3099|true|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Anatomy|Body Part, Organ, or Organ Component|General Exam|3102,3107|true|false|false|C0024109|Lung|Lungs
Event|Event|General Exam|3109,3114|true|false|false|||Clear
Finding|Idea or Concept|General Exam|3109,3114|true|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|General Exam|3118,3130|true|false|false|||auscultation
Procedure|Diagnostic Procedure|General Exam|3118,3130|true|false|false|C0004339|Auscultation|auscultation
Event|Event|General Exam|3147,3154|true|false|false|||wheezes
Finding|Sign or Symptom|General Exam|3147,3154|true|false|false|C0043144|Wheezing|wheezes
Event|Event|General Exam|3156,3161|true|false|false|||rales
Finding|Finding|General Exam|3156,3161|true|false|false|C0034642;C0240859|Basilar Rales;Rales|rales
Event|Event|General Exam|3164,3171|true|false|false|||rhonchi
Finding|Finding|General Exam|3164,3171|true|false|false|C0035508|Rhonchi|rhonchi
Event|Activity|General Exam|3186,3190|false|false|false|C0871208|Rating (action)|rate
Event|Event|General Exam|3186,3190|false|false|false|||rate
Finding|Idea or Concept|General Exam|3186,3190|false|false|false|C1549480|Amount type - Rate|rate
Event|Event|General Exam|3195,3201|true|false|false|||rhythm
Finding|Finding|General Exam|3195,3201|true|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|General Exam|3195,3201|true|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Event|Event|General Exam|3222,3229|true|false|false|||murmurs
Finding|Finding|General Exam|3222,3229|true|false|false|C0018808|Heart murmur|murmurs
Event|Event|General Exam|3231,3235|true|false|false|||rubs
Finding|Finding|General Exam|3231,3235|true|false|false|C0232267|Pericardial friction rub|rubs
Event|Event|General Exam|3238,3245|true|false|false|||gallops
Anatomy|Body Location or Region|General Exam|3248,3255|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|General Exam|3248,3255|false|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Event|Event|General Exam|3248,3255|false|false|false|||Abdomen
Finding|Finding|General Exam|3248,3255|false|false|false|C0941288|Abdomen problem|Abdomen
Disorder|Disease or Syndrome|General Exam|3257,3261|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|General Exam|3257,3261|false|false|false|||soft
Anatomy|Body Part, Organ, or Organ Component|General Exam|3278,3283|false|false|false|C0021853|Intestines|bowel
Finding|Finding|General Exam|3278,3290|false|false|false|C0232693|Bowel sounds|bowel sounds
Event|Event|General Exam|3284,3290|false|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|General Exam|3284,3290|false|false|false|C0037709||sounds
Finding|Finding|General Exam|3291,3298|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|General Exam|3291,3298|false|false|false|C0150312;C0449450|Present;Presentation|present
Disorder|Disease or Syndrome|General Exam|3300,3303|false|false|false|C0034155;C1268935|Congenital Thrombotic Thrombocytopenic Purpura;Purpura, Thrombotic Thrombocytopenic|TTP
Drug|Amino Acid, Peptide, or Protein|General Exam|3300,3303|false|false|false|C1506603;C4723973|ZFP36 protein, human;thiamine triphosphorate|TTP
Drug|Biologically Active Substance|General Exam|3300,3303|false|false|false|C1506603;C4723973|ZFP36 protein, human;thiamine triphosphorate|TTP
Drug|Organic Chemical|General Exam|3300,3303|false|false|false|C1506603;C4723973|ZFP36 protein, human;thiamine triphosphorate|TTP
Drug|Vitamin|General Exam|3300,3303|false|false|false|C1506603;C4723973|ZFP36 protein, human;thiamine triphosphorate|TTP
Event|Event|General Exam|3300,3303|false|false|false|||TTP
Finding|Gene or Genome|General Exam|3300,3303|false|false|false|C1413036;C1421571;C3539814|ADAMTS13 gene;ZFP36 gene;ZFP36 wt Allele|TTP
Anatomy|Body Location or Region|General Exam|3307,3310|true|false|false|C0230178|Structure of right lower quadrant of abdomen|RLQ
Attribute|Clinical Attribute|General Exam|3317,3321|true|false|false|C4318566|Deep Resection Margin|deep
Procedure|Diagnostic Procedure|General Exam|3317,3331|true|false|false|C0278328|Deep palpation|deep palpation
Event|Event|General Exam|3322,3331|true|false|false|||palpation
Procedure|Diagnostic Procedure|General Exam|3322,3331|true|false|false|C0030247|Palpation|palpation
Finding|Sign or Symptom|General Exam|3341,3359|true|false|false|C0234246|Rebound tenderness|rebound tenderness
Event|Event|General Exam|3349,3359|true|false|false|||tenderness
Finding|Mental Process|General Exam|3349,3359|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|General Exam|3349,3359|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Event|Event|General Exam|3363,3371|true|false|false|||guarding
Finding|Finding|General Exam|3363,3371|true|false|false|C0427198|Protective muscle spasm|guarding
Event|Event|General Exam|3373,3375|true|false|false|||no
Event|Event|General Exam|3377,3389|true|false|false|||organomegaly
Finding|Finding|General Exam|3377,3389|true|false|false|C4054315|Organomegaly|organomegaly
Disorder|Congenital Abnormality|General Exam|3392,3395|true|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Event|Event|General Exam|3392,3395|true|false|false|||Ext
Finding|Gene or Genome|General Exam|3392,3395|true|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Event|Event|General Exam|3397,3401|false|false|false|||Warm
Finding|Finding|General Exam|3397,3401|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|General Exam|3397,3401|false|false|false|C0687712|warming process|Warm
Finding|Finding|General Exam|3403,3407|true|false|false|C5575035|Well (answer to question)|well
Event|Event|General Exam|3408,3416|true|false|false|||perfused
Drug|Food|General Exam|3421,3427|true|false|false|C5890763||pulses
Event|Event|General Exam|3421,3427|true|false|false|||pulses
Finding|Physiologic Function|General Exam|3421,3427|true|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|General Exam|3421,3427|true|false|false|C0034107|Pulse taking|pulses
Disorder|Anatomical Abnormality|General Exam|3432,3440|true|false|false|C0149651|Clubbing|clubbing
Event|Event|General Exam|3432,3440|true|false|false|||clubbing
Event|Event|General Exam|3442,3450|true|false|false|||cyanosis
Finding|Sign or Symptom|General Exam|3442,3450|true|false|false|C0010520|Cyanosis|cyanosis
Attribute|Clinical Attribute|General Exam|3455,3460|true|false|false|C1717255||edema
Event|Event|General Exam|3455,3460|true|false|false|||edema
Finding|Pathologic Function|General Exam|3455,3460|true|false|false|C0013604|Edema|edema
Attribute|Clinical Attribute|General Exam|3485,3495|false|false|false|C2598148||Laboratory
Finding|Functional Concept|General Exam|3485,3495|false|false|false|C1548427;C1571737;C3244292|Diagnostic Service Section ID - Laboratory;Laboratory domain;Referral type - Laboratory|Laboratory
Finding|Intellectual Product|General Exam|3485,3495|false|false|false|C1548427;C1571737;C3244292|Diagnostic Service Section ID - Laboratory;Laboratory domain;Referral type - Laboratory|Laboratory
Lab|Laboratory or Test Result|General Exam|3485,3495|false|false|false|C4283904|Laboratory observation|Laboratory
Lab|Laboratory or Test Result|General Exam|3485,3504|false|false|false|C0587081|Laboratory test finding|Laboratory Findings
Attribute|Clinical Attribute|General Exam|3496,3504|false|false|false|C2926606||Findings
Event|Event|General Exam|3496,3504|false|false|false|||Findings
Finding|Functional Concept|General Exam|3496,3504|false|false|false|C2607943|findings aspects|Findings
Disorder|Disease or Syndrome|General Exam|3518,3523|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3518,3523|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3518,3523|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|3524,3527|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|3534,3537|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|3534,3537|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|3534,3537|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|3544,3547|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|3544,3547|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|3544,3547|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|3544,3547|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|3553,3556|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|3553,3556|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|3564,3567|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|3564,3567|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|3564,3567|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|3564,3567|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|3564,3567|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|3571,3574|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|3571,3574|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|3571,3574|false|false|false|||MCH
Finding|Gene or Genome|General Exam|3571,3574|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|3571,3574|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|3571,3574|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|General Exam|3580,3584|false|false|false|||MCHC
Procedure|Laboratory Procedure|General Exam|3580,3584|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|3599,3602|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|3619,3624|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3619,3624|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3619,3624|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Antibiotic|General Exam|3641,3646|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|General Exam|3641,3646|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|General Exam|3641,3646|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|General Exam|3651,3654|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|Eos
Event|Event|General Exam|3651,3654|false|false|false|||Eos
Finding|Gene or Genome|General Exam|3651,3654|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|Eos
Disorder|Disease or Syndrome|General Exam|3681,3686|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3681,3686|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3681,3686|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|General Exam|3703,3708|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3703,3708|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3703,3708|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|3703,3716|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|3703,3716|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|3703,3716|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|3709,3716|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|3709,3716|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|3709,3716|false|false|false|C0017725|glucose|Glucose
Event|Event|General Exam|3709,3716|false|false|false|||Glucose
Lab|Laboratory or Test Result|General Exam|3709,3716|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|3709,3716|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|General Exam|3762,3766|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|3762,3766|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|General Exam|3762,3766|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|General Exam|3791,3796|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3791,3796|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3791,3796|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|3797,3800|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|General Exam|3797,3800|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|General Exam|3797,3800|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|General Exam|3797,3800|false|false|false|||ALT
Finding|Gene or Genome|General Exam|3797,3800|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|General Exam|3797,3800|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|General Exam|3797,3800|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|General Exam|3797,3800|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|General Exam|3804,3807|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|General Exam|3804,3807|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|3804,3807|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|General Exam|3804,3807|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|General Exam|3804,3807|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|General Exam|3804,3807|false|false|false|||AST
Finding|Gene or Genome|General Exam|3804,3807|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|3811,3818|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|General Exam|3811,3818|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Disorder|Disease or Syndrome|General Exam|3846,3851|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3846,3851|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3846,3851|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|3852,3858|false|false|false|C0023764|lipase|Lipase
Drug|Enzyme|General Exam|3852,3858|false|false|false|C0023764|lipase|Lipase
Drug|Pharmacologic Substance|General Exam|3852,3858|false|false|false|C0023764|lipase|Lipase
Procedure|Laboratory Procedure|General Exam|3852,3858|false|false|false|C0373670|Lipase measurement|Lipase
Disorder|Disease or Syndrome|General Exam|3874,3879|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3874,3879|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3874,3879|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|3874,3887|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|General Exam|3880,3887|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|General Exam|3880,3887|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|General Exam|3880,3887|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|General Exam|3880,3887|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|General Exam|3880,3887|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|General Exam|3880,3887|false|false|false|||Calcium
Finding|Physiologic Function|General Exam|3880,3887|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|General Exam|3880,3887|false|false|false|C0201925|Calcium measurement|Calcium
Disorder|Disease or Syndrome|General Exam|3923,3928|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3923,3928|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3923,3928|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|3923,3936|false|false|false|C3824990|lactate in blood (lab test)|BLOOD Lactate
Drug|Organic Chemical|General Exam|3929,3936|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Drug|Pharmacologic Substance|General Exam|3929,3936|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Event|Event|General Exam|3929,3936|false|false|false|||Lactate
Procedure|Laboratory Procedure|General Exam|3929,3936|false|false|false|C0202115|Lactic acid measurement|Lactate
Disorder|Disease or Syndrome|General Exam|3953,3958|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3953,3958|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3953,3958|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|3959,3962|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|3967,3970|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|3967,3970|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|3967,3970|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|3977,3980|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|3977,3980|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|3977,3980|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|3977,3980|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|3987,3990|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|3987,3990|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|3998,4001|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|3998,4001|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|3998,4001|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|3998,4001|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|3998,4001|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|4005,4008|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|4005,4008|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|4005,4008|false|false|false|||MCH
Finding|Gene or Genome|General Exam|4005,4008|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|4005,4008|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|4005,4008|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|General Exam|4014,4018|false|false|false|||MCHC
Procedure|Laboratory Procedure|General Exam|4014,4018|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|4033,4036|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|4053,4058|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4053,4058|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4053,4058|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|4053,4066|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|4053,4066|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|4053,4066|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|4059,4066|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|4059,4066|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|4059,4066|false|false|false|C0017725|glucose|Glucose
Event|Event|General Exam|4059,4066|false|false|false|||Glucose
Lab|Laboratory or Test Result|General Exam|4059,4066|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|4059,4066|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|General Exam|4110,4114|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|4110,4114|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|General Exam|4110,4114|false|false|false|C0202059|Bicarbonate measurement|HCO3
Finding|Body Substance|General Exam|4139,4144|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|4139,4144|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|4139,4144|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Finding|General Exam|4139,4150|false|false|false|C0278030|Color of urine|URINE Color
Drug|Biomedical or Dental Material|General Exam|4145,4150|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|Color
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|4145,4150|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|Color
Event|Event|General Exam|4145,4150|false|false|false|||Color
Drug|Organic Chemical|General Exam|4151,4156|false|false|false|C4047917|Cereal plant straw|Straw
Finding|Idea or Concept|General Exam|4164,4169|false|false|false|C1550016|Remote control command - Clear|Clear
Finding|Body Substance|General Exam|4189,4194|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|4189,4194|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|4189,4194|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Disorder|Disease or Syndrome|General Exam|4189,4200|false|false|false|C0018965|Hematuria|URINE Blood
Disorder|Disease or Syndrome|General Exam|4195,4200|false|false|false|C0851353|Blood and lymphatic system disorders|Blood
Event|Event|General Exam|4195,4200|false|false|false|||Blood
Finding|Body Substance|General Exam|4195,4200|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Drug|Biologically Active Substance|General Exam|4204,4211|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|Nitrite
Drug|Inorganic Chemical|General Exam|4204,4211|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|Nitrite
Drug|Pharmacologic Substance|General Exam|4204,4211|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|Nitrite
Event|Event|General Exam|4212,4215|false|false|false|||NEG
Finding|Finding|General Exam|4212,4215|false|false|false|C5848551|Neg - answer|NEG
Drug|Amino Acid, Peptide, or Protein|General Exam|4216,4223|false|false|false|C0033684|Proteins|Protein
Drug|Biologically Active Substance|General Exam|4216,4223|false|false|false|C0033684|Proteins|Protein
Event|Event|General Exam|4216,4223|false|false|false|||Protein
Finding|Conceptual Entity|General Exam|4216,4223|false|false|false|C1521746|Protein Info|Protein
Procedure|Laboratory Procedure|General Exam|4216,4223|false|false|false|C0202202|Protein measurement|Protein
Event|Event|General Exam|4224,4227|false|false|false|||NEG
Finding|Finding|General Exam|4224,4227|false|false|false|C5848551|Neg - answer|NEG
Drug|Biologically Active Substance|General Exam|4229,4236|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|4229,4236|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|4229,4236|false|false|false|C0017725|glucose|Glucose
Event|Event|General Exam|4229,4236|false|false|false|||Glucose
Lab|Laboratory or Test Result|General Exam|4229,4236|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|4229,4236|false|false|false|C0337438|Glucose measurement|Glucose
Event|Event|General Exam|4237,4240|false|false|false|||NEG
Finding|Finding|General Exam|4237,4240|false|false|false|C5848551|Neg - answer|NEG
Drug|Organic Chemical|General Exam|4241,4247|false|false|false|C0022634|Ketones|Ketone
Event|Event|General Exam|4248,4251|false|false|false|||NEG
Finding|Finding|General Exam|4248,4251|false|false|false|C5848551|Neg - answer|NEG
Finding|Finding|General Exam|4260,4263|false|false|false|C5848551|Neg - answer|NEG
Finding|Finding|General Exam|4272,4275|false|false|false|C5848551|Neg - answer|NEG
Disorder|Disease or Syndrome|General Exam|4289,4292|false|false|false|C0011860|Diabetes Mellitus, Non-Insulin-Dependent|MOD
Event|Event|General Exam|4289,4292|false|false|false|||MOD
Finding|Body Substance|General Exam|4305,4310|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|4305,4310|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|4305,4310|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Lab|Laboratory or Test Result|General Exam|4305,4314|false|false|false|C0221752;C2188659|Red blood cells urine positive|URINE RBC
Anatomy|Cell|General Exam|4311,4314|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|4311,4314|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|4311,4314|false|false|false|C0014792|Erythrocytes|RBC
Anatomy|Cell|General Exam|4318,4321|false|false|false|C0023516|Leukocytes|WBC
Drug|Food|General Exam|4336,4341|true|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|Yeast
Drug|Immunologic Factor|General Exam|4336,4341|true|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|Yeast
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|4336,4341|true|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|Yeast
Drug|Pharmacologic Substance|General Exam|4336,4341|true|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|Yeast
Disorder|Disease or Syndrome|General Exam|4347,4350|true|false|false|C0267963|Exocrine pancreatic insufficiency|Epi
Drug|Amino Acid, Peptide, or Protein|General Exam|4347,4350|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Biologically Active Substance|General Exam|4347,4350|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Hormone|General Exam|4347,4350|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Organic Chemical|General Exam|4347,4350|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Pharmacologic Substance|General Exam|4347,4350|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Event|Event|General Exam|4347,4350|true|false|false|||Epi
Finding|Gene or Genome|General Exam|4347,4350|true|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|Epi
Finding|Intellectual Product|General Exam|4347,4350|true|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|Epi
Procedure|Diagnostic Procedure|General Exam|4347,4350|true|false|false|C0162734;C3641909|Echo-Planar Imaging;Electronic Portal Imaging|Epi
Event|Event|General Exam|4354,4366|true|false|false|||Microbiology
Finding|Functional Concept|General Exam|4354,4366|true|false|false|C0025953;C1571921;C4049106|Microbiological;Microbiology - Laboratory Class;Microbiology Diagnostic Service Section ID|Microbiology
Finding|Intellectual Product|General Exam|4354,4366|true|false|false|C0025953;C1571921;C4049106|Microbiological;Microbiology - Laboratory Class;Microbiology Diagnostic Service Section ID|Microbiology
Procedure|Laboratory Procedure|General Exam|4354,4366|true|false|false|C0085672|Microbiology procedure|Microbiology
Finding|Body Substance|General Exam|4368,4373|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|4368,4373|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|4368,4373|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Procedure|Laboratory Procedure|General Exam|4368,4381|false|false|false|C0430404|Urine culture|URINE CULTURE
Drug|Biomedical or Dental Material|General Exam|4374,4381|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|General Exam|4374,4381|false|false|false|||CULTURE
Finding|Functional Concept|General Exam|4374,4381|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|General Exam|4374,4381|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|General Exam|4374,4381|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Event|Event|General Exam|4383,4388|false|false|false|||Final
Finding|Idea or Concept|General Exam|4383,4388|false|false|false|C1546485|Diagnosis Type - Final|Final
Disorder|Disease or Syndrome|General Exam|4418,4423|false|false|false|C0851353|Blood and lymphatic system disorders|Blood
Event|Event|General Exam|4418,4423|false|false|false|||Blood
Finding|Body Substance|General Exam|4418,4423|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Procedure|Laboratory Procedure|General Exam|4418,4431|false|false|false|C0200949|Blood culture|Blood Culture
Drug|Biomedical or Dental Material|General Exam|4424,4431|false|false|false|C1706355|Culture Dose Form|Culture
Event|Event|General Exam|4424,4431|false|false|false|||Culture
Finding|Functional Concept|General Exam|4424,4431|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|Culture
Finding|Idea or Concept|General Exam|4424,4431|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|Culture
Procedure|Laboratory Procedure|General Exam|4424,4431|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|Culture
Event|Event|General Exam|4440,4446|true|false|false|||growth
Finding|Finding|General Exam|4440,4446|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|growth
Finding|Organ or Tissue Function|General Exam|4440,4446|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|growth
Finding|Organism Function|General Exam|4440,4446|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|growth
Finding|Physiologic Function|General Exam|4440,4446|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|growth
Phenomenon|Phenomenon or Process|General Exam|4440,4446|true|false|false|C2911660|Growth action|growth
Event|Event|General Exam|4452,4457|true|false|false|||final
Finding|Idea or Concept|General Exam|4452,4457|true|false|false|C1546485|Diagnosis Type - Final|final
Finding|Finding|General Exam|4461,4465|true|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|General Exam|4461,4465|true|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|General Exam|4461,4465|true|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|General Exam|4470,4479|true|false|false|||discharge
Finding|Body Substance|General Exam|4470,4479|true|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|General Exam|4470,4479|true|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|General Exam|4470,4479|true|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|General Exam|4470,4479|true|false|false|C0030685|Patient Discharge|discharge
Event|Event|General Exam|4482,4489|false|false|false|||Imaging
Finding|Finding|General Exam|4482,4489|false|false|false|C0740845|Imaging problem|Imaging
Procedure|Diagnostic Procedure|General Exam|4482,4489|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|Imaging
Anatomy|Body Part, Organ, or Organ Component|General Exam|4491,4497|false|false|false|C0030797|Pelvis|Pelvic
Attribute|Clinical Attribute|General Exam|4507,4515|false|false|false|C2926606||FINDINGS
Event|Event|General Exam|4507,4515|false|false|false|||FINDINGS
Finding|Functional Concept|General Exam|4507,4515|false|false|false|C2607943|findings aspects|FINDINGS
Anatomy|Body Part, Organ, or Organ Component|General Exam|4538,4544|false|false|false|C0042149;C1519876;C4266525|Mouse Uterus;Pelvis>Uterus;Uterus|uterus
Anatomy|Tissue|General Exam|4538,4544|false|false|false|C0042149;C1519876;C4266525|Mouse Uterus;Pelvis>Uterus;Uterus|uterus
Disorder|Disease or Syndrome|General Exam|4538,4544|false|false|false|C0042131;C0496919|Neoplasm of uncertain or unknown behavior of uterus;Uterine Diseases|uterus
Disorder|Neoplastic Process|General Exam|4538,4544|false|false|false|C0042131;C0496919|Neoplasm of uncertain or unknown behavior of uterus;Uterine Diseases|uterus
Procedure|Diagnostic Procedure|General Exam|4538,4544|false|false|false|C0869889|examination of uterus|uterus
Event|Event|General Exam|4545,4553|false|false|false|||measures
Finding|Functional Concept|General Exam|4545,4553|false|false|false|C1879489|Measures (attribute)|measures
Event|Event|General Exam|4591,4604|true|false|false|||heterogeneous
Attribute|Clinical Attribute|General Exam|4608,4618|true|false|false|C0550215||appearance
Event|Event|General Exam|4608,4618|true|false|false|||appearance
Procedure|Health Care Activity|General Exam|4608,4618|true|false|false|C2051406|patient appearance regarding mental status exam|appearance
Disorder|Neoplastic Process|General Exam|4637,4645|true|false|false|C0023267;C0042133|Fibroid Tumor;Uterine Fibroids|fibroids
Event|Event|General Exam|4637,4645|true|false|false|||fibroids
Event|Event|General Exam|4646,4650|true|false|false|||seen
Event|Event|General Exam|4665,4669|false|false|false|||exam
Finding|Functional Concept|General Exam|4665,4669|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|General Exam|4665,4669|false|false|false|C0582103|Medical Examination|exam
Finding|Idea or Concept|General Exam|4689,4695|false|false|false|C1550462|Observation Interpretation - better|better
Event|Event|General Exam|4696,4706|false|false|false|||evaluation
Finding|Idea or Concept|General Exam|4696,4706|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|General Exam|4696,4706|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Anatomy|Body Part, Organ, or Organ Component|General Exam|4714,4720|false|false|false|C0042149;C1519876;C4266525|Mouse Uterus;Pelvis>Uterus;Uterus|uterus
Anatomy|Tissue|General Exam|4714,4720|false|false|false|C0042149;C1519876;C4266525|Mouse Uterus;Pelvis>Uterus;Uterus|uterus
Disorder|Disease or Syndrome|General Exam|4714,4720|false|false|false|C0042131;C0496919|Neoplasm of uncertain or unknown behavior of uterus;Uterine Diseases|uterus
Disorder|Neoplastic Process|General Exam|4714,4720|false|false|false|C0042131;C0496919|Neoplasm of uncertain or unknown behavior of uterus;Uterine Diseases|uterus
Procedure|Diagnostic Procedure|General Exam|4714,4720|false|false|false|C0869889|examination of uterus|uterus
Anatomy|Body Part, Organ, or Organ Component|General Exam|4725,4731|false|false|false|C0001575;C0229243;C4522151|Adnexa;Ocular adnexa structure;Uterine adnexae structure|adnexa
Event|Event|General Exam|4750,4756|false|false|false|||stripe
Finding|Functional Concept|General Exam|4776,4780|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|General Exam|4776,4786|false|false|false|C0227874|Structure of left ovary|left ovary
Anatomy|Body Part, Organ, or Organ Component|General Exam|4781,4786|false|false|false|C0029939;C0227898;C4266530|Both ovaries;Ovary;Pelvis>Ovary|ovary
Disorder|Disease or Syndrome|General Exam|4781,4786|false|false|false|C0029928;C0496920|Neoplasm of uncertain or unknown behavior of ovary;Ovarian Diseases|ovary
Disorder|Neoplastic Process|General Exam|4781,4786|false|false|false|C0029928;C0496920|Neoplasm of uncertain or unknown behavior of ovary;Ovarian Diseases|ovary
Event|Event|General Exam|4781,4786|false|false|false|||ovary
Event|Event|General Exam|4787,4795|false|false|false|||measures
Finding|Functional Concept|General Exam|4821,4826|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|General Exam|4821,4832|false|false|false|C0227873|Structure of right ovary|right ovary
Anatomy|Body Part, Organ, or Organ Component|General Exam|4827,4832|false|false|false|C0029939;C0227898;C4266530|Both ovaries;Ovary;Pelvis>Ovary|ovary
Disorder|Disease or Syndrome|General Exam|4827,4832|false|false|false|C0029928;C0496920|Neoplasm of uncertain or unknown behavior of ovary;Ovarian Diseases|ovary
Disorder|Neoplastic Process|General Exam|4827,4832|false|false|false|C0029928;C0496920|Neoplasm of uncertain or unknown behavior of ovary;Ovarian Diseases|ovary
Event|Event|General Exam|4833,4841|false|false|false|||measures
Finding|Finding|General Exam|4880,4889|false|false|false|C4697723|Echogenic|echogenic
Event|Event|General Exam|4890,4895|false|false|false|||focus
Finding|Functional Concept|General Exam|4890,4895|false|false|false|C1285542|Has focus|focus
Finding|Functional Concept|General Exam|4907,4912|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|General Exam|4907,4918|false|false|false|C0227873|Structure of right ovary|right ovary
Anatomy|Body Part, Organ, or Organ Component|General Exam|4913,4918|false|false|false|C0029939;C0227898;C4266530|Both ovaries;Ovary;Pelvis>Ovary|ovary
Disorder|Disease or Syndrome|General Exam|4913,4918|false|false|false|C0029928;C0496920|Neoplasm of uncertain or unknown behavior of ovary;Ovarian Diseases|ovary
Disorder|Neoplastic Process|General Exam|4913,4918|false|false|false|C0029928;C0496920|Neoplasm of uncertain or unknown behavior of ovary;Ovarian Diseases|ovary
Event|Event|General Exam|4919,4928|false|false|false|||measuring
Finding|Finding|General Exam|4944,4950|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|General Exam|4944,4950|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Disorder|Anatomical Abnormality|General Exam|4959,4975|false|false|false|C0333145|Hemorrhagic cyst|hemorrhagic cyst
Disorder|Anatomical Abnormality|General Exam|4971,4975|false|false|false|C0010709|Cyst|cyst
Event|Event|General Exam|4971,4975|false|false|false|||cyst
Finding|Body Substance|General Exam|4971,4975|false|false|false|C1546594;C1550626|SpecimenType - Cyst|cyst
Finding|Intellectual Product|General Exam|4971,4975|false|false|false|C1546594;C1550626|SpecimenType - Cyst|cyst
Anatomy|Body Part, Organ, or Organ Component|General Exam|4977,4989|false|false|false|C0227898|Both ovaries|Both ovaries
Anatomy|Body Part, Organ, or Organ Component|General Exam|4982,4989|false|false|false|C0029939;C0227898|Both ovaries;Ovary|ovaries
Event|Event|General Exam|4990,5001|false|false|false|||demonstrate
Anatomy|Body Part, Organ, or Organ Component|General Exam|5010,5018|false|false|false|C0003842|Arteries|arterial
Anatomy|Body Part, Organ, or Organ Component|General Exam|5023,5029|false|false|false|C0042449|Veins|venous
Event|Event|General Exam|5030,5039|false|false|false|||waveforms
Phenomenon|Natural Phenomenon or Process|General Exam|5030,5039|false|false|false|C0450448|Waveforms|waveforms
Event|Event|Impression|5064,5072|true|false|false|||evidence
Finding|Idea or Concept|Impression|5064,5072|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Impression|5064,5075|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Anatomy|Body Part, Organ, or Organ Component|Impression|5076,5083|true|false|false|C0205065|Ovarian|ovarian
Disorder|Anatomical Abnormality|Impression|5076,5091|true|false|false|C0149952|Ovarian Torsion|ovarian torsion
Event|Event|Impression|5084,5091|true|false|false|||torsion
Finding|Pathologic Function|Impression|5084,5091|true|false|false|C0040480;C1265748|Musculoskeletal torsion (function);Torsion (malposition)|torsion
Finding|Physiologic Function|Impression|5084,5091|true|false|false|C0040480;C1265748|Musculoskeletal torsion (function);Torsion (malposition)|torsion
Finding|Functional Concept|Impression|5104,5109|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|Impression|5110,5117|false|false|false|C0205065|Ovarian|ovarian
Disorder|Anatomical Abnormality|Impression|5118,5134|false|false|false|C0333145|Hemorrhagic cyst|hemorrhagic cyst
Disorder|Anatomical Abnormality|Impression|5130,5134|false|false|false|C0010709|Cyst|cyst
Event|Event|Impression|5130,5134|false|false|false|||cyst
Finding|Body Substance|Impression|5130,5134|false|false|false|C1546594;C1550626|SpecimenType - Cyst|cyst
Finding|Intellectual Product|Impression|5130,5134|false|false|false|C1546594;C1550626|SpecimenType - Cyst|cyst
Attribute|Clinical Attribute|Impression|5139,5145|false|false|false|C1644645||CT abd
Anatomy|Body Location or Region|Impression|5142,5145|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|abd
Disorder|Cell or Molecular Dysfunction|Impression|5142,5145|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|abd
Anatomy|Body Part, Organ, or Organ Component|Impression|5146,5152|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Anatomy|Body Space or Junction|Impression|5146,5152|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Disorder|Neoplastic Process|Impression|5146,5152|false|false|false|C0153663|Malignant neoplasm of pelvis|pelvis
Event|Event|Impression|5146,5152|false|false|false|||pelvis
Finding|Finding|Impression|5146,5152|false|false|false|C0812455|Pelvis problem|pelvis
Event|Event|Impression|5154,5155|false|false|false|||/
Drug|Indicator, Reagent, or Diagnostic Aid|Impression|5157,5165|false|false|false|C0009924|Contrast Media|contrast
Event|Event|Impression|5157,5165|false|false|false|||contrast
Event|Event|Impression|5193,5203|false|false|false|||granulomas
Finding|Pathologic Function|Impression|5193,5203|false|false|false|C0018188|Granuloma|granulomas
Anatomy|Body Location or Region|Impression|5212,5216|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Impression|5212,5216|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Impression|5212,5216|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Impression|5212,5216|false|false|false|C0740941|Lung Problem|lung
Drug|Chemical Viewed Functionally|Impression|5217,5222|false|false|false|C0178499|Base|bases
Event|Event|Impression|5217,5222|false|false|false|||bases
Event|Event|Impression|5227,5233|false|false|false|||stable
Finding|Intellectual Product|Impression|5227,5233|false|false|false|C1547311|Patient Condition Code - Stable|stable
Finding|Finding|Impression|5247,5250|true|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Impression|5247,5250|true|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Anatomy|Body Part, Organ, or Organ Component|Impression|5257,5266|true|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Impression|5257,5266|true|false|false|C2707265||pulmonary
Finding|Finding|Impression|5257,5266|true|false|false|C4522268|Pulmonary (intended site)|pulmonary
Event|Event|Impression|5268,5274|true|false|false|||nodule
Disorder|Disease or Syndrome|Impression|5277,5290|false|false|false|C0521530|Lung consolidation|consolidation
Event|Event|Impression|5277,5290|false|false|false|||consolidation
Event|Event|Impression|5295,5303|false|false|false|||effusion
Finding|Body Substance|Impression|5295,5303|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|Impression|5295,5303|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|Impression|5295,5303|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Anatomy|Body Part, Organ, or Organ Component|Impression|5309,5316|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|Impression|5309,5316|false|false|false|C1314974|Cardiac attachment|cardiac
Anatomy|Body Location or Region|Impression|5309,5321|false|false|false|C0225811|Structure of apex of heart|cardiac apex
Anatomy|Cell Component|Impression|5317,5321|false|false|false|C3890171|dinoflagellate apex|apex
Drug|Amino Acid, Peptide, or Protein|Impression|5317,5321|false|false|false|C0140145|APEX1 protein, human|apex
Drug|Enzyme|Impression|5317,5321|false|false|false|C0140145|APEX1 protein, human|apex
Finding|Gene or Genome|Impression|5317,5321|false|false|false|C1332102|APEX1 gene|apex
Event|Event|Impression|5332,5338|false|false|false|||normal
Event|Event|Impression|5340,5346|false|false|false|||limits
Finding|Functional Concept|Impression|5340,5346|false|false|false|C0439801|Limited (extensiveness)|limits
Drug|Organic Chemical|Impression|5350,5358|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|Complete
Drug|Pharmacologic Substance|Impression|5350,5358|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|Complete
Drug|Vitamin|Impression|5350,5358|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|Complete
Finding|Functional Concept|Impression|5350,5358|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|Complete
Finding|Idea or Concept|Impression|5350,5358|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|Complete
Event|Event|Impression|5359,5369|false|false|false|||evaluation
Finding|Idea or Concept|Impression|5359,5369|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|Impression|5359,5369|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Finding|Functional Concept|Impression|5377,5392|false|false|false|C1512911|Intraabdominal Route of Administration|intra-abdominal
Anatomy|Body Part, Organ, or Organ Component|Impression|5393,5400|false|false|false|C0042779;C1285145|Structure of viscus;Viscera|viscera
Event|Event|Impression|5404,5411|false|false|false|||limited
Event|Event|Impression|5434,5443|false|false|false|||technique
Finding|Functional Concept|Impression|5434,5443|false|false|false|C0449851|Techniques|technique
Anatomy|Body Part, Organ, or Organ Component|Impression|5458,5463|true|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|Impression|5458,5463|true|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|Impression|5458,5463|true|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|Impression|5458,5463|true|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|Impression|5458,5463|true|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|Impression|5458,5463|true|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|Impression|5458,5463|true|false|false|||liver
Finding|Finding|Impression|5458,5463|true|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|Impression|5458,5463|true|false|false|C0872387|Procedures on liver|liver
Event|Event|Impression|5472,5483|true|false|false|||homogeneous
Event|Event|Impression|5499,5505|true|false|false|||lesion
Finding|Finding|Impression|5499,5505|true|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|Impression|5499,5505|true|false|false|C0221198;C1546698|Lesion|lesion
Finding|Functional Concept|Impression|5534,5541|true|false|false|C0521378|Biliary|biliary
Event|Event|Impression|5550,5560|false|false|false|||dilatation
Finding|Finding|Impression|5550,5560|false|false|false|C0012359;C0700124|Dilated;Pathological Dilatation|dilatation
Finding|Pathologic Function|Impression|5550,5560|false|false|false|C0012359;C0700124|Dilated;Pathological Dilatation|dilatation
Procedure|Therapeutic or Preventive Procedure|Impression|5550,5560|false|false|false|C1322279|Dilate procedure|dilatation
Event|Event|Impression|5564,5574|false|false|false|||identified
Anatomy|Body Part, Organ, or Organ Component|Impression|5581,5592|false|false|false|C0016976;C1524055;C4071903|Abdomen>Gallbladder;Gallbladder;Gallbladder (MMHCC)|gallbladder
Anatomy|Tissue|Impression|5581,5592|false|false|false|C0016976;C1524055;C4071903|Abdomen>Gallbladder;Gallbladder;Gallbladder (MMHCC)|gallbladder
Procedure|Health Care Activity|Impression|5581,5592|false|false|false|C2032932|examination of gallbladder|gallbladder
Anatomy|Body Part, Organ, or Organ Component|Impression|5594,5600|false|false|false|C0037993;C4037984|Abdomen>Spleen;Spleen|spleen
Disorder|Neoplastic Process|Impression|5594,5600|false|false|false|C0153470|Malignant neoplasm of spleen|spleen
Event|Event|Impression|5594,5600|false|false|false|||spleen
Finding|Finding|Impression|5594,5600|false|false|false|C0812414|Spleen problem|spleen
Procedure|Therapeutic or Preventive Procedure|Impression|5594,5600|false|false|false|C0869677|Procedures on Spleen|spleen
Anatomy|Body Part, Organ, or Organ Component|Impression|5606,5614|false|false|false|C0030274;C4037927|Abdomen>Pancreas;Pancreas|pancreas
Disorder|Disease or Syndrome|Impression|5606,5614|false|false|false|C0030286;C0347284|Benign tumor of pancreas;Pancreatic Diseases|pancreas
Disorder|Neoplastic Process|Impression|5606,5614|false|false|false|C0030286;C0347284|Benign tumor of pancreas;Pancreatic Diseases|pancreas
Drug|Organic Chemical|Impression|5606,5614|false|false|false|C0771711|pancreas extract|pancreas
Drug|Pharmacologic Substance|Impression|5606,5614|false|false|false|C0771711|pancreas extract|pancreas
Event|Event|Impression|5606,5614|false|false|false|||pancreas
Finding|Finding|Impression|5606,5614|false|false|false|C0813176|Pancreas problem|pancreas
Procedure|Health Care Activity|Impression|5606,5614|false|false|false|C0869826|Procedures on Pancreas|pancreas
Event|Event|Impression|5616,5622|false|false|false|||appear
Finding|Finding|Impression|5623,5643|false|false|false|C0442816||within normal limits
Event|Event|Impression|5637,5643|false|false|false|||limits
Finding|Functional Concept|Impression|5637,5643|false|false|false|C0439801|Limited (extensiveness)|limits
Anatomy|Body Part, Organ, or Organ Component|Impression|5649,5656|true|false|false|C0001625|Adrenal Glands|adrenal
Finding|Finding|Impression|5649,5656|true|false|false|C0521428|Adrenal|adrenal
Anatomy|Body Part, Organ, or Organ Component|Impression|5649,5663|true|false|false|C0001625|Adrenal Glands|adrenal glands
Anatomy|Body Part, Organ, or Organ Component|Impression|5657,5663|true|false|false|C1285092|Gland|glands
Event|Event|Impression|5668,5677|true|false|false|||symmetric
Finding|Conceptual Entity|Impression|5668,5677|true|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Finding|Impression|5668,5677|true|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Event|Event|Impression|5693,5699|true|false|false|||nodule
Anatomy|Body Part, Organ, or Organ Component|Impression|5705,5712|true|false|false|C0022646;C0227665|Both kidneys;Kidney|kidneys
Event|Event|Impression|5720,5731|true|false|false|||homogeneous
Event|Event|Impression|5747,5753|true|false|false|||lesion
Finding|Finding|Impression|5747,5753|true|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|Impression|5747,5753|true|false|false|C0221198;C1546698|Lesion|lesion
Disorder|Disease or Syndrome|Impression|5757,5771|true|false|false|C0020295|Hydronephrosis|hydronephrosis
Event|Event|Impression|5757,5771|true|false|false|||hydronephrosis
Anatomy|Body Location or Region|Impression|5777,5786|false|false|false|C0000726|Abdomen|abdominal
Anatomy|Body Part, Organ, or Organ Component|Impression|5777,5792|false|false|false|C0003484;C4037989|Abdomen>Aorta.abdominal;Abdominal aorta structure|abdominal aorta
Procedure|Health Care Activity|Impression|5777,5792|false|false|false|C2228415|examination of abdominal aorta|abdominal aorta
Anatomy|Body Part, Organ, or Organ Component|Impression|5787,5792|false|false|false|C0003483;C4037978|Aorta;Chest+Abdomen>Aorta|aorta
Procedure|Health Care Activity|Impression|5787,5792|false|false|false|C0869784|Procedure on aorta|aorta
Event|Event|Impression|5797,5811|false|false|false|||non-aneurysmal
Event|Event|Impression|5838,5844|false|false|false|||course
Finding|Functional Concept|Impression|5850,5856|false|false|false|C1522484;C1561503;C1705190|Precision - second;Second Suffix;metastatic qualifier|second
Finding|Idea or Concept|Impression|5850,5856|false|false|false|C1522484;C1561503;C1705190|Precision - second;Second Suffix;metastatic qualifier|second
Finding|Intellectual Product|Impression|5850,5856|false|false|false|C1522484;C1561503;C1705190|Precision - second;Second Suffix;metastatic qualifier|second
Event|Event|Impression|5868,5876|false|false|false|||portions
Anatomy|Body Part, Organ, or Organ Component|Impression|5884,5892|false|false|false|C0013303|Duodenum|duodenum
Disorder|Neoplastic Process|Impression|5884,5892|false|false|false|C0153426;C0496869|Benign neoplasm of duodenum;Malignant neoplasm of duodenum|duodenum
Event|Event|Impression|5909,5918|false|false|false|||thickened
Event|Event|Impression|5940,5955|false|false|false|||underdistension
Anatomy|Body Location or Region|Impression|5960,5971|true|false|false|C0021852;C4319010|Abdomen>Small bowel;Intestines, Small|small bowel
Anatomy|Body Part, Organ, or Organ Component|Impression|5960,5971|true|false|false|C0021852;C4319010|Abdomen>Small bowel;Intestines, Small|small bowel
Disorder|Disease or Syndrome|Impression|5960,5983|true|false|false|C0235329|Small bowel obstruction|small bowel obstruction
Anatomy|Body Part, Organ, or Organ Component|Impression|5966,5971|true|false|false|C0021853|Intestines|bowel
Disorder|Disease or Syndrome|Impression|5966,5983|true|false|false|C0021843|Intestinal Obstruction|bowel obstruction
Event|Event|Impression|5972,5983|true|false|false|||obstruction
Finding|Finding|Impression|5972,5983|true|false|false|C0028778|Obstruction|obstruction
Event|Event|Impression|5988,5998|true|false|false|||identified
Anatomy|Body Part, Organ, or Organ Component|Impression|6004,6012|false|false|false|C0003617;C4037994|Abdomen+Pelvis>Appendix;Appendix|appendix
Disorder|Neoplastic Process|Impression|6004,6012|false|false|false|C0348899;C0496779;C0496860|Benign neoplasm of appendix;Malignant neoplasm of appendix;Neoplasm of uncertain or unknown behavior of appendix|appendix
Event|Event|Impression|6004,6012|false|false|false|||appendix
Finding|Intellectual Product|Impression|6004,6012|false|false|false|C1552860|appendix - HTML link|appendix
Procedure|Therapeutic or Preventive Procedure|Impression|6004,6012|false|false|false|C0869813|Procedure on appendix|appendix
Finding|Finding|Impression|6016,6020|false|false|false|C5575035|Well (answer to question)|well
Event|Event|Impression|6021,6031|false|false|false|||visualized
Attribute|Clinical Attribute|Impression|6050,6060|false|false|false|C0550215||appearance
Event|Event|Impression|6050,6060|false|false|false|||appearance
Procedure|Health Care Activity|Impression|6050,6060|false|false|false|C2051406|patient appearance regarding mental status exam|appearance
Finding|Functional Concept|Impression|6074,6078|true|false|false|C0332296|Free of (attribute)|free
Finding|Pathologic Function|Impression|6074,6084|true|false|false|C0013687|effusion|free fluid
Drug|Substance|Impression|6079,6084|true|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|Impression|6079,6084|true|false|false|||fluid
Finding|Intellectual Product|Impression|6079,6084|true|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|Impression|6088,6092|true|false|false|||free
Finding|Functional Concept|Impression|6088,6092|true|false|false|C0332296|Free of (attribute)|free
Drug|Inorganic Chemical|Impression|6093,6096|true|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|Impression|6093,6096|true|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|Impression|6093,6096|true|false|false|C0001861;C3536832|Air (substance);air|air
Event|Event|Impression|6093,6096|true|false|false|||air
Finding|Finding|Impression|6093,6096|true|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|Impression|6093,6096|true|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|Impression|6093,6096|true|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Attribute|Clinical Attribute|Impression|6102,6111|true|false|false|C0882057||CT PELVIS
Procedure|Diagnostic Procedure|Impression|6102,6111|true|false|false|C0412628|Computed tomography of pelvis|CT PELVIS
Anatomy|Body Part, Organ, or Organ Component|Impression|6105,6111|true|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|PELVIS
Anatomy|Body Space or Junction|Impression|6105,6111|true|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|PELVIS
Disorder|Neoplastic Process|Impression|6105,6111|true|false|false|C0153663|Malignant neoplasm of pelvis|PELVIS
Event|Event|Impression|6105,6111|true|false|false|||PELVIS
Finding|Finding|Impression|6105,6111|true|false|false|C0812455|Pelvis problem|PELVIS
Finding|Functional Concept|Impression|6120,6131|true|false|false|C1522726|Intravenous Route of Administration|INTRAVENOUS
Drug|Indicator, Reagent, or Diagnostic Aid|Impression|6120,6140|true|false|false|C4072741|IV contrast|INTRAVENOUS CONTRAST
Drug|Indicator, Reagent, or Diagnostic Aid|Impression|6132,6140|true|false|false|C0009924|Contrast Media|CONTRAST
Event|Event|Impression|6132,6140|true|false|false|||CONTRAST
Finding|Idea or Concept|Impression|6146,6153|false|false|false|C1555582|Initial (abbreviation)|Initial
Event|Event|Impression|6162,6174|false|false|false|||demonstrated
Drug|Biomedical or Dental Material|Impression|6177,6182|false|false|false|C0302909;C1378566|Solid Dose Form;solid substance|solid
Drug|Substance|Impression|6177,6182|false|false|false|C0302909;C1378566|Solid Dose Form;solid substance|solid
Event|Event|Impression|6183,6187|false|false|false|||mass
Finding|Finding|Impression|6183,6187|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|Impression|6183,6187|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|Impression|6183,6187|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Disorder|Congenital Abnormality|Impression|6193,6204|false|false|false|C0000768|Congenital Abnormality|abnormality
Event|Event|Impression|6193,6204|false|false|false|||abnormality
Finding|Finding|Impression|6193,6204|false|false|false|C1704258|Abnormality|abnormality
Anatomy|Body Part, Organ, or Organ Component|Impression|6212,6217|false|false|false|C0007531|Cecum|cecal
Event|Event|Impression|6218,6221|false|false|false|||tip
Finding|Gene or Genome|Impression|6218,6221|false|false|false|C1705504;C1823282;C1825626;C1825978|ITFG1 gene;KAT5 wt Allele;METTL8 gene;TIPRL gene|tip
Procedure|Therapeutic or Preventive Procedure|Impression|6218,6221|false|false|false|C0673828|TIP regimen|tip
Event|Event|Impression|6223,6232|false|false|false|||measuring
Event|Event|Impression|6286,6296|false|false|false|||concerning
Anatomy|Body Part, Organ, or Organ Component|Impression|6303,6308|false|false|false|C0007531|Cecum|cecal
Finding|Finding|Impression|6303,6313|false|true|false|C3670817|Cecal mass|cecal mass
Event|Event|Impression|6309,6313|false|false|false|||mass
Finding|Finding|Impression|6309,6313|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|Impression|6309,6313|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|Impression|6309,6313|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Event|Event|Impression|6315,6325|false|false|false|||rescanning
Finding|Functional Concept|Impression|6331,6338|false|false|false|C0439801;C3542948|Limited (extensiveness);Limited component (foundation metadata concept)|limited
Finding|Intellectual Product|Impression|6331,6338|false|false|false|C0439801;C3542948|Limited (extensiveness);Limited component (foundation metadata concept)|limited
Anatomy|Body Part, Organ, or Organ Component|Impression|6351,6357|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Anatomy|Body Space or Junction|Impression|6351,6357|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Disorder|Neoplastic Process|Impression|6351,6357|false|false|false|C0153663|Malignant neoplasm of pelvis|pelvis
Event|Event|Impression|6351,6357|false|false|false|||pelvis
Finding|Finding|Impression|6351,6357|false|false|false|C0812455|Pelvis problem|pelvis
Event|Event|Impression|6378,6385|false|false|false|||passage
Procedure|Laboratory Procedure|Impression|6378,6385|false|false|false|C1709474|Passage tissue culture technique|passage
Anatomy|Body Space or Junction|Impression|6389,6393|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Impression|6389,6393|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Impression|6389,6393|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Impression|6389,6393|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Drug|Indicator, Reagent, or Diagnostic Aid|Impression|6394,6402|false|false|false|C0009924|Contrast Media|contrast
Event|Event|Impression|6394,6402|false|false|false|||contrast
Event|Event|Impression|6404,6414|false|false|false|||confirming
Finding|Finding|Impression|6404,6414|false|false|false|C0750484|Confirmation|confirming
Event|Event|Impression|6420,6427|false|false|false|||finding
Finding|Finding|Impression|6420,6427|false|false|false|C0037088;C0243095;C2825141|Experimental Finding;Finding;Signs and Symptoms|finding
Finding|Sign or Symptom|Impression|6420,6427|false|false|false|C0037088;C0243095;C2825141|Experimental Finding;Finding;Signs and Symptoms|finding
Event|Event|Impression|6432,6445|false|false|false|||demonstrating
Event|Event|Impression|6453,6457|false|false|false|||mass
Finding|Finding|Impression|6453,6457|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|Impression|6453,6457|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|Impression|6453,6457|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Event|Event|Impression|6463,6473|false|false|false|||thickening
Finding|Finding|Impression|6463,6473|false|false|false|C0205400|Thickened|thickening
Anatomy|Body Part, Organ, or Organ Component|Impression|6491,6496|false|false|false|C0007531|Cecum|cecal
Anatomy|Body Part, Organ, or Organ Component|Impression|6491,6501|false|false|false|C0734005|Wall of cecum|cecal wall
Anatomy|Body Part, Organ, or Organ Component|Impression|6525,6533|true|false|false|C0003617;C4037994|Abdomen+Pelvis>Appendix;Appendix|appendix
Disorder|Neoplastic Process|Impression|6525,6533|true|false|false|C0348899;C0496779;C0496860|Benign neoplasm of appendix;Malignant neoplasm of appendix;Neoplasm of uncertain or unknown behavior of appendix|appendix
Event|Event|Impression|6525,6533|true|false|false|||appendix
Finding|Intellectual Product|Impression|6525,6533|true|false|false|C1552860|appendix - HTML link|appendix
Procedure|Therapeutic or Preventive Procedure|Impression|6525,6533|true|false|false|C0869813|Procedure on appendix|appendix
Event|Event|Impression|6537,6543|true|false|false|||normal
Finding|Functional Concept|Impression|6571,6583|true|false|false|C0333348|Inflammatory|inflammatory
Event|Event|Impression|6584,6590|true|false|false|||change
Finding|Functional Concept|Impression|6584,6590|true|false|false|C0392747|Changing|change
Procedure|Therapeutic or Preventive Procedure|Impression|6584,6590|true|false|false|C4319952|Change - procedure|change
Anatomy|Body Part, Organ, or Organ Component|Impression|6615,6620|true|false|false|C0009368;C4071907|Abdomen+Pelvis>Colon;Colon structure (body structure)|colon
Disorder|Disease or Syndrome|Impression|6615,6620|true|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Disorder|Neoplastic Process|Impression|6615,6620|true|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Event|Event|Impression|6615,6620|true|false|false|||colon
Finding|Finding|Impression|6615,6620|true|false|false|C0750873|COLON PROBLEM|colon
Event|Event|Impression|6624,6630|true|false|false|||normal
Event|Event|Impression|6639,6647|true|false|false|||evidence
Finding|Idea or Concept|Impression|6639,6647|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Impression|6639,6650|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Event|Event|Impression|6652,6663|true|false|false|||obstruction
Finding|Finding|Impression|6652,6663|true|false|false|C0028778|Obstruction|obstruction
Event|Event|Impression|6668,6680|true|false|false|||inflammation
Finding|Pathologic Function|Impression|6668,6680|true|false|false|C0021368|Inflammation|inflammation
Procedure|Health Care Activity|Impression|6686,6694|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Procedure|Therapeutic or Preventive Procedure|Impression|6686,6694|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Procedure|Therapeutic or Preventive Procedure|Impression|6686,6706|false|false|false|C0677554||surgical anastomosis
Anatomy|Body Space or Junction|Impression|6695,6706|false|false|false|C0500470|Anatomical anastomosis|anastomosis
Disorder|Acquired Abnormality|Impression|6695,6706|false|false|false|C0332853|Anastomosis|anastomosis
Event|Event|Impression|6695,6706|false|false|false|||anastomosis
Procedure|Therapeutic or Preventive Procedure|Impression|6695,6706|false|false|false|C0677554||anastomosis
Anatomy|Body Location or Region|Impression|6718,6723|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|Impression|6718,6723|false|false|false|C2003888|Lower (action)|lower
Anatomy|Cell Component|Impression|6724,6731|false|false|false|C1660780|midline cell component|midline
Anatomy|Body Part, Organ, or Organ Component|Impression|6733,6739|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Anatomy|Body Space or Junction|Impression|6733,6739|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Disorder|Neoplastic Process|Impression|6733,6739|false|false|false|C0153663|Malignant neoplasm of pelvis|pelvis
Finding|Finding|Impression|6733,6739|false|false|false|C0812455|Pelvis problem|pelvis
Event|Event|Impression|6749,6761|false|false|false|||unremarkable
Anatomy|Body Part, Organ, or Organ Component|Impression|6775,6781|true|false|false|C0030797|Pelvis|pelvic
Finding|Body Substance|Impression|6775,6792|true|false|false|C0237041|pelvic free fluid|pelvic free fluid
Finding|Functional Concept|Impression|6782,6786|true|false|false|C0332296|Free of (attribute)|free
Finding|Pathologic Function|Impression|6782,6792|true|false|false|C0013687|effusion|free fluid
Drug|Substance|Impression|6787,6792|true|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|Impression|6787,6792|true|false|false|||fluid
Finding|Intellectual Product|Impression|6787,6792|true|false|false|C1546638|Fluid Specimen Code|fluid
Anatomy|Body Part, Organ, or Organ Component|Impression|6798,6804|false|false|false|C0042149;C1519876;C4266525|Mouse Uterus;Pelvis>Uterus;Uterus|uterus
Anatomy|Tissue|Impression|6798,6804|false|false|false|C0042149;C1519876;C4266525|Mouse Uterus;Pelvis>Uterus;Uterus|uterus
Disorder|Disease or Syndrome|Impression|6798,6804|false|false|false|C0042131;C0496919|Neoplasm of uncertain or unknown behavior of uterus;Uterine Diseases|uterus
Disorder|Neoplastic Process|Impression|6798,6804|false|false|false|C0042131;C0496919|Neoplasm of uncertain or unknown behavior of uterus;Uterine Diseases|uterus
Event|Event|Impression|6798,6804|false|false|false|||uterus
Procedure|Diagnostic Procedure|Impression|6798,6804|false|false|false|C0869889|examination of uterus|uterus
Anatomy|Body Part, Organ, or Organ Component|Impression|6810,6816|false|false|false|C0001575;C0229243;C4522151|Adnexa;Ocular adnexa structure;Uterine adnexae structure|adnexa
Event|Event|Impression|6818,6824|false|false|false|||appear
Finding|Finding|Impression|6825,6845|false|false|false|C0442816||within normal limits
Event|Event|Impression|6839,6845|false|false|false|||limits
Finding|Functional Concept|Impression|6839,6845|false|false|false|C0439801|Limited (extensiveness)|limits
Anatomy|Body Part, Organ, or Organ Component|Impression|6851,6858|false|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|Impression|6851,6858|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Event|Event|Impression|6851,6858|false|false|false|||bladder
Procedure|Therapeutic or Preventive Procedure|Impression|6851,6858|false|false|false|C0872388|Procedures on bladder|bladder
Event|Event|Impression|6871,6880|false|false|false|||distended
Finding|Finding|Impression|6871,6880|false|false|false|C0700124|Dilated|distended
Event|Event|Impression|6900,6912|false|false|false|||unremarkable
Procedure|Therapeutic or Preventive Procedure|Impression|6932,6940|true|false|false|C1293134|Enlargement procedure|enlarged
Anatomy|Body Part, Organ, or Organ Component|Impression|6941,6947|true|false|false|C0030797|Pelvis|pelvic
Anatomy|Body Location or Region|Impression|6952,6960|true|false|false|C0018246|Inguinal region|inguinal
Anatomy|Body Part, Organ, or Organ Component|Impression|6952,6972|true|false|false|C0729596|Inguinal lymph node group|inguinal lymph nodes
Finding|Body Substance|Impression|6961,6966|true|false|false|C0024202|Lymph|lymph
Anatomy|Body Part, Organ, or Organ Component|Impression|6961,6972|true|false|false|C0024204|lymph nodes|lymph nodes
Disorder|Neoplastic Process|Impression|6961,6972|true|false|false|C0154054|benign neoplasm of lymph nodes|lymph nodes
Event|Event|Impression|6977,6987|false|false|false|||identified
Anatomy|Body Part, Organ, or Organ Component|Impression|6990,6997|false|false|false|C0262950;C4520924|Bone Tissue, Human;Skeletal bone|OSSEOUS
Anatomy|Tissue|Impression|6990,6997|false|false|false|C0262950;C4520924|Bone Tissue, Human;Skeletal bone|OSSEOUS
Event|Event|Impression|6998,7008|false|false|false|||STRUCTURES
Anatomy|Body Part, Organ, or Organ Component|Impression|7013,7017|true|false|false|C0262950;C1442209|Skeletal bone;XXX bone|bone
Finding|Body Substance|Impression|7013,7017|true|false|false|C1546560;C1550616|Specimen Type - Bone|bone
Finding|Intellectual Product|Impression|7013,7017|true|false|false|C1546560;C1550616|Specimen Type - Bone|bone
Finding|Individual Behavior|Impression|7018,7029|true|false|false|C0233520|Destructive behavior|destructive
Event|Event|Impression|7030,7036|true|false|false|||lesion
Finding|Finding|Impression|7030,7036|true|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|Impression|7030,7036|true|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|Impression|7040,7045|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Disorder|Injury or Poisoning|Impression|7046,7054|true|false|false|C0016658|Fracture|fracture
Event|Event|Impression|7046,7054|true|false|false|||fracture
Event|Event|Impression|7060,7070|false|false|false|||identified
Attribute|Clinical Attribute|Impression|7090,7098|false|false|false|C2926606||Findings
Event|Event|Impression|7090,7098|false|false|false|||Findings
Finding|Functional Concept|Impression|7090,7098|false|false|false|C2607943|findings aspects|Findings
Event|Event|Impression|7099,7109|false|false|false|||consistent
Finding|Idea or Concept|Impression|7099,7109|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|Impression|7099,7114|false|false|false|C0332290|Consistent with|consistent with
Anatomy|Body Part, Organ, or Organ Component|Impression|7122,7127|false|false|false|C0007531|Cecum|cecal
Finding|Finding|Impression|7122,7132|false|false|false|C3670817|Cecal mass|cecal mass
Event|Event|Impression|7128,7132|false|false|false|||mass
Finding|Finding|Impression|7128,7132|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|Impression|7128,7132|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|Impression|7128,7132|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Event|Event|Impression|7137,7147|false|false|false|||thickening
Finding|Finding|Impression|7137,7147|false|false|false|C0205400|Thickened|thickening
Anatomy|Body Part, Organ, or Organ Component|Impression|7156,7161|false|false|false|C0007531|Cecum|cecal
Event|Event|Impression|7162,7165|false|false|false|||tip
Finding|Gene or Genome|Impression|7162,7165|false|false|false|C1705504;C1823282;C1825626;C1825978|ITFG1 gene;KAT5 wt Allele;METTL8 gene;TIPRL gene|tip
Procedure|Therapeutic or Preventive Procedure|Impression|7162,7165|false|false|false|C0673828|TIP regimen|tip
Disorder|Neoplastic Process|Impression|7181,7189|false|false|false|C0027651;C1882062|Neoplasms;Neoplastic disease|neoplasm
Event|Event|Impression|7181,7189|false|false|false|||neoplasm
Finding|Finding|Impression|7191,7199|false|false|false|C0741302|atypia morphology|Atypical
Disorder|Disease or Syndrome|Impression|7200,7210|false|false|false|C0009450|Communicable Diseases|infectious
Event|Event|Impression|7200,7210|false|false|false|||infectious
Anatomy|Body Part, Organ, or Organ Component|Impression|7212,7219|false|false|false|C1184743|bony process|process
Drug|Pharmacologic Substance|Impression|7212,7219|false|false|false|C1951340|Process Pharmacologic Substance|process
Event|Event|Impression|7212,7219|false|false|false|||process
Finding|Functional Concept|Impression|7212,7219|false|false|false|C4521054|Process (qualifier value)|process
Phenomenon|Phenomenon or Process|Impression|7212,7219|false|false|false|C1522240|Process|process
Event|Event|Impression|7220,7227|false|false|false|||causing
Attribute|Clinical Attribute|Impression|7233,7243|false|false|false|C0550215||appearance
Event|Event|Impression|7233,7243|false|false|false|||appearance
Procedure|Health Care Activity|Impression|7233,7243|false|false|false|C2051406|patient appearance regarding mental status exam|appearance
Event|Event|Impression|7247,7251|false|false|false|||felt
Event|Event|Impression|7257,7263|false|false|false|||likely
Finding|Finding|Impression|7257,7263|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Impression|7257,7263|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Functional Concept|Impression|7280,7292|false|false|false|C0333348|Inflammatory|inflammatory
Event|Event|Impression|7293,7302|false|false|false|||stranding
Event|Event|Impression|7314,7325|false|false|false|||colonoscopy
Procedure|Diagnostic Procedure|Impression|7314,7325|false|false|true|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Procedure|Health Care Activity|Impression|7314,7325|false|false|true|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Event|Event|Impression|7339,7349|false|false|false|||evaluation
Finding|Idea or Concept|Impression|7339,7349|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|Impression|7339,7349|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Anatomy|Body Part, Organ, or Organ Component|Impression|7363,7371|true|false|false|C0003617;C4037994|Abdomen+Pelvis>Appendix;Appendix|appendix
Disorder|Neoplastic Process|Impression|7363,7371|true|false|false|C0348899;C0496779;C0496860|Benign neoplasm of appendix;Malignant neoplasm of appendix;Neoplasm of uncertain or unknown behavior of appendix|appendix
Event|Event|Impression|7363,7371|true|false|false|||appendix
Finding|Intellectual Product|Impression|7363,7371|true|false|false|C1552860|appendix - HTML link|appendix
Procedure|Therapeutic or Preventive Procedure|Impression|7363,7371|true|false|false|C0869813|Procedure on appendix|appendix
Event|Event|Impression|7376,7381|true|false|false|||signs
Finding|Finding|Impression|7376,7381|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|Impression|7376,7381|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Event|Event|Impression|7385,7397|true|false|false|||inflammation
Finding|Pathologic Function|Impression|7385,7397|true|false|false|C0021368|Inflammation|inflammation
Finding|Gene or Genome|Impression|7415,7420|true|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Anatomy|Body Part, Organ, or Organ Component|Impression|7415,7426|true|false|false|C0021851|Large Intestine|large bowel
Finding|Pathologic Function|Impression|7415,7438|true|false|false|C0460048|Large bowel obstruction|large bowel obstruction
Anatomy|Body Part, Organ, or Organ Component|Impression|7421,7426|true|false|false|C0021853|Intestines|bowel
Disorder|Disease or Syndrome|Impression|7421,7438|true|false|false|C0021843|Intestinal Obstruction|bowel obstruction
Event|Event|Impression|7427,7438|true|false|false|||obstruction
Finding|Finding|Impression|7427,7438|true|false|false|C0028778|Obstruction|obstruction
Event|Event|Impression|7454,7464|false|false|false|||thickening
Finding|Finding|Impression|7454,7464|false|false|false|C0205400|Thickened|thickening
Anatomy|Body Part, Organ, or Organ Component|Impression|7468,7476|false|false|false|C0013303|Duodenum|duodenum
Disorder|Neoplastic Process|Impression|7468,7476|false|false|false|C0153426;C0496869|Benign neoplasm of duodenum;Malignant neoplasm of duodenum|duodenum
Finding|Finding|Impression|7477,7483|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Impression|7477,7483|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Drug|Organic Chemical|Impression|7484,7491|false|true|false|C0163712|Relate - vinyl resin|related
Event|Event|Impression|7484,7491|false|false|false|||related
Finding|Finding|Impression|7484,7491|false|true|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Finding|Functional Concept|Impression|7484,7491|false|true|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Event|Event|Impression|7496,7511|false|false|false|||underdistention
Event|Event|Impression|7516,7527|false|false|false|||Colonoscopy
Procedure|Diagnostic Procedure|Impression|7516,7527|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|Colonoscopy
Procedure|Health Care Activity|Impression|7516,7527|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|Colonoscopy
Anatomy|Body Space or Junction|Findings|7546,7551|false|false|false|C0524461|Structure of lumen of body system|Lumen
Event|Event|Findings|7553,7561|false|false|false|||Evidence
Finding|Idea or Concept|Findings|7553,7561|false|false|false|C3887511|Evidence|Evidence
Finding|Functional Concept|Findings|7553,7564|false|false|false|C0332120|Evidence of (contextual qualifier)|Evidence of
Drug|Amino Acid, Peptide, or Protein|Findings|7576,7579|false|false|false|C0082420|Endoglin, human|end
Drug|Immunologic Factor|Findings|7576,7579|false|false|false|C0082420|Endoglin, human|end
Event|Event|Findings|7576,7579|false|false|false|||end
Finding|Functional Concept|Findings|7576,7579|false|false|false|C1366583;C1561490;C1704837|ENG gene;ENG wt Allele;end - ActRelationshipCheckpoint|end
Finding|Gene or Genome|Findings|7576,7579|false|false|false|C1366583;C1561490;C1704837|ENG gene;ENG wt Allele;end - ActRelationshipCheckpoint|end
Drug|Amino Acid, Peptide, or Protein|Findings|7583,7586|false|false|false|C0082420|Endoglin, human|end
Drug|Immunologic Factor|Findings|7583,7586|false|false|false|C0082420|Endoglin, human|end
Event|Event|Findings|7583,7586|false|false|false|||end
Finding|Functional Concept|Findings|7583,7586|false|false|false|C1366583;C1561490;C1704837|ENG gene;ENG wt Allele;end - ActRelationshipCheckpoint|end
Finding|Gene or Genome|Findings|7583,7586|false|false|false|C1366583;C1561490;C1704837|ENG gene;ENG wt Allele;end - ActRelationshipCheckpoint|end
Anatomy|Body Space or Junction|Findings|7592,7603|false|false|false|C0500470|Anatomical anastomosis|anastomosis
Disorder|Acquired Abnormality|Findings|7592,7603|false|false|false|C0332853|Anastomosis|anastomosis
Event|Event|Findings|7592,7603|false|false|false|||anastomosis
Procedure|Therapeutic or Preventive Procedure|Findings|7592,7603|false|false|false|C0677554||anastomosis
Event|Event|Findings|7608,7612|false|false|false|||seen
Anatomy|Body Part, Organ, or Organ Component|Findings|7620,7627|false|false|false|C0227391|Sigmoid colon|sigmoid
Anatomy|Body Part, Organ, or Organ Component|Findings|7620,7633|false|false|false|C0227391|Sigmoid colon|sigmoid colon
Disorder|Neoplastic Process|Findings|7620,7633|false|false|false|C0153436;C0496864|Benign neoplasm of sigmoid colon;Malignant neoplasm of sigmoid colon|sigmoid colon
Anatomy|Body Part, Organ, or Organ Component|Findings|7628,7633|false|false|false|C0009368;C4071907|Abdomen+Pelvis>Colon;Colon structure (body structure)|colon
Disorder|Disease or Syndrome|Findings|7628,7633|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Disorder|Neoplastic Process|Findings|7628,7633|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Finding|Finding|Findings|7628,7633|false|false|false|C0750873|COLON PROBLEM|colon
Disorder|Anatomical Abnormality|Findings|7638,7648|false|false|false|C0333056|protrusion|Protruding
Event|Event|Findings|7638,7648|false|false|false|||Protruding
Finding|Finding|Findings|7649,7656|false|false|false|C0221198|Lesion|Lesions
Finding|Pathologic Function|Findings|7659,7668|false|false|false|C0041582;C3887532|Ulcer;Ulceration|ulcerated
Event|Event|Findings|7674,7678|false|false|false|||mass
Finding|Finding|Findings|7674,7678|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|Findings|7674,7678|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|Findings|7674,7678|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Event|Event|Findings|7682,7691|false|false|false|||malignant
Attribute|Clinical Attribute|Findings|7693,7703|false|false|false|C0550215||appearance
Event|Event|Findings|7693,7703|false|false|false|||appearance
Procedure|Health Care Activity|Findings|7693,7703|false|false|false|C2051406|patient appearance regarding mental status exam|appearance
Event|Event|Findings|7708,7713|false|false|false|||found
Anatomy|Body Part, Organ, or Organ Component|Findings|7721,7726|false|false|false|C0007531|Cecum|cecum
Disorder|Neoplastic Process|Findings|7721,7726|false|false|false|C0153437;C0496859|Benign neoplasm of cecum;Malignant neoplasm of cecum|cecum
Finding|Conceptual Entity|Findings|7732,7737|false|false|false|C1710028|Scope|scope
Event|Event|Findings|7738,7747|false|false|false|||traversed
Event|Event|Findings|7753,7759|false|false|false|||lesion
Finding|Finding|Findings|7753,7759|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|Findings|7753,7759|false|false|false|C0221198;C1546698|Lesion|lesion
Disorder|Disease or Syndrome|Findings|7761,7765|false|false|false|C0009443;C0024117|Chronic Obstructive Airway Disease;Common Cold|Cold
Drug|Organic Chemical|Findings|7761,7765|false|false|false|C0719425|Cold brand of chlorpheniramine-phenylpropanolamine|Cold
Drug|Pharmacologic Substance|Findings|7761,7765|false|false|false|C0719425|Cold brand of chlorpheniramine-phenylpropanolamine|Cold
Event|Event|Findings|7761,7765|false|false|false|||Cold
Finding|Organism Function|Findings|7761,7765|false|false|false|C0234192|Cold Sensation|Cold
Phenomenon|Natural Phenomenon or Process|Findings|7761,7765|false|false|false|C0009264|Cold Temperature|Cold
Procedure|Therapeutic or Preventive Procedure|Findings|7761,7765|false|false|false|C0010412|Cold Therapy|Cold
Event|Event|Findings|7774,7782|false|false|false|||biopsies
Procedure|Diagnostic Procedure|Findings|7774,7782|false|false|false|C0005558|Biopsy|biopsies
Event|Event|Findings|7802,7811|false|false|false|||histology
Finding|Functional Concept|Findings|7802,7811|false|false|false|C4048239;C4321399|Histology aspects;PATH.HISTO|histology
Finding|Intellectual Product|Findings|7802,7811|false|false|false|C4048239;C4321399|Histology aspects;PATH.HISTO|histology
Procedure|Laboratory Procedure|Findings|7802,7811|false|false|false|C0344441|Histologic test|histology
Anatomy|Body Part, Organ, or Organ Component|Findings|7820,7825|false|false|false|C0007531|Cecum|cecum
Disorder|Neoplastic Process|Findings|7820,7825|false|false|false|C0153437;C0496859|Benign neoplasm of cecum;Malignant neoplasm of cecum|cecum
Finding|Finding|Findings|7840,7847|false|false|false|C0221198|Lesion|Lesions
Disorder|Anatomical Abnormality|Findings|7848,7868|false|false|false|C1265782|Multiple diverticula|Multiple diverticula
Finding|Finding|Findings|7848,7868|false|false|false|C2238327||Multiple diverticula
Disorder|Anatomical Abnormality|Findings|7857,7868|false|false|false|C0012817|Diverticulum|diverticula
Event|Event|Findings|7857,7868|false|false|false|||diverticula
Event|Event|Findings|7880,7888|false|false|false|||openings
Event|Event|Findings|7895,7899|false|false|false|||seen
Finding|Functional Concept|Findings|7907,7917|false|false|false|C1547177|Sequencing - Descending|descending
Anatomy|Body Part, Organ, or Organ Component|Findings|7907,7923|false|false|false|C0227389|Descending colon|descending colon
Disorder|Neoplastic Process|Findings|7907,7923|false|false|false|C0153435;C0496863|Benign neoplasm of descending colon;Malignant neoplasm of descending colon|descending colon
Anatomy|Body Part, Organ, or Organ Component|Findings|7918,7923|false|false|false|C0009368;C4071907|Abdomen+Pelvis>Colon;Colon structure (body structure)|colon
Disorder|Disease or Syndrome|Findings|7918,7923|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Disorder|Neoplastic Process|Findings|7918,7923|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Event|Event|Findings|7918,7923|false|false|false|||colon
Finding|Finding|Findings|7918,7923|false|false|false|C0750873|COLON PROBLEM|colon
Event|Event|Findings|7927,7937|false|false|false|||Impression
Finding|Intellectual Product|Findings|7927,7937|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|Impression
Finding|Mental Process|Findings|7927,7937|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|Impression
Event|Event|Findings|7939,7943|false|false|false|||Mass
Finding|Finding|Findings|7939,7943|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|Mass
Finding|Gene or Genome|Findings|7939,7943|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|Mass
Finding|Intellectual Product|Findings|7939,7943|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|Mass
Anatomy|Body Part, Organ, or Organ Component|Findings|7951,7956|false|false|false|C0007531|Cecum|cecum
Disorder|Neoplastic Process|Findings|7951,7956|false|false|false|C0153437;C0496859|Benign neoplasm of cecum;Malignant neoplasm of cecum|cecum
Event|Event|Findings|7958,7964|false|false|false|||biopsy
Finding|Finding|Findings|7958,7964|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Finding|Intellectual Product|Findings|7958,7964|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Procedure|Diagnostic Procedure|Findings|7958,7964|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Procedure|Health Care Activity|Findings|7958,7964|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Disorder|Disease or Syndrome|Findings|7966,7980|false|false|false|C1510475|Diverticulosis|Diverticulosis
Event|Event|Findings|7966,7980|false|false|false|||Diverticulosis
Finding|Functional Concept|Findings|7988,7998|false|false|false|C1547177|Sequencing - Descending|descending
Anatomy|Body Part, Organ, or Organ Component|Findings|7988,8004|false|false|false|C0227389|Descending colon|descending colon
Disorder|Neoplastic Process|Findings|7988,8004|false|false|false|C0153435;C0496863|Benign neoplasm of descending colon;Malignant neoplasm of descending colon|descending colon
Anatomy|Body Part, Organ, or Organ Component|Findings|7999,8004|false|false|false|C0009368;C4071907|Abdomen+Pelvis>Colon;Colon structure (body structure)|colon
Disorder|Disease or Syndrome|Findings|7999,8004|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Disorder|Neoplastic Process|Findings|7999,8004|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Event|Event|Findings|7999,8004|false|false|false|||colon
Finding|Finding|Findings|7999,8004|false|false|false|C0750873|COLON PROBLEM|colon
Drug|Amino Acid, Peptide, or Protein|Findings|8014,8017|false|false|false|C0082420|Endoglin, human|end
Drug|Immunologic Factor|Findings|8014,8017|false|false|false|C0082420|Endoglin, human|end
Event|Event|Findings|8014,8017|false|false|false|||end
Finding|Functional Concept|Findings|8014,8017|false|false|false|C1366583;C1561490;C1704837|ENG gene;ENG wt Allele;end - ActRelationshipCheckpoint|end
Finding|Gene or Genome|Findings|8014,8017|false|false|false|C1366583;C1561490;C1704837|ENG gene;ENG wt Allele;end - ActRelationshipCheckpoint|end
Drug|Amino Acid, Peptide, or Protein|Findings|8021,8024|false|false|false|C0082420|Endoglin, human|end
Drug|Immunologic Factor|Findings|8021,8024|false|false|false|C0082420|Endoglin, human|end
Event|Event|Findings|8021,8024|false|false|false|||end
Finding|Functional Concept|Findings|8021,8024|false|false|false|C1366583;C1561490;C1704837|ENG gene;ENG wt Allele;end - ActRelationshipCheckpoint|end
Finding|Gene or Genome|Findings|8021,8024|false|false|false|C1366583;C1561490;C1704837|ENG gene;ENG wt Allele;end - ActRelationshipCheckpoint|end
Anatomy|Body Space or Junction|Findings|8029,8040|false|false|false|C0500470|Anatomical anastomosis|anastomosis
Disorder|Acquired Abnormality|Findings|8029,8040|false|false|false|C0332853|Anastomosis|anastomosis
Event|Event|Findings|8029,8040|false|false|false|||anastomosis
Procedure|Therapeutic or Preventive Procedure|Findings|8029,8040|false|false|false|C0677554||anastomosis
Anatomy|Body Part, Organ, or Organ Component|Findings|8048,8055|false|false|false|C0227391|Sigmoid colon|sigmoid
Anatomy|Body Part, Organ, or Organ Component|Findings|8057,8062|false|false|false|C0009368;C4071907|Abdomen+Pelvis>Colon;Colon structure (body structure)|colon
Disorder|Disease or Syndrome|Findings|8057,8062|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Disorder|Neoplastic Process|Findings|8057,8062|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Event|Event|Findings|8057,8062|false|false|false|||colon
Finding|Finding|Findings|8057,8062|false|false|false|C0750873|COLON PROBLEM|colon
Event|Event|Findings|8080,8091|false|false|false|||colonoscopy
Procedure|Diagnostic Procedure|Findings|8080,8091|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Procedure|Health Care Activity|Findings|8080,8091|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Anatomy|Body Part, Organ, or Organ Component|Findings|8095,8100|false|false|false|C0007531|Cecum|cecum
Disorder|Neoplastic Process|Findings|8095,8100|false|false|false|C0153437;C0496859|Benign neoplasm of cecum;Malignant neoplasm of cecum|cecum
Anatomy|Body Location or Region|Findings|8105,8119|false|false|false|C0227327|Distal part of ileum|terminal ileum
Anatomy|Body Part, Organ, or Organ Component|Findings|8114,8119|false|false|false|C0020885|ileum|ileum
Disorder|Neoplastic Process|Findings|8114,8119|false|false|false|C0153428|Malignant neoplasm of ileum|ileum
Event|Event|Findings|8123,8132|false|false|false|||PATHOLOGY
Finding|Functional Concept|Findings|8123,8132|false|false|false|C0205469;C0677042|Pathological aspects;Pathology processes|PATHOLOGY
Finding|Pathologic Function|Findings|8123,8132|false|false|false|C0205469;C0677042|Pathological aspects;Pathology processes|PATHOLOGY
Procedure|Laboratory Procedure|Findings|8123,8132|false|false|false|C0919386|Pathology procedure|PATHOLOGY
Anatomy|Body Part, Organ, or Organ Component|Diagnosis|8147,8152|false|false|false|C0007531|Cecum|Cecal
Finding|Finding|Diagnosis|8147,8157|false|false|false|C3670817|Cecal mass|Cecal mass
Event|Event|Diagnosis|8153,8157|false|false|false|||mass
Finding|Finding|Diagnosis|8153,8157|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|Diagnosis|8153,8157|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|Diagnosis|8153,8157|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Anatomy|Tissue|Diagnosis|8160,8167|false|false|false|C0026724|Mucous Membrane|mucosal
Event|Event|Diagnosis|8168,8176|false|false|false|||biopsies
Procedure|Diagnostic Procedure|Diagnosis|8168,8176|false|false|false|C0005558|Biopsy|biopsies
Anatomy|Body Part, Organ, or Organ Component|Diagnosis|8179,8186|false|false|false|C0009368|Colon structure (body structure)|Colonic
Anatomy|Body Part, Organ, or Organ Component|Diagnosis|8179,8193|false|false|false|C0227349|Colonic mucous membrane|Colonic mucosa
Anatomy|Tissue|Diagnosis|8187,8193|false|false|false|C0026724|Mucous Membrane|mucosa
Finding|Intellectual Product|Diagnosis|8187,8193|false|false|false|C1561514||mucosa
Finding|Functional Concept|Diagnosis|8205,8213|false|false|false|C0475224|Ischemic|ischemic
Finding|Finding|Diagnosis|8205,8220|false|false|false|C2826576|Ischemic Change|ischemic change
Event|Event|Diagnosis|8214,8220|false|false|false|||change
Finding|Functional Concept|Diagnosis|8214,8220|false|false|false|C0392747|Changing|change
Procedure|Therapeutic or Preventive Procedure|Diagnosis|8214,8220|false|false|false|C4319952|Change - procedure|change
Event|Event|Diagnosis|8225,8233|false|false|false|||abundant
Event|Event|Diagnosis|8246,8256|false|false|false|||ulceration
Finding|Pathologic Function|Diagnosis|8246,8256|false|false|false|C0041582;C3887532|Ulcer;Ulceration|ulceration
Event|Event|Diagnosis|8258,8265|false|false|false|||exudate
Finding|Body Substance|Diagnosis|8258,8265|false|false|false|C0015388;C1546629|Exudate|exudate
Finding|Intellectual Product|Diagnosis|8258,8265|false|false|false|C0015388;C1546629|Exudate|exudate
Event|Event|Diagnosis|8271,8282|false|false|false|||granulation
Finding|Finding|Diagnosis|8271,8282|false|false|false|C0518864|Granulation finding|granulation
Procedure|Laboratory Procedure|Diagnosis|8271,8282|false|false|false|C4281706|Granulation procedure|granulation
Anatomy|Tissue|Diagnosis|8271,8289|false|false|false|C0018180|Granulation Tissue|granulation tissue
Finding|Finding|Diagnosis|8271,8289|false|false|false|C3806379|Granulation of tissue|granulation tissue
Anatomy|Tissue|Diagnosis|8283,8289|false|false|false|C0040300|Body tissue|tissue
Finding|Intellectual Product|Diagnosis|8283,8289|false|false|false|C1547928|Tissue Specimen Code|tissue
Event|Event|Diagnosis|8291,8300|false|false|false|||formation
Finding|Functional Concept|Diagnosis|8291,8300|false|false|false|C1522492|Formation|formation
Phenomenon|Biologic Function|Diagnosis|8291,8300|false|false|false|C0220781|Anabolism|formation
Disorder|Neoplastic Process|Diagnosis|8305,8314|true|false|false|C0007097|Carcinoma|carcinoma
Event|Event|Diagnosis|8305,8314|true|false|false|||carcinoma
Disorder|Congenital Abnormality|Diagnosis|8318,8327|true|false|false|C0334044|Dysplasia|dysplasia
Event|Event|Diagnosis|8318,8327|true|false|false|||dysplasia
Event|Event|Diagnosis|8353,8359|false|false|false|||levels
Event|Event|Diagnosis|8364,8372|false|false|false|||examined
Finding|Body Substance|Hospital Course|8407,8414|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|8407,8414|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|8407,8414|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|8424,8428|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|Hospital Course|8424,8428|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Event|Event|Hospital Course|8429,8432|false|false|false|||old
Event|Event|Hospital Course|8445,8452|false|false|false|||history
Finding|Conceptual Entity|Hospital Course|8445,8452|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|8445,8452|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Hospital Course|8445,8452|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Idea or Concept|Hospital Course|8453,8464|false|false|false|C0750502|Significant|significant
Event|Event|Hospital Course|8465,8468|false|false|false|||for
Disorder|Disease or Syndrome|Hospital Course|8470,8484|false|false|false|C0012813|Diverticulitis|diverticulitis
Event|Event|Hospital Course|8470,8484|false|false|false|||diverticulitis
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8489,8496|false|false|false|C0227391|Sigmoid colon|sigmoid
Event|Event|Hospital Course|8497,8506|false|false|false|||resection
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8497,8506|false|false|false|C0015252;C0728940|Excision;removal technique|resection
Event|Event|Hospital Course|8519,8528|false|false|false|||presented
Anatomy|Body Location or Region|Hospital Course|8535,8544|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|Hospital Course|8535,8549|false|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|Hospital Course|8545,8549|false|false|false|C2598155||pain
Event|Event|Hospital Course|8545,8549|false|false|false|||pain
Finding|Functional Concept|Hospital Course|8545,8549|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|8545,8549|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|8558,8563|false|false|false|||found
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8572,8577|false|false|false|C0007531|Cecum|cecal
Finding|Finding|Hospital Course|8572,8582|false|false|false|C3670817|Cecal mass|cecal mass
Event|Event|Hospital Course|8578,8582|false|false|false|||mass
Finding|Finding|Hospital Course|8578,8582|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|Hospital Course|8578,8582|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|Hospital Course|8578,8582|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Anatomy|Body Location or Region|Hospital Course|8592,8601|false|false|false|C0000726|Abdomen|Abdominal
Finding|Sign or Symptom|Hospital Course|8592,8606|false|false|false|C0000737|Abdominal Pain|Abdominal pain
Attribute|Clinical Attribute|Hospital Course|8602,8606|false|false|false|C2598155||pain
Event|Event|Hospital Course|8602,8606|false|false|false|||pain
Finding|Functional Concept|Hospital Course|8602,8606|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|8602,8606|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Idea or Concept|Hospital Course|8612,8623|false|false|false|C0750501|most likely|most likely
Finding|Finding|Hospital Course|8617,8623|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Hospital Course|8617,8623|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Drug|Organic Chemical|Hospital Course|8624,8631|false|false|false|C0163712|Relate - vinyl resin|related
Event|Event|Hospital Course|8624,8631|false|false|false|||related
Finding|Finding|Hospital Course|8624,8631|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Finding|Functional Concept|Hospital Course|8624,8631|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8647,8654|false|false|false|C0205065|Ovarian|ovarian
Disorder|Anatomical Abnormality|Hospital Course|8656,8660|false|false|false|C0010709|Cyst|cyst
Event|Event|Hospital Course|8656,8660|false|false|false|||cyst
Finding|Body Substance|Hospital Course|8656,8660|false|false|false|C1546594;C1550626|SpecimenType - Cyst|cyst
Finding|Intellectual Product|Hospital Course|8656,8660|false|false|false|C1546594;C1550626|SpecimenType - Cyst|cyst
Finding|Body Substance|Hospital Course|8674,8681|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|8674,8681|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|8674,8681|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|8686,8697|true|false|false|C0750502|Significant|significant
Attribute|Clinical Attribute|Hospital Course|8698,8702|true|false|false|C2598155||pain
Event|Event|Hospital Course|8698,8702|true|false|false|||pain
Finding|Functional Concept|Hospital Course|8698,8702|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|8698,8702|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|8717,8725|true|false|false|||relieved
Drug|Organic Chemical|Hospital Course|8731,8739|true|false|false|C0728755|Dilaudid|dilaudid
Drug|Pharmacologic Substance|Hospital Course|8731,8739|true|false|false|C0728755|Dilaudid|dilaudid
Event|Event|Hospital Course|8731,8739|true|false|false|||dilaudid
Event|Event|Hospital Course|8760,8766|false|false|false|||course
Attribute|Clinical Attribute|Hospital Course|8788,8792|false|false|false|C2598155||pain
Event|Event|Hospital Course|8788,8792|false|false|false|||pain
Finding|Functional Concept|Hospital Course|8788,8792|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|8788,8792|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|8793,8801|false|false|false|||resolved
Finding|Finding|Hospital Course|8809,8812|false|false|false|C5939094|Own|own
Event|Event|Hospital Course|8831,8839|true|false|false|||required
Attribute|Clinical Attribute|Hospital Course|8845,8849|true|false|false|C2598155||pain
Event|Event|Hospital Course|8845,8849|true|false|false|||pain
Finding|Functional Concept|Hospital Course|8845,8849|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|8845,8849|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|Hospital Course|8850,8861|true|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Hospital Course|8850,8861|true|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Hospital Course|8850,8861|true|false|false|||medications
Finding|Intellectual Product|Hospital Course|8850,8861|true|false|false|C4284232|Medications|medications
Event|Event|Hospital Course|8864,8873|true|false|false|||Bloodwork
Event|Event|Hospital Course|8878,8885|true|false|false|||imaging
Finding|Finding|Hospital Course|8878,8885|true|false|false|C0740845|Imaging problem|imaging
Procedure|Diagnostic Procedure|Hospital Course|8878,8885|true|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|imaging
Event|Event|Hospital Course|8895,8905|true|false|false|||suggestive
Finding|Functional Concept|Hospital Course|8895,8905|true|false|false|C0332299|Suggestive of|suggestive
Finding|Functional Concept|Hospital Course|8895,8908|true|false|false|C0332299|Suggestive of|suggestive of
Finding|Functional Concept|Hospital Course|8914,8929|true|false|false|C1512911|Intraabdominal Route of Administration|intra-abdominal
Disorder|Disease or Syndrome|Hospital Course|8914,8939|true|false|false|C1112209|Abdominal Infection|intra-abdominal infection
Disorder|Disease or Syndrome|Hospital Course|8930,8939|true|false|false|C0009450|Communicable Diseases|infection
Event|Event|Hospital Course|8930,8939|true|false|false|||infection
Finding|Pathologic Function|Hospital Course|8930,8939|true|false|false|C3714514|Infection|infection
Finding|Body Substance|Hospital Course|8946,8953|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|8946,8953|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|8946,8953|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|8958,8965|false|false|false|||advised
Event|Event|Hospital Course|8970,8976|false|false|false|||follow
Event|Event|Hospital Course|9002,9011|false|false|false|||regarding
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9016,9023|false|false|false|C0205065|Ovarian|ovarian
Disorder|Disease or Syndrome|Hospital Course|9016,9028|false|false|false|C0029927|Ovarian Cysts|ovarian cyst
Disorder|Anatomical Abnormality|Hospital Course|9024,9028|false|false|false|C0010709|Cyst|cyst
Event|Event|Hospital Course|9024,9028|false|false|false|||cyst
Finding|Body Substance|Hospital Course|9024,9028|false|false|false|C1546594;C1550626|SpecimenType - Cyst|cyst
Finding|Intellectual Product|Hospital Course|9024,9028|false|false|false|C1546594;C1550626|SpecimenType - Cyst|cyst
Event|Event|Hospital Course|9039,9043|false|false|false|||need
Finding|Functional Concept|Hospital Course|9039,9043|false|false|false|C0686904|Patient need for (contextual qualifier)|need
Finding|Functional Concept|Hospital Course|9039,9047|false|false|false|C0686904|Patient need for (contextual qualifier)|need for
Finding|Idea or Concept|Hospital Course|9048,9057|false|false|false|C0549178|Continuous|continued
Event|Event|Hospital Course|9058,9065|false|false|false|||therapy
Finding|Finding|Hospital Course|9058,9065|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|Hospital Course|9058,9065|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9058,9065|false|false|false|C0087111|Therapeutic procedure|therapy
Finding|Finding|Hospital Course|9071,9074|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|Hospital Course|9071,9074|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Drug|Pharmacologic Substance|Hospital Course|9071,9098|false|false|false|C0086736|Oral Contraceptives, Low-Dose|low dose oral contraceptive
Event|Event|Hospital Course|9075,9079|false|false|false|||dose
Anatomy|Body Space or Junction|Hospital Course|9080,9084|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|9080,9084|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|9080,9084|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|9080,9084|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Drug|Pharmacologic Substance|Hospital Course|9080,9098|false|false|false|C0009905|Contraceptives, Oral|oral contraceptive
Finding|Finding|Hospital Course|9080,9098|false|false|false|C0029151|Uses oral contraception (finding)|oral contraceptive
Drug|Pharmacologic Substance|Hospital Course|9085,9098|false|false|false|C0009871|Contraceptive Agents|contraceptive
Event|Event|Hospital Course|9085,9098|false|false|false|||contraceptive
Finding|Finding|Hospital Course|9085,9098|false|false|false|C0344225|Encounter due to presence of intrauterine contraceptive device|contraceptive
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9110,9115|false|false|false|C0007531|Cecum|Cecal
Finding|Finding|Hospital Course|9110,9120|false|false|false|C3670817|Cecal mass|Cecal Mass
Event|Event|Hospital Course|9116,9120|false|false|false|||Mass
Finding|Finding|Hospital Course|9116,9120|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|Mass
Finding|Gene or Genome|Hospital Course|9116,9120|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|Mass
Finding|Intellectual Product|Hospital Course|9116,9120|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|Mass
Event|Event|Hospital Course|9133,9139|false|false|false|||workup
Finding|Body Substance|Hospital Course|9148,9155|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|9148,9155|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|9148,9155|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Anatomy|Body Location or Region|Hospital Course|9158,9167|false|false|false|C0000726|Abdomen|abdominal
Attribute|Clinical Attribute|Hospital Course|9169,9173|false|false|false|C2598155||pain
Event|Event|Hospital Course|9169,9173|false|false|false|||pain
Finding|Functional Concept|Hospital Course|9169,9173|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|9169,9173|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|9177,9179|false|false|false|||CT
Anatomy|Body Location or Region|Hospital Course|9187,9194|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|abdomen
Disorder|Neoplastic Process|Hospital Course|9187,9194|false|false|false|C0153662|Malignant neoplasm of abdomen|abdomen
Finding|Finding|Hospital Course|9187,9194|false|false|false|C0941288|Abdomen problem|abdomen
Anatomy|Body Location or Region|Hospital Course|9187,9198|false|false|false|C0000726|Abdomen|abdomen and
Anatomy|Body Location or Region|Hospital Course|9187,9205|false|false|false|C1508499|Abdominopelvic structure|abdomen and pelvis
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9199,9205|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Anatomy|Body Space or Junction|Hospital Course|9199,9205|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Disorder|Neoplastic Process|Hospital Course|9199,9205|false|false|false|C0153663|Malignant neoplasm of pelvis|pelvis
Finding|Finding|Hospital Course|9199,9205|false|false|false|C0812455|Pelvis problem|pelvis
Event|Event|Hospital Course|9206,9214|false|false|false|||revealed
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9222,9227|false|false|false|C0007531|Cecum|cecal
Finding|Finding|Hospital Course|9222,9232|false|false|false|C3670817|Cecal mass|cecal mass
Event|Event|Hospital Course|9228,9232|false|false|false|||mass
Finding|Finding|Hospital Course|9228,9232|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|Hospital Course|9228,9232|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|Hospital Course|9228,9232|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Disorder|Neoplastic Process|Hospital Course|9249,9259|false|false|false|C0006826;C1306459|Malignant Neoplasms;Primary malignant neoplasm|malignancy
Event|Event|Hospital Course|9249,9259|false|false|false|||malignancy
Event|Event|Hospital Course|9274,9289|false|false|false|||hospitalization
Procedure|Health Care Activity|Hospital Course|9274,9289|false|false|false|C0019993|Hospitalization|hospitalization
Event|Event|Hospital Course|9305,9316|false|false|false|||colonoscopy
Procedure|Diagnostic Procedure|Hospital Course|9305,9316|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Procedure|Health Care Activity|Hospital Course|9305,9316|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Procedure|Diagnostic Procedure|Hospital Course|9305,9328|false|false|false|C0372088;C0810150|Colonoscopy and Biopsy;Colonoscopy through stoma; with biopsy, single or multiple|colonoscopy with biopsy
Event|Event|Hospital Course|9322,9328|false|false|false|||biopsy
Finding|Finding|Hospital Course|9322,9328|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Finding|Intellectual Product|Hospital Course|9322,9328|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Procedure|Diagnostic Procedure|Hospital Course|9322,9328|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Procedure|Health Care Activity|Hospital Course|9322,9328|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Event|Event|Hospital Course|9336,9340|false|false|false|||mass
Finding|Finding|Hospital Course|9336,9340|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|Hospital Course|9336,9340|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|Hospital Course|9336,9340|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Event|Event|Hospital Course|9352,9362|false|false|false|||instructed
Event|Event|Hospital Course|9366,9372|false|false|false|||follow
Finding|Classification|Hospital Course|9385,9395|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|9385,9395|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|Hospital Course|9396,9414|false|false|false|||gastroenterologist
Event|Event|Hospital Course|9430,9437|false|false|false|||results
Event|Event|Hospital Course|9446,9452|false|false|false|||biopsy
Finding|Finding|Hospital Course|9446,9452|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Finding|Intellectual Product|Hospital Course|9446,9452|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Procedure|Diagnostic Procedure|Hospital Course|9446,9452|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Procedure|Health Care Activity|Hospital Course|9446,9452|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Finding|Intellectual Product|Hospital Course|9460,9464|false|false|false|C1561540|Transaction counts and value totals - week|week
Event|Event|Hospital Course|9471,9477|true|false|false|||biopsy
Finding|Finding|Hospital Course|9471,9477|true|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Finding|Intellectual Product|Hospital Course|9471,9477|true|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Procedure|Diagnostic Procedure|Hospital Course|9471,9477|true|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Procedure|Health Care Activity|Hospital Course|9471,9477|true|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Event|Event|Hospital Course|9483,9491|false|false|false|||negative
Finding|Classification|Hospital Course|9483,9491|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|9483,9491|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|9483,9491|false|false|false|C5237010|Expression Negative|negative
Finding|Finding|Hospital Course|9483,9495|false|false|false|C0205160|Negative|negative for
Disorder|Neoplastic Process|Hospital Course|9496,9506|true|false|false|C0006826;C1306459|Malignant Neoplasms;Primary malignant neoplasm|malignancy
Event|Event|Hospital Course|9496,9506|true|false|false|||malignancy
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9517,9524|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|Anxiety
Event|Event|Hospital Course|9517,9524|false|false|false|||Anxiety
Finding|Sign or Symptom|Hospital Course|9517,9524|false|false|false|C0860603|Anxiety symptoms|Anxiety
Event|Event|Hospital Course|9527,9534|false|false|false|||Patient
Finding|Body Substance|Hospital Course|9527,9534|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|9527,9534|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|9527,9534|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Hospital Course|9539,9548|false|false|false|||continued
Finding|Idea or Concept|Hospital Course|9552,9556|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|9552,9556|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|9552,9556|false|false|false|C1553498|home health encounter|home
Event|Event|Hospital Course|9557,9564|false|false|false|||regimen
Finding|Intellectual Product|Hospital Course|9557,9564|false|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9557,9564|false|false|false|C0040808|Treatment Protocols|regimen
Drug|Organic Chemical|Hospital Course|9568,9574|false|false|false|C0284660|Zoloft|zoloft
Drug|Pharmacologic Substance|Hospital Course|9568,9574|false|false|false|C0284660|Zoloft|zoloft
Drug|Organic Chemical|Hospital Course|9580,9586|false|false|false|C0699194|Ativan|ativan
Drug|Pharmacologic Substance|Hospital Course|9580,9586|false|false|false|C0699194|Ativan|ativan
Event|Event|Hospital Course|9580,9586|false|false|false|||ativan
Disorder|Disease or Syndrome|Hospital Course|9596,9600|false|false|false|C0017168|Gastroesophageal reflux disease|Gerd
Event|Event|Hospital Course|9596,9600|false|false|false|||Gerd
Finding|Body Substance|Hospital Course|9603,9610|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|9603,9610|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|9603,9610|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Hospital Course|9611,9620|false|false|false|||continued
Drug|Organic Chemical|Hospital Course|9624,9634|false|false|false|C0028978|omeprazole|omeprazole
Drug|Pharmacologic Substance|Hospital Course|9624,9634|false|false|false|C0028978|omeprazole|omeprazole
Event|Event|Hospital Course|9624,9634|false|false|false|||omeprazole
Drug|Organic Chemical|Hospital Course|9636,9642|false|false|false|C0592278|Zantac|zantac
Drug|Pharmacologic Substance|Hospital Course|9636,9642|false|false|false|C0592278|Zantac|zantac
Event|Event|Hospital Course|9636,9642|false|false|false|||zantac
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9643,9646|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9643,9646|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|9643,9646|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|9643,9646|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|9643,9646|false|false|false|C1332410|BID gene|BID
Finding|Classification|Hospital Course|9652,9662|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|9652,9662|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|Hospital Course|9663,9670|false|false|false|||regimen
Finding|Intellectual Product|Hospital Course|9663,9670|false|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9663,9670|false|false|false|C0040808|Treatment Protocols|regimen
Attribute|Clinical Attribute|Hospital Course|9677,9688|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|9677,9688|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|9677,9688|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|9677,9688|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|9677,9701|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|Hospital Course|9692,9701|false|false|false|||Admission
Procedure|Health Care Activity|Hospital Course|9692,9701|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Food|Hospital Course|9704,9708|false|false|false|C3257082;C4521129|Fish (substance);Fish extract|Fish
Drug|Organic Chemical|Hospital Course|9704,9708|false|false|false|C3257082;C4521129|Fish (substance);Fish extract|Fish
Event|Event|Hospital Course|9704,9708|false|false|false|||Fish
Finding|Gene or Genome|Hospital Course|9704,9708|false|false|false|C1822711;C3274826|SH3PXD2A gene;SH3PXD2A wt Allele|Fish
Procedure|Molecular Biology Research Technique|Hospital Course|9704,9708|false|false|false|C0162789|Fluorescent in Situ Hybridization|Fish
Drug|Organic Chemical|Hospital Course|9704,9712|false|false|false|C0016157|fish oils|Fish Oil
Drug|Pharmacologic Substance|Hospital Course|9704,9712|false|false|false|C0016157|fish oils|Fish Oil
Drug|Biomedical or Dental Material|Hospital Course|9709,9712|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|Oil
Drug|Food|Hospital Course|9709,9712|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|Oil
Drug|Organic Chemical|Hospital Course|9709,9712|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|Oil
Drug|Pharmacologic Substance|Hospital Course|9709,9712|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|Oil
Disorder|Congenital Abnormality|Hospital Course|9722,9725|false|false|false|C1855179|CATARACT, ANTERIOR POLAR|Cap
Drug|Biomedical or Dental Material|Hospital Course|9722,9725|false|false|false|C0006935|capsule (pharmacologic)|Cap
Event|Event|Hospital Course|9722,9725|false|false|false|||Cap
Finding|Gene or Genome|Hospital Course|9722,9725|false|false|false|C1416891;C1418551;C1419093;C1422073;C1422760;C2985259;C4522312|BRD4 gene;BRD4 wt Allele;CAP1 gene;HACD1 gene;LNPEP gene;SERPINB6 gene;SORBS1 gene|Cap
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9722,9725|false|false|false|C0278651;C0280547;C1879916|CAP Regimen;cisplatin/cyclophosphamide/doxorubicin protocol;cyclophosphamide/doxorubicin/prednisone protocol|Cap
Drug|Organic Chemical|Hospital Course|9729,9734|false|false|false|C0939679|Axert|Axert
Drug|Pharmacologic Substance|Hospital Course|9729,9734|false|false|false|C0939679|Axert|Axert
Drug|Biomedical or Dental Material|Hospital Course|9743,9746|false|false|false|C0039225|Tablet Dosage Form|Tab
Drug|Biomedical or Dental Material|Hospital Course|9751,9757|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Functional Concept|Hospital Course|9761,9769|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|9764,9769|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|9764,9769|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Event|Event|Hospital Course|9789,9795|false|false|false|||repeat
Finding|Idea or Concept|Hospital Course|9819,9822|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|9819,9822|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|Hospital Course|9826,9833|false|false|false|C1170371|Lexapro|Lexapro
Drug|Pharmacologic Substance|Hospital Course|9826,9833|false|false|false|C1170371|Lexapro|Lexapro
Drug|Biomedical or Dental Material|Hospital Course|9840,9843|false|false|false|C0039225|Tablet Dosage Form|Tab
Drug|Organic Chemical|Hospital Course|9853,9868|false|false|false|C0008318|cholecalciferol|Cholecalciferol
Drug|Pharmacologic Substance|Hospital Course|9853,9868|false|false|false|C0008318|cholecalciferol|Cholecalciferol
Drug|Vitamin|Hospital Course|9853,9868|false|false|false|C0008318|cholecalciferol|Cholecalciferol
Event|Event|Hospital Course|9853,9868|false|false|false|||Cholecalciferol
Drug|Organic Chemical|Hospital Course|9853,9881|false|false|false|C0008318|cholecalciferol|Cholecalciferol (Vitamin D3)
Drug|Pharmacologic Substance|Hospital Course|9853,9881|false|false|false|C0008318|cholecalciferol|Cholecalciferol (Vitamin D3)
Drug|Vitamin|Hospital Course|9853,9881|false|false|false|C0008318|cholecalciferol|Cholecalciferol (Vitamin D3)
Drug|Organic Chemical|Hospital Course|9870,9877|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|Hospital Course|9870,9877|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|Hospital Course|9870,9877|false|false|false|C0042890|Vitamins|Vitamin
Drug|Organic Chemical|Hospital Course|9870,9880|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|Vitamin D3
Drug|Pharmacologic Substance|Hospital Course|9870,9880|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|Vitamin D3
Drug|Vitamin|Hospital Course|9870,9880|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|Vitamin D3
Drug|Biomedical or Dental Material|Hospital Course|9893,9896|false|false|false|C0039225|Tablet Dosage Form|Tab
Event|Event|Hospital Course|9893,9896|false|false|false|||Tab
Drug|Organic Chemical|Hospital Course|9900,9909|false|false|false|C0024002|lorazepam|lorazepam
Drug|Pharmacologic Substance|Hospital Course|9900,9909|false|false|false|C0024002|lorazepam|lorazepam
Drug|Biomedical or Dental Material|Hospital Course|9917,9920|false|false|false|C0039225|Tablet Dosage Form|Tab
Finding|Gene or Genome|Hospital Course|9924,9927|false|false|false|C1422467|CIAO3 gene|prn
Drug|Organic Chemical|Hospital Course|9931,9941|false|false|false|C0028978|omeprazole|Omeprazole
Drug|Pharmacologic Substance|Hospital Course|9931,9941|false|false|false|C0028978|omeprazole|Omeprazole
Disorder|Congenital Abnormality|Hospital Course|9948,9951|false|false|false|C1855179|CATARACT, ANTERIOR POLAR|Cap
Drug|Biomedical or Dental Material|Hospital Course|9948,9951|false|false|false|C0006935|capsule (pharmacologic)|Cap
Event|Event|Hospital Course|9948,9951|false|false|false|||Cap
Finding|Gene or Genome|Hospital Course|9948,9951|false|false|false|C1416891;C1418551;C1419093;C1422073;C1422760;C2985259;C4522312|BRD4 gene;BRD4 wt Allele;CAP1 gene;HACD1 gene;LNPEP gene;SERPINB6 gene;SORBS1 gene|Cap
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9948,9951|false|false|false|C0278651;C0280547;C1879916|CAP Regimen;cisplatin/cyclophosphamide/doxorubicin protocol;cyclophosphamide/doxorubicin/prednisone protocol|Cap
Event|Event|Hospital Course|9961,9968|false|false|false|||Release
Finding|Functional Concept|Hospital Course|9961,9968|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|9961,9968|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9961,9968|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9969,9972|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9969,9972|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|9969,9972|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|9969,9972|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|9969,9972|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|9976,9984|false|false|false|C0040610|tramadol|tramadol
Drug|Pharmacologic Substance|Hospital Course|9976,9984|false|false|false|C0040610|tramadol|tramadol
Event|Event|Hospital Course|9976,9984|false|false|false|||tramadol
Procedure|Laboratory Procedure|Hospital Course|9976,9984|false|false|false|C1266765|Tramadol measurement (procedure)|tramadol
Drug|Biomedical or Dental Material|Hospital Course|9991,9994|false|false|false|C0039225|Tablet Dosage Form|Tab
Event|Event|Hospital Course|10018,10024|false|false|false|||needed
Attribute|Clinical Attribute|Hospital Course|10029,10033|false|false|false|C2598155||pain
Event|Event|Hospital Course|10029,10033|false|false|false|||pain
Finding|Functional Concept|Hospital Course|10029,10033|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|10029,10033|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|Hospital Course|10037,10046|false|false|false|C0030049|oxycodone|oxycodone
Drug|Pharmacologic Substance|Hospital Course|10037,10046|false|false|false|C0030049|oxycodone|oxycodone
Event|Event|Hospital Course|10037,10046|false|false|false|||oxycodone
Procedure|Laboratory Procedure|Hospital Course|10037,10046|false|false|false|C0524222|Oxycodone measurement|oxycodone
Drug|Biomedical or Dental Material|Hospital Course|10052,10055|false|false|false|C0039225|Tablet Dosage Form|Tab
Drug|Biomedical or Dental Material|Hospital Course|10062,10068|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|10062,10068|false|false|false|||Tablet
Finding|Functional Concept|Hospital Course|10072,10080|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|10075,10080|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|10075,10080|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Gene or Genome|Hospital Course|10085,10088|false|false|false|C1422467|CIAO3 gene|prn
Event|Event|Hospital Course|10092,10098|false|false|false|||needed
Attribute|Clinical Attribute|Hospital Course|10103,10107|false|false|false|C2598155||pain
Event|Event|Hospital Course|10103,10107|false|false|false|||pain
Finding|Functional Concept|Hospital Course|10103,10107|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|10103,10107|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|Hospital Course|10111,10123|false|false|false|C0301532|Multivitamin preparation|Multivitamin
Drug|Pharmacologic Substance|Hospital Course|10111,10123|false|false|false|C0301532|Multivitamin preparation|Multivitamin
Drug|Vitamin|Hospital Course|10111,10123|false|false|false|C0301532|Multivitamin preparation|Multivitamin
Disorder|Congenital Abnormality|Hospital Course|10124,10127|false|false|false|C1855179|CATARACT, ANTERIOR POLAR|Cap
Drug|Biomedical or Dental Material|Hospital Course|10124,10127|false|false|false|C0006935|capsule (pharmacologic)|Cap
Event|Event|Hospital Course|10124,10127|false|false|false|||Cap
Finding|Gene or Genome|Hospital Course|10124,10127|false|false|false|C1416891;C1418551;C1419093;C1422073;C1422760;C2985259;C4522312|BRD4 gene;BRD4 wt Allele;CAP1 gene;HACD1 gene;LNPEP gene;SERPINB6 gene;SORBS1 gene|Cap
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10124,10127|false|false|false|C0278651;C0280547;C1879916|CAP Regimen;cisplatin/cyclophosphamide/doxorubicin protocol;cyclophosphamide/doxorubicin/prednisone protocol|Cap
Drug|Organic Chemical|Hospital Course|10131,10137|false|false|false|C0592278|Zantac|Zantac
Drug|Pharmacologic Substance|Hospital Course|10131,10137|false|false|false|C0592278|Zantac|Zantac
Drug|Organic Chemical|Hospital Course|10131,10141|false|false|false|C0724451|Zantac 150|Zantac 150
Drug|Pharmacologic Substance|Hospital Course|10131,10141|false|false|false|C0724451|Zantac 150|Zantac 150
Disorder|Congenital Abnormality|Hospital Course|10145,10148|false|false|false|C1855179|CATARACT, ANTERIOR POLAR|Cap
Drug|Biomedical or Dental Material|Hospital Course|10145,10148|false|false|false|C0006935|capsule (pharmacologic)|Cap
Event|Event|Hospital Course|10145,10148|false|false|false|||Cap
Finding|Gene or Genome|Hospital Course|10145,10148|false|false|false|C1416891;C1418551;C1419093;C1422073;C1422760;C2985259;C4522312|BRD4 gene;BRD4 wt Allele;CAP1 gene;HACD1 gene;LNPEP gene;SERPINB6 gene;SORBS1 gene|Cap
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10145,10148|false|false|false|C0278651;C0280547;C1879916|CAP Regimen;cisplatin/cyclophosphamide/doxorubicin protocol;cyclophosphamide/doxorubicin/prednisone protocol|Cap
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10151,10158|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|10151,10158|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|10151,10158|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Finding|Functional Concept|Hospital Course|10162,10170|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|10165,10170|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|10165,10170|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Idea or Concept|Hospital Course|10179,10182|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|10179,10182|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|Hospital Course|10186,10197|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Hospital Course|10186,10197|false|false|false|C0082607|fluticasone|Fluticasone
Event|Event|Hospital Course|10186,10197|false|false|false|||Fluticasone
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10215,10220|false|false|false|C0028429||Nasal
Drug|Biomedical or Dental Material|Hospital Course|10215,10220|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Organic Chemical|Hospital Course|10215,10220|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Pharmacologic Substance|Hospital Course|10215,10220|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Finding|Finding|Hospital Course|10215,10220|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Finding|Functional Concept|Hospital Course|10215,10220|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Drug|Pharmacologic Substance|Hospital Course|10215,10226|false|false|false|C2608294|Nasal Spray brand of phenylephrine|Nasal Spray
Drug|Biomedical or Dental Material|Hospital Course|10221,10226|false|false|false|C1154182|Spray Dosage Form|Spray
Event|Activity|Hospital Course|10221,10226|false|false|false|C2003858|Spray (action)|Spray
Event|Event|Hospital Course|10221,10226|false|false|false|||Spray
Finding|Functional Concept|Hospital Course|10221,10226|false|false|false|C4521772|Spray (administration method)|Spray
Drug|Biomedical or Dental Material|Hospital Course|10228,10232|false|false|false|C0038960|Suspensions|Susp
Event|Event|Hospital Course|10228,10232|false|false|false|||Susp
Finding|Molecular Function|Hospital Course|10228,10232|false|false|false|C1150157|SUMO-specific protease activity|Susp
Disorder|Mental or Behavioral Dysfunction|Hospital Course|10237,10243|false|false|false|C0233601|Spraying behavior|sprays
Drug|Biomedical or Dental Material|Hospital Course|10237,10243|false|false|false|C1154182|Spray Dosage Form|sprays
Event|Event|Hospital Course|10237,10243|false|false|false|||sprays
Finding|Intellectual Product|Hospital Course|10268,10272|false|false|false|C1720594|Then - dosing instruction fragment|then
Drug|Biomedical or Dental Material|Hospital Course|10275,10280|false|false|false|C1154182|Spray Dosage Form|spray
Event|Activity|Hospital Course|10275,10280|false|false|false|C2003858|Spray (action)|spray
Event|Event|Hospital Course|10275,10280|false|false|false|||spray
Finding|Functional Concept|Hospital Course|10275,10280|false|false|false|C4521772|Spray (administration method)|spray
Drug|Biologically Active Substance|Hospital Course|10287,10294|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|Hospital Course|10287,10294|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|Hospital Course|10287,10294|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|Hospital Course|10287,10294|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|Hospital Course|10287,10294|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|Hospital Course|10287,10294|false|false|false|||Calcium
Finding|Physiologic Function|Hospital Course|10287,10294|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|Hospital Course|10287,10294|false|false|false|C0201925|Calcium measurement|Calcium
Drug|Organic Chemical|Hospital Course|10287,10302|false|false|false|C0108101|calcium citrate|Calcium Citrate
Drug|Pharmacologic Substance|Hospital Course|10287,10302|false|false|false|C0108101|calcium citrate|Calcium Citrate
Drug|Organic Chemical|Hospital Course|10295,10302|false|false|false|C0008857;C0376259|Citrates;citrate|Citrate
Drug|Pharmacologic Substance|Hospital Course|10295,10302|false|false|false|C0008857;C0376259|Citrates;citrate|Citrate
Event|Event|Hospital Course|10295,10302|false|false|false|||Citrate
Procedure|Laboratory Procedure|Hospital Course|10295,10302|false|false|false|C0201956|Citrate measurement|Citrate
Drug|Biomedical or Dental Material|Hospital Course|10312,10315|false|false|false|C0039225|Tablet Dosage Form|Tab
Event|Event|Hospital Course|10336,10343|false|false|false|||started
Finding|Gene or Genome|Hospital Course|10352,10355|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Event|Event|Hospital Course|10361,10370|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|10361,10370|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|10361,10370|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|10361,10370|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|10361,10370|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|10361,10382|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|10371,10382|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|10371,10382|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|10371,10382|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|10371,10382|false|false|false|C4284232|Medications|Medications
Event|Event|Hospital Course|10387,10392|false|false|false|||omega
Finding|Intellectual Product|Hospital Course|10387,10392|false|false|false|C1719844|Omega|omega
Drug|Biologically Active Substance|Hospital Course|10387,10394|false|false|false|C0015689|omega-3 fatty acids|omega-3
Drug|Organic Chemical|Hospital Course|10387,10394|false|false|false|C0015689|omega-3 fatty acids|omega-3
Drug|Pharmacologic Substance|Hospital Course|10387,10394|false|false|false|C0015689|omega-3 fatty acids|omega-3
Drug|Biologically Active Substance|Hospital Course|10387,10406|false|false|false|C0015689|omega-3 fatty acids|omega-3 fatty acids
Drug|Organic Chemical|Hospital Course|10387,10406|false|false|false|C0015689|omega-3 fatty acids|omega-3 fatty acids
Drug|Pharmacologic Substance|Hospital Course|10387,10406|false|false|false|C0015689|omega-3 fatty acids|omega-3 fatty acids
Drug|Organic Chemical|Hospital Course|10395,10406|false|false|false|C0015684|Fatty Acids|fatty acids
Drug|Chemical|Hospital Course|10401,10406|false|false|false|C0001128|Acids|acids
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10411,10418|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|10411,10418|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|10411,10418|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10432,10439|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|10432,10439|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|10432,10439|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Drug|Organic Chemical|Hospital Course|10464,10469|false|false|false|C0939679|Axert|Axert
Drug|Pharmacologic Substance|Hospital Course|10464,10469|false|false|false|C0939679|Axert|Axert
Drug|Biomedical or Dental Material|Hospital Course|10478,10484|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|10478,10484|false|false|false|||Tablet
Drug|Biomedical or Dental Material|Hospital Course|10498,10504|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|10498,10504|false|false|false|||Tablet
Event|Event|Hospital Course|10505,10507|false|false|false|||PO
Finding|Intellectual Product|Hospital Course|10508,10512|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|Hospital Course|10508,10518|false|false|false|C3537736|Once A Day|once a day
Finding|Idea or Concept|Hospital Course|10515,10518|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|10515,10518|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Hospital Course|10523,10529|false|false|false|||needed
Disorder|Disease or Syndrome|Hospital Course|10534,10542|false|false|false|C0149931|Migraine Disorders|migraine
Event|Event|Hospital Course|10534,10542|false|false|false|||migraine
Drug|Organic Chemical|Hospital Course|10549,10561|false|false|false|C1099456|escitalopram|escitalopram
Drug|Pharmacologic Substance|Hospital Course|10549,10561|false|false|false|C1099456|escitalopram|escitalopram
Event|Event|Hospital Course|10549,10561|false|false|false|||escitalopram
Drug|Biomedical or Dental Material|Hospital Course|10568,10574|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|10588,10594|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|10588,10594|false|false|false|||Tablet
Drug|Organic Chemical|Hospital Course|10619,10634|false|false|false|C0008318|cholecalciferol|cholecalciferol
Drug|Pharmacologic Substance|Hospital Course|10619,10634|false|false|false|C0008318|cholecalciferol|cholecalciferol
Drug|Vitamin|Hospital Course|10619,10634|false|false|false|C0008318|cholecalciferol|cholecalciferol
Event|Event|Hospital Course|10619,10634|false|false|false|||cholecalciferol
Drug|Organic Chemical|Hospital Course|10619,10647|false|false|false|C0008318|cholecalciferol|cholecalciferol (vitamin D3)
Drug|Pharmacologic Substance|Hospital Course|10619,10647|false|false|false|C0008318|cholecalciferol|cholecalciferol (vitamin D3)
Drug|Vitamin|Hospital Course|10619,10647|false|false|false|C0008318|cholecalciferol|cholecalciferol (vitamin D3)
Drug|Organic Chemical|Hospital Course|10636,10643|false|false|false|C0042890|Vitamins|vitamin
Drug|Pharmacologic Substance|Hospital Course|10636,10643|false|false|false|C0042890|Vitamins|vitamin
Drug|Vitamin|Hospital Course|10636,10643|false|false|false|C0042890|Vitamins|vitamin
Event|Event|Hospital Course|10636,10643|false|false|false|||vitamin
Drug|Organic Chemical|Hospital Course|10636,10646|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Drug|Pharmacologic Substance|Hospital Course|10636,10646|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Drug|Vitamin|Hospital Course|10636,10646|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10659,10666|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|10659,10666|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|10659,10666|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10681,10688|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|10681,10688|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|10681,10688|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Event|Event|Hospital Course|10689,10691|false|false|false|||PO
Finding|Intellectual Product|Hospital Course|10692,10696|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|Hospital Course|10692,10702|false|false|false|C3537736|Once A Day|once a day
Finding|Idea or Concept|Hospital Course|10699,10702|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|10699,10702|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|Hospital Course|10709,10718|false|false|false|C0024002|lorazepam|lorazepam
Drug|Pharmacologic Substance|Hospital Course|10709,10718|false|false|false|C0024002|lorazepam|lorazepam
Event|Event|Hospital Course|10709,10718|false|false|false|||lorazepam
Drug|Biomedical or Dental Material|Hospital Course|10726,10732|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|10733,10736|false|false|false|||Sig
Drug|Biomedical or Dental Material|Hospital Course|10746,10752|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|10746,10752|false|false|false|||Tablet
Event|Event|Hospital Course|10776,10782|false|false|false|||needed
Disorder|Mental or Behavioral Dysfunction|Hospital Course|10787,10794|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Event|Event|Hospital Course|10787,10794|false|false|false|||anxiety
Finding|Sign or Symptom|Hospital Course|10787,10794|false|false|false|C0860603|Anxiety symptoms|anxiety
Drug|Organic Chemical|Hospital Course|10801,10811|false|false|false|C0028978|omeprazole|omeprazole
Drug|Pharmacologic Substance|Hospital Course|10801,10811|false|false|false|C0028978|omeprazole|omeprazole
Event|Event|Hospital Course|10801,10811|false|false|false|||omeprazole
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10818,10825|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|10818,10825|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|10818,10825|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Attribute|Clinical Attribute|Hospital Course|10827,10834|false|false|false|C1545665|Views delayed|Delayed
Drug|Biomedical or Dental Material|Hospital Course|10827,10842|false|false|false|C1707664|Delayed Release Dosage Form|Delayed Release
Event|Event|Hospital Course|10835,10842|false|false|false|||Release
Finding|Functional Concept|Hospital Course|10835,10842|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|10835,10842|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10835,10842|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Event|Event|Hospital Course|10849,10852|false|false|false|||Sig
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10863,10870|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|10863,10870|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|10863,10870|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Attribute|Clinical Attribute|Hospital Course|10872,10879|false|false|false|C1545665|Views delayed|Delayed
Drug|Biomedical or Dental Material|Hospital Course|10872,10887|false|false|false|C1707664|Delayed Release Dosage Form|Delayed Release
Event|Event|Hospital Course|10880,10887|false|false|false|||Release
Finding|Functional Concept|Hospital Course|10880,10887|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|10880,10887|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10880,10887|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Disorder|Mental or Behavioral Dysfunction|Hospital Course|10897,10900|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10897,10900|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|10897,10900|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|10897,10900|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|10897,10900|false|false|false|C1332410|BID gene|BID
Finding|Finding|Hospital Course|10902,10909|false|false|false|C4035627|2 times|2 times
Disorder|Disease or Syndrome|Hospital Course|10904,10909|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|Hospital Course|10912,10915|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|10912,10915|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|Hospital Course|10923,10935|false|false|false|C0301532|Multivitamin preparation|multivitamin
Drug|Pharmacologic Substance|Hospital Course|10923,10935|false|false|false|C0301532|Multivitamin preparation|multivitamin
Drug|Vitamin|Hospital Course|10923,10935|false|false|false|C0301532|Multivitamin preparation|multivitamin
Event|Event|Hospital Course|10923,10935|false|false|false|||multivitamin
Drug|Pharmacologic Substance|Hospital Course|10923,10946|false|false|false|C0978787|Multivitamin tablet|multivitamin     Tablet
Drug|Biomedical or Dental Material|Hospital Course|10940,10946|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|10940,10946|false|false|false|||Tablet
Drug|Biomedical or Dental Material|Hospital Course|10960,10966|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|10960,10966|false|false|false|||Tablet
Drug|Organic Chemical|Hospital Course|10991,11001|false|false|false|C0034665|ranitidine|ranitidine
Drug|Pharmacologic Substance|Hospital Course|10991,11001|false|false|false|C0034665|ranitidine|ranitidine
Event|Event|Hospital Course|10991,11001|false|false|false|||ranitidine
Drug|Organic Chemical|Hospital Course|10991,11005|false|false|false|C0700466|ranitidine hydrochloride|ranitidine HCl
Drug|Pharmacologic Substance|Hospital Course|10991,11005|false|false|false|C0700466|ranitidine hydrochloride|ranitidine HCl
Disorder|Neoplastic Process|Hospital Course|11002,11005|false|false|false|C0023443|Hairy Cell Leukemia|HCl
Drug|Immunologic Factor|Hospital Course|11002,11005|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Inorganic Chemical|Hospital Course|11002,11005|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Pharmacologic Substance|Hospital Course|11002,11005|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Event|Event|Hospital Course|11002,11005|false|false|false|||HCl
Drug|Biomedical or Dental Material|Hospital Course|11013,11019|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|11033,11039|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|11033,11039|false|false|false|||Tablet
Disorder|Mental or Behavioral Dysfunction|Hospital Course|11043,11046|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11043,11046|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|11043,11046|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|11043,11046|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|11043,11046|false|false|false|C1332410|BID gene|BID
Disorder|Disease or Syndrome|Hospital Course|11051,11056|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|Hospital Course|11059,11062|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|11059,11062|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|Hospital Course|11070,11081|false|false|false|C0082607|fluticasone|fluticasone
Drug|Pharmacologic Substance|Hospital Course|11070,11081|false|false|false|C0082607|fluticasone|fluticasone
Event|Event|Hospital Course|11070,11081|false|false|false|||fluticasone
Drug|Biomedical or Dental Material|Hospital Course|11099,11104|false|false|false|C1154182|Spray Dosage Form|Spray
Event|Activity|Hospital Course|11099,11104|false|false|false|C2003858|Spray (action)|Spray
Event|Event|Hospital Course|11099,11104|false|false|false|||Spray
Finding|Functional Concept|Hospital Course|11099,11104|false|false|false|C4521772|Spray (administration method)|Spray
Drug|Biomedical or Dental Material|Hospital Course|11099,11116|false|false|false|C1710170|SPRAY, SUSPENSION|Spray, Suspension
Drug|Biomedical or Dental Material|Hospital Course|11106,11116|false|false|false|C0038960;C1382107|Suspension substance;Suspensions|Suspension
Drug|Substance|Hospital Course|11106,11116|false|false|false|C0038960;C1382107|Suspension substance;Suspensions|Suspension
Event|Event|Hospital Course|11106,11116|false|false|false|||Suspension
Finding|Functional Concept|Hospital Course|11106,11116|false|false|false|C1705537|Suspension (action)|Suspension
Drug|Biomedical or Dental Material|Hospital Course|11131,11136|false|false|false|C1154182|Spray Dosage Form|Spray
Event|Activity|Hospital Course|11131,11136|false|false|false|C2003858|Spray (action)|Spray
Event|Event|Hospital Course|11131,11136|false|false|false|||Spray
Finding|Functional Concept|Hospital Course|11131,11136|false|false|false|C4521772|Spray (administration method)|Spray
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11137,11142|false|false|false|C0028429||Nasal
Drug|Biomedical or Dental Material|Hospital Course|11137,11142|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Organic Chemical|Hospital Course|11137,11142|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Pharmacologic Substance|Hospital Course|11137,11142|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Finding|Finding|Hospital Course|11137,11142|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Finding|Functional Concept|Hospital Course|11137,11142|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Event|Event|Hospital Course|11143,11148|false|false|false|||DAILY
Drug|Biologically Active Substance|Hospital Course|11164,11171|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Element, Ion, or Isotope|Hospital Course|11164,11171|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Inorganic Chemical|Hospital Course|11164,11171|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Pharmacologic Substance|Hospital Course|11164,11171|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Vitamin|Hospital Course|11164,11171|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Event|Event|Hospital Course|11164,11171|false|false|false|||calcium
Finding|Physiologic Function|Hospital Course|11164,11171|false|false|false|C4553026|Calcium metabolic function|calcium
Procedure|Laboratory Procedure|Hospital Course|11164,11171|false|false|false|C0201925|Calcium measurement|calcium
Drug|Inorganic Chemical|Hospital Course|11164,11181|false|false|false|C0006681|calcium carbonate|calcium carbonate
Drug|Pharmacologic Substance|Hospital Course|11164,11181|false|false|false|C0006681|calcium carbonate|calcium carbonate
Drug|Element, Ion, or Isotope|Hospital Course|11172,11181|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|carbonate
Drug|Organic Chemical|Hospital Course|11172,11181|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|carbonate
Drug|Pharmacologic Substance|Hospital Course|11172,11181|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|carbonate
Event|Event|Hospital Course|11172,11181|false|false|false|||carbonate
Drug|Biologically Active Substance|Hospital Course|11189,11196|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Element, Ion, or Isotope|Hospital Course|11189,11196|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Inorganic Chemical|Hospital Course|11189,11196|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Pharmacologic Substance|Hospital Course|11189,11196|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Vitamin|Hospital Course|11189,11196|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Event|Event|Hospital Course|11189,11196|false|false|false|||calcium
Finding|Physiologic Function|Hospital Course|11189,11196|false|false|false|C4553026|Calcium metabolic function|calcium
Procedure|Laboratory Procedure|Hospital Course|11189,11196|false|false|false|C0201925|Calcium measurement|calcium
Drug|Biomedical or Dental Material|Hospital Course|11208,11214|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|11208,11214|false|false|false|||Tablet
Drug|Biomedical or Dental Material|Hospital Course|11229,11235|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|11236,11238|false|false|false|||PO
Finding|Intellectual Product|Hospital Course|11239,11243|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|Hospital Course|11239,11249|false|false|false|C3537736|Once A Day|once a day
Finding|Idea or Concept|Hospital Course|11246,11249|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|11246,11249|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Hospital Course|11256,11265|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|11256,11265|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|11256,11265|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|11256,11265|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|11256,11265|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|11256,11277|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|11256,11277|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|11266,11277|false|false|false|C2926604||Disposition
Event|Event|Hospital Course|11266,11277|false|false|false|||Disposition
Procedure|Health Care Activity|Hospital Course|11266,11277|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|Hospital Course|11279,11283|false|false|false|||Home
Finding|Idea or Concept|Hospital Course|11279,11283|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|11279,11283|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|11279,11283|false|false|false|C1553498|home health encounter|Home
Event|Event|Hospital Course|11286,11295|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|11286,11295|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|11286,11295|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|11286,11295|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|11286,11295|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|11286,11305|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|11296,11305|false|false|false|C0945731||Diagnosis
Event|Event|Hospital Course|11296,11305|false|false|false|||Diagnosis
Finding|Classification|Hospital Course|11296,11305|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|11296,11305|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|11296,11305|false|false|false|C0011900|Diagnosis|Diagnosis
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11307,11312|false|false|false|C0007531|Cecum|Cecal
Finding|Finding|Hospital Course|11307,11317|false|false|false|C3670817|Cecal mass|Cecal Mass
Event|Event|Hospital Course|11313,11317|false|false|false|||Mass
Finding|Finding|Hospital Course|11313,11317|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|Mass
Finding|Gene or Genome|Hospital Course|11313,11317|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|Mass
Finding|Intellectual Product|Hospital Course|11313,11317|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|Mass
Disorder|Acquired Abnormality|Hospital Course|11318,11342|false|false|false|C0473311|Hemorrhagic cyst of ovary|Hemorrhagic ovarian cyst
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11330,11337|false|false|false|C0205065|Ovarian|ovarian
Disorder|Disease or Syndrome|Hospital Course|11330,11342|false|false|false|C0029927|Ovarian Cysts|ovarian cyst
Disorder|Anatomical Abnormality|Hospital Course|11338,11342|false|false|false|C0010709|Cyst|cyst
Event|Event|Hospital Course|11338,11342|false|false|false|||cyst
Finding|Body Substance|Hospital Course|11338,11342|false|false|false|C1546594;C1550626|SpecimenType - Cyst|cyst
Finding|Intellectual Product|Hospital Course|11338,11342|false|false|false|C1546594;C1550626|SpecimenType - Cyst|cyst
Finding|Mental Process|Discharge Condition|11367,11373|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|11367,11380|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|11367,11380|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|11374,11380|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|11374,11380|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|11382,11387|false|false|false|||Clear
Finding|Idea or Concept|Discharge Condition|11382,11387|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|Discharge Condition|11392,11400|false|false|false|||coherent
Finding|Finding|Discharge Condition|11392,11400|false|false|false|C4068804|Coherent|coherent
Event|Event|Discharge Condition|11402,11407|false|false|false|||Level
Attribute|Clinical Attribute|Discharge Condition|11402,11424|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|11402,11424|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|Discharge Condition|11411,11424|false|false|false|||Consciousness
Finding|Finding|Discharge Condition|11411,11424|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|11411,11424|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|11426,11431|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|11426,11431|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|11426,11431|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|Discharge Condition|11426,11431|false|false|false|||Alert
Finding|Finding|Discharge Condition|11426,11431|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|11426,11431|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|11426,11431|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|Discharge Condition|11436,11447|false|false|false|||interactive
Finding|Functional Concept|Discharge Condition|11436,11447|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|11449,11457|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|11449,11457|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|11449,11457|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|11458,11464|false|false|false|C5889824||Status
Event|Event|Discharge Condition|11458,11464|false|false|false|||Status
Finding|Idea or Concept|Discharge Condition|11458,11464|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|11466,11476|false|false|false|||Ambulatory
Finding|Functional Concept|Discharge Condition|11466,11476|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|Discharge Condition|11466,11476|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|Discharge Condition|11466,11476|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|Discharge Condition|11466,11476|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|Discharge Condition|11479,11490|false|false|false|||Independent
Finding|Finding|Discharge Condition|11479,11490|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|Discharge Condition|11479,11490|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Gene or Genome|Discharge Instructions|11519,11523|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Event|Event|Discharge Instructions|11543,11551|false|false|false|||admitted
Finding|Idea or Concept|Discharge Instructions|11559,11567|false|false|false|C1547192|Organization unit type - Hospital|hospital
Anatomy|Body Location or Region|Discharge Instructions|11572,11581|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|Discharge Instructions|11572,11586|false|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|Discharge Instructions|11582,11586|false|true|false|C2598155||pain
Event|Event|Discharge Instructions|11582,11586|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|11582,11586|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|11582,11586|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Mental Process|Discharge Instructions|11598,11603|false|false|false|C0039869||think
Event|Event|Discharge Instructions|11608,11615|false|false|false|||related
Disorder|Acquired Abnormality|Discharge Instructions|11621,11645|false|false|false|C0473311|Hemorrhagic cyst of ovary|hemorrhagic ovarian cyst
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|11633,11640|false|false|false|C0205065|Ovarian|ovarian
Disorder|Disease or Syndrome|Discharge Instructions|11633,11645|false|false|false|C0029927|Ovarian Cysts|ovarian cyst
Disorder|Anatomical Abnormality|Discharge Instructions|11641,11645|false|false|false|C0010709|Cyst|cyst
Event|Event|Discharge Instructions|11641,11645|false|false|false|||cyst
Finding|Body Substance|Discharge Instructions|11641,11645|false|false|false|C1546594;C1550626|SpecimenType - Cyst|cyst
Finding|Intellectual Product|Discharge Instructions|11641,11645|false|false|false|C1546594;C1550626|SpecimenType - Cyst|cyst
Event|Event|Discharge Instructions|11658,11665|false|false|false|||treated
Drug|Hazardous or Poisonous Substance|Discharge Instructions|11671,11681|false|false|false|C0002771;C4722089|Analgesics;Analgesics [TC]|analgesics
Drug|Organic Chemical|Discharge Instructions|11671,11681|false|false|false|C0002771;C4722089|Analgesics;Analgesics [TC]|analgesics
Drug|Pharmacologic Substance|Discharge Instructions|11671,11681|false|false|false|C0002771;C4722089|Analgesics;Analgesics [TC]|analgesics
Event|Event|Discharge Instructions|11671,11681|false|false|false|||analgesics
Attribute|Clinical Attribute|Discharge Instructions|11692,11696|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|11692,11696|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|11692,11696|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|11692,11696|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Discharge Instructions|11697,11705|false|false|false|||resolved
Disorder|Congenital Abnormality|Discharge Instructions|11724,11727|false|false|false|C0041207|Truncus Arteriosus, Persistent|CAT
Drug|Amino Acid, Peptide, or Protein|Discharge Instructions|11724,11727|false|false|false|C0008169;C1443200;C3530118|CAT protein, human;Cat hair antigen;Chloramphenicol O-Acetyltransferase|CAT
Drug|Enzyme|Discharge Instructions|11724,11727|false|false|false|C0008169;C1443200;C3530118|CAT protein, human;Cat hair antigen;Chloramphenicol O-Acetyltransferase|CAT
Drug|Immunologic Factor|Discharge Instructions|11724,11727|false|false|false|C0008169;C1443200;C3530118|CAT protein, human;Cat hair antigen;Chloramphenicol O-Acetyltransferase|CAT
Event|Event|Discharge Instructions|11724,11727|false|false|false|||CAT
Finding|Gene or Genome|Discharge Instructions|11724,11727|false|false|false|C1151515;C1366498;C1413138;C4050461;C4758039|CAT gene;Chloramphenicol Acetyl Transferase Gene;Chronic Obstructive Pulmonary Disease Assessment Test scale;Cutaneous Assessment Tool;catalase activity|CAT
Finding|Intellectual Product|Discharge Instructions|11724,11727|false|false|false|C1151515;C1366498;C1413138;C4050461;C4758039|CAT gene;Chloramphenicol Acetyl Transferase Gene;Chronic Obstructive Pulmonary Disease Assessment Test scale;Cutaneous Assessment Tool;catalase activity|CAT
Finding|Molecular Function|Discharge Instructions|11724,11727|false|false|false|C1151515;C1366498;C1413138;C4050461;C4758039|CAT gene;Chloramphenicol Acetyl Transferase Gene;Chronic Obstructive Pulmonary Disease Assessment Test scale;Cutaneous Assessment Tool;catalase activity|CAT
Procedure|Diagnostic Procedure|Discharge Instructions|11724,11727|false|false|false|C0040405;C0280589;C2097305|X-Ray Computed Tomography;allergy testing cat;cytarabine/thioguanine protocol|CAT
Procedure|Laboratory Procedure|Discharge Instructions|11724,11727|false|false|false|C0040405;C0280589;C2097305|X-Ray Computed Tomography;allergy testing cat;cytarabine/thioguanine protocol|CAT
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|11724,11727|false|false|false|C0040405;C0280589;C2097305|X-Ray Computed Tomography;allergy testing cat;cytarabine/thioguanine protocol|CAT
Finding|Intellectual Product|Discharge Instructions|11724,11732|false|false|false|C1547980|CAT Scan Section ID|CAT scan
Procedure|Diagnostic Procedure|Discharge Instructions|11724,11732|false|false|false|C0040405|X-Ray Computed Tomography|CAT scan
Event|Event|Discharge Instructions|11728,11732|false|false|false|||scan
Procedure|Diagnostic Procedure|Discharge Instructions|11728,11732|false|false|false|C0034606;C0441633|Radionuclide Imaging;Scanning|scan
Event|Event|Discharge Instructions|11733,11740|false|false|false|||showing
Finding|Finding|Discharge Instructions|11741,11747|false|false|false|C0577559|Mass of body structure|a mass
Event|Event|Discharge Instructions|11743,11747|false|false|false|||mass
Finding|Finding|Discharge Instructions|11743,11747|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|Discharge Instructions|11743,11747|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|Discharge Instructions|11743,11747|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|11755,11760|false|false|false|C0007531|Cecum|cecum
Disorder|Neoplastic Process|Discharge Instructions|11755,11760|false|false|false|C0153437;C0496859|Benign neoplasm of cecum;Malignant neoplasm of cecum|cecum
Event|Event|Discharge Instructions|11780,11791|false|false|false|||colonoscopy
Procedure|Diagnostic Procedure|Discharge Instructions|11780,11791|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Procedure|Health Care Activity|Discharge Instructions|11780,11791|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Event|Event|Discharge Instructions|11795,11801|false|false|false|||biopsy
Event|Event|Discharge Instructions|11807,11811|false|false|false|||mass
Finding|Finding|Discharge Instructions|11807,11811|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|Discharge Instructions|11807,11811|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|Discharge Instructions|11807,11811|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Event|Event|Discharge Instructions|11828,11834|false|false|false|||follow
Event|Event|Discharge Instructions|11849,11867|false|false|false|||gastroenterologist
Event|Event|Discharge Instructions|11887,11890|false|false|false|||see
Event|Event|Discharge Instructions|11896,11908|false|false|false|||gynecologist
Event|Event|Discharge Instructions|11923,11927|false|false|false|||need
Finding|Functional Concept|Discharge Instructions|11923,11927|false|false|false|C0686904|Patient need for (contextual qualifier)|need
Event|Event|Discharge Instructions|11932,11939|false|false|false|||restart
Anatomy|Body Space or Junction|Discharge Instructions|11945,11949|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Discharge Instructions|11945,11949|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Discharge Instructions|11945,11949|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Discharge Instructions|11945,11949|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Drug|Pharmacologic Substance|Discharge Instructions|11945,11963|false|false|false|C0009905|Contraceptives, Oral|oral contraceptive
Finding|Finding|Discharge Instructions|11945,11963|false|false|false|C0029151|Uses oral contraception (finding)|oral contraceptive
Drug|Pharmacologic Substance|Discharge Instructions|11950,11963|false|false|false|C0009871|Contraceptive Agents|contraceptive
Event|Event|Discharge Instructions|11950,11963|false|false|false|||contraceptive
Finding|Finding|Discharge Instructions|11950,11963|false|false|false|C0344225|Encounter due to presence of intrauterine contraceptive device|contraceptive
Event|Event|Discharge Instructions|11977,11981|true|false|false|||make
Event|Event|Discharge Instructions|11986,11993|true|false|false|||changes
Finding|Functional Concept|Discharge Instructions|11986,11993|true|false|false|C0392747|Changing|changes
Finding|Idea or Concept|Discharge Instructions|12002,12006|true|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Discharge Instructions|12002,12006|true|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Discharge Instructions|12002,12006|true|false|false|C1553498|home health encounter|home
Attribute|Clinical Attribute|Discharge Instructions|12007,12018|true|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|12007,12018|true|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Discharge Instructions|12007,12018|true|false|false|||medications
Finding|Intellectual Product|Discharge Instructions|12007,12018|true|false|false|C4284232|Medications|medications
Procedure|Health Care Activity|Discharge Instructions|12023,12031|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|12032,12044|false|false|false|C3263700||Instructions
Event|Event|Discharge Instructions|12032,12044|false|false|false|||Instructions
Finding|Intellectual Product|Discharge Instructions|12032,12044|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

