 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
_|27,28
_|28,29
_|29,30
No|31,33
:|33,34
_|37,38
_|38,39
_|39,40
<EOL>|40,41
<EOL>|42,43
Admission|43,52
Date|53,57
:|57,58
_|60,61
_|61,62
_|62,63
Discharge|77,86
Date|87,91
:|91,92
_|95,96
_|96,97
_|97,98
<EOL>|98,99
<EOL>|100,101
Date|101,105
of|106,108
Birth|109,114
:|114,115
_|117,118
_|118,119
_|119,120
Sex|133,136
:|136,137
F|140,141
<EOL>|141,142
<EOL>|143,144
Service|144,151
:|151,152
MEDICINE|153,161
<EOL>|161,162
<EOL>|163,164
Allergies|164,173
:|173,174
<EOL>|175,176
meropenem|176,185
<EOL>|185,186
<EOL>|187,188
Attending|188,197
:|197,198
_|199,200
_|200,201
_|201,202
<EOL>|202,203
<EOL>|204,205
_|205,206
_|206,207
_|207,208
Complaint|209,218
:|218,219
<EOL>|219,220
Hypercarbic|220,231
Respiratory|232,243
Failure|244,251
<EOL>|251,252
<EOL>|253,254
Major|254,259
Surgical|260,268
or|269,271
Invasive|272,280
Procedure|281,290
:|290,291
<EOL>|291,292
Mechanical|292,302
Intubation|303,313
,|313,314
Arterial|315,323
-|324,325
Line|325,329
,|329,330
Central|331,338
Venous|339,345
Access|346,352
<EOL>|353,354
Line|354,358
<EOL>|358,359
<EOL>|360,361
History|361,368
of|369,371
Present|372,379
Illness|380,387
:|387,388
<EOL>|388,389
This|389,393
is|394,396
an|397,399
_|400,401
_|401,402
_|402,403
year|404,408
old|409,412
woman|413,418
,|418,419
recently|420,428
hospitalized|429,441
for|442,445
C|446,447
.|447,448
<EOL>|449,450
Difficile|450,459
sepsis|460,466
and|467,470
shock|471,476
,|476,477
complicated|478,489
by|490,492
readmission|493,504
<EOL>|505,506
hypoxia|506,513
/|513,514
hypercarbia|514,525
(|526,527
_|527,528
_|528,529
_|529,530
)|530,531
who|532,535
presents|536,544
with|545,549
respiratory|550,561
<EOL>|562,563
distress|563,571
and|572,575
respiratory|576,587
failure|588,595
.|595,596
<EOL>|596,597
.|597,598
<EOL>|598,599
The|599,602
patient|603,610
had|611,614
reportedly|615,625
been|626,630
doing|631,636
well|637,641
_|642,643
_|643,644
_|644,645
rehab|646,651
until|652,657
today|658,663
<EOL>|664,665
when|665,669
she|670,673
was|674,677
noted|678,683
to|684,686
have|687,691
an|692,694
altered|695,702
(|703,704
depressed|704,713
)|713,714
mental|715,721
status|722,728
,|728,729
<EOL>|730,731
tachypnea|731,740
,|740,741
and|742,745
dyspnea|746,753
.|753,754
EMS|756,759
was|760,763
called|764,770
who|771,774
found|775,780
the|781,784
patient|785,792
_|793,794
_|794,795
_|795,796
<EOL>|797,798
extremis|798,806
,|806,807
intubation|808,818
was|819,822
attempted|823,832
x2|833,835
and|836,839
failed|840,846
.|846,847
A|849,850
_|851,852
_|852,853
_|853,854
airway|855,861
<EOL>|862,863
was|863,866
placed|867,873
and|874,877
the|878,881
patient|882,889
was|890,893
transported|894,905
to|906,908
_|909,910
_|910,911
_|911,912
emergency|913,922
<EOL>|923,924
department|924,934
.|934,935
There|937,942
were|943,947
no|948,950
reports|951,958
of|959,961
increased|962,971
coughing|972,980
or|981,983
<EOL>|984,985
stooling|985,993
from|994,998
_|999,1000
_|1000,1001
_|1001,1002
.|1002,1003
<EOL>|1003,1004
.|1004,1005
<EOL>|1005,1006
The|1006,1009
patient|1010,1017
has|1018,1021
had|1022,1025
a|1026,1027
complicated|1028,1039
medical|1040,1047
course|1048,1054
_|1055,1056
_|1056,1057
_|1057,1058
the|1059,1062
past|1063,1067
<EOL>|1068,1069
month|1069,1074
-|1075,1076
<EOL>|1077,1078
.|1078,1079
<EOL>|1079,1080
_|1080,1081
_|1081,1082
_|1082,1083
brief|1084,1089
,|1089,1090
the|1091,1094
patient|1095,1102
was|1103,1106
initially|1107,1116
discharge|1117,1126
on|1127,1129
_|1130,1131
_|1131,1132
_|1132,1133
after|1134,1139
<EOL>|1140,1141
a|1141,1142
14|1143,1145
hosptilazation|1146,1160
for|1161,1164
c|1165,1166
.|1166,1167
diff|1167,1171
colitis|1172,1179
complicated|1180,1191
by|1192,1194
sepsis|1195,1201
and|1202,1205
<EOL>|1206,1207
hypercarbic|1207,1218
respiratory|1219,1230
failure|1231,1238
requiring|1239,1248
intubation|1249,1259
.|1259,1260
On|1262,1264
the|1265,1268
<EOL>|1269,1270
day|1270,1273
following|1274,1283
discharge|1284,1293
from|1294,1298
that|1299,1303
admission|1304,1313
,|1313,1314
the|1315,1318
patient|1319,1326
was|1327,1330
<EOL>|1331,1332
noted|1332,1337
to|1338,1340
be|1341,1343
complaining|1344,1355
of|1356,1358
worsening|1359,1368
SOB|1369,1372
and|1373,1376
ABG|1377,1380
at|1381,1383
_|1384,1385
_|1385,1386
_|1386,1387
<EOL>|1388,1389
was|1389,1392
7.4|1393,1396
/|1396,1397
_|1397,1398
_|1398,1399
_|1399,1400
.|1400,1401
She|1402,1405
was|1406,1409
re-admitted|1410,1421
to|1422,1424
_|1425,1426
_|1426,1427
_|1427,1428
on|1429,1431
_|1432,1433
_|1433,1434
_|1434,1435
to|1436,1438
the|1439,1442
MICU|1443,1447
<EOL>|1448,1449
and|1449,1452
intially|1453,1461
reuqired|1462,1470
biPAP|1471,1476
for|1477,1480
HD1|1481,1484
-|1484,1485
2|1485,1486
.|1486,1487
Her|1488,1491
oxygen|1492,1498
requirement|1499,1510
on|1511,1513
<EOL>|1514,1515
d|1515,1516
/|1516,1517
c|1517,1518
was|1519,1522
2L|1523,1525
NC|1526,1528
.|1528,1529
The|1532,1535
etiology|1536,1544
of|1545,1547
her|1548,1551
hypercarbic|1552,1563
respiratory|1564,1575
<EOL>|1576,1577
failure|1577,1584
was|1585,1588
felt|1589,1593
to|1594,1596
be|1597,1599
_|1600,1601
_|1601,1602
_|1602,1603
hypoventilation|1604,1619
from|1620,1624
somnolence|1625,1635
<EOL>|1636,1637
related|1637,1644
to|1645,1647
oversedation|1648,1660
with|1661,1665
zyprexa|1666,1673
which|1674,1679
was|1680,1683
held|1684,1688
on|1689,1691
<EOL>|1692,1693
discharge|1693,1702
.|1702,1703
A|1704,1705
CTA|1706,1709
chest|1710,1715
was|1716,1719
negative|1720,1728
for|1729,1732
PE|1733,1735
and|1736,1739
showed|1740,1746
no|1747,1749
clear|1750,1755
<EOL>|1756,1757
evidence|1757,1765
of|1766,1768
pneumonia|1769,1778
.|1778,1779
She|1781,1784
was|1785,1788
initially|1789,1798
started|1799,1806
on|1807,1809
HCAP|1810,1814
<EOL>|1815,1816
antibiotics|1816,1827
with|1828,1832
vanc|1833,1837
/|1837,1838
cefepime|1838,1846
which|1847,1852
were|1853,1857
stopped|1858,1865
on|1866,1868
HD|1869,1871
4|1872,1873
prior|1874,1879
<EOL>|1880,1881
to|1881,1883
discharge|1884,1893
given|1894,1899
that|1900,1904
all|1905,1908
cultures|1909,1917
were|1918,1922
negative|1923,1931
and|1932,1935
there|1936,1941
was|1942,1945
<EOL>|1946,1947
no|1947,1949
consolidation|1950,1963
on|1964,1966
imaging|1967,1974
.|1974,1975
<EOL>|1976,1977
.|1977,1978
<EOL>|1978,1979
_|1979,1980
_|1980,1981
_|1981,1982
the|1983,1986
ED|1987,1989
,|1989,1990
initial|1991,1998
VS|1999,2001
were|2002,2006
:|2006,2007
HR|2008,2010
:|2010,2011
82|2012,2014
BP|2015,2017
:|2017,2018
94|2019,2021
systolic|2022,2030
Resp|2031,2035
:|2035,2036
No|2037,2039
<EOL>|2040,2041
spontaneous|2041,2052
respirations|2053,2065
O|2066,2067
(|2067,2068
2|2068,2069
)|2069,2070
Sat|2070,2073
:|2073,2074
100|2075,2078
;|2078,2079
Initial|2081,2088
labs|2089,2093
<EOL>|2094,2095
demonstrated|2095,2107
hct|2108,2111
22.0|2112,2116
,|2116,2117
wbc|2118,2121
16.0|2122,2126
,|2126,2127
creatinine|2128,2138
0.3|2139,2142
,|2142,2143
BIN|2144,2147
18|2148,2150
,|2150,2151
lipase|2152,2158
<EOL>|2159,2160
148|2160,2163
and|2164,2167
lactate|2168,2175
0.9|2176,2179
.|2179,2180
A|2181,2182
cxr|2183,2186
demonstrated|2187,2199
bilateral|2200,2209
pleural|2210,2217
<EOL>|2218,2219
effusions|2219,2228
with|2229,2233
R|2234,2235
>|2235,2236
L|2236,2237
.|2237,2238
A|2241,2242
UA|2243,2245
demonstrated|2246,2258
large|2259,2264
leuks|2265,2270
,|2270,2271
positive|2272,2280
<EOL>|2281,2282
nitrites|2282,2290
and|2291,2294
104|2295,2298
wbc|2299,2302
.|2302,2303
Due|2305,2308
respiratory|2309,2320
failure|2321,2328
the|2329,2332
patient|2333,2340
was|2341,2344
<EOL>|2345,2346
intubated|2346,2355
.|2355,2356
<EOL>|2358,2359
.|2359,2360
<EOL>|2360,2361
An|2361,2363
initial|2364,2371
ABG|2372,2375
was|2376,2379
7.|2380,2382
_|2382,2383
_|2383,2384
_|2384,2385
/|2385,2386
128|2386,2389
which|2390,2395
was|2396,2399
7.|2400,2402
_|2402,2403
_|2403,2404
_|2404,2405
/|2405,2406
395|2406,2409
post|2410,2414
<EOL>|2415,2416
intubation|2416,2426
.|2426,2427
The|2429,2432
patient|2433,2440
was|2441,2444
given|2445,2450
vancomycin|2451,2461
and|2462,2465
cefepime|2466,2474
for|2475,2478
<EOL>|2479,2480
coverage|2480,2488
of|2489,2491
both|2492,2496
a|2497,2498
urinary|2499,2506
and|2507,2510
pulmonary|2511,2520
source|2521,2527
.|2527,2528
Post|2529,2533
intubation|2534,2544
<EOL>|2545,2546
her|2546,2549
BP|2550,2552
dropped|2553,2560
to|2561,2563
the|2564,2567
_|2568,2569
_|2569,2570
_|2570,2571
.|2571,2572
She|2573,2576
was|2577,2580
started|2581,2588
on|2589,2591
levophed|2592,2600
and|2601,2604
<EOL>|2605,2606
phenylephrine|2606,2619
through|2620,2627
her|2628,2631
existing|2632,2640
PICC|2641,2645
line|2646,2650
.|2650,2651
Given|2652,2657
her|2658,2661
altered|2662,2669
<EOL>|2670,2671
mental|2671,2677
status|2678,2684
on|2685,2687
arrival|2688,2695
,|2695,2696
a|2697,2698
head|2699,2703
CT|2704,2706
was|2707,2710
performed|2711,2720
which|2721,2726
showed|2727,2733
<EOL>|2734,2735
no|2735,2737
acute|2738,2743
findings|2744,2752
.|2752,2753
Vitals|2754,2760
on|2761,2763
transfer|2764,2772
were|2773,2777
:|2777,2778
36.3|2779,2783
66|2784,2786
118|2787,2790
107|2791,2794
/|2794,2795
58|2795,2797
<EOL>|2798,2799
99|2799,2801
%|2801,2802
.|2802,2803
<EOL>|2804,2805
.|2805,2806
<EOL>|2806,2807
Vent|2807,2811
settings|2812,2820
were|2821,2825
:|2825,2826
fio2|2827,2831
60|2832,2834
%|2834,2835
RR|2836,2838
18|2839,2841
Vt|2842,2844
400|2845,2848
peep|2849,2853
5.|2854,2856
Sedation|2857,2865
with|2866,2870
<EOL>|2871,2872
midazolam|2872,2881
and|2882,2885
fentanyl|2886,2894
.|2894,2895
She|2896,2899
was|2900,2903
transferred|2904,2915
on|2916,2918
levophed|2919,2927
alone|2928,2933
w|2934,2935
/|2935,2936
<EOL>|2937,2938
MAPs|2938,2942
>|2942,2943
70|2944,2946
.|2946,2947
<EOL>|2947,2948
.|2948,2949
<EOL>|2952,2953
On|2953,2955
arrival|2956,2963
to|2964,2966
the|2967,2970
MICU|2971,2975
,|2975,2976
vitals|2978,2984
were|2985,2989
:|2989,2990
36.2|2991,2995
106|2996,2999
/|2999,3000
58|3000,3002
77|3003,3005
18|3006,3008
(|3009,3010
vented|3010,3016
)|3016,3017
<EOL>|3018,3019
100|3019,3022
%|3022,3023
on|3024,3026
40|3027,3029
%|3029,3030
FiO2|3031,3035
.|3035,3036
The|3038,3041
patient|3042,3049
was|3050,3053
on|3054,3056
a|3057,3058
levophed|3059,3067
drip|3068,3072
,|3072,3073
was|3074,3077
not|3078,3081
<EOL>|3082,3083
sedated|3083,3090
,|3090,3091
was|3092,3095
unresponsive|3096,3108
to|3109,3111
verbal|3112,3118
and|3119,3122
painful|3123,3130
stimuli|3131,3138
,|3138,3139
was|3140,3143
<EOL>|3144,3145
thought|3145,3152
to|3153,3155
have|3156,3160
a|3161,3162
brief|3163,3168
episode|3169,3176
of|3177,3179
decerebrate|3180,3191
posturing|3192,3201
with|3202,3206
<EOL>|3207,3208
the|3208,3211
upper|3212,3217
extremities|3218,3229
.|3229,3230
<EOL>|3230,3231
.|3231,3232
<EOL>|3233,3234
Review|3234,3240
of|3241,3243
systems|3244,3251
:|3251,3252
Unable|3254,3260
to|3261,3263
Obtain|3264,3270
<EOL>|3270,3271
<EOL>|3271,3272
<EOL>|3273,3274
Past|3274,3278
Medical|3279,3286
History|3287,3294
:|3294,3295
<EOL>|3295,3296
Anemia|3296,3302
<EOL>|3304,3305
Borderline|3305,3315
cholesterol|3316,3327
<EOL>|3329,3330
Recurrent|3330,3339
C.|3340,3342
Diff|3343,3347
<EOL>|3349,3350
Flatulence|3350,3360
<EOL>|3362,3363
Heart|3363,3368
Murmur|3369,3375
<EOL>|3377,3378
Hypertension|3378,3390
<EOL>|3392,3393
Hypothyroidism|3393,3407
<EOL>|3409,3410
Mitral|3410,3416
Regurgitation|3417,3430
<EOL>|3432,3433
Osteoporosis|3433,3445
<EOL>|3447,3448
Pneumonia|3448,3457
<EOL>|3459,3460
Sinusitis|3460,3469
<EOL>|3471,3472
Sjogren|3472,3479
<EOL>|3481,3482
<EOL>|3483,3484
Social|3484,3490
History|3491,3498
:|3498,3499
<EOL>|3499,3500
_|3500,3501
_|3501,3502
_|3502,3503
<EOL>|3503,3504
Family|3504,3510
History|3511,3518
:|3518,3519
<EOL>|3519,3520
Long|3520,3524
history|3525,3532
of|3533,3535
hypertension|3536,3548
_|3549,3550
_|3550,3551
_|3551,3552
her|3553,3556
family|3557,3563
.|3563,3564
Father|3566,3572
's|3572,3574
family|3575,3581
has|3582,3585
<EOL>|3586,3587
a|3587,3588
history|3589,3596
of|3597,3599
multiple|3600,3608
cancers|3609,3616
.|3616,3617
She|3619,3622
has|3623,3626
a|3627,3628
grandfather|3629,3640
with|3641,3645
a|3646,3647
<EOL>|3648,3649
history|3649,3656
of|3657,3659
stomach|3660,3667
cancer|3668,3674
and|3675,3678
an|3679,3681
uncle|3682,3687
with|3688,3692
a|3693,3694
history|3695,3702
of|3703,3705
throat|3706,3712
<EOL>|3713,3714
cancer|3714,3720
.|3720,3721
No|3723,3725
history|3726,3733
of|3734,3736
colon|3737,3742
cancers|3743,3750
.|3750,3751
Father|3752,3758
had|3759,3762
stroke|3763,3769
.|3769,3770
No|3771,3773
<EOL>|3774,3775
family|3775,3781
h|3782,3783
/|3783,3784
o|3784,3785
MI|3786,3788
.|3788,3789
Mother|3790,3796
had|3797,3800
a|3801,3802
heart|3803,3808
valve|3809,3814
replaced|3815,3823
.|3823,3824
<EOL>|3824,3825
<EOL>|3825,3826
<EOL>|3827,3828
Physical|3828,3836
Exam|3837,3841
:|3841,3842
<EOL>|3842,3843
ADMISSION|3843,3852
PHYSICAL|3853,3861
EXAM|3862,3866
:|3866,3867
<EOL>|3868,3869
36.2|3869,3873
106|3874,3877
/|3877,3878
58|3878,3880
77|3881,3883
18|3884,3886
(|3887,3888
vented|3888,3894
)|3894,3895
100|3896,3899
%|3899,3900
on|3901,3903
40|3904,3906
%|3906,3907
FiO2|3908,3912
<EOL>|3914,3915
General|3915,3922
:|3922,3923
Intubated|3924,3933
,|3933,3934
unresponsive|3935,3947
,|3947,3948
pale|3949,3953
,|3953,3954
very|3955,3959
thin|3960,3964
<EOL>|3966,3967
HEENT|3967,3972
:|3972,3973
Sclera|3974,3980
anicteric|3981,3990
,|3990,3991
MMM|3992,3995
,|3995,3996
oropharynx|3997,4007
clear|4008,4013
,|4013,4014
pupils|4015,4021
<EOL>|4022,4023
constricted|4023,4034
and|4035,4038
sluggish|4039,4047
b|4048,4049
/|4049,4050
l|4050,4051
;|4051,4052
there|4053,4058
is|4059,4061
a|4062,4063
dobhoff|4064,4071
and|4072,4075
an|4076,4078
NGT|4079,4082
<EOL>|4083,4084
present|4084,4091
<EOL>|4093,4094
Neck|4094,4098
:|4098,4099
supple|4100,4106
,|4106,4107
JVP|4108,4111
not|4112,4115
elevated|4116,4124
,|4124,4125
no|4126,4128
LAD|4129,4132
<EOL>|4134,4135
CV|4135,4137
:|4137,4138
Regular|4139,4146
rate|4147,4151
and|4152,4155
rhythm|4156,4162
,|4162,4163
normal|4164,4170
S1|4171,4173
+|4174,4175
S2|4176,4178
,|4178,4179
there|4180,4185
is|4186,4188
a|4189,4190
_|4191,4192
_|4192,4193
_|4193,4194
SEM|4195,4198
<EOL>|4199,4200
best|4200,4204
heard|4205,4210
over|4211,4215
the|4216,4219
LSB|4220,4223
.|4223,4224
There|4226,4231
is|4232,4234
a|4235,4236
midline|4237,4244
catheter|4245,4253
present|4254,4261
_|4262,4263
_|4263,4264
_|4264,4265
<EOL>|4266,4267
the|4267,4270
R|4271,4272
arm|4273,4276
<EOL>|4276,4277
Lungs|4277,4282
:|4282,4283
Bilateral|4284,4293
crackles|4294,4302
R|4303,4304
>|4305,4306
L|4307,4308
,|4308,4309
no|4310,4312
spontaneous|4313,4324
respirations|4325,4337
;|4337,4338
<EOL>|4339,4340
there|4340,4345
is|4346,4348
an|4349,4351
ETT|4352,4355
_|4356,4357
_|4357,4358
_|4358,4359
place|4360,4365
.|4365,4366
<EOL>|4366,4367
Abdomen|4367,4374
:|4374,4375
soft|4376,4380
,|4380,4381
non-distended|4382,4395
,|4395,4396
bowel|4397,4402
sounds|4403,4409
present|4410,4417
,|4417,4418
no|4419,4421
<EOL>|4422,4423
organomegaly|4423,4435
<EOL>|4437,4438
GU|4438,4440
:|4440,4441
Foley|4442,4447
present|4448,4455
;|4455,4456
there|4457,4462
is|4463,4465
a|4466,4467
candidal|4468,4476
rash|4477,4481
_|4482,4483
_|4483,4484
_|4484,4485
the|4486,4489
groin|4490,4495
area|4496,4500
,|4500,4501
<EOL>|4502,4503
there|4503,4508
is|4509,4511
powder|4512,4518
c|4519,4520
/|4520,4521
w|4521,4522
miconazole|4523,4533
powder|4534,4540
present|4541,4548
over|4549,4553
the|4554,4557
same|4558,4562
<EOL>|4563,4564
distribution|4564,4576
<EOL>|4578,4579
Ext|4579,4582
:|4582,4583
warm|4584,4588
,|4588,4589
well|4590,4594
perfused|4595,4603
,|4603,4604
2|4605,4606
+|4606,4607
pulses|4608,4614
,|4614,4615
no|4616,4618
clubbing|4619,4627
,|4627,4628
cyanosis|4629,4637
or|4638,4640
<EOL>|4641,4642
edema|4642,4647
<EOL>|4649,4650
Neuro|4650,4655
:|4655,4656
Unable|4657,4663
to|4664,4666
fully|4667,4672
evaluate|4673,4681
due|4682,4685
to|4686,4688
unresponsiveness|4689,4705
.|4705,4706
The|4708,4711
<EOL>|4712,4713
patient|4713,4720
has|4721,4724
1|4725,4726
+|4726,4727
DTRs|4728,4732
bilaterally|4733,4744
_|4745,4746
_|4746,4747
_|4747,4748
all|4749,4752
extremities|4753,4764
;|4764,4765
<EOL>|4766,4767
decerebration|4767,4780
briefly|4781,4788
noted|4789,4794
_|4795,4796
_|4796,4797
_|4797,4798
the|4799,4802
upper|4803,4808
extremities|4809,4820
.|4820,4821
<EOL>|4823,4824
.|4824,4825
<EOL>|4825,4826
DISCHARGE|4826,4835
PHYSICAL|4836,4844
EXAM|4845,4849
:|4849,4850
*|4851,4852
*|4852,4853
*|4853,4854
*|4854,4855
<EOL>|4855,4856
<EOL>|4857,4858
Pertinent|4858,4867
Results|4868,4875
:|4875,4876
<EOL>|4876,4877
ADMISSION|4877,4886
LABS|4887,4891
:|4891,4892
<EOL>|4892,4893
<EOL>|4893,4894
_|4894,4895
_|4895,4896
_|4896,4897
11|4898,4900
:|4900,4901
43AM|4901,4905
BLOOD|4906,4911
WBC|4912,4915
-|4915,4916
16|4916,4918
.|4918,4919
0|4919,4920
*|4920,4921
RBC|4922,4925
-|4925,4926
2|4926,4927
.|4927,4928
84|4928,4930
*|4930,4931
Hgb|4932,4935
-|4935,4936
8|4936,4937
.|4937,4938
4|4938,4939
*|4939,4940
Hct|4941,4944
-|4944,4945
29|4945,4947
.|4947,4948
0|4948,4949
*|4949,4950
<EOL>|4951,4952
MCV|4952,4955
-|4955,4956
102|4956,4959
*|4959,4960
MCH|4961,4964
-|4964,4965
29.7|4965,4969
MCHC|4970,4974
-|4974,4975
29|4975,4977
.|4977,4978
1|4978,4979
*|4979,4980
RDW|4981,4984
-|4984,4985
16|4985,4987
.|4987,4988
4|4988,4989
*|4989,4990
Plt|4991,4994
_|4995,4996
_|4996,4997
_|4997,4998
<EOL>|4998,4999
_|4999,5000
_|5000,5001
_|5001,5002
11|5003,5005
:|5005,5006
43AM|5006,5010
BLOOD|5011,5016
_|5017,5018
_|5018,5019
_|5019,5020
PTT|5021,5024
-|5024,5025
38|5025,5027
.|5027,5028
4|5028,5029
*|5029,5030
_|5031,5032
_|5032,5033
_|5033,5034
<EOL>|5034,5035
_|5035,5036
_|5036,5037
_|5037,5038
11|5039,5041
:|5041,5042
43AM|5042,5046
BLOOD|5047,5052
_|5053,5054
_|5054,5055
_|5055,5056
02|5057,5059
:|5059,5060
46AM|5060,5064
BLOOD|5065,5070
Glucose|5071,5078
-|5078,5079
96|5079,5081
UreaN|5082,5087
-|5087,5088
12|5088,5090
Creat|5091,5096
-|5096,5097
0.4|5097,5100
Na|5101,5103
-|5103,5104
135|5104,5107
<EOL>|5108,5109
K|5109,5110
-|5110,5111
3|5111,5112
.|5112,5113
1|5113,5114
*|5114,5115
Cl|5116,5118
-|5118,5119
107|5119,5122
HCO3|5123,5127
-|5127,5128
23|5128,5130
AnGap|5131,5136
-|5136,5137
8|5137,5138
<EOL>|5138,5139
_|5139,5140
_|5140,5141
_|5141,5142
11|5143,5145
:|5145,5146
43AM|5146,5150
BLOOD|5151,5156
CK|5157,5159
(|5159,5160
CPK|5160,5163
)|5163,5164
-|5164,5165
28|5165,5167
*|5167,5168
<EOL>|5168,5169
_|5169,5170
_|5170,5171
_|5171,5172
11|5173,5175
:|5175,5176
43AM|5176,5180
BLOOD|5181,5186
Lipase|5187,5193
-|5193,5194
148|5194,5197
*|5197,5198
<EOL>|5198,5199
_|5199,5200
_|5200,5201
_|5201,5202
11|5203,5205
:|5205,5206
43AM|5206,5210
BLOOD|5211,5216
CK|5217,5219
-|5219,5220
MB|5220,5222
-|5222,5223
6|5223,5224
cTropnT|5225,5232
-|5232,5233
0|5233,5234
.|5234,5235
02|5235,5237
*|5237,5238
<EOL>|5238,5239
_|5239,5240
_|5240,5241
_|5241,5242
02|5243,5245
:|5245,5246
46AM|5246,5250
BLOOD|5251,5256
Calcium|5257,5264
-|5264,5265
8|5265,5266
.|5266,5267
1|5267,5268
*|5268,5269
Phos|5270,5274
-|5274,5275
3.2|5275,5278
Mg|5279,5281
-|5281,5282
1.8|5282,5285
Iron|5286,5290
-|5290,5291
17|5291,5293
*|5293,5294
<EOL>|5294,5295
_|5295,5296
_|5296,5297
_|5297,5298
02|5299,5301
:|5301,5302
46AM|5302,5306
BLOOD|5307,5312
calTIBC|5313,5320
-|5320,5321
222|5321,5324
*|5324,5325
VitB12|5326,5332
-|5332,5333
726|5333,5336
Folate|5337,5343
-|5343,5344
15.3|5344,5348
<EOL>|5349,5350
Ferritn|5350,5357
-|5357,5358
101|5358,5361
TRF|5362,5365
-|5365,5366
171|5366,5369
*|5369,5370
<EOL>|5370,5371
_|5371,5372
_|5372,5373
_|5373,5374
11|5375,5377
:|5377,5378
43AM|5378,5382
BLOOD|5383,5388
ASA|5389,5392
-|5392,5393
NEG|5393,5396
Ethanol|5397,5404
-|5404,5405
NEG|5405,5408
Acetmnp|5409,5416
-|5416,5417
NEG|5417,5420
<EOL>|5421,5422
Bnzodzp|5422,5429
-|5429,5430
NEG|5430,5433
Barbitr|5434,5441
-|5441,5442
NEG|5442,5445
Tricycl|5446,5453
-|5453,5454
NEG|5454,5457
<EOL>|5457,5458
_|5458,5459
_|5459,5460
_|5460,5461
11|5462,5464
:|5464,5465
44AM|5465,5469
BLOOD|5470,5475
pO2|5476,5479
-|5479,5480
128|5480,5483
*|5483,5484
pCO2|5485,5489
-|5489,5490
70|5490,5492
*|5492,5493
pH|5494,5496
-|5496,5497
7|5497,5498
.|5498,5499
22|5499,5501
*|5501,5502
calTCO2|5503,5510
-|5510,5511
30|5511,5513
<EOL>|5514,5515
Base|5515,5519
XS|5520,5522
-|5522,5523
0|5523,5524
Comment|5525,5532
-|5532,5533
GREEN|5533,5538
TOP|5539,5542
<EOL>|5542,5543
_|5543,5544
_|5544,5545
_|5545,5546
11|5547,5549
:|5549,5550
44AM|5550,5554
BLOOD|5555,5560
Glucose|5561,5568
-|5568,5569
132|5569,5572
*|5572,5573
Lactate|5574,5581
-|5581,5582
0.9|5582,5585
Na|5586,5588
-|5588,5589
130|5589,5592
*|5592,5593
K|5594,5595
-|5595,5596
3.6|5596,5599
<EOL>|5600,5601
Cl|5601,5603
-|5603,5604
98|5604,5606
<EOL>|5606,5607
_|5607,5608
_|5608,5609
_|5609,5610
11|5611,5613
:|5613,5614
44AM|5614,5618
BLOOD|5619,5624
Hgb|5625,5628
-|5628,5629
8|5629,5630
.|5630,5631
8|5631,5632
*|5632,5633
calcHCT|5634,5641
-|5641,5642
26|5642,5644
O2|5645,5647
Sat|5648,5651
-|5651,5652
96|5652,5654
COHgb|5655,5660
-|5660,5661
3|5661,5662
<EOL>|5663,5664
MetHgb|5664,5670
-|5670,5671
0|5671,5672
<EOL>|5672,5673
_|5673,5674
_|5674,5675
_|5675,5676
12|5677,5679
:|5679,5680
30PM|5680,5684
URINE|5685,5690
Color|5691,5696
-|5696,5697
Yellow|5697,5703
Appear|5704,5710
-|5710,5711
Hazy|5711,5715
Sp|5716,5718
_|5719,5720
_|5720,5721
_|5721,5722
<EOL>|5722,5723
_|5723,5724
_|5724,5725
_|5725,5726
12|5727,5729
:|5729,5730
30PM|5730,5734
URINE|5735,5740
Blood|5741,5746
-|5746,5747
MOD|5747,5750
Nitrite|5751,5758
-|5758,5759
POS|5759,5762
Protein|5763,5770
-|5770,5771
100|5771,5774
<EOL>|5775,5776
Glucose|5776,5783
-|5783,5784
NEG|5784,5787
Ketone|5788,5794
-|5794,5795
NEG|5795,5798
Bilirub|5799,5806
-|5806,5807
NEG|5807,5810
Urobiln|5811,5818
-|5818,5819
NEG|5819,5822
pH|5823,5825
-|5825,5826
6.5|5826,5829
Leuks|5830,5835
-|5835,5836
LG|5836,5838
<EOL>|5838,5839
_|5839,5840
_|5840,5841
_|5841,5842
12|5843,5845
:|5845,5846
30PM|5846,5850
URINE|5851,5856
RBC|5857,5860
-|5860,5861
18|5861,5863
*|5863,5864
WBC|5865,5868
-|5868,5869
104|5869,5872
*|5872,5873
Bacteri|5874,5881
-|5881,5882
MOD|5882,5885
Yeast|5886,5891
-|5891,5892
NONE|5892,5896
<EOL>|5897,5898
Epi|5898,5901
-|5901,5902
0|5902,5903
TransE|5904,5910
-|5910,5911
2|5911,5912
<EOL>|5912,5913
_|5913,5914
_|5914,5915
_|5915,5916
12|5917,5919
:|5919,5920
30PM|5920,5924
URINE|5925,5930
CastHy|5931,5937
-|5937,5938
3|5938,5939
*|5939,5940
<EOL>|5940,5941
_|5941,5942
_|5942,5943
_|5943,5944
12|5945,5947
:|5947,5948
30PM|5948,5952
URINE|5953,5958
CastHy|5959,5965
-|5965,5966
3|5966,5967
*|5967,5968
<EOL>|5968,5969
_|5969,5970
_|5970,5971
_|5971,5972
12|5973,5975
:|5975,5976
30PM|5976,5980
URINE|5981,5986
Mucous|5987,5993
-|5993,5994
RARE|5994,5998
<EOL>|5998,5999
<EOL>|5999,6000
DISCHARGE|6000,6009
LABS|6010,6014
:|6014,6015
*|6016,6017
*|6017,6018
*|6018,6019
*|6019,6020
<EOL>|6020,6021
<EOL>|6021,6022
MICROBIOLOGY|6022,6034
:|6034,6035
<EOL>|6036,6037
<EOL>|6037,6038
-|6038,6039
Urine|6039,6044
culture|6045,6052
(|6053,6054
_|6054,6055
_|6055,6056
_|6056,6057
)|6057,6058
:|6058,6059
PSEUDOMONAS|6060,6071
AERUGINOSA|6072,6082
.|6082,6083
>|6084,6085
100,000|6085,6092
<EOL>|6093,6094
ORGANISMS|6094,6103
/|6103,6104
ML|6104,6106
.|6106,6107
.|6107,6108
<EOL>|6109,6110
SENSITIVITIES|6110,6123
:|6123,6124
MIC|6125,6128
expressed|6129,6138
_|6139,6140
_|6140,6141
_|6141,6142
MCG|6143,6146
/|6146,6147
ML|6147,6149
<EOL>|6149,6150
AMIKACIN|6155,6163
-|6163,6164
-|6164,6165
-|6165,6166
-|6166,6167
-|6167,6168
-|6168,6169
-|6169,6170
-|6170,6171
-|6171,6172
-|6172,6173
-|6173,6174
-|6174,6175
-|6175,6176
-|6176,6177
<|6180,6181
=|6181,6182
2|6182,6183
S|6184,6185
<EOL>|6185,6186
CEFEPIME|6191,6199
-|6199,6200
-|6200,6201
-|6201,6202
-|6202,6203
-|6203,6204
-|6204,6205
-|6205,6206
-|6206,6207
-|6207,6208
-|6208,6209
-|6209,6210
-|6210,6211
-|6211,6212
-|6212,6213
<|6216,6217
=|6217,6218
1|6218,6219
S|6220,6221
<EOL>|6221,6222
CEFTAZIDIME|6227,6238
-|6238,6239
-|6239,6240
-|6240,6241
-|6241,6242
-|6242,6243
-|6243,6244
-|6244,6245
-|6245,6246
-|6246,6247
-|6247,6248
-|6248,6249
<|6252,6253
=|6253,6254
1|6254,6255
S|6256,6257
<EOL>|6257,6258
CIPROFLOXACIN|6263,6276
-|6276,6277
-|6277,6278
-|6278,6279
-|6279,6280
-|6280,6281
-|6281,6282
-|6282,6283
-|6283,6284
-|6284,6285
2|6290,6291
I|6292,6293
<EOL>|6293,6294
GENTAMICIN|6299,6309
-|6309,6310
-|6310,6311
-|6311,6312
-|6312,6313
-|6313,6314
-|6314,6315
-|6315,6316
-|6316,6317
-|6317,6318
-|6318,6319
-|6319,6320
-|6320,6321
=|6323,6324
>|6324,6325
16|6325,6327
R|6328,6329
<EOL>|6329,6330
MEROPENEM|6335,6344
-|6344,6345
-|6345,6346
-|6346,6347
-|6347,6348
-|6348,6349
-|6349,6350
-|6350,6351
-|6351,6352
-|6352,6353
-|6353,6354
-|6354,6355
-|6355,6356
-|6356,6357
1|6362,6363
S|6364,6365
<EOL>|6365,6366
PIPERACILLIN|6371,6383
/|6383,6384
TAZO|6384,6388
-|6388,6389
-|6389,6390
-|6390,6391
-|6391,6392
-|6392,6393
S|6400,6401
<EOL>|6401,6402
TOBRAMYCIN|6407,6417
-|6417,6418
-|6418,6419
-|6419,6420
-|6420,6421
-|6421,6422
-|6422,6423
-|6423,6424
-|6424,6425
-|6425,6426
-|6426,6427
-|6427,6428
-|6428,6429
8|6434,6435
I|6436,6437
<EOL>|6437,6438
<EOL>|6438,6439
-|6439,6440
Blood|6440,6445
culture|6446,6453
(|6454,6455
_|6455,6456
_|6456,6457
_|6457,6458
)|6458,6459
:|6459,6460
LACTOBACILLUS|6461,6474
SPECIES|6475,6482
.|6482,6483
Isolated|6484,6492
from|6493,6497
<EOL>|6498,6499
only|6499,6503
one|6504,6507
set|6508,6511
_|6512,6513
_|6513,6514
_|6514,6515
the|6516,6519
previous|6520,6528
five|6529,6533
days|6534,6538
.|6538,6539
<EOL>|6540,6541
SENSITIVITIES|6541,6554
:|6554,6555
MIC|6556,6559
expressed|6560,6569
_|6570,6571
_|6571,6572
_|6572,6573
MCG|6574,6577
/|6577,6578
ML|6578,6580
<EOL>|6580,6581
AMPICILLIN|6586,6596
-|6596,6597
-|6597,6598
-|6598,6599
-|6599,6600
-|6600,6601
-|6601,6602
-|6602,6603
-|6603,6604
-|6604,6605
-|6605,6606
-|6606,6607
-|6607,6608
1|6613,6614
S|6615,6616
<EOL>|6616,6617
GENTAMICIN|6622,6632
-|6632,6633
-|6633,6634
-|6634,6635
-|6635,6636
-|6636,6637
-|6637,6638
-|6638,6639
-|6639,6640
-|6640,6641
-|6641,6642
-|6642,6643
-|6643,6644
2|6649,6650
S|6651,6652
<EOL>|6652,6653
PENICILLIN|6658,6668
G|6669,6670
-|6670,6671
-|6671,6672
-|6672,6673
-|6673,6674
-|6674,6675
-|6675,6676
-|6676,6677
-|6677,6678
-|6678,6679
-|6679,6680
0.5|6683,6686
S|6687,6688
<EOL>|6688,6689
<EOL>|6689,6690
-|6690,6691
Sputum|6691,6697
culture|6698,6705
_|6706,6707
_|6707,6708
_|6708,6709
,|6709,6710
endotracheal|6711,6723
source|6724,6730
)|6730,6731
:|6731,6732
<EOL>|6733,6734
GRAM|6737,6741
STAIN|6742,6747
:|6747,6748
>|6749,6750
25|6750,6752
PMNs|6753,6757
and|6758,6761
<|6762,6763
10|6763,6765
epithelial|6766,6776
cells|6777,6782
/|6782,6783
100X|6783,6787
field|6788,6793
.|6793,6794
<EOL>|6795,6796
2|6802,6803
+|6803,6804
_|6807,6808
_|6808,6809
_|6809,6810
per|6811,6814
1000X|6815,6820
FIELD|6821,6826
)|6826,6827
:|6827,6828
BUDDING|6831,6838
YEAST|6839,6844
WITH|6845,6849
<EOL>|6850,6851
PSEUDOHYPHAE|6851,6863
.|6863,6864
<EOL>|6865,6866
1|6872,6873
+|6873,6874
(|6878,6879
<|6879,6880
1|6880,6881
per|6882,6885
1000X|6886,6891
FIELD|6892,6897
)|6897,6898
:|6898,6899
GRAM|6902,6906
POSITIVE|6907,6915
COCCI|6916,6921
.|6921,6922
<EOL>|6923,6924
_|6960,6961
_|6961,6962
_|6962,6963
PAIRS|6964,6969
AND|6970,6973
SINGLY|6974,6980
.|6980,6981
<EOL>|6982,6983
RESPIRATORY|6986,6997
CULTURE|6998,7005
(|7006,7007
Final|7007,7012
_|7013,7014
_|7014,7015
_|7015,7016
:|7016,7017
<EOL>|7018,7019
MODERATE|7025,7033
GROWTH|7034,7040
Commensal|7041,7050
Respiratory|7051,7062
Flora|7063,7068
.|7068,7069
<EOL>|7070,7071
YEAST|7077,7082
.|7082,7083
SPARSE|7084,7090
GROWTH|7091,7097
.|7097,7098
<EOL>|7099,7100
LEGIONELLA|7103,7113
CULTURE|7114,7121
(|7122,7123
Preliminary|7123,7134
)|7134,7135
:|7135,7136
NO|7140,7142
LEGIONELLA|7143,7153
ISOLATED|7154,7162
.|7162,7163
<EOL>|7164,7165
<EOL>|7165,7166
-|7166,7167
Urine|7167,7172
culture|7173,7180
_|7181,7182
_|7182,7183
_|7183,7184
,|7184,7185
foley|7186,7191
)|7191,7192
:|7192,7193
YEAST|7194,7199
.|7199,7200
10,000|7201,7207
-|7207,7208
100,000|7208,7215
<EOL>|7216,7217
ORGANISMS|7217,7226
/|7226,7227
ML|7227,7229
.|7229,7230
<EOL>|7230,7231
<EOL>|7231,7232
-|7232,7233
Blood|7233,7238
culture|7239,7246
_|7247,7248
_|7248,7249
_|7249,7250
,|7250,7251
final|7252,7257
)|7257,7258
:|7258,7259
NEGATIVE|7260,7268
<EOL>|7268,7269
-|7269,7270
Blood|7270,7275
culture|7276,7283
_|7284,7285
_|7285,7286
_|7286,7287
,|7287,7288
final|7289,7294
)|7294,7295
:|7295,7296
NEGATIVE|7297,7305
<EOL>|7305,7306
-|7306,7307
Blood|7307,7312
culture|7313,7320
_|7321,7322
_|7322,7323
_|7323,7324
,|7324,7325
pending|7326,7333
)|7333,7334
:|7334,7335
NO|7336,7338
GROWTH|7339,7345
TO|7346,7348
DATE|7349,7353
<EOL>|7353,7354
<EOL>|7355,7356
AP|7356,7358
CHEST|7359,7364
X-RAY|7365,7370
(|7371,7372
_|7372,7373
_|7373,7374
_|7374,7375
)|7375,7376
:|7376,7377
<EOL>|7378,7379
1.|7379,7381
Bilateral|7382,7391
pleural|7392,7399
effusion|7400,7408
,|7408,7409
right|7410,7415
greater|7416,7423
than|7424,7428
left|7429,7433
.|7433,7434
<EOL>|7435,7436
Underlying|7436,7446
<EOL>|7447,7448
consolidation|7448,7461
can|7462,7465
not|7465,7468
be|7469,7471
completely|7472,7482
excluded|7483,7491
.|7491,7492
<EOL>|7493,7494
2.|7494,7496
Endotracheal|7497,7509
tube|7510,7514
terminates|7515,7525
1.8|7526,7529
cm|7530,7532
above|7533,7538
the|7539,7542
carina|7543,7549
.|7549,7550
<EOL>|7551,7552
Recommend|7552,7561
<EOL>|7562,7563
repositioning|7563,7576
.|7576,7577
<EOL>|7578,7579
3.|7579,7581
NG|7582,7584
tube|7585,7589
terminates|7590,7600
_|7601,7602
_|7602,7603
_|7603,7604
stomach|7605,7612
with|7613,7617
sidehole|7618,7626
_|7627,7628
_|7628,7629
_|7629,7630
distal|7631,7637
<EOL>|7638,7639
esophagus|7639,7648
.|7648,7649
<EOL>|7650,7651
3.|7651,7653
Right|7654,7659
PICC|7660,7664
terminates|7665,7675
_|7676,7677
_|7677,7678
_|7678,7679
the|7680,7683
axilla|7684,7690
.|7690,7691
<EOL>|7692,7693
<EOL>|7693,7694
CT|7694,7696
HEAD|7697,7701
WITHOUT|7702,7709
CONTRAST|7710,7718
(|7719,7720
_|7720,7721
_|7721,7722
_|7722,7723
)|7723,7724
:|7724,7725
There|7726,7731
is|7732,7734
no|7735,7737
evidence|7738,7746
of|7747,7749
<EOL>|7750,7751
hemorrhage|7751,7761
,|7761,7762
edema|7763,7768
,|7768,7769
infarction|7770,7780
,|7780,7781
or|7782,7784
mass|7785,7789
effect|7790,7796
.|7796,7797
The|7798,7801
ventricles|7802,7812
<EOL>|7813,7814
and|7814,7817
sulci|7818,7823
are|7824,7827
prominent|7828,7837
,|7837,7838
suggesting|7839,7849
age|7850,7853
-|7853,7854
related|7854,7861
involutional|7862,7874
<EOL>|7875,7876
changes|7876,7883
or|7884,7886
atrophy|7887,7894
.|7894,7895
Periventricular|7896,7911
white|7912,7917
matter|7918,7924
hypodensities|7925,7938
<EOL>|7939,7940
are|7940,7943
compatible|7944,7954
with|7955,7959
chronic|7960,7967
small|7968,7973
vessel|7974,7980
ischemic|7981,7989
disease|7990,7997
.|7997,7998
Basal|7999,8004
<EOL>|8005,8006
cisterns|8006,8014
appear|8015,8021
patent|8022,8028
,|8028,8029
and|8030,8033
there|8034,8039
is|8040,8042
preservation|8043,8055
of|8056,8058
gray|8059,8063
-|8063,8064
white|8064,8069
<EOL>|8070,8071
matter|8071,8077
differentiation|8078,8093
.|8093,8094
No|8095,8097
fracture|8098,8106
is|8107,8109
identified|8110,8120
.|8120,8121
There|8122,8127
is|8128,8130
<EOL>|8131,8132
fluid|8132,8137
within|8138,8144
the|8145,8148
nasal|8149,8154
cavity|8155,8161
,|8161,8162
likely|8163,8169
secondary|8170,8179
to|8180,8182
intubated|8183,8192
<EOL>|8193,8194
state|8194,8199
.|8199,8200
Atherosclerotic|8202,8217
mural|8218,8223
calcifications|8224,8238
of|8239,8241
the|8242,8245
internal|8246,8254
<EOL>|8255,8256
carotid|8256,8263
arteries|8264,8272
are|8273,8276
present|8277,8284
.|8284,8285
The|8286,8289
visualized|8290,8300
paranasal|8301,8310
sinuses|8311,8318
,|8318,8319
<EOL>|8320,8321
mastoid|8321,8328
air|8329,8332
cells|8333,8338
,|8338,8339
and|8340,8343
middle|8344,8350
ear|8351,8354
cavities|8355,8363
are|8364,8367
otherwise|8368,8377
clear|8378,8383
.|8383,8384
<EOL>|8385,8386
Bilateral|8386,8395
ocular|8396,8402
lenses|8403,8409
have|8410,8414
been|8415,8419
replaced|8420,8428
.|8428,8429
IMPRESSION|8430,8440
:|8440,8441
No|8442,8444
<EOL>|8445,8446
intracranial|8446,8458
hemorrhage|8459,8469
or|8470,8472
mass|8473,8477
effect|8478,8484
.|8484,8485
<EOL>|8486,8487
<EOL>|8487,8488
TTE|8488,8491
(|8492,8493
_|8493,8494
_|8494,8495
_|8495,8496
)|8496,8497
:|8497,8498
The|8499,8502
left|8503,8507
atrium|8508,8514
is|8515,8517
normal|8518,8524
_|8525,8526
_|8526,8527
_|8527,8528
size|8529,8533
.|8533,8534
There|8535,8540
is|8541,8543
mild|8544,8548
<EOL>|8549,8550
(|8550,8551
non-obstructive|8551,8566
)|8566,8567
focal|8568,8573
hypertrophy|8574,8585
of|8586,8588
the|8589,8592
basal|8593,8598
septum|8599,8605
.|8605,8606
The|8607,8610
<EOL>|8611,8612
left|8612,8616
ventricular|8617,8628
cavity|8629,8635
size|8636,8640
is|8641,8643
normal|8644,8650
.|8650,8651
Left|8652,8656
ventricular|8657,8668
<EOL>|8669,8670
systolic|8670,8678
function|8679,8687
is|8688,8690
hyperdynamic|8691,8703
(|8704,8705
EF|8705,8707
=|8708,8709
75|8710,8712
%|8712,8713
)|8713,8714
.|8714,8715
Right|8716,8721
ventricular|8722,8733
<EOL>|8734,8735
chamber|8735,8742
size|8743,8747
and|8748,8751
free|8752,8756
wall|8757,8761
motion|8762,8768
are|8769,8772
normal|8773,8779
.|8779,8780
The|8781,8784
aortic|8785,8791
valve|8792,8797
<EOL>|8798,8799
leaflets|8799,8807
(|8808,8809
3|8809,8810
)|8810,8811
are|8812,8815
mildly|8816,8822
thickened|8823,8832
.|8832,8833
There|8834,8839
is|8840,8842
mild|8843,8847
aortic|8848,8854
valve|8855,8860
<EOL>|8861,8862
stenosis|8862,8870
(|8871,8872
valve|8872,8877
area|8878,8882
1.2|8883,8886
-|8886,8887
1.9|8887,8890
cm2|8890,8893
)|8893,8894
.|8894,8895
Trace|8896,8901
aortic|8902,8908
regurgitation|8909,8922
is|8923,8925
<EOL>|8926,8927
seen|8927,8931
.|8931,8932
The|8933,8936
mitral|8937,8943
valve|8944,8949
leaflets|8950,8958
are|8959,8962
mildly|8963,8969
thickened|8970,8979
.|8979,8980
There|8981,8986
is|8987,8989
<EOL>|8990,8991
severe|8991,8997
mitral|8998,9004
annular|9005,9012
calcification|9013,9026
.|9026,9027
Moderate|9028,9036
(|9037,9038
2|9038,9039
+|9039,9040
)|9040,9041
mitral|9042,9048
<EOL>|9049,9050
regurgitation|9050,9063
is|9064,9066
seen|9067,9071
.|9071,9072
[|9073,9074
Due|9074,9077
to|9078,9080
acoustic|9081,9089
shadowing|9090,9099
,|9099,9100
the|9101,9104
severity|9105,9113
<EOL>|9114,9115
of|9115,9117
mitral|9118,9124
regurgitation|9125,9138
may|9139,9142
be|9143,9145
significantly|9146,9159
UNDERestimated|9160,9174
.|9174,9175
]|9175,9176
<EOL>|9177,9178
There|9178,9183
is|9184,9186
mild|9187,9191
pulmonary|9192,9201
artery|9202,9208
systolic|9209,9217
hypertension|9218,9230
.|9230,9231
There|9232,9237
is|9238,9240
<EOL>|9241,9242
no|9242,9244
pericardial|9245,9256
effusion|9257,9265
.|9265,9266
<EOL>|9267,9268
<EOL>|9268,9269
Compared|9269,9277
with|9278,9282
the|9283,9286
prior|9287,9292
study|9293,9298
dated|9299,9304
_|9305,9306
_|9306,9307
_|9307,9308
(|9309,9310
images|9310,9316
reviewed|9317,9325
)|9325,9326
,|9326,9327
<EOL>|9328,9329
findings|9329,9337
are|9338,9341
similar|9342,9349
.|9349,9350
<EOL>|9352,9353
<EOL>|9353,9354
AP|9354,9356
UPRIGHT|9357,9364
CHEST|9365,9370
X-RAY|9371,9376
(|9377,9378
_|9378,9379
_|9379,9380
_|9380,9381
)|9381,9382
:|9382,9383
Compared|9384,9392
to|9393,9395
the|9396,9399
most|9400,9404
recent|9405,9411
<EOL>|9412,9413
study|9413,9418
,|9418,9419
there|9420,9425
is|9426,9428
improvement|9429,9440
_|9441,9442
_|9442,9443
_|9443,9444
the|9445,9448
mild|9449,9453
pulmonary|9454,9463
edema|9464,9469
and|9470,9473
<EOL>|9474,9475
decrease|9475,9483
_|9484,9485
_|9485,9486
_|9486,9487
the|9488,9491
small|9492,9497
left|9498,9502
pleural|9503,9510
effusion|9511,9519
.|9519,9520
Moderate|9521,9529
right|9530,9535
<EOL>|9536,9537
pleural|9537,9544
effusion|9545,9553
and|9554,9557
bibasilar|9558,9567
atelectasis|9568,9579
are|9580,9583
stable|9584,9590
.|9590,9591
<EOL>|9592,9593
<EOL>|9593,9594
AP|9594,9596
UPRIGHT|9597,9604
CHEST|9605,9610
X-RAY|9611,9616
(|9617,9618
_|9618,9619
_|9619,9620
_|9620,9621
)|9621,9622
:|9622,9623
Cardiac|9624,9631
size|9632,9636
is|9637,9639
normal|9640,9646
.|9646,9647
Lines|9648,9653
<EOL>|9654,9655
and|9655,9658
tubes|9659,9664
are|9665,9668
_|9669,9670
_|9670,9671
_|9671,9672
the|9673,9676
standard|9677,9685
position|9686,9694
.|9694,9695
Large|9696,9701
right|9702,9707
and|9708,9711
moderate|9712,9720
<EOL>|9721,9722
left|9722,9726
pleural|9727,9734
effusions|9735,9744
are|9745,9748
grossly|9749,9756
unchanged|9757,9766
allowing|9767,9775
the|9776,9779
<EOL>|9780,9781
differences|9781,9792
_|9793,9794
_|9794,9795
_|9795,9796
positioning|9797,9808
of|9809,9811
the|9812,9815
patient|9816,9823
.|9823,9824
Right|9825,9830
upper|9831,9836
lobe|9837,9841
<EOL>|9842,9843
opacity|9843,9850
has|9851,9854
improved|9855,9863
consistent|9864,9874
with|9875,9879
improving|9880,9889
atelectasis|9890,9901
.|9901,9902
<EOL>|9903,9904
Pleural|9904,9911
effusions|9912,9921
are|9922,9925
associated|9926,9936
with|9937,9941
atelectasis|9942,9953
,|9953,9954
larger|9955,9961
on|9962,9964
the|9965,9968
<EOL>|9969,9970
right|9970,9975
side|9976,9980
.|9980,9981
There|9982,9987
is|9988,9990
mild|9991,9995
vascular|9996,10004
congestion|10005,10015
.|10015,10016
<EOL>|10017,10018
<EOL>|10019,10020
Brief|10020,10025
Hospital|10026,10034
Course|10035,10041
:|10041,10042
<EOL>|10042,10043
HOSPITAL|10043,10051
COURSE|10052,10058
:|10058,10059
<EOL>|10059,10060
This|10060,10064
is|10065,10067
an|10068,10070
_|10071,10072
_|10072,10073
_|10073,10074
year|10075,10079
old|10080,10083
woman|10084,10089
,|10089,10090
recently|10091,10099
hospitalized|10100,10112
for|10113,10116
C|10117,10118
.|10118,10119
<EOL>|10120,10121
Difficile|10121,10130
sepsis|10131,10137
and|10138,10141
shock|10142,10147
,|10147,10148
complicated|10149,10160
by|10161,10163
readmission|10164,10175
<EOL>|10176,10177
hypoxia|10177,10184
/|10184,10185
hypercarbia|10185,10196
(|10197,10198
_|10198,10199
_|10199,10200
_|10200,10201
)|10201,10202
p|10203,10204
/|10204,10205
w|10205,10206
hypercarbic|10207,10218
respiratory|10219,10230
<EOL>|10231,10232
failure|10232,10239
and|10240,10243
urinary|10244,10251
tract|10252,10257
infection|10258,10267
.|10267,10268
<EOL>|10269,10270
.|10270,10271
<EOL>|10271,10272
#|10272,10273
Hypercarbic|10274,10285
Respiratory|10286,10297
Failure|10298,10305
:|10305,10306
Etiology|10307,10315
likely|10316,10322
<EOL>|10323,10324
multifactorial|10324,10338
,|10338,10339
primarily|10340,10349
respiratory|10350,10361
muscle|10362,10368
weakness|10369,10377
and|10378,10381
pulm|10382,10386
<EOL>|10387,10388
edema|10388,10393
with|10394,10398
pleural|10399,10406
effusions|10407,10416
as|10417,10419
noted|10420,10425
on|10426,10428
admission|10429,10438
x-ray|10439,10444
(|10445,10446
has|10446,10449
<EOL>|10450,10451
history|10451,10458
of|10459,10461
2|10462,10463
+|10463,10464
mitral|10465,10471
regurg|10472,10478
)|10478,10479
.|10479,10480
She|10481,10484
remained|10485,10493
intubated|10494,10503
for|10504,10507
most|10508,10512
of|10513,10515
<EOL>|10516,10517
her|10517,10520
MICU|10521,10525
stay|10526,10530
due|10531,10534
to|10535,10537
pulmonary|10538,10547
edema|10548,10553
and|10554,10557
respiratory|10558,10569
muscle|10570,10576
<EOL>|10577,10578
weakness|10578,10586
with|10587,10591
a|10592,10593
poor|10594,10598
negative|10599,10607
inspiratory|10608,10619
force|10620,10625
(|10626,10627
NIF|10627,10630
)|10630,10631
.|10631,10632
Her|10633,10636
NIF|10637,10640
<EOL>|10641,10642
gradually|10642,10651
improved|10652,10660
with|10661,10665
optimization|10666,10678
of|10679,10681
her|10682,10685
nutrition|10686,10695
and|10696,10699
<EOL>|10700,10701
supportive|10701,10711
care|10712,10716
.|10716,10717
Her|10718,10721
pulmonary|10722,10731
edema|10732,10737
was|10738,10741
addressed|10742,10751
with|10752,10756
<EOL>|10757,10758
aggressive|10758,10768
diuresis|10769,10777
with|10778,10782
IV|10783,10785
and|10786,10789
PO|10790,10792
Lasix|10793,10798
boluses|10799,10806
(|10807,10808
responds|10808,10816
well|10817,10821
<EOL>|10822,10823
to|10823,10825
Lasix|10826,10831
10mg|10832,10836
IV|10837,10839
)|10839,10840
.|10840,10841
With|10842,10846
treatment|10847,10856
of|10857,10859
these|10860,10865
issues|10866,10872
,|10872,10873
she|10874,10877
was|10878,10881
able|10882,10886
<EOL>|10887,10888
to|10888,10890
be|10891,10893
successfully|10894,10906
extubated|10907,10916
to|10917,10919
nasal|10920,10925
cannula|10926,10933
on|10934,10936
_|10937,10938
_|10938,10939
_|10939,10940
.|10940,10941
She|10942,10945
<EOL>|10946,10947
was|10947,10950
started|10951,10958
on|10959,10961
Lisinopril|10962,10972
5mg|10973,10976
daily|10977,10982
for|10983,10986
afterload|10987,10996
reduction|10997,11006
_|11007,11008
_|11008,11009
_|11009,11010
<EOL>|11011,11012
setting|11012,11019
of|11020,11022
her|11023,11026
2|11027,11028
+|11028,11029
MR|11030,11032
which|11033,11038
may|11039,11042
have|11043,11047
been|11048,11052
causing|11053,11060
the|11061,11064
pulmonary|11065,11074
<EOL>|11075,11076
edema|11076,11081
.|11081,11082
She|11083,11086
may|11087,11090
require|11091,11098
further|11099,11106
PRN|11107,11110
doses|11111,11116
of|11117,11119
Lasix|11120,11125
at|11126,11128
rehab|11129,11134
;|11134,11135
if|11136,11138
<EOL>|11139,11140
so|11140,11142
would|11143,11148
try|11149,11152
Lasix|11153,11158
20mg|11159,11163
PO|11164,11166
PRN|11167,11170
.|11170,11171
Consider|11172,11180
increasing|11181,11191
lisinopril|11192,11202
<EOL>|11203,11204
to|11204,11206
10mg|11207,11211
for|11212,11215
better|11216,11222
afterload|11223,11232
reduction|11233,11242
pressure|11243,11251
tolerating|11252,11262
.|11262,11263
<EOL>|11263,11264
.|11264,11265
<EOL>|11265,11266
#|11266,11267
Pseudomonas|11268,11279
UTI|11280,11283
:|11283,11284
Patient|11285,11292
grew|11293,11297
out|11298,11301
Pseudomonas|11302,11313
sensitive|11314,11323
to|11324,11326
<EOL>|11327,11328
everything|11328,11338
but|11339,11342
Gentamicin|11343,11353
on|11354,11356
_|11357,11358
_|11358,11359
_|11359,11360
urine|11361,11366
culture|11367,11374
.|11374,11375
She|11376,11379
was|11380,11383
<EOL>|11384,11385
initially|11385,11394
started|11395,11402
on|11403,11405
double|11406,11412
coverage|11413,11421
with|11422,11426
Cipro|11427,11432
/|11432,11433
Cefepime|11433,11441
while|11442,11447
<EOL>|11448,11449
cultures|11449,11457
pending|11458,11465
,|11465,11466
then|11467,11471
narrowed|11472,11480
to|11481,11483
Cefepime|11484,11492
alone|11493,11498
,|11498,11499
then|11500,11504
<EOL>|11505,11506
broadened|11506,11515
to|11516,11518
Meropenam|11519,11528
per|11529,11532
ID|11533,11535
recs|11536,11540
.|11540,11541
There|11542,11547
was|11548,11551
concern|11552,11559
that|11560,11564
<EOL>|11565,11566
Meropenam|11566,11575
caused|11576,11582
a|11583,11584
drug|11585,11589
rash|11590,11594
so|11595,11597
she|11598,11601
was|11602,11605
then|11606,11610
switched|11611,11619
to|11620,11622
IV|11623,11625
<EOL>|11626,11627
Zosyn|11627,11632
.|11632,11633
She|11634,11637
completed|11638,11647
Zosyn|11648,11653
course|11654,11660
on|11661,11663
_|11664,11665
_|11665,11666
_|11666,11667
,|11667,11668
received|11669,11677
total|11678,11683
of|11684,11686
10|11687,11689
<EOL>|11690,11691
days|11691,11695
antibiotics|11696,11707
for|11708,11711
complicated|11712,11723
UTI|11724,11727
.|11727,11728
<EOL>|11729,11730
.|11730,11731
<EOL>|11731,11732
#|11732,11733
RASH|11734,11738
:|11738,11739
pt|11740,11742
noted|11743,11748
to|11749,11751
have|11752,11756
red|11757,11760
macular|11761,11768
rash|11769,11773
on|11774,11776
extremities|11777,11788
after|11789,11794
<EOL>|11795,11796
starting|11796,11804
meropenam|11805,11814
,|11814,11815
initially|11816,11825
presumed|11826,11834
to|11835,11837
be|11838,11840
meropenam|11841,11850
drug|11851,11855
rash|11856,11860
<EOL>|11861,11862
so|11862,11864
meropenam|11865,11874
was|11875,11878
stopped|11879,11886
.|11886,11887
However|11888,11895
this|11896,11900
was|11901,11904
later|11905,11910
believed|11911,11919
to|11920,11922
be|11923,11925
<EOL>|11926,11927
more|11927,11931
consistent|11932,11942
with|11943,11947
contact|11948,11955
dermatitis|11956,11966
vs|11967,11969
.|11969,11970
eczema|11971,11977
.|11977,11978
<EOL>|11979,11980
Triamcinolone|11980,11993
cream|11994,11999
was|12000,12003
started|12004,12011
and|12012,12015
rash|12016,12020
improved|12021,12029
.|12029,12030
<EOL>|12031,12032
.|12032,12033
<EOL>|12033,12034
#|12034,12035
C|12036,12037
Diff|12038,12042
Colitis|12043,12050
:|12050,12051
Patient|12052,12059
was|12060,12063
recently|12064,12072
admitted|12073,12081
for|12082,12085
C.|12086,12088
diff|12089,12093
<EOL>|12094,12095
colitis|12095,12102
with|12103,12107
sepsis|12108,12114
.|12114,12115
Repeat|12116,12122
C|12123,12124
Diff|12125,12129
PCR|12130,12133
was|12134,12137
negative|12138,12146
during|12147,12153
last|12154,12158
<EOL>|12159,12160
hospitalization|12160,12175
.|12175,12176
She|12177,12180
completed|12181,12190
her|12191,12194
PO|12195,12197
vancomycin|12198,12208
course|12209,12215
on|12216,12218
<EOL>|12219,12220
_|12220,12221
_|12221,12222
_|12222,12223
.|12223,12224
Her|12225,12228
PO|12229,12231
vancomycin|12232,12242
was|12243,12246
continued|12247,12256
during|12257,12263
hospitalization|12264,12279
<EOL>|12280,12281
because|12281,12288
of|12289,12291
concurrent|12292,12302
treatment|12303,12312
with|12313,12317
broad|12318,12323
-|12323,12324
spectrum|12324,12332
antibiotics|12333,12344
<EOL>|12345,12346
(|12346,12347
zosyn|12347,12352
)|12352,12353
for|12354,12357
pseudomonas|12358,12369
UTI|12370,12373
.|12373,12374
Her|12375,12378
zosyn|12379,12384
was|12385,12388
completed|12389,12398
on|12399,12401
_|12402,12403
_|12403,12404
_|12404,12405
,|12405,12406
<EOL>|12407,12408
should|12408,12414
continued|12415,12424
PO|12425,12427
vanco|12428,12433
until|12434,12439
_|12440,12441
_|12441,12442
_|12442,12443
.|12443,12444
<EOL>|12445,12446
.|12446,12447
<EOL>|12447,12448
#|12448,12449
Anemia|12450,12456
:|12456,12457
Patient|12458,12465
with|12466,12470
guaiac|12471,12477
positive|12478,12486
stools|12487,12493
during|12494,12500
last|12501,12505
<EOL>|12506,12507
admission|12507,12516
,|12516,12517
new|12518,12521
from|12522,12526
past|12527,12531
admission|12532,12541
.|12541,12542
Hct|12543,12546
stable|12547,12553
_|12554,12555
_|12555,12556
_|12556,12557
high|12558,12562
_|12563,12564
_|12564,12565
_|12565,12566
<EOL>|12567,12568
throughout|12568,12578
hospitalization|12579,12594
;|12594,12595
she|12596,12599
did|12600,12603
receive|12604,12611
one|12612,12615
unit|12616,12620
pRBC|12621,12625
for|12626,12629
<EOL>|12630,12631
colloid|12631,12638
pressure|12639,12647
support|12648,12655
.|12655,12656
<EOL>|12656,12657
.|12657,12658
<EOL>|12658,12659
#|12659,12660
Hypothyroidism|12661,12675
:|12675,12676
Continued|12677,12686
on|12687,12689
levothyroxine|12690,12703
50|12704,12706
mcg|12707,12710
daily|12711,12716
.|12716,12717
<EOL>|12717,12718
.|12718,12719
<EOL>|12719,12720
#|12720,12721
GERD|12722,12726
:|12726,12727
Patient|12728,12735
previously|12736,12746
on|12747,12749
omeprazole|12750,12760
last|12761,12765
hospitalization|12766,12781
,|12781,12782
<EOL>|12783,12784
which|12784,12789
was|12790,12793
stopped|12794,12801
after|12802,12807
C.|12808,12810
diff|12811,12815
came|12816,12820
back|12821,12825
positive|12826,12834
,|12834,12835
and|12836,12839
she|12840,12843
was|12844,12847
<EOL>|12848,12849
transitioned|12849,12861
to|12862,12864
H2|12865,12867
blocker|12868,12875
for|12876,12879
GI|12880,12882
prophylaxis|12883,12894
which|12895,12900
was|12901,12904
held|12905,12909
_|12910,12911
_|12911,12912
_|12912,12913
<EOL>|12914,12915
setting|12915,12922
of|12923,12925
delirium|12926,12934
.|12934,12935
Famotidine|12936,12946
was|12947,12950
restarted|12951,12960
at|12961,12963
20mg|12964,12968
BID|12969,12972
once|12973,12977
<EOL>|12978,12979
she|12979,12982
was|12983,12986
no|12987,12989
longer|12990,12996
delirious|12997,13006
.|13006,13007
<EOL>|13008,13009
<EOL>|13009,13010
#|13010,13011
EKG|13012,13015
Changes|13016,13023
:|13023,13024
Patient|13025,13032
had|13033,13036
lateral|13037,13044
STE|13045,13048
and|13049,13052
mildly|13053,13059
elevated|13060,13068
<EOL>|13069,13070
troponin|13070,13078
x3|13079,13081
(|13082,13083
CK|13083,13085
/|13085,13086
MB|13086,13088
flat|13089,13093
)|13093,13094
on|13094,13096
admission|13097,13106
,|13106,13107
felt|13108,13112
likely|13113,13119
due|13120,13123
to|13124,13126
blunt|13127,13132
<EOL>|13133,13134
injury|13134,13140
_|13141,13142
_|13142,13143
_|13143,13144
compressions|13145,13157
_|13158,13159
_|13159,13160
_|13160,13161
ED|13162,13164
vs|13165,13167
.|13167,13168
demand|13169,13175
ischemia|13176,13184
.|13184,13185
<EOL>|13186,13187
.|13187,13188
<EOL>|13188,13189
#|13189,13190
A-line|13191,13197
:|13197,13198
patient|13199,13206
had|13207,13210
femoral|13211,13218
A-line|13219,13225
placed|13226,13232
_|13233,13234
_|13234,13235
_|13235,13236
ED|13237,13239
_|13240,13241
_|13241,13242
_|13242,13243
setting|13244,13251
of|13252,13254
<EOL>|13255,13256
her|13256,13259
hypotension|13260,13271
.|13271,13272
This|13273,13277
was|13278,13281
discontinued|13282,13294
_|13295,13296
_|13296,13297
_|13297,13298
ICU|13299,13302
and|13303,13306
replaced|13307,13315
with|13316,13320
<EOL>|13321,13322
PICC|13322,13326
.|13326,13327
She|13328,13331
had|13332,13335
one|13336,13339
set|13340,13343
of|13344,13346
BCx|13347,13350
which|13351,13356
grew|13357,13361
Lactobacillus|13362,13375
,|13375,13376
likely|13377,13383
<EOL>|13384,13385
skin|13385,13389
contaminant|13390,13401
.|13401,13402
Other|13403,13408
surveillance|13409,13421
cx|13422,13424
negative|13425,13433
.|13433,13434
<EOL>|13435,13436
.|13436,13437
<EOL>|13437,13438
TRANSITIONAL|13438,13450
ISSUES|13451,13457
:|13457,13458
<EOL>|13458,13459
-|13459,13460
Code|13461,13465
:|13465,13466
Full|13467,13471
<EOL>|13471,13472
-|13472,13473
Labs|13474,13478
:|13478,13479
She|13480,13483
should|13484,13490
have|13491,13495
a|13496,13497
daily|13498,13503
chem|13504,13508
7|13509,13510
for|13511,13514
phos|13515,13519
repletions|13520,13530
and|13531,13534
<EOL>|13535,13536
while|13536,13541
being|13542,13547
diuresed|13548,13556
<EOL>|13556,13557
-|13557,13558
Nutrition|13559,13568
:|13568,13569
Tube|13570,13574
Feeds|13575,13580
+|13581,13582
soft|13583,13587
diet|13588,13592
and|13593,13596
thin|13597,13601
liqiuds|13602,13609
<EOL>|13609,13610
<EOL>|13611,13612
Medications|13612,13623
on|13624,13626
Admission|13627,13636
:|13636,13637
<EOL>|13637,13638
1.|13638,13640
fluticasone|13641,13652
50|13653,13655
mcg|13656,13659
/|13659,13660
actuation|13660,13669
Spray|13670,13675
,|13675,13676
Suspension|13677,13687
_|13688,13689
_|13689,13690
_|13690,13691
puffs|13692,13697
BID|13698,13701
<EOL>|13702,13703
2.|13703,13705
levothyroxine|13706,13719
50|13720,13722
mcg|13723,13726
Tablet|13727,13733
Sig|13734,13737
:|13737,13738
One|13739,13742
(|13743,13744
1|13744,13745
)|13745,13746
Tablet|13747,13753
PO|13754,13756
DAILY|13757,13762
<EOL>|13764,13765
3.|13765,13767
acetaminophen|13768,13781
325|13782,13785
mg|13786,13788
Tablet|13789,13795
Sig|13796,13799
:|13799,13800
_|13801,13802
_|13802,13803
_|13803,13804
Tablets|13805,13812
q4hr|13814,13818
prn|13819,13822
<EOL>|13822,13823
4.|13823,13825
polyvinyl|13826,13835
alcohol|13836,13843
1.4|13844,13847
%|13848,13849
Drops|13850,13855
1every|13856,13862
four|13863,13867
(|13868,13869
4|13869,13870
)|13870,13871
hours|13872,13877
prn|13878,13881
<EOL>|13881,13882
5.|13882,13884
insulin|13885,13892
lispro|13893,13899
100|13900,13903
unit|13904,13908
/|13908,13909
mL|13909,13911
Solution|13912,13920
SS|13921,13923
TID|13924,13927
Sliding|13928,13935
scale|13936,13941
<EOL>|13942,13943
units|13943,13948
<EOL>|13949,13950
Subcutaneous|13950,13962
three|13963,13968
times|13969,13974
a|13975,13976
day|13977,13980
:|13980,13981
150|13982,13985
-|13985,13986
200|13986,13989
-|13990,13991
2|13992,13993
units|13994,13999
;|13999,14000
201|14001,14004
-|14004,14005
250|14005,14008
-|14009,14010
4|14011,14012
<EOL>|14013,14014
units|14014,14019
;|14019,14020
251|14021,14024
-|14024,14025
300|14025,14028
-|14029,14030
6|14031,14032
units|14033,14038
;|14038,14039
301|14040,14043
-|14043,14044
350|14044,14047
-|14048,14049
8|14050,14051
units|14052,14057
;|14057,14058
351|14059,14062
-|14062,14063
400|14063,14066
-|14067,14068
10|14069,14071
units|14072,14077
;|14077,14078
<EOL>|14079,14080
<EOL>|14080,14081
over|14081,14085
400|14086,14089
-|14090,14091
10|14092,14094
units|14095,14100
and|14101,14104
call|14105,14109
MD|14110,14112
.|14112,14113
<EOL>|14115,14116
6.|14116,14118
miconazole|14119,14129
nitrate|14130,14137
2|14138,14139
%|14140,14141
Powder|14142,14148
1|14149,14150
TID|14151,14154
prn|14155,14158
rash|14159,14163
<EOL>|14163,14164
7.|14164,14166
vancomycin|14167,14177
125|14178,14181
mg|14182,14184
Capsule|14185,14192
1|14193,14194
PO|14195,14197
Q6H|14198,14201
for|14202,14205
7|14206,14207
days|14208,14212
<EOL>|14212,14213
8.|14213,14215
heparin|14216,14223
(|14224,14225
porcine|14225,14232
)|14232,14233
5,000|14234,14239
unit|14240,14244
/|14244,14245
mL|14245,14247
Solution|14248,14256
5000|14257,14261
(|14262,14263
5000|14263,14267
)|14267,14268
TID|14269,14272
<EOL>|14272,14273
9.|14273,14275
albuterol|14276,14285
sulfate|14286,14293
2.5|14294,14297
mg|14298,14300
/|14301,14302
3|14302,14303
mL|14304,14306
(|14307,14308
0.083|14308,14313
%|14314,14315
)|14315,14316
Solution|14317,14325
1|14326,14327
q4hr|14328,14332
prn|14333,14336
<EOL>|14337,14338
SOB|14338,14341
<EOL>|14341,14342
10.|14342,14345
ipratropium|14346,14357
bromide|14358,14365
0.02|14366,14370
%|14371,14372
Solution|14373,14381
1|14382,14383
q6hr|14384,14388
prn|14389,14392
SOB|14393,14396
<EOL>|14396,14397
<EOL>|14398,14399
Discharge|14399,14408
Medications|14409,14420
:|14420,14421
<EOL>|14421,14422
1.|14422,14424
Vancomycin|14425,14435
Oral|14436,14440
Liquid|14441,14447
_|14448,14449
_|14449,14450
_|14450,14451
mg|14452,14454
PO|14455,14457
Q6H|14458,14461
Duration|14462,14470
:|14470,14471
12|14472,14474
Days|14475,14479
<EOL>|14480,14481
Last|14481,14485
day|14486,14489
=|14490,14491
_|14492,14493
_|14493,14494
_|14494,14495
<EOL>|14496,14497
2.|14497,14499
Fluticasone|14500,14511
Propionate|14512,14522
110mcg|14523,14529
2|14530,14531
PUFF|14532,14536
IH|14537,14539
BID|14540,14543
<EOL>|14544,14545
3.|14545,14547
Levothyroxine|14548,14561
Sodium|14562,14568
50|14569,14571
mcg|14572,14575
PO|14576,14578
DAILY|14579,14584
<EOL>|14585,14586
4.|14586,14588
Triamcinolone|14589,14602
Acetonide|14603,14612
0.025|14613,14618
%|14618,14619
Cream|14620,14625
1|14626,14627
Appl|14628,14632
TP|14633,14635
BID|14636,14639
<EOL>|14640,14641
pls|14641,14644
apply|14645,14650
thin|14651,14655
layer|14656,14661
to|14662,14664
rash|14665,14669
<EOL>|14670,14671
5.|14671,14673
Miconazole|14674,14684
Powder|14685,14691
2|14692,14693
%|14693,14694
1|14695,14696
Appl|14697,14701
TP|14702,14704
TID|14705,14708
<EOL>|14709,14710
to|14710,14712
groin|14713,14718
rash|14719,14723
<EOL>|14724,14725
6.|14725,14727
Insulin|14728,14735
SC|14736,14738
<EOL>|14739,14740
Sliding|14746,14753
Scale|14754,14759
<EOL>|14759,14760
<EOL>|14760,14761
Fingerstick|14761,14772
QACHS|14773,14778
<EOL>|14778,14779
Insulin|14779,14786
SC|14787,14789
Sliding|14790,14797
Scale|14798,14803
using|14804,14809
lispro|14810,14816
Insulin|14817,14824
<EOL>|14824,14825
7.|14825,14827
Lisinopril|14828,14838
5|14839,14840
mg|14841,14843
PO|14844,14846
DAILY|14847,14852
<EOL>|14853,14854
HOLD|14854,14858
for|14859,14862
SBP|14863,14866
<|14866,14867
100|14867,14870
<EOL>|14871,14872
8.|14872,14874
Famotidine|14875,14885
20|14886,14888
mg|14889,14891
PO|14892,14894
Q12H|14895,14899
<EOL>|14900,14901
9.|14901,14903
Heparin|14904,14911
5000|14912,14916
UNIT|14917,14921
SC|14922,14924
TID|14925,14928
<EOL>|14929,14930
10.|14930,14933
polyvinyl|14934,14943
alcohol|14944,14951
*|14952,14953
NF|14953,14955
*|14955,14956
1.4|14957,14960
%|14961,14962
_|14963,14964
_|14964,14965
_|14965,14966
q4|14967,14969
hours|14970,14975
PRN|14976,14979
dry|14980,14983
eyes|14984,14988
<EOL>|14989,14990
11|14990,14992
.|14992,14993
Docusate|14994,15002
Sodium|15003,15009
(|15010,15011
Liquid|15011,15017
)|15017,15018
100|15019,15022
mg|15023,15025
PO|15026,15028
BID|15029,15032
<EOL>|15033,15034
12.|15034,15037
Furosemide|15038,15048
20|15049,15051
mg|15052,15054
PO|15055,15057
DAILY|15058,15063
<EOL>|15064,15065
as|15065,15067
needed|15068,15074
for|15075,15078
volume|15079,15085
overload|15086,15094
,|15094,15095
please|15096,15102
check|15103,15108
electrolytes|15109,15121
<EOL>|15122,15123
13.|15123,15126
Albuterol|15127,15136
0.083|15137,15142
%|15142,15143
Neb|15144,15147
Soln|15148,15152
1|15153,15154
NEB|15155,15158
IH|15159,15161
Q6H|15162,15165
:|15165,15166
PRN|15166,15169
wheeze|15170,15176
<EOL>|15177,15178
14.|15178,15181
Ipratropium|15182,15193
Bromide|15194,15201
Neb|15202,15205
1|15206,15207
NEB|15208,15211
IH|15212,15214
Q6H|15215,15218
:|15218,15219
PRN|15219,15222
wheeze|15223,15229
<EOL>|15230,15231
<EOL>|15231,15232
<EOL>|15233,15234
Discharge|15234,15243
Disposition|15244,15255
:|15255,15256
<EOL>|15256,15257
Extended|15257,15265
Care|15266,15270
<EOL>|15270,15271
<EOL>|15272,15273
Facility|15273,15281
:|15281,15282
<EOL>|15282,15283
_|15283,15284
_|15284,15285
_|15285,15286
<EOL>|15286,15287
<EOL>|15288,15289
Discharge|15289,15298
Diagnosis|15299,15308
:|15308,15309
<EOL>|15309,15310
ACUTE|15310,15315
ISSUES|15316,15322
:|15322,15323
<EOL>|15323,15324
1.|15324,15326
Hypercarbic|15327,15338
respiratory|15339,15350
failure|15351,15358
<EOL>|15358,15359
2.|15359,15361
Sepsis|15362,15368
due|15369,15372
to|15373,15375
urinary|15376,15383
source|15384,15390
<EOL>|15390,15391
3.|15391,15393
Recurrent|15394,15403
C.|15404,15406
difficile|15407,15416
colitis|15417,15424
<EOL>|15424,15425
<EOL>|15425,15426
CHRONIC|15426,15433
ISSUES|15434,15440
:|15440,15441
<EOL>|15442,15443
1.|15443,15445
Hypothyroidism|15446,15460
<EOL>|15460,15461
2.|15461,15463
Chronic|15464,15471
anemia|15472,15478
<EOL>|15478,15479
3.|15479,15481
Mitral|15482,15488
regurgitation|15489,15502
<EOL>|15502,15503
4.|15503,15505
Osteoporosis|15506,15518
<EOL>|15518,15519
5.|15519,15521
Sjogren|15522,15529
syndrome|15530,15538
<EOL>|15538,15539
<EOL>|15539,15540
<EOL>|15541,15542
Discharge|15542,15551
Condition|15552,15561
:|15561,15562
<EOL>|15562,15563
Mental|15563,15569
Status|15570,15576
:|15576,15577
Clear|15578,15583
and|15584,15587
coherent|15588,15596
.|15596,15597
<EOL>|15597,15598
Level|15598,15603
of|15604,15606
Consciousness|15607,15620
:|15620,15621
Alert|15622,15627
and|15628,15631
interactive|15632,15643
.|15643,15644
<EOL>|15644,15645
Activity|15645,15653
Status|15654,15660
:|15660,15661
Out|15662,15665
of|15666,15668
Bed|15669,15672
with|15673,15677
assistance|15678,15688
to|15689,15691
chair|15692,15697
or|15698,15700
<EOL>|15701,15702
wheelchair|15702,15712
.|15712,15713
<EOL>|15713,15714
<EOL>|15714,15715
<EOL>|15716,15717
Discharge|15717,15726
Instructions|15727,15739
:|15739,15740
<EOL>|15740,15741
Dear|15741,15745
Ms.|15746,15749
_|15750,15751
_|15751,15752
_|15752,15753
,|15753,15754
<EOL>|15755,15756
<EOL>|15756,15757
It|15757,15759
was|15760,15763
a|15764,15765
pleasure|15766,15774
participating|15775,15788
_|15789,15790
_|15790,15791
_|15791,15792
your|15793,15797
care|15798,15802
at|15803,15805
_|15806,15807
_|15807,15808
_|15808,15809
<EOL>|15810,15811
_|15811,15812
_|15812,15813
_|15813,15814
.|15814,15815
You|15816,15819
were|15820,15824
admitted|15825,15833
to|15834,15836
the|15837,15840
hospital|15841,15849
with|15850,15854
<EOL>|15855,15856
respiratory|15856,15867
failure|15868,15875
requiring|15876,15885
intubation|15886,15896
and|15897,15900
mechanical|15901,15911
<EOL>|15912,15913
ventilation|15913,15924
.|15924,15925
This|15926,15930
was|15931,15934
likely|15935,15941
due|15942,15945
to|15946,15948
a|15949,15950
combination|15951,15962
of|15963,15965
severe|15966,15972
<EOL>|15973,15974
weakness|15974,15982
caused|15983,15989
by|15990,15992
chronic|15993,16000
illness|16001,16008
,|16008,16009
pleural|16010,16017
effusions|16018,16027
and|16028,16031
<EOL>|16032,16033
pulmonary|16033,16042
edema|16043,16048
(|16049,16050
fluid|16050,16055
_|16056,16057
_|16057,16058
_|16058,16059
the|16060,16063
lungs|16064,16069
)|16069,16070
.|16070,16071
You|16072,16075
were|16076,16080
also|16081,16085
found|16086,16091
to|16092,16094
<EOL>|16095,16096
have|16096,16100
a|16101,16102
urinary|16103,16110
tract|16111,16116
infection|16117,16126
causing|16127,16134
sepsis|16135,16141
(|16142,16143
bloodstream|16143,16154
<EOL>|16155,16156
infection|16156,16165
)|16165,16166
,|16166,16167
which|16168,16173
likely|16174,16180
also|16181,16185
contributed|16186,16197
to|16198,16200
your|16201,16205
respiratory|16206,16217
<EOL>|16218,16219
failure|16219,16226
.|16226,16227
You|16228,16231
were|16232,16236
treated|16237,16244
with|16245,16249
antibiotics|16250,16261
,|16261,16262
your|16263,16267
symptoms|16268,16276
and|16277,16280
<EOL>|16281,16282
breathing|16282,16291
improved|16292,16300
,|16300,16301
and|16302,16305
you|16306,16309
were|16310,16314
successfully|16315,16327
extubated|16328,16337
on|16338,16340
_|16341,16342
_|16342,16343
_|16343,16344
.|16344,16345
<EOL>|16346,16347
You|16347,16350
will|16351,16355
be|16356,16358
discharged|16359,16369
to|16370,16372
rehab|16373,16378
where|16379,16384
you|16385,16388
will|16389,16393
receive|16394,16401
intensive|16402,16411
<EOL>|16412,16413
physical|16413,16421
therapy|16422,16429
and|16430,16433
your|16434,16438
nutrition|16439,16448
will|16449,16453
be|16454,16456
optimized|16457,16466
to|16467,16469
help|16470,16474
<EOL>|16475,16476
you|16476,16479
continue|16480,16488
regaining|16489,16498
strength|16499,16507
.|16507,16508
<EOL>|16509,16510
.|16510,16511
<EOL>|16511,16512
When|16512,16516
you|16517,16520
are|16521,16524
discharged|16525,16535
from|16536,16540
rehab|16541,16546
,|16546,16547
you|16548,16551
will|16552,16556
need|16557,16561
to|16562,16564
follow|16565,16571
up|16572,16574
<EOL>|16575,16576
with|16576,16580
your|16581,16585
primary|16586,16593
care|16594,16598
doctor|16599,16605
_|16606,16607
_|16607,16608
_|16608,16609
.|16609,16610
<EOL>|16611,16612
.|16612,16613
<EOL>|16613,16614
We|16614,16616
made|16617,16621
the|16622,16625
following|16626,16635
changes|16636,16643
to|16644,16646
your|16647,16651
medications|16652,16663
:|16663,16664
<EOL>|16665,16666
1.|16666,16668
STARTED|16669,16676
famotidine|16677,16687
20mg|16688,16692
by|16693,16695
mouth|16696,16701
twice|16702,16707
daily|16708,16713
for|16714,16717
heartburn|16718,16727
<EOL>|16727,16728
2.|16728,16730
STARTED|16731,16738
triamcinolone|16739,16752
acetonide|16753,16762
0.025|16763,16768
%|16768,16769
cream|16770,16775
three|16776,16781
times|16782,16787
<EOL>|16788,16789
daily|16789,16794
for|16795,16798
rash|16799,16803
<EOL>|16803,16804
3.|16804,16806
RESTARTED|16807,16816
lisinopril|16817,16827
5mg|16828,16831
by|16832,16834
mouth|16835,16840
daily|16841,16846
for|16847,16850
high|16851,16855
blood|16856,16861
<EOL>|16862,16863
pressure|16863,16871
and|16872,16875
heart|16876,16881
failure|16882,16889
<EOL>|16889,16890
4.|16890,16892
STARTED|16893,16900
docusate|16901,16909
(|16910,16911
Colace|16911,16917
)|16917,16918
100mg|16919,16924
by|16925,16927
mouth|16928,16933
twice|16934,16939
daily|16940,16945
for|16946,16949
<EOL>|16950,16951
constipation|16951,16963
<EOL>|16963,16964
5.|16964,16966
CONTINUED|16967,16976
vancomycin|16977,16987
oral|16988,16992
liquid|16993,16999
_|17000,17001
_|17001,17002
_|17002,17003
by|17004,17006
mouth|17007,17012
every|17013,17018
6|17019,17020
hours|17021,17026
<EOL>|17027,17028
(|17028,17029
last|17029,17033
day|17034,17037
=|17038,17039
_|17040,17041
_|17041,17042
_|17042,17043
<EOL>|17044,17045
6.|17045,17047
START|17048,17053
lasix|17054,17059
po|17060,17062
20mg|17063,17067
daily|17068,17073
prn|17074,17077
volume|17078,17084
overload|17085,17093
<EOL>|17093,17094
<EOL>|17095,17096
Followup|17096,17104
Instructions|17105,17117
:|17117,17118
<EOL>|17118,17119
_|17119,17120
_|17120,17121
_|17121,17122
<EOL>|17122,17123

