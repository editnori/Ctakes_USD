 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|32,36
No|37,39
:|39,40
_|43,44
_|44,45
_|45,46
<EOL>|46,47
<EOL>|48,49
Admission|49,58
Date|59,63
:|63,64
_|66,67
_|67,68
_|68,69
Discharge|83,92
Date|93,97
:|97,98
_|101,102
_|102,103
_|103,104
<EOL>|104,105
<EOL>|106,107
Date|107,111
of|112,114
Birth|115,120
:|120,121
_|123,124
_|124,125
_|125,126
Sex|139,142
:|142,143
F|146,147
<EOL>|147,148
<EOL>|149,150
Service|150,157
:|157,158
SURGERY|159,166
<EOL>|166,167
<EOL>|168,169
IV|181,183
Dye|184,187
,|187,188
Iodine|189,195
Containing|196,206
<EOL>|206,207
<EOL>|208,209
Attending|209,218
:|218,219
_|220,221
_|221,222
_|222,223
.|223,224
<EOL>|224,225
<EOL>|226,227
nausea|244,250
,|250,251
vomiting|252,260
x|261,262
1|263,264
day|265,268
<EOL>|268,269
<EOL>|270,271
Major|271,276
Surgical|277,285
or|286,288
Invasive|289,297
Procedure|298,307
:|307,308
<EOL>|308,309
none|309,313
<EOL>|313,314
<EOL>|315,316
_|344,345
_|345,346
_|346,347
s|348,349
/|349,350
p|350,351
sigmoid|352,359
colectomy|360,369
for|370,373
recurrent|374,383
diverticulitis|384,398
on|399,401
_|402,403
_|403,404
_|404,405
<EOL>|406,407
discharged|407,417
home|418,422
on|423,425
_|426,427
_|427,428
_|428,429
after|430,435
tolerating|436,446
a|447,448
low|449,452
residue|453,460
diet|461,465
<EOL>|466,467
and|467,470
po|471,473
antibiotics|474,485
for|486,489
a|490,491
wound|492,497
infection|498,507
.|507,508
She|510,513
returned|514,522
one|523,526
week|527,531
<EOL>|532,533
after|533,538
discharge|539,548
with|549,553
1|554,555
day|556,559
of|560,562
intense|563,570
nausea|571,577
and|578,581
emesis|582,588
<EOL>|589,590
(|590,591
non-bloody|591,601
,|601,602
non-biliary|603,614
)|614,615
.|615,616
The|618,621
nausea|622,628
is|629,631
associated|632,642
with|643,647
a|648,649
<EOL>|650,651
slight|651,657
increase|658,666
in|667,669
epigastric|670,680
abdominal|681,690
pain|691,695
without|696,703
any|704,707
<EOL>|708,709
significant|709,720
tenderness|721,731
on|732,734
exam|735,739
.|739,740
<EOL>|741,742
<EOL>|743,744
diverticulitis|766,780
s|781,782
/|782,783
p|783,784
lap|785,788
sigmoid|789,796
colectomy|797,806
c|807,808
/|808,809
b|809,810
wound|811,816
infection|817,826
<EOL>|827,828
Migraines|828,837
<EOL>|837,838
Left|838,842
finger|843,849
cellulitis|850,860
<EOL>|860,861
<EOL>|862,863
:|877,878
<EOL>|878,879
_|879,880
_|880,881
_|881,882
<EOL>|882,883
:|897,898
<EOL>|898,899
father|899,905
with|906,910
h|911,912
/|912,913
o|913,914
colitis|915,922
<EOL>|922,923
<EOL>|924,925
afebrile|940,948
,|948,949
vital|950,955
signs|956,961
within|962,968
normal|969,975
limits|976,982
<EOL>|982,983
NAD|983,986
,|986,987
talkative|988,997
<EOL>|997,998
EOM|998,1001
full|1002,1006
,|1006,1007
PERRL|1008,1013
,|1013,1014
anicteric|1015,1024
sclera|1025,1031
<EOL>|1031,1032
Chest|1032,1037
clear|1038,1043
<EOL>|1043,1044
RRR|1044,1047
,|1047,1048
no|1049,1051
murmurs|1052,1059
<EOL>|1059,1060
Abdomen|1060,1067
soft|1068,1072
,|1072,1073
round|1074,1079
,|1079,1080
non-tender|1081,1091
,|1091,1092
non-distended|1093,1106
with|1107,1111
6cm|1112,1115
of|1116,1118
open|1119,1123
<EOL>|1124,1125
transverse|1125,1135
incision|1136,1144
through|1145,1152
the|1153,1156
subcutis|1157,1165
with|1166,1170
intact|1171,1177
deep|1178,1182
<EOL>|1183,1184
fascia|1184,1190
;|1190,1191
no|1192,1194
erythema|1195,1203
or|1204,1206
induration|1207,1217
;|1217,1218
minimal|1219,1226
serous|1227,1233
output|1234,1240
.|1240,1241
<EOL>|1243,1244
_|1244,1245
_|1245,1246
_|1246,1247
without|1248,1255
edema|1256,1261
,|1261,1262
2|1263,1264
+|1264,1265
DP|1266,1268
pulses|1269,1275
<EOL>|1275,1276
<EOL>|1277,1278
Pertinent|1278,1287
Results|1288,1295
:|1295,1296
<EOL>|1296,1297
CT|1297,1299
ABDOMEN|1300,1307
W|1308,1309
/|1309,1310
O|1310,1311
CONTRAST|1312,1320
_|1322,1323
_|1323,1324
_|1324,1325
6|1326,1327
:|1327,1328
_|1328,1329
_|1329,1330
_|1330,1331
BDOMEN|1331,1337
W|1338,1339
/|1339,1340
O|1340,1341
CONTRAST|1342,1350
;|1350,1351
CT|1352,1354
PELVIS|1355,1361
W|1362,1363
/|1363,1364
O|1364,1365
CONTRAST|1366,1374
<EOL>|1374,1375
<EOL>|1375,1376
Reason|1376,1382
:|1382,1383
r|1384,1385
/|1385,1386
o|1386,1387
abscess|1388,1395
-|1395,1396
NO|1396,1398
IV|1399,1401
contrast|1402,1410
,|1410,1411
PO|1412,1414
only|1415,1419
<EOL>|1420,1421
Field|1421,1426
of|1427,1429
view|1430,1434
:|1434,1435
40|1436,1438
<EOL>|1438,1439
<EOL>|1439,1440
UNDERLYING|1440,1450
MEDICAL|1451,1458
CONDITION|1459,1468
:|1468,1469
<EOL>|1469,1470
_|1470,1471
_|1471,1472
_|1472,1473
year|1474,1478
old|1479,1482
woman|1483,1488
with|1489,1493
h|1494,1495
/|1495,1496
o|1496,1497
divertic|1498,1506
s|1507,1508
/|1508,1509
p|1509,1510
colectomy|1511,1520
here|1521,1525
with|1526,1530
<EOL>|1531,1532
elevated|1532,1540
WBC|1541,1544
and|1545,1548
nausea|1549,1555
<EOL>|1556,1557
REASON|1557,1563
FOR|1564,1567
THIS|1568,1572
EXAMINATION|1573,1584
:|1584,1585
<EOL>|1585,1586
r|1586,1587
/|1587,1588
o|1588,1589
abscess|1590,1597
-|1597,1598
NO|1598,1600
IV|1601,1603
contrast|1604,1612
,|1612,1613
PO|1614,1616
only|1617,1621
<EOL>|1622,1623
CONTRAINDICATIONS|1623,1640
for|1641,1644
IV|1645,1647
CONTRAST|1648,1656
:|1656,1657
RF|1658,1660
<EOL>|1660,1661
<EOL>|1661,1662
INDICATION|1662,1672
:|1672,1673
_|1674,1675
_|1675,1676
_|1676,1677
woman|1678,1683
with|1684,1688
elevated|1689,1697
white|1698,1703
blood|1704,1709
cell|1710,1714
<EOL>|1715,1716
count|1716,1721
and|1722,1725
nausea|1726,1732
,|1732,1733
history|1734,1741
of|1742,1744
recent|1745,1751
colectomy|1752,1761
for|1762,1765
recurrent|1766,1775
<EOL>|1776,1777
diverticulitis|1777,1791
.|1791,1792
<EOL>|1792,1793
<EOL>|1793,1794
COMPARISON|1794,1804
:|1804,1805
CT|1806,1808
abdomen|1809,1816
and|1817,1820
pelvis|1821,1827
of|1828,1830
_|1831,1832
_|1832,1833
_|1833,1834
.|1834,1835
<EOL>|1835,1836
<EOL>|1836,1837
TECHNIQUE|1837,1846
:|1846,1847
MDCT|1848,1852
acquired|1853,1861
axial|1862,1867
images|1868,1874
were|1875,1879
obtained|1880,1888
through|1889,1896
the|1897,1900
<EOL>|1901,1902
abdomen|1902,1909
and|1910,1913
pelvis|1914,1920
after|1921,1926
the|1927,1930
administration|1931,1945
of|1946,1948
oral|1949,1953
contrast|1954,1962
.|1962,1963
No|1964,1966
<EOL>|1967,1968
intravenous|1968,1979
contrast|1980,1988
was|1989,1992
administered|1993,2005
.|2005,2006
Multiplanar|2007,2018
reformatted|2019,2030
<EOL>|2031,2032
images|2032,2038
were|2039,2043
also|2044,2048
obtained|2049,2057
.|2057,2058
<EOL>|2058,2059
<EOL>|2059,2060
:|2068,2069
<EOL>|2070,2071
<EOL>|2071,2072
The|2072,2075
lung|2076,2080
bases|2081,2086
are|2087,2090
clear|2091,2096
.|2096,2097
A|2098,2099
4|2100,2101
-|2101,2102
mm|2102,2104
calcified|2105,2114
granuloma|2115,2124
in|2125,2127
the|2128,2131
<EOL>|2132,2133
right|2133,2138
lung|2139,2143
base|2144,2148
is|2149,2151
unchanged|2152,2161
.|2161,2162
Limited|2163,2170
images|2171,2177
of|2178,2180
the|2181,2184
heart|2185,2190
are|2191,2194
<EOL>|2195,2196
unremarkable|2196,2208
.|2208,2209
There|2210,2215
is|2216,2218
no|2219,2221
pericardial|2222,2233
effusion|2234,2242
.|2242,2243
<EOL>|2243,2244
<EOL>|2244,2245
In|2245,2247
the|2248,2251
abdomen|2252,2259
,|2259,2260
the|2261,2264
liver|2265,2270
,|2270,2271
gallbladder|2272,2283
,|2283,2284
spleen|2285,2291
,|2291,2292
kidneys|2293,2300
,|2300,2301
adrenal|2302,2309
<EOL>|2310,2311
glands|2311,2317
,|2317,2318
pancreas|2319,2327
,|2327,2328
stomach|2329,2336
,|2336,2337
and|2338,2341
intra-abdominal|2342,2357
loops|2358,2363
of|2364,2366
small|2367,2372
<EOL>|2373,2374
and|2374,2377
large|2378,2383
bowel|2384,2389
are|2390,2393
unremarkable|2394,2406
.|2406,2407
There|2408,2413
is|2414,2416
no|2417,2419
mesenteric|2420,2430
<EOL>|2431,2432
lymphadenopathy|2432,2447
.|2447,2448
There|2449,2454
is|2455,2457
no|2458,2460
free|2461,2465
fluid|2466,2471
or|2472,2474
free|2475,2479
air|2480,2483
in|2484,2486
the|2487,2490
<EOL>|2491,2492
abdomen|2492,2499
.|2499,2500
Immediately|2501,2512
adjacent|2513,2521
to|2522,2524
the|2525,2528
left|2529,2533
common|2534,2540
iliac|2541,2546
artery|2547,2553
,|2553,2554
<EOL>|2555,2556
is|2556,2558
a|2559,2560
linear|2561,2567
focus|2568,2573
of|2574,2576
hyper|2577,2582
-|2582,2583
attenuating|2583,2594
material|2595,2603
,|2603,2604
with|2605,2609
the|2610,2613
<EOL>|2614,2615
appearance|2615,2625
of|2626,2628
suture|2629,2635
material|2636,2644
,|2644,2645
largely|2646,2653
unchanged|2654,2663
from|2664,2668
the|2669,2672
prior|2673,2678
<EOL>|2679,2680
examination|2680,2691
.|2691,2692
<EOL>|2692,2693
<EOL>|2693,2694
In|2694,2696
the|2697,2700
pelvis|2701,2707
,|2707,2708
suture|2709,2715
material|2716,2724
is|2725,2727
seen|2728,2732
in|2733,2735
the|2736,2739
distal|2740,2746
sigmoid|2747,2754
<EOL>|2755,2756
colon|2756,2761
,|2761,2762
unchanged|2763,2772
in|2773,2775
appearance|2776,2786
from|2787,2791
prior|2792,2797
examination|2798,2809
and|2810,2813
<EOL>|2814,2815
consistent|2815,2825
with|2826,2830
colonic|2831,2838
anastomosis|2839,2850
.|2850,2851
There|2852,2857
is|2858,2860
no|2861,2863
evidence|2864,2872
of|2873,2875
<EOL>|2876,2877
stricture|2877,2886
or|2887,2889
obstruction|2890,2901
at|2902,2904
this|2905,2909
site|2910,2914
.|2914,2915
There|2916,2921
is|2922,2924
no|2925,2927
local|2928,2933
fluid|2934,2939
<EOL>|2940,2941
collection|2941,2951
to|2952,2954
indicate|2955,2963
abscess|2964,2971
.|2971,2972
There|2973,2978
are|2979,2982
no|2983,2985
signs|2986,2991
of|2992,2994
<EOL>|2995,2996
inflammation|2996,3008
.|3008,3009
The|3010,3013
intrapelvic|3014,3025
loops|3026,3031
of|3032,3034
small|3035,3040
and|3041,3044
large|3045,3050
bowel|3051,3056
are|3057,3060
<EOL>|3061,3062
unremarkable|3062,3074
,|3074,3075
containing|3076,3086
air|3087,3090
and|3091,3094
stool|3095,3100
in|3101,3103
a|3104,3105
normal|3106,3112
pattern|3113,3120
<EOL>|3121,3122
without|3122,3129
bowel|3130,3135
dilatation|3136,3146
.|3146,3147
The|3148,3151
appendix|3152,3160
is|3161,3163
visualized|3164,3174
and|3175,3178
is|3179,3181
<EOL>|3182,3183
normal|3183,3189
.|3189,3190
The|3191,3194
urinary|3195,3202
bladder|3203,3210
,|3210,3211
uterus|3212,3218
,|3218,3219
and|3220,3223
adnexa|3224,3230
are|3231,3234
<EOL>|3235,3236
unremarkable|3236,3248
.|3248,3249
There|3250,3255
are|3256,3259
no|3260,3262
abnormally|3263,3273
enlarged|3274,3282
lymph|3283,3288
nodes|3289,3294
in|3295,3297
<EOL>|3298,3299
the|3299,3302
pelvis|3303,3309
.|3309,3310
A|3311,3312
fat|3313,3316
-|3316,3317
containing|3317,3327
left|3328,3332
inguinal|3333,3341
hernia|3342,3348
is|3349,3351
unchanged|3352,3361
.|3361,3362
<EOL>|3362,3363
<EOL>|3363,3364
Examination|3364,3375
of|3376,3378
soft|3379,3383
tissues|3384,3391
reveals|3392,3399
stranding|3400,3409
and|3410,3413
subcutaneous|3414,3426
<EOL>|3427,3428
air|3428,3431
of|3432,3434
the|3435,3438
soft|3439,3443
tissues|3444,3451
along|3452,3457
the|3458,3461
midline|3462,3469
lower|3470,3475
anterior|3476,3484
<EOL>|3485,3486
abdominal|3486,3495
wall|3496,3500
,|3500,3501
slightly|3502,3510
larger|3511,3517
in|3518,3520
size|3521,3525
than|3526,3530
on|3531,3533
the|3534,3537
prior|3538,3543
<EOL>|3544,3545
examination|3545,3556
of|3557,3559
approximately|3560,3573
2|3574,3575
weeks|3576,3581
ago|3582,3585
.|3585,3586
Additionally|3587,3599
,|3599,3600
a|3601,3602
small|3603,3608
<EOL>|3609,3610
focus|3610,3615
of|3616,3618
fluid|3619,3624
attenuating|3625,3636
material|3637,3645
now|3646,3649
extends|3650,3657
from|3658,3662
the|3663,3666
<EOL>|3667,3668
abdominal|3668,3677
wall|3678,3682
musculature|3683,3694
through|3695,3702
the|3703,3706
subcutaneous|3707,3719
tissues|3720,3727
,|3727,3728
and|3729,3732
<EOL>|3733,3734
appears|3734,3741
to|3742,3744
drain|3745,3750
into|3751,3755
an|3756,3758
external|3759,3767
collecting|3768,3778
device|3779,3785
.|3785,3786
No|3787,3789
discrete|3790,3798
<EOL>|3799,3800
fluid|3800,3805
collection|3806,3816
is|3817,3819
identified|3820,3830
to|3831,3833
indicate|3834,3842
abscess|3843,3850
formation|3851,3860
,|3860,3861
or|3862,3864
<EOL>|3865,3866
that|3866,3870
would|3871,3876
be|3877,3879
amenable|3880,3888
to|3889,3891
drainage|3892,3900
.|3900,3901
However|3902,3909
,|3909,3910
this|3911,3915
appearance|3916,3926
<EOL>|3927,3928
suggests|3928,3936
continued|3937,3946
cellulitis|3947,3957
.|3957,3958
<EOL>|3958,3959
<EOL>|3959,3960
Examination|3960,3971
of|3972,3974
osseous|3975,3982
structures|3983,3993
reveals|3994,4001
mild|4002,4006
degenerative|4007,4019
<EOL>|4020,4021
disease|4021,4028
at|4029,4031
L5|4032,4034
-|4034,4035
S1|4035,4037
and|4038,4041
are|4042,4045
otherwise|4046,4055
unremarkable|4056,4068
.|4068,4069
<EOL>|4069,4070
<EOL>|4070,4071
1.|4083,4085
Stable|4086,4092
appearance|4093,4103
of|4104,4106
sigmoid|4107,4114
colon|4115,4120
anastomosis|4121,4132
without|4133,4140
<EOL>|4141,4142
obstruction|4142,4153
or|4154,4156
abscess|4157,4164
formation|4165,4174
.|4174,4175
<EOL>|4175,4176
2.|4176,4178
Stranding|4179,4188
and|4189,4192
subcutaneous|4193,4205
air|4206,4209
along|4210,4215
the|4216,4219
lower|4220,4225
abdominal|4226,4235
wall|4236,4240
<EOL>|4241,4242
in|4242,4244
the|4245,4248
midline|4249,4256
,|4256,4257
indicating|4258,4268
cellulitis|4269,4279
,|4279,4280
but|4281,4284
without|4285,4292
discrete|4293,4301
or|4302,4304
<EOL>|4305,4306
drainable|4306,4315
fluid|4316,4321
collection|4322,4332
<EOL>|4332,4333
<EOL>|4333,4334
The|4334,4337
study|4338,4343
and|4344,4347
the|4348,4351
report|4352,4358
were|4359,4363
reviewed|4364,4372
by|4373,4375
the|4376,4379
staff|4380,4385
radiologist|4386,4397
.|4397,4398
<EOL>|4398,4399
_|4399,4400
_|4400,4401
_|4401,4402
.|4402,4403
_|4404,4405
_|4405,4406
_|4406,4407
<EOL>|4407,4408
_|4408,4409
_|4409,4410
_|4410,4411
.|4411,4412
_|4413,4414
_|4414,4415
_|4415,4416
<EOL>|4416,4417
_|4417,4418
_|4418,4419
_|4419,4420
.|4420,4421
_|4422,4423
_|4423,4424
_|4424,4425
:|4425,4426
SUN|4427,4430
_|4431,4432
_|4432,4433
_|4433,4434
9|4435,4436
:|4436,4437
36|4437,4439
AM|4440,4442
<EOL>|4442,4443
_|4443,4444
_|4444,4445
_|4445,4446
_|4446,4447
_|4447,4448
_|4448,4449
_|4449,4450
_|4450,4451
_|4451,4452
_|4452,4453
_|4453,4454
_|4454,4455
_|4455,4456
_|4456,4457
_|4457,4458
_|4458,4459
_|4459,4460
_|4460,4461
_|4461,4462
_|4462,4463
_|4463,4464
_|4464,4465
_|4465,4466
_|4466,4467
_|4467,4468
_|4468,4469
_|4469,4470
_|4470,4471
_|4471,4472
_|4472,4473
_|4473,4474
_|4474,4475
_|4475,4476
_|4476,4477
_|4477,4478
_|4478,4479
_|4479,4480
_|4480,4481
_|4481,4482
_|4482,4483
_|4483,4484
_|4484,4485
_|4485,4486
_|4486,4487
<EOL>|4487,4488
<EOL>|4488,4489
_|4489,4490
_|4490,4491
_|4491,4492
03|4493,4495
:|4495,4496
45AM|4496,4500
URINE|4501,4506
COLOR|4508,4513
-|4513,4514
Straw|4514,4519
APPEAR|4520,4526
-|4526,4527
Clear|4527,4532
SP|4533,4535
_|4536,4537
_|4537,4538
_|4538,4539
<EOL>|4539,4540
_|4540,4541
_|4541,4542
_|4542,4543
03|4544,4546
:|4546,4547
45AM|4547,4551
URINE|4552,4557
BLOOD|4559,4564
-|4564,4565
NEG|4565,4568
NITRITE|4569,4576
-|4576,4577
NEG|4577,4580
PROTEIN|4581,4588
-|4588,4589
NEG|4589,4592
<EOL>|4593,4594
GLUCOSE|4594,4601
-|4601,4602
NEG|4602,4605
KETONE|4606,4612
-|4612,4613
NEG|4613,4616
BILIRUBIN|4617,4626
-|4626,4627
NEG|4627,4630
UROBILNGN|4631,4640
-|4640,4641
NEG|4641,4644
PH|4645,4647
-|4647,4648
7.0|4648,4651
<EOL>|4652,4653
LEUK|4653,4657
-|4657,4658
NEG|4658,4661
<EOL>|4661,4662
_|4662,4663
_|4663,4664
_|4664,4665
02|4666,4668
:|4668,4669
20AM|4669,4673
GLUCOSE|4676,4683
-|4683,4684
124|4684,4687
*|4687,4688
UREA|4689,4693
N|4694,4695
-|4695,4696
20|4696,4698
CREAT|4699,4704
-|4704,4705
1|4705,4706
.|4706,4707
4|4707,4708
*|4708,4709
SODIUM|4710,4716
-|4716,4717
138|4717,4720
<EOL>|4721,4722
POTASSIUM|4722,4731
-|4731,4732
4.8|4732,4735
CHLORIDE|4736,4744
-|4744,4745
98|4745,4747
TOTAL|4748,4753
CO2|4754,4757
-|4757,4758
30|4758,4760
ANION|4761,4766
GAP|4767,4770
-|4770,4771
15|4771,4773
<EOL>|4773,4774
_|4774,4775
_|4775,4776
_|4776,4777
02|4778,4780
:|4780,4781
20AM|4781,4785
estGFR|4788,4794
-|4794,4795
Using|4795,4800
this|4801,4805
<EOL>|4805,4806
_|4806,4807
_|4807,4808
_|4808,4809
02|4810,4812
:|4812,4813
20AM|4813,4817
ALT|4820,4823
(|4823,4824
SGPT|4824,4828
)|4828,4829
-|4829,4830
38|4830,4832
AST|4833,4836
(|4836,4837
SGOT|4837,4841
)|4841,4842
-|4842,4843
20|4843,4845
ALK|4846,4849
PHOS|4850,4854
-|4854,4855
107|4855,4858
TOT|4859,4862
<EOL>|4863,4864
BILI|4864,4868
-|4868,4869
0.6|4869,4872
<EOL>|4872,4873
_|4873,4874
_|4874,4875
_|4875,4876
02|4877,4879
:|4879,4880
20AM|4880,4884
LIPASE|4887,4893
-|4893,4894
62|4894,4896
*|4896,4897
<EOL>|4897,4898
_|4898,4899
_|4899,4900
_|4900,4901
02|4902,4904
:|4904,4905
20AM|4905,4909
WBC|4912,4915
-|4915,4916
15|4916,4918
.|4918,4919
4|4919,4920
*|4920,4921
#|4921,4922
RBC|4923,4926
-|4926,4927
3|4927,4928
.|4928,4929
17|4929,4931
*|4931,4932
HGB|4933,4936
-|4936,4937
9|4937,4938
.|4938,4939
4|4939,4940
*|4940,4941
HCT|4942,4945
-|4945,4946
28|4946,4948
.|4948,4949
2|4949,4950
*|4950,4951
<EOL>|4952,4953
MCV|4953,4956
-|4956,4957
89|4957,4959
MCH|4960,4963
-|4963,4964
29.7|4964,4968
MCHC|4969,4973
-|4973,4974
33.4|4974,4978
RDW|4979,4982
-|4982,4983
13.7|4983,4987
<EOL>|4987,4988
_|4988,4989
_|4989,4990
_|4990,4991
02|4992,4994
:|4994,4995
20AM|4995,4999
NEUTS|5002,5007
-|5007,5008
85|5008,5010
.|5010,5011
8|5011,5012
*|5012,5013
LYMPHS|5014,5020
-|5020,5021
10|5021,5023
.|5023,5024
0|5024,5025
*|5025,5026
MONOS|5027,5032
-|5032,5033
2.5|5033,5036
EOS|5037,5040
-|5040,5041
1.2|5041,5044
<EOL>|5045,5046
BASOS|5046,5051
-|5051,5052
0.5|5052,5055
<EOL>|5055,5056
_|5056,5057
_|5057,5058
_|5058,5059
02|5060,5062
:|5062,5063
20AM|5063,5067
PLT|5070,5073
COUNT|5074,5079
-|5079,5080
730|5080,5083
*|5083,5084
#|5084,5085
<EOL>|5085,5086
<EOL>|5087,5088
GI|5111,5113
:|5113,5114
Admitted|5115,5123
in|5124,5126
early|5127,5132
morning|5133,5140
on|5141,5143
_|5144,5145
_|5145,5146
_|5146,5147
the|5148,5151
pt|5152,5154
was|5155,5158
made|5159,5163
NPO|5164,5167
with|5168,5172
<EOL>|5173,5174
IVF|5174,5177
resuscitation|5178,5191
.|5191,5192
A|5194,5195
abdominal|5196,5205
/|5205,5206
pelvic|5206,5212
CT|5213,5215
was|5216,5219
done|5220,5224
and|5225,5228
<EOL>|5229,5230
demonstrated|5230,5242
a|5243,5244
stable|5245,5251
sigmoid|5252,5259
anastomosis|5260,5271
without|5272,5279
any|5280,5283
fluid|5284,5289
<EOL>|5290,5291
collections|5291,5302
or|5303,5305
free|5306,5310
air|5311,5314
.|5314,5315
Over|5317,5321
the|5322,5325
first|5326,5331
night|5332,5337
her|5338,5341
urine|5342,5347
output|5348,5354
<EOL>|5355,5356
increased|5356,5365
and|5366,5369
a|5370,5371
foley|5372,5377
was|5378,5381
not|5382,5385
placed|5386,5392
.|5392,5393
Due|5395,5398
to|5399,5401
her|5402,5405
constant|5406,5414
loose|5415,5420
<EOL>|5421,5422
stools|5422,5428
,|5428,5429
toxin|5430,5435
screens|5436,5443
of|5444,5446
C|5447,5448
.|5448,5449
diff|5449,5453
were|5454,5458
sent|5459,5463
and|5464,5467
returned|5468,5476
negative|5477,5485
.|5485,5486
<EOL>|5487,5488
By|5489,5491
HD2|5492,5495
,|5495,5496
the|5497,5500
nausea|5501,5507
persisted|5508,5517
an|5518,5520
a|5521,5522
GI|5523,5525
consult|5526,5533
was|5534,5537
obtained|5538,5546
.|5546,5547
The|5549,5552
<EOL>|5553,5554
GI|5554,5556
service|5557,5564
believed|5565,5573
the|5574,5577
nausea|5578,5584
to|5585,5587
be|5588,5590
related|5591,5598
to|5599,5601
baseline|5602,5610
reflux|5611,5617
<EOL>|5618,5619
exacerbated|5619,5630
by|5631,5633
her|5634,5637
postop|5638,5644
course|5645,5651
,|5651,5652
including|5653,5662
a|5663,5664
wound|5665,5670
infection|5671,5680
.|5680,5681
<EOL>|5683,5684
Per|5684,5687
their|5688,5693
recommendations|5694,5709
,|5709,5710
she|5711,5714
was|5715,5718
started|5719,5726
on|5727,5729
an|5730,5732
antacid|5733,5740
and|5741,5744
<EOL>|5745,5746
upon|5746,5750
discharge|5751,5760
she|5761,5764
will|5765,5769
follow|5770,5776
up|5777,5779
with|5780,5784
a|5785,5786
gastroenterologist|5787,5805
to|5806,5808
<EOL>|5809,5810
determine|5810,5819
her|5820,5823
H|5824,5825
.|5825,5826
pylori|5826,5832
status|5833,5839
.|5839,5840
Prior|5843,5848
to|5849,5851
discharge|5852,5861
,|5861,5862
she|5863,5866
was|5867,5870
<EOL>|5871,5872
tolerating|5872,5882
a|5883,5884
low|5885,5888
residue|5889,5896
diet|5897,5901
and|5902,5905
able|5906,5910
to|5911,5913
hydrate|5914,5921
herself|5922,5929
.|5929,5930
<EOL>|5932,5933
<EOL>|5934,5935
Discharge|5935,5944
Medications|5945,5956
:|5956,5957
<EOL>|5957,5958
1.|5958,5960
Escitalopram|5961,5973
10|5974,5976
mg|5977,5979
Tablet|5980,5986
Sig|5987,5990
:|5990,5991
One|5992,5995
(|5996,5997
1|5997,5998
)|5998,5999
Tablet|6000,6006
PO|6007,6009
DAILY|6010,6015
<EOL>|6016,6017
(|6017,6018
Daily|6018,6023
)|6023,6024
.|6024,6025
<EOL>|6025,6026
Disp|6026,6030
:|6030,6031
*|6031,6032
0|6032,6033
Tablet|6034,6040
(|6040,6041
s|6041,6042
)|6042,6043
*|6043,6044
Refills|6045,6052
:|6052,6053
*|6053,6054
0|6054,6055
*|6055,6056
<EOL>|6056,6057
2.|6057,6059
Pantoprazole|6060,6072
40|6073,6075
mg|6076,6078
Tablet|6079,6085
,|6085,6086
Delayed|6087,6094
Release|6095,6102
(|6103,6104
E.C|6104,6107
.|6107,6108
)|6108,6109
Sig|6110,6113
:|6113,6114
One|6115,6118
<EOL>|6119,6120
(|6120,6121
1|6121,6122
)|6122,6123
Tablet|6124,6130
,|6130,6131
Delayed|6132,6139
Release|6140,6147
(|6148,6149
E.C|6149,6152
.|6152,6153
)|6153,6154
PO|6155,6157
Q12H|6158,6162
(|6163,6164
every|6164,6169
12|6170,6172
hours|6173,6178
)|6178,6179
.|6179,6180
<EOL>|6180,6181
Disp|6181,6185
:|6185,6186
*|6186,6187
60|6187,6189
Tablet|6190,6196
,|6196,6197
Delayed|6198,6205
Release|6206,6213
(|6214,6215
E.C|6215,6218
.|6218,6219
)|6219,6220
(|6220,6221
s|6221,6222
)|6222,6223
*|6223,6224
Refills|6225,6232
:|6232,6233
*|6233,6234
2|6234,6235
*|6235,6236
<EOL>|6236,6237
3.|6237,6239
Ranitidine|6240,6250
HCl|6251,6254
150|6255,6258
mg|6259,6261
Tablet|6262,6268
Sig|6269,6272
:|6272,6273
One|6274,6277
(|6278,6279
1|6279,6280
)|6280,6281
Tablet|6282,6288
PO|6289,6291
HS|6292,6294
(|6295,6296
at|6296,6298
<EOL>|6299,6300
bedtime|6300,6307
)|6307,6308
.|6308,6309
<EOL>|6309,6310
Disp|6310,6314
:|6314,6315
*|6315,6316
30|6316,6318
Tablet|6319,6325
(|6325,6326
s|6326,6327
)|6327,6328
*|6328,6329
Refills|6330,6337
:|6337,6338
*|6338,6339
2|6339,6340
*|6340,6341
<EOL>|6341,6342
4.|6342,6344
Fluticasone|6345,6356
50|6357,6359
mcg|6360,6363
/|6363,6364
Actuation|6364,6373
Spray|6374,6379
,|6379,6380
Suspension|6381,6391
Sig|6392,6395
:|6395,6396
One|6397,6400
(|6401,6402
1|6402,6403
)|6403,6404
<EOL>|6405,6406
Spray|6406,6411
Nasal|6412,6417
DAILY|6418,6423
(|6424,6425
Daily|6425,6430
)|6430,6431
.|6431,6432
<EOL>|6432,6433
Disp|6433,6437
:|6437,6438
*|6438,6439
0|6439,6440
*|6441,6442
Refills|6443,6450
:|6450,6451
*|6451,6452
0|6452,6453
*|6453,6454
<EOL>|6454,6455
<EOL>|6455,6456
<EOL>|6457,6458
Discharge|6458,6467
Disposition|6468,6479
:|6479,6480
<EOL>|6480,6481
Home|6481,6485
With|6486,6490
Service|6491,6498
<EOL>|6498,6499
<EOL>|6500,6501
Facility|6501,6509
:|6509,6510
<EOL>|6510,6511
_|6511,6512
_|6512,6513
_|6513,6514
<EOL>|6514,6515
<EOL>|6516,6517
Discharge|6517,6526
Diagnosis|6527,6536
:|6536,6537
<EOL>|6537,6538
nausea|6538,6544
and|6545,6548
vomiting|6549,6557
<EOL>|6557,6558
<EOL>|6558,6559
<EOL>|6560,6561
Followup|6582,6590
Instructions|6591,6603
:|6603,6604
<EOL>|6604,6605
_|6605,6606
_|6606,6607
_|6607,6608
<EOL>|6608,6609

