 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|29,33
No|34,36
:|36,37
_|40,41
_|41,42
_|42,43
<EOL>|43,44
<EOL>|45,46
Admission|46,55
Date|56,60
:|60,61
_|63,64
_|64,65
_|65,66
Discharge|80,89
Date|90,94
:|94,95
_|98,99
_|99,100
_|100,101
<EOL>|101,102
<EOL>|103,104
Date|104,108
of|109,111
Birth|112,117
:|117,118
_|120,121
_|121,122
_|122,123
Sex|136,139
:|139,140
F|143,144
<EOL>|144,145
<EOL>|146,147
Service|147,154
:|154,155
MEDICINE|156,164
<EOL>|164,165
<EOL>|166,167
Patient|179,186
recorded|187,195
as|196,198
having|199,205
No|206,208
Known|209,214
Allergies|215,224
to|225,227
Drugs|228,233
<EOL>|233,234
<EOL>|235,236
Attending|236,245
:|245,246
_|247,248
_|248,249
_|249,250
<EOL>|250,251
<EOL>|252,253
CP|270,272
<EOL>|272,273
<EOL>|274,275
Major|275,280
Surgical|281,289
or|290,292
Invasive|293,301
Procedure|302,311
:|311,312
<EOL>|312,313
None|313,317
<EOL>|317,318
<EOL>|318,319
<EOL>|320,321
_|349,350
_|350,351
_|351,352
yo|353,355
F|356,357
with|358,362
hx|363,365
CAD|366,369
(|370,371
BMS|371,374
x|375,376
1|377,378
_|379,380
_|380,381
_|381,382
,|382,383
_|384,385
_|385,386
_|386,387
2|388,389
in|390,392
_|393,394
_|394,395
_|395,396
and|397,400
_|401,402
_|402,403
_|403,404
to|405,407
LAD|408,411
)|411,412
,|412,413
<EOL>|414,415
poorly|415,421
controlled|422,432
type|433,437
2|438,439
IDDM|440,444
,|444,445
HTN|446,449
presented|450,459
to|460,462
PCP|463,466
's|466,468
office|469,475
<EOL>|476,477
this|477,481
AM|482,484
reporting|485,494
episode|495,502
of|503,505
CP|506,508
last|509,513
night|514,519
.|519,520
Over|521,525
the|526,529
past|530,534
week|535,539
<EOL>|540,541
patient|541,548
's|548,550
jan|551,554
_|554,555
_|555,556
_|556,557
duties|558,564
have|565,569
increased|570,579
and|580,583
has|584,587
felt|588,592
weak|593,597
and|598,601
<EOL>|602,603
fatigued|603,611
.|611,612
Admits|613,619
to|620,622
radiation|623,632
to|633,635
R|636,637
arm|638,641
.|641,642
At|643,645
approx|646,652
10pm|653,657
last|658,662
<EOL>|663,664
night|664,669
,|669,670
patient|671,678
felt|679,683
faint|684,689
and|690,693
c|694,695
/|695,696
o|696,697
_|698,699
_|699,700
_|700,701
chest|702,707
tightness|708,717
,|717,718
<EOL>|719,720
relieved|720,728
by|729,731
took|732,736
2|737,738
NTG|739,742
.|742,743
Denies|744,750
any|751,754
associated|755,765
SOB|766,769
,|769,770
Diaphoresis|771,782
.|782,783
<EOL>|784,785
Patient|785,792
c|793,794
/|794,795
o|795,796
perisistent|797,808
_|809,810
_|810,811
_|811,812
CP|813,815
Today|816,821
and|822,825
feels|826,831
mildly|832,838
SOB|839,842
.|842,843
<EOL>|845,846
In|846,848
the|849,852
ER|853,855
,|855,856
patient|857,864
's|864,866
VS|867,869
were|870,874
97.2|875,879
,|879,880
99|881,883
,|883,884
145|885,888
/|888,889
97|889,891
,|891,892
15|893,895
,|895,896
100|897,900
%|900,901
2L|902,904
NC|905,907
.|907,908
<EOL>|909,910
Patient|910,917
had|918,921
CP|922,924
relief|925,931
to|932,934
2|935,936
SL|937,939
NTG|940,943
.|943,944
On|945,947
transfer|948,956
to|957,959
floor|960,965
,|965,966
patient|967,974
<EOL>|975,976
has|976,979
no|980,982
chest|983,988
pain|989,993
.|993,994
<EOL>|996,997
.|997,998
<EOL>|1000,1001
Patient|1001,1008
denies|1009,1015
any|1016,1019
N|1020,1021
,|1021,1022
V|1023,1024
,|1024,1025
D|1026,1027
,|1027,1028
CP|1029,1031
,|1031,1032
SOB|1033,1036
currently|1037,1046
.|1046,1047
All|1048,1051
other|1052,1057
ROS|1058,1061
<EOL>|1062,1063
negative|1063,1071
unless|1072,1078
otherwise|1079,1088
specified|1089,1098
<EOL>|1099,1100
<EOL>|1100,1101
<EOL>|1102,1103
asthma|1125,1131
,|1131,1132
emphysema|1133,1142
,|1142,1143
chronic|1144,1151
bronchitis|1152,1162
,|1162,1163
HTN|1164,1167
,|1167,1168
CAD|1169,1172
(|1173,1174
MIx2|1174,1178
,|1178,1179
2|1180,1181
<EOL>|1181,1182
cardiac|1182,1189
stents|1190,1196
_|1197,1198
_|1198,1199
_|1199,1200
,|1200,1201
migraines|1202,1211
,|1211,1212
GERD|1213,1217
,|1217,1218
DM|1219,1221
(|1222,1223
takes|1223,1228
pills|1229,1234
and|1235,1238
<EOL>|1238,1239
insulin|1239,1246
)|1246,1247
,|1247,1248
Anemia|1249,1255
,|1255,1256
neuropathy|1257,1267
,|1267,1268
anxiety|1269,1276
<EOL>|1276,1277
<EOL>|1277,1278
<EOL>|1279,1280
:|1294,1295
<EOL>|1295,1296
_|1296,1297
_|1297,1298
_|1298,1299
<EOL>|1299,1300
:|1314,1315
<EOL>|1315,1316
parents|1316,1323
not|1324,1327
known|1328,1333
.|1333,1334
daughter|1335,1343
htn|1344,1347
<EOL>|1349,1350
<EOL>|1350,1351
<EOL>|1352,1353
Physical|1353,1361
_|1362,1363
_|1363,1364
_|1364,1365
:|1365,1366
<EOL>|1366,1367
VS|1367,1369
-|1370,1371
98.3|1372,1376
,|1376,1377
142|1378,1381
/|1381,1382
77|1382,1384
,|1384,1385
89|1386,1388
,|1388,1389
16|1390,1392
,|1392,1393
93|1394,1396
%|1396,1397
RA|1397,1399
<EOL>|1401,1402
Gen|1402,1405
:|1405,1406
WDWN|1407,1411
middle|1412,1418
aged|1419,1423
male|1424,1428
in|1429,1431
NAD|1432,1435
.|1435,1436
Oriented|1437,1445
x3|1446,1448
.|1448,1449
Mood|1450,1454
,|1454,1455
affect|1456,1462
<EOL>|1463,1464
appropriate|1464,1475
.|1475,1476
<EOL>|1478,1479
HEENT|1479,1484
:|1484,1485
NCAT|1486,1490
.|1490,1491
Sclera|1492,1498
anicteric|1499,1508
.|1508,1509
PERRL|1510,1515
,|1515,1516
EOMI|1517,1521
.|1521,1522
Conjunctiva|1523,1534
were|1535,1539
<EOL>|1540,1541
pink|1541,1545
,|1545,1546
no|1547,1549
pallor|1550,1556
or|1557,1559
cyanosis|1560,1568
of|1569,1571
the|1572,1575
oral|1576,1580
mucosa|1581,1587
.|1587,1588
No|1589,1591
xanthalesma|1592,1603
.|1603,1604
<EOL>|1606,1607
<EOL>|1607,1608
Neck|1608,1612
:|1612,1613
No|1614,1616
JVD|1617,1620
<EOL>|1622,1623
CV|1623,1625
:|1625,1626
RR|1627,1629
,|1629,1630
normal|1631,1637
S1|1638,1640
,|1640,1641
S2|1642,1644
.|1644,1645
No|1646,1648
m|1649,1650
/|1650,1651
r|1651,1652
/|1652,1653
g|1653,1654
.|1654,1655
No|1656,1658
thrills|1659,1666
,|1666,1667
lifts|1668,1673
.|1673,1674
No|1675,1677
S3|1678,1680
or|1681,1683
S4|1684,1686
.|1686,1687
<EOL>|1688,1689
<EOL>|1690,1691
Chest|1691,1696
:|1696,1697
CTAB|1698,1702
,|1702,1703
no|1704,1706
crackles|1707,1715
,|1715,1716
wheezes|1717,1724
or|1725,1727
rhonchi|1728,1735
.|1735,1736
<EOL>|1738,1739
Abd|1739,1742
:|1742,1743
Soft|1744,1748
,|1748,1749
NTND|1750,1754
.|1754,1755
No|1756,1758
HSM|1759,1762
or|1763,1765
tenderness|1766,1776
.|1776,1777
Abd|1778,1781
aorta|1782,1787
not|1788,1791
enlarged|1792,1800
by|1801,1803
<EOL>|1804,1805
palpation|1805,1814
.|1814,1815
No|1816,1818
abdominial|1819,1829
bruits|1830,1836
.|1836,1837
<EOL>|1839,1840
Ext|1840,1843
:|1843,1844
No|1845,1847
c|1848,1849
/|1849,1850
c|1850,1851
/|1851,1852
e|1852,1853
.|1853,1854
No|1855,1857
femoral|1858,1865
bruits|1866,1872
.|1872,1873
<EOL>|1875,1876
Skin|1876,1880
:|1880,1881
No|1882,1884
stasis|1885,1891
dermatitis|1892,1902
,|1902,1903
ulcers|1904,1910
,|1910,1911
scars|1912,1917
,|1917,1918
or|1919,1921
xanthomas|1922,1931
.|1931,1932
<EOL>|1934,1935
.|1935,1936
<EOL>|1938,1939
Pulses|1939,1945
:|1945,1946
<EOL>|1948,1949
Right|1949,1954
:|1954,1955
Carotid|1956,1963
2|1964,1965
+|1965,1966
DP|1967,1969
2|1970,1971
+|1971,1972
_|1973,1974
_|1974,1975
_|1975,1976
2|1977,1978
+|1978,1979
<EOL>|1981,1982
Left|1982,1986
:|1986,1987
Carotid|1988,1995
2|1996,1997
+|1997,1998
DP|1999,2001
2|2002,2003
+|2003,2004
_|2005,2006
_|2006,2007
_|2007,2008
2|2009,2010
+|2010,2011
<EOL>|2013,2014
<EOL>|2014,2015
<EOL>|2016,2017
Pertinent|2017,2026
Results|2027,2034
:|2034,2035
<EOL>|2035,2036
_|2036,2037
_|2037,2038
_|2038,2039
Stress|2040,2046
<EOL>|2046,2047
INTERPRETATION|2047,2061
:|2061,2062
This|2063,2067
_|2068,2069
_|2069,2070
_|2070,2071
yo|2072,2074
Type|2075,2079
II|2080,2082
IDDM|2083,2087
woman|2088,2093
with|2094,2098
a|2099,2100
h|2101,2102
/|2102,2103
o|2103,2104
MI|2105,2107
and|2108,2111
<EOL>|2112,2113
stent|2113,2118
in|2119,2121
_|2122,2123
_|2123,2124
_|2124,2125
was|2126,2129
referred|2130,2138
for|2139,2142
evaluation|2143,2153
of|2154,2156
chest|2157,2162
pain|2163,2167
.|2167,2168
The|2169,2172
<EOL>|2173,2174
patient|2174,2181
was|2182,2185
<EOL>|2186,2187
infused|2187,2194
with|2195,2199
0.142|2200,2205
mg|2205,2207
/|2207,2208
kg|2208,2210
/|2210,2211
min|2211,2214
of|2215,2217
persantine|2218,2228
over|2229,2233
4|2234,2235
minutes|2236,2243
.|2243,2244
During|2245,2251
<EOL>|2252,2253
<EOL>|2253,2254
infusion|2254,2262
,|2262,2263
the|2264,2267
patient|2268,2275
reported|2276,2284
_|2285,2286
_|2286,2287
_|2287,2288
mid-sternal|2289,2300
chest|2301,2306
"|2307,2308
pressure|2308,2316
"|2316,2317
<EOL>|2318,2319
which|2319,2324
<EOL>|2325,2326
was|2326,2329
increased|2330,2339
slightly|2340,2348
with|2349,2353
inspiration|2354,2365
.|2365,2366
This|2367,2371
symptom|2372,2379
was|2380,2383
<EOL>|2384,2385
relieved|2385,2393
after|2394,2399
<EOL>|2400,2401
125mg|2401,2406
of|2407,2409
IV|2410,2412
aminophylline|2413,2426
was|2427,2430
given|2431,2436
post-isotope|2437,2449
injection|2450,2459
.|2459,2460
No|2461,2463
<EOL>|2464,2465
significant|2465,2476
ST|2477,2479
segment|2480,2487
changes|2488,2495
were|2496,2500
noted|2501,2506
.|2506,2507
The|2508,2511
rhythm|2512,2518
was|2519,2522
sinus|2523,2528
<EOL>|2529,2530
without|2530,2537
<EOL>|2538,2539
ectopy|2539,2545
.|2545,2546
Hemodynamic|2547,2558
response|2559,2567
to|2568,2570
infusion|2571,2579
was|2580,2583
appropriate|2584,2595
.|2595,2596
<EOL>|2597,2598
<EOL>|2600,2601
IMPRESSION|2601,2611
:|2611,2612
Possible|2613,2621
anginal|2622,2629
type|2630,2634
symptoms|2635,2643
in|2644,2646
the|2647,2650
absence|2651,2658
of|2659,2661
<EOL>|2662,2663
ischemic|2663,2671
<EOL>|2672,2673
EKG|2673,2676
changes|2677,2684
.|2684,2685
Nuclear|2686,2693
report|2694,2700
sent|2701,2705
separately|2706,2716
.|2716,2717
<EOL>|2718,2719
<EOL>|2719,2720
<EOL>|2721,2722
IMPRESSION|2722,2732
:|2732,2733
Normal|2734,2740
myocardial|2741,2751
perfusion|2752,2761
and|2762,2765
function|2766,2774
(|2775,2776
EF|2776,2778
57|2779,2781
%|2781,2782
)|2782,2783
<EOL>|2784,2785
<EOL>|2785,2786
_|2786,2787
_|2787,2788
_|2788,2789
06|2790,2792
:|2792,2793
25AM|2793,2797
BLOOD|2798,2803
WBC|2804,2807
-|2807,2808
7.5|2808,2811
RBC|2812,2815
-|2815,2816
3|2816,2817
.|2817,2818
94|2818,2820
*|2820,2821
Hgb|2822,2825
-|2825,2826
13.0|2826,2830
Hct|2831,2834
-|2834,2835
36.1|2835,2839
<EOL>|2840,2841
MCV|2841,2844
-|2844,2845
92|2845,2847
MCH|2848,2851
-|2851,2852
32|2852,2854
.|2854,2855
9|2855,2856
*|2856,2857
MCHC|2858,2862
-|2862,2863
36|2863,2865
.|2865,2866
0|2866,2867
*|2867,2868
RDW|2869,2872
-|2872,2873
13.1|2873,2877
Plt|2878,2881
_|2882,2883
_|2883,2884
_|2884,2885
<EOL>|2885,2886
_|2886,2887
_|2887,2888
_|2888,2889
07|2890,2892
:|2892,2893
00AM|2893,2897
BLOOD|2898,2903
WBC|2904,2907
-|2907,2908
7.1|2908,2911
RBC|2912,2915
-|2915,2916
3|2916,2917
.|2917,2918
84|2918,2920
*|2920,2921
Hgb|2922,2925
-|2925,2926
12.9|2926,2930
Hct|2931,2934
-|2934,2935
35|2935,2937
.|2937,2938
3|2938,2939
*|2939,2940
<EOL>|2941,2942
MCV|2942,2945
-|2945,2946
92|2946,2948
MCH|2949,2952
-|2952,2953
33|2953,2955
.|2955,2956
7|2956,2957
*|2957,2958
MCHC|2959,2963
-|2963,2964
36|2964,2966
.|2966,2967
6|2967,2968
*|2968,2969
RDW|2970,2973
-|2973,2974
12.1|2974,2978
Plt|2979,2982
_|2983,2984
_|2984,2985
_|2985,2986
<EOL>|2986,2987
_|2987,2988
_|2988,2989
_|2989,2990
05|2991,2993
:|2993,2994
30AM|2994,2998
BLOOD|2999,3004
WBC|3005,3008
-|3008,3009
8.1|3009,3012
RBC|3013,3016
-|3016,3017
3|3017,3018
.|3018,3019
76|3019,3021
*|3021,3022
Hgb|3023,3026
-|3026,3027
12.6|3027,3031
Hct|3032,3035
-|3035,3036
34|3036,3038
.|3038,3039
9|3039,3040
*|3040,3041
<EOL>|3042,3043
MCV|3043,3046
-|3046,3047
93|3047,3049
MCH|3050,3053
-|3053,3054
33|3054,3056
.|3056,3057
6|3057,3058
*|3058,3059
MCHC|3060,3064
-|3064,3065
36|3065,3067
.|3067,3068
2|3068,3069
*|3069,3070
RDW|3071,3074
-|3074,3075
13.2|3075,3079
Plt|3080,3083
_|3084,3085
_|3085,3086
_|3086,3087
<EOL>|3087,3088
_|3088,3089
_|3089,3090
_|3090,3091
06|3092,3094
:|3094,3095
25AM|3095,3099
BLOOD|3100,3105
Plt|3106,3109
_|3110,3111
_|3111,3112
_|3112,3113
<EOL>|3113,3114
_|3114,3115
_|3115,3116
_|3116,3117
07|3118,3120
:|3120,3121
00AM|3121,3125
BLOOD|3126,3131
Plt|3132,3135
_|3136,3137
_|3137,3138
_|3138,3139
<EOL>|3139,3140
_|3140,3141
_|3141,3142
_|3142,3143
05|3144,3146
:|3146,3147
30AM|3147,3151
BLOOD|3152,3157
Plt|3158,3161
_|3162,3163
_|3163,3164
_|3164,3165
<EOL>|3165,3166
_|3166,3167
_|3167,3168
_|3168,3169
06|3170,3172
:|3172,3173
25AM|3173,3177
BLOOD|3178,3183
Glucose|3184,3191
-|3191,3192
68|3192,3194
*|3194,3195
UreaN|3196,3201
-|3201,3202
17|3202,3204
Creat|3205,3210
-|3210,3211
0.8|3211,3214
Na|3215,3217
-|3217,3218
141|3218,3221
<EOL>|3222,3223
K|3223,3224
-|3224,3225
4.0|3225,3228
Cl|3229,3231
-|3231,3232
102|3232,3235
HCO3|3236,3240
-|3240,3241
32|3241,3243
AnGap|3244,3249
-|3249,3250
11|3250,3252
<EOL>|3252,3253
_|3253,3254
_|3254,3255
_|3255,3256
07|3257,3259
:|3259,3260
00AM|3260,3264
BLOOD|3265,3270
Glucose|3271,3278
-|3278,3279
90|3279,3281
UreaN|3282,3287
-|3287,3288
18|3288,3290
Creat|3291,3296
-|3296,3297
0.7|3297,3300
Na|3301,3303
-|3303,3304
139|3304,3307
<EOL>|3308,3309
K|3309,3310
-|3310,3311
4.1|3311,3314
Cl|3315,3317
-|3317,3318
101|3318,3321
HCO3|3322,3326
-|3326,3327
31|3327,3329
AnGap|3330,3335
-|3335,3336
11|3336,3338
<EOL>|3338,3339
_|3339,3340
_|3340,3341
_|3341,3342
05|3343,3345
:|3345,3346
30AM|3346,3350
BLOOD|3351,3356
Glucose|3357,3364
-|3364,3365
178|3365,3368
*|3368,3369
UreaN|3370,3375
-|3375,3376
22|3376,3378
*|3378,3379
Creat|3380,3385
-|3385,3386
0.8|3386,3389
Na|3390,3392
-|3392,3393
136|3393,3396
<EOL>|3397,3398
K|3398,3399
-|3399,3400
3.9|3400,3403
Cl|3404,3406
-|3406,3407
101|3407,3410
HCO3|3411,3415
-|3415,3416
24|3416,3418
AnGap|3419,3424
-|3424,3425
15|3425,3427
<EOL>|3427,3428
<EOL>|3429,3430
Patient|3453,3460
is|3461,3463
a|3464,3465
_|3466,3467
_|3467,3468
_|3468,3469
y|3470,3471
/|3471,3472
o|3472,3473
F|3474,3475
with|3476,3480
a|3481,3482
history|3483,3490
of|3491,3493
CAD|3494,3497
with|3498,3502
BMS|3503,3506
x|3507,3508
1|3509,3510
_|3511,3512
_|3512,3513
_|3513,3514
,|3514,3515
<EOL>|3516,3517
_|3517,3518
_|3518,3519
_|3519,3520
2|3521,3522
in|3523,3525
_|3526,3527
_|3527,3528
_|3528,3529
and|3530,3533
_|3534,3535
_|3535,3536
_|3536,3537
to|3538,3540
LAD|3541,3544
,|3544,3545
DM|3546,3548
,|3548,3549
HTN|3550,3553
,|3553,3554
Hypercholesterolemia|3555,3575
who|3576,3579
<EOL>|3580,3581
presents|3581,3589
with|3590,3594
atypical|3595,3603
chest|3604,3609
pain|3610,3614
.|3614,3615
<EOL>|3617,3618
.|3618,3619
<EOL>|3621,3622
#|3622,3623
.|3623,3624
CAD|3625,3628
:|3628,3629
Pt|3630,3632
with|3633,3637
hx|3638,3640
CAD|3641,3644
,|3644,3645
poorly|3646,3652
controlled|3653,3663
DM|3664,3666
,|3666,3667
episode|3668,3675
of|3676,3678
CP|3679,3681
<EOL>|3682,3683
prior|3683,3688
to|3689,3691
admission|3692,3701
concerning|3702,3712
for|3713,3716
angina|3717,3723
.|3723,3724
Patient|3726,3733
's|3733,3735
EKG|3736,3739
showed|3740,3746
<EOL>|3747,3748
TWI|3748,3751
in|3752,3754
AVL|3755,3758
that|3759,3763
is|3764,3766
nonspecific|3767,3778
.|3778,3779
Patient|3780,3787
ruled|3788,3793
out|3794,3797
for|3798,3801
MI|3802,3804
.|3804,3805
<EOL>|3807,3808
Patient|3808,3815
's|3815,3817
CP|3818,3820
that|3821,3825
was|3826,3829
likely|3830,3836
of|3837,3839
noncardiac|3840,3850
origin|3851,3857
,|3857,3858
given|3859,3864
the|3865,3868
<EOL>|3869,3870
multiple|3870,3878
episodes|3879,3887
of|3888,3890
waxing|3891,3897
and|3898,3901
waning|3902,3908
CP|3909,3911
with|3912,3916
rest|3917,3921
and|3922,3925
or|3926,3928
<EOL>|3929,3930
exertion|3930,3938
,|3938,3939
and|3940,3943
lack|3944,3948
of|3949,3951
EKG|3952,3955
changes|3956,3963
and|3964,3967
negative|3968,3976
cardiac|3977,3984
enzymes|3985,3992
.|3992,3993
<EOL>|3995,3996
Patient|3996,4003
had|4004,4007
a|4008,4009
nuclear|4010,4017
stress|4018,4024
as|4025,4027
an|4028,4030
inpatient|4031,4040
and|4041,4044
was|4045,4048
negative|4049,4057
<EOL>|4058,4059
for|4059,4062
any|4063,4066
perfusion|4067,4076
defects|4077,4084
.|4084,4085
<EOL>|4087,4088
-|4088,4089
Continue|4090,4098
ASA|4099,4102
,|4102,4103
Plavix|4104,4110
<EOL>|4112,4113
-|4113,4114
Contine|4115,4122
ACE|4123,4126
,|4126,4127
BB|4128,4130
<EOL>|4132,4133
-|4133,4134
Continue|4135,4143
Statin|4144,4150
<EOL>|4152,4153
.|4153,4154
<EOL>|4156,4157
#|4157,4158
.|4158,4159
Pump|4160,4164
:|4164,4165
Euvolemic|4166,4175
on|4176,4178
exam|4179,4183
.|4183,4184
<EOL>|4186,4187
.|4187,4188
<EOL>|4190,4191
#|4191,4192
.|4192,4193
Rhythm|4194,4200
:|4200,4201
NSR|4202,4205
.|4205,4206
<EOL>|4208,4209
.|4209,4210
<EOL>|4212,4213
#|4213,4214
HTN|4215,4218
:|4218,4219
SBP|4220,4223
120|4224,4227
-|4227,4228
140s|4228,4232
on|4233,4235
discharge|4236,4245
.|4245,4246
Concern|4248,4255
that|4256,4260
patient|4261,4268
may|4269,4272
be|4273,4275
<EOL>|4276,4277
non|4277,4280
compliant|4281,4290
with|4291,4295
medication|4296,4306
regimen|4307,4314
.|4314,4315
Patient|4317,4324
had|4325,4328
dropped|4329,4336
SBP|4337,4340
<EOL>|4341,4342
into|4342,4346
_|4347,4348
_|4348,4349
_|4349,4350
on|4351,4353
admission|4354,4363
once|4364,4368
home|4369,4373
medications|4374,4385
were|4386,4390
administered|4391,4403
.|4403,4404
<EOL>|4406,4407
Her|4407,4410
does|4411,4415
of|4416,4418
BB|4419,4421
and|4422,4425
Imdur|4426,4431
have|4432,4436
been|4437,4441
decreased|4442,4451
,|4451,4452
SBPs|4453,4457
have|4458,4462
been|4463,4467
<EOL>|4468,4469
controlled|4469,4479
,|4479,4480
but|4481,4484
may|4485,4488
need|4489,4493
outpatient|4494,4504
titration|4505,4514
.|4514,4515
<EOL>|4517,4518
-|4518,4519
Continue|4520,4528
BP|4529,4531
meds|4532,4536
.|4536,4537
<EOL>|4538,4539
.|4539,4540
<EOL>|4542,4543
#|4543,4544
.|4544,4545
DM|4546,4548
-|4549,4550
HbA1c|4551,4556
10.0|4557,4561
on|4562,4564
_|4565,4566
_|4566,4567
_|4567,4568
.|4568,4569
Poorly|4570,4576
controlled|4577,4587
.|4587,4588
Currently|4589,4598
on|4599,4601
<EOL>|4602,4603
Levemir|4603,4610
50|4611,4613
units|4614,4619
sq|4620,4622
in|4623,4625
AM|4626,4628
,|4628,4629
60|4630,4632
in|4633,4635
_|4636,4637
_|4637,4638
_|4638,4639
,|4639,4640
Metformin|4641,4650
500|4651,4654
mg|4655,4657
tid|4658,4661
,|4661,4662
<EOL>|4663,4664
although|4664,4672
not|4673,4676
compliant|4677,4686
with|4687,4691
this|4692,4696
.|4696,4697
<EOL>|4699,4700
-|4700,4701
Continue|4702,4710
metformin|4711,4720
<EOL>|4722,4723
-|4723,4724
Continue|4725,4733
Lantus|4734,4740
50u|4741,4744
qAM|4745,4748
/|4748,4749
60u|4749,4752
qHS|4753,4756
<EOL>|4758,4759
.|4759,4760
<EOL>|4762,4763
#|4763,4764
.|4764,4765
hyperlipidemia|4766,4780
-|4781,4782
Continue|4783,4791
Lipitor|4792,4799
80|4800,4802
mg|4803,4805
qday|4806,4810
.|4810,4811
<EOL>|4813,4814
<EOL>|4814,4815
<EOL>|4816,4817
Medications|4817,4828
on|4829,4831
Admission|4832,4841
:|4841,4842
<EOL>|4842,4843
Advair|4843,4849
250|4850,4853
/|4853,4854
50|4854,4856
daily|4857,4862
<EOL>|4864,4865
Albuterol|4865,4874
Aerosol|4875,4882
prn|4883,4886
<EOL>|4888,4889
ASA|4889,4892
325mg|4893,4898
daily|4899,4904
<EOL>|4906,4907
Atenolol|4907,4915
100mg|4916,4921
qday|4922,4926
<EOL>|4928,4929
Insulin|4929,4936
levimir|4937,4944
50|4945,4947
units|4948,4953
AM|4954,4956
;|4956,4957
60|4958,4960
units|4961,4966
_|4967,4968
_|4968,4969
_|4969,4970
,|4970,4971
<EOL>|4973,4974
Isosorbide|4974,4984
Mononitrate|4985,4996
120mg|4997,5002
daily|5003,5008
<EOL>|5010,5011
Lisinopril|5011,5021
10mg|5022,5026
daily|5027,5032
<EOL>|5034,5035
Metformin|5035,5044
500|5045,5048
mg|5049,5051
TID|5052,5055
,|5055,5056
<EOL>|5058,5059
Nitroglycerin|5059,5072
SL|5073,5075
<EOL>|5077,5078
Omeprazole|5078,5088
40|5089,5091
mg|5092,5094
daily|5095,5100
<EOL>|5102,5103
Plavix|5103,5109
75|5110,5112
mg|5113,5115
daily|5116,5121
,|5121,5122
<EOL>|5124,5125
Potassium|5125,5134
chloride|5135,5143
20|5144,5146
mEq|5147,5150
<EOL>|5152,5153
Simvastatin|5153,5164
80|5165,5167
mg|5168,5170
<EOL>|5172,5173
<EOL>|5173,5174
<EOL>|5175,5176
Discharge|5176,5185
Medications|5186,5197
:|5197,5198
<EOL>|5198,5199
1.|5199,5201
Fluticasone|5202,5213
-|5213,5214
Salmeterol|5214,5224
250|5225,5228
-|5228,5229
50|5229,5231
mcg|5232,5235
/|5235,5236
Dose|5236,5240
Disk|5241,5245
with|5246,5250
Device|5251,5257
Sig|5258,5261
:|5261,5262
<EOL>|5263,5264
One|5264,5267
(|5268,5269
1|5269,5270
)|5270,5271
Disk|5272,5276
with|5277,5281
Device|5282,5288
Inhalation|5289,5299
BID|5300,5303
(|5304,5305
2|5305,5306
times|5307,5312
a|5313,5314
day|5315,5318
)|5318,5319
.|5319,5320
<EOL>|5322,5323
2.|5323,5325
Aspirin|5326,5333
325|5334,5337
mg|5338,5340
Tablet|5341,5347
Sig|5348,5351
:|5351,5352
One|5353,5356
(|5357,5358
1|5358,5359
)|5359,5360
Tablet|5361,5367
PO|5368,5370
DAILY|5371,5376
(|5377,5378
Daily|5378,5383
)|5383,5384
.|5384,5385
<EOL>|5387,5388
3.|5388,5390
Albuterol|5391,5400
90|5401,5403
mcg|5404,5407
/|5407,5408
Actuation|5408,5417
Aerosol|5418,5425
Sig|5426,5429
:|5429,5430
_|5431,5432
_|5432,5433
_|5433,5434
Puffs|5435,5440
Inhalation|5441,5451
<EOL>|5452,5453
Q6H|5453,5456
(|5457,5458
every|5458,5463
6|5464,5465
hours|5466,5471
)|5471,5472
as|5473,5475
needed|5476,5482
.|5482,5483
<EOL>|5485,5486
4.|5486,5488
Clopidogrel|5489,5500
75|5501,5503
mg|5504,5506
Tablet|5507,5513
Sig|5514,5517
:|5517,5518
One|5519,5522
(|5523,5524
1|5524,5525
)|5525,5526
Tablet|5527,5533
PO|5534,5536
DAILY|5537,5542
<EOL>|5543,5544
(|5544,5545
Daily|5545,5550
)|5550,5551
.|5551,5552
<EOL>|5554,5555
5.|5555,5557
Simvastatin|5558,5569
40|5570,5572
mg|5573,5575
Tablet|5576,5582
Sig|5583,5586
:|5586,5587
Two|5588,5591
(|5592,5593
2|5593,5594
)|5594,5595
Tablet|5596,5602
PO|5603,5605
DAILY|5606,5611
<EOL>|5612,5613
(|5613,5614
Daily|5614,5619
)|5619,5620
.|5620,5621
<EOL>|5623,5624
6.|5624,5626
Omeprazole|5627,5637
20|5638,5640
mg|5641,5643
Capsule|5644,5651
,|5651,5652
Delayed|5653,5660
Release|5661,5668
(|5668,5669
E.C|5669,5672
.|5672,5673
)|5673,5674
Sig|5675,5678
:|5678,5679
Two|5680,5683
(|5684,5685
2|5685,5686
)|5686,5687
<EOL>|5688,5689
Capsule|5689,5696
,|5696,5697
Delayed|5698,5705
Release|5706,5713
(|5713,5714
E.C|5714,5717
.|5717,5718
)|5718,5719
PO|5720,5722
DAILY|5723,5728
(|5729,5730
Daily|5730,5735
)|5735,5736
.|5736,5737
<EOL>|5739,5740
7.|5740,5742
Oxycodone|5743,5752
-|5752,5753
Acetaminophen|5753,5766
_|5767,5768
_|5768,5769
_|5769,5770
mg|5771,5773
Tablet|5774,5780
Sig|5781,5784
:|5784,5785
_|5786,5787
_|5787,5788
_|5788,5789
Tablets|5790,5797
PO|5798,5800
<EOL>|5801,5802
Q6H|5802,5805
(|5806,5807
every|5807,5812
6|5813,5814
hours|5815,5820
)|5820,5821
as|5822,5824
needed|5825,5831
.|5831,5832
<EOL>|5834,5835
8.|5835,5837
Levemir|5838,5845
100|5846,5849
unit|5850,5854
/|5854,5855
mL|5855,5857
Solution|5858,5866
Sig|5867,5870
:|5870,5871
One|5872,5875
(|5876,5877
1|5877,5878
)|5878,5879
Subcutaneous|5881,5893
twice|5894,5899
<EOL>|5900,5901
a|5901,5902
day|5903,5906
:|5906,5907
50units|5908,5915
qAM|5916,5919
,|5919,5920
60|5921,5923
qPM|5924,5927
.|5927,5928
<EOL>|5930,5931
9.|5931,5933
Metformin|5934,5943
500|5944,5947
mg|5948,5950
Tablet|5951,5957
Sig|5958,5961
:|5961,5962
One|5963,5966
(|5967,5968
1|5968,5969
)|5969,5970
Tablet|5971,5977
PO|5978,5980
three|5981,5986
times|5987,5992
a|5993,5994
<EOL>|5995,5996
day|5996,5999
.|5999,6000
<EOL>|6002,6003
10.|6003,6006
Potassium|6007,6016
Chloride|6017,6025
10|6026,6028
mEq|6029,6032
Capsule|6033,6040
,|6040,6041
Sustained|6042,6051
Release|6052,6059
Sig|6060,6063
:|6063,6064
<EOL>|6065,6066
Two|6066,6069
(|6070,6071
2|6071,6072
)|6072,6073
Capsule|6074,6081
,|6081,6082
Sustained|6083,6092
Release|6093,6100
PO|6101,6103
once|6104,6108
a|6109,6110
day|6111,6114
.|6114,6115
<EOL>|6117,6118
11.|6118,6121
Nitroglycerin|6122,6135
0.4|6136,6139
mg|6140,6142
Tablet|6143,6149
,|6149,6150
Sublingual|6151,6161
Sig|6162,6165
:|6165,6166
One|6167,6170
(|6171,6172
1|6172,6173
)|6173,6174
tablet|6175,6181
<EOL>|6182,6183
Sublingual|6183,6193
q5min|6194,6199
as|6200,6202
needed|6203,6209
for|6210,6213
chest|6214,6219
pain|6220,6224
:|6224,6225
Sit|6226,6229
down|6230,6234
prior|6235,6240
to|6241,6243
<EOL>|6244,6245
taking|6245,6251
.|6251,6252
Take|6253,6257
one|6258,6261
tab|6262,6265
every|6266,6271
5|6272,6273
minutes|6274,6281
until|6282,6287
chest|6288,6293
pain|6294,6298
resolves|6299,6307
.|6307,6308
<EOL>|6309,6310
If|6310,6312
pain|6313,6317
not|6318,6321
resolved|6322,6330
,|6330,6331
please|6332,6338
call|6339,6343
EMS|6344,6347
.|6347,6348
<EOL>|6350,6351
12.|6351,6354
Lisinopril|6355,6365
5|6366,6367
mg|6368,6370
Tablet|6371,6377
Sig|6378,6381
:|6381,6382
One|6383,6386
(|6387,6388
1|6388,6389
)|6389,6390
Tablet|6391,6397
PO|6398,6400
DAILY|6401,6406
(|6407,6408
Daily|6408,6413
)|6413,6414
.|6414,6415
<EOL>|6415,6416
Disp|6416,6420
:|6420,6421
*|6421,6422
30|6422,6424
Tablet|6425,6431
(|6431,6432
s|6432,6433
)|6433,6434
*|6434,6435
Refills|6436,6443
:|6443,6444
*|6444,6445
2|6445,6446
*|6446,6447
<EOL>|6447,6448
13.|6448,6451
Metoprolol|6452,6462
Tartrate|6463,6471
25|6472,6474
mg|6475,6477
Tablet|6478,6484
Sig|6485,6488
:|6488,6489
1.5|6490,6493
Tablets|6494,6501
PO|6502,6504
BID|6505,6508
(|6509,6510
2|6510,6511
<EOL>|6512,6513
times|6513,6518
a|6519,6520
day|6521,6524
)|6524,6525
.|6525,6526
<EOL>|6526,6527
Disp|6527,6531
:|6531,6532
*|6532,6533
90|6533,6535
Tablet|6536,6542
(|6542,6543
s|6543,6544
)|6544,6545
*|6545,6546
Refills|6547,6554
:|6554,6555
*|6555,6556
2|6556,6557
*|6557,6558
<EOL>|6558,6559
14.|6559,6562
Isosorbide|6563,6573
Mononitrate|6574,6585
30|6586,6588
mg|6589,6591
Tablet|6592,6598
Sustained|6599,6608
Release|6609,6616
24|6617,6619
hr|6620,6622
<EOL>|6623,6624
Sig|6624,6627
:|6627,6628
One|6629,6632
(|6633,6634
1|6634,6635
)|6635,6636
Tablet|6637,6643
Sustained|6644,6653
Release|6654,6661
24|6662,6664
hr|6665,6667
PO|6668,6670
DAILY|6671,6676
(|6677,6678
Daily|6678,6683
)|6683,6684
.|6684,6685
<EOL>|6685,6686
Disp|6686,6690
:|6690,6691
*|6691,6692
30|6692,6694
Tablet|6695,6701
Sustained|6702,6711
Release|6712,6719
24|6720,6722
hr|6723,6725
(|6725,6726
s|6726,6727
)|6727,6728
*|6728,6729
Refills|6730,6737
:|6737,6738
*|6738,6739
2|6739,6740
*|6740,6741
<EOL>|6741,6742
<EOL>|6742,6743
<EOL>|6744,6745
Discharge|6745,6754
Disposition|6755,6766
:|6766,6767
<EOL>|6767,6768
Home|6768,6772
<EOL>|6772,6773
<EOL>|6774,6775
Discharge|6775,6784
Diagnosis|6785,6794
:|6794,6795
<EOL>|6795,6796
Primary|6796,6803
<EOL>|6803,6804
-|6804,6805
Atypical|6806,6814
Chest|6815,6820
pain|6821,6825
<EOL>|6825,6826
-|6826,6827
Coronary|6828,6836
artery|6837,6843
disase|6844,6850
<EOL>|6850,6851
Secondary|6851,6860
<EOL>|6860,6861
-|6861,6862
Hypertension|6863,6875
<EOL>|6875,6876
-|6876,6877
Diabetes|6878,6886
,|6886,6887
insulin|6888,6895
dependent|6896,6905
<EOL>|6905,6906
<EOL>|6906,6907
<EOL>|6908,6909
Afebrile|6930,6938
,|6938,6939
Chest|6940,6945
pain|6946,6950
free|6951,6955
,|6955,6956
stable|6957,6963
.|6963,6964
<EOL>|6966,6967
<EOL>|6967,6968
<EOL>|6969,6970
You|6994,6997
were|6998,7002
hospitalized|7003,7015
because|7016,7023
you|7024,7027
had|7028,7031
chest|7032,7037
pain|7038,7042
.|7042,7043
You|7045,7048
did|7049,7052
not|7053,7056
<EOL>|7057,7058
have|7058,7062
a|7063,7064
heart|7065,7070
attack|7071,7077
.|7077,7078
Your|7080,7084
chest|7085,7090
pain|7091,7095
resolved|7096,7104
.|7104,7105
Your|7107,7111
blood|7112,7117
<EOL>|7118,7119
pressure|7119,7127
was|7128,7131
a|7132,7133
little|7134,7140
low|7141,7144
on|7145,7147
the|7148,7151
regimen|7152,7159
you|7160,7163
had|7164,7167
previously|7168,7178
been|7179,7183
<EOL>|7184,7185
taking|7185,7191
at|7192,7194
home|7195,7199
.|7199,7200
Several|7202,7209
of|7210,7212
your|7213,7217
doses|7218,7223
have|7224,7228
been|7229,7233
changed|7234,7241
:|7241,7242
<EOL>|7242,7243
<EOL>|7243,7244
We|7244,7246
made|7247,7251
the|7252,7255
following|7256,7265
changes|7266,7273
to|7274,7276
your|7277,7281
medications|7282,7293
:|7293,7294
<EOL>|7294,7295
1|7295,7296
.|7296,7297
We|7298,7300
changed|7301,7308
your|7309,7313
imdur|7314,7319
to|7320,7322
30mg|7323,7327
daily|7328,7333
<EOL>|7333,7334
2|7334,7335
.|7335,7336
We|7337,7339
changed|7340,7347
your|7348,7352
lisinopril|7353,7363
to|7364,7366
5mg|7367,7370
daily|7371,7376
<EOL>|7376,7377
3|7377,7378
.|7378,7379
We|7380,7382
discontinued|7383,7395
your|7396,7400
atenolol|7401,7409
.|7409,7410
<EOL>|7410,7411
4|7411,7412
.|7412,7413
We|7414,7416
started|7417,7424
metoprolol|7425,7435
37.5|7436,7440
mg|7440,7442
,|7442,7443
twice|7444,7449
daily|7450,7455
.|7455,7456
<EOL>|7458,7459
<EOL>|7459,7460
You|7460,7463
had|7464,7467
a|7468,7469
stress|7470,7476
test|7477,7481
that|7482,7486
was|7487,7490
normal|7491,7497
.|7497,7498
Please|7500,7506
continue|7507,7515
to|7516,7518
<EOL>|7519,7520
adhere|7520,7526
to|7527,7529
a|7530,7531
healthy|7532,7539
diet|7540,7544
and|7545,7548
exercise|7549,7557
daily|7558,7563
.|7563,7564
<EOL>|7566,7567
<EOL>|7567,7568
If|7568,7570
you|7571,7574
experience|7575,7585
any|7586,7589
additional|7590,7600
chest|7601,7606
pain|7607,7611
,|7611,7612
shortness|7613,7622
of|7623,7625
<EOL>|7626,7627
breath|7627,7633
,|7633,7634
nausea|7635,7641
,|7641,7642
vomiting|7643,7651
,|7651,7652
please|7653,7659
call|7660,7664
your|7665,7669
PCP|7670,7673
or|7674,7676
return|7677,7683
to|7684,7686
the|7687,7690
<EOL>|7691,7692
ER|7692,7694
.|7694,7695
<EOL>|7697,7698
<EOL>|7699,7700
Followup|7700,7708
Instructions|7709,7721
:|7721,7722
<EOL>|7722,7723
_|7723,7724
_|7724,7725
_|7725,7726
<EOL>|7726,7727

