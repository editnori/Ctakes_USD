CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Pharmaceutical Preparations|Drug|false|false||MEDICINEnull|Medicine|Title|false|false||MEDICINEnull|Dyes|Drug|false|false||Dyenull|Iodine, Homeopathic preparation|Drug|false|false||Iodine
null|iodine|Drug|false|false||Iodine
null|iodine|Drug|false|false||Iodine
null|iodine|Drug|false|false||Iodinenull|Containing (qualifier value)|Finding|false|false||Containingnull|Contain (action)|Event|false|false||Containingnull|Contrast Media|Drug|false|false|C1254021;C0162867|Contrast Medianull|Contrast Media|Drug|false|false||Contrastnull|Contrast|Modifier|false|false||Contrastnull|Communications Media|Finding|false|false|C1254021;C0162867|Media
null|PAMS Media|Finding|false|false|C1254021;C0162867|Medianull|Tunica Media|Anatomy|false|false|C0677540;C0009458;C0009924;C0524222|Media
null|Media layer|Anatomy|false|false|C0677540;C0009458;C0009924;C0524222|Medianull|oxycodone|Drug|false|false||Oxycodone
null|oxycodone|Drug|false|false||Oxycodonenull|Oxycodone measurement|Procedure|false|false|C1254021;C0162867|Oxycodonenull|cilostazol|Drug|false|false||cilostazol
null|cilostazol|Drug|false|false||cilostazolnull|varenicline|Drug|false|false||Varenicline
null|varenicline|Drug|false|false||Vareniclinenull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Chest Pain|Finding|false|false|C1527391;C0817096|Chest painnull|null|Attribute|false|false|C1527391;C0817096|Chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|Chestnull|Chest|Anatomy|false|false|C0008031;C2926613;C0741025;C1549543;C0030193|Chest
null|Anterior thoracic region|Anatomy|false|false|C0008031;C2926613;C0741025;C1549543;C0030193|Chestnull|Administration Method - Pain|Finding|false|false|C1527391;C0817096|pain
null|Pain|Finding|false|false|C1527391;C0817096|painnull|null|Attribute|false|false||painnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Transaction counts and value totals - year|Finding|false|false||year
null|Precision - year|Finding|false|false||yearnull|year|Time|false|false||yearnull|Old|Time|false|false||oldnull|Females|Subject|false|false||female
null|Woman|Subject|false|false||femalenull|Female, Self-Report|Modifier|false|false||female
null|Female Phenotype|Modifier|false|false||femalenull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Peripheral Vascular Diseases|Disorder|false|false||PVDnull|Pomalidomide/Bortezomib/Dexamethasone Regimen|Procedure|false|false||PVDnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|Chest Pain|Finding|false|false|C1527391;C0817096|chest painnull|null|Attribute|false|false|C1527391;C0817096|chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0741025;C2926613;C0008031|chest
null|Anterior thoracic region|Anatomy|false|false|C0741025;C2926613;C0008031|chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Dyspnea|Finding|false|false||shortness of breathnull|null|Attribute|false|false||shortness of breathnull|Breath|Finding|false|false||breathnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Report (document)|Finding|false|false||reportsnull|Reporting|Procedure|false|false||reportsnull|5 minutes Office visit|Procedure|false|false||5 minutesnull|5 minutes|Time|false|false||5 minutesnull|Minute of time|Time|false|false||minutesnull|Minute Unit of Plane Angle|LabModifier|false|false||minutes
null|Minute (diminutive)|LabModifier|false|false||minutes
null|Small|LabModifier|false|false||minutesnull|Several|LabModifier|false|false||severalnull|More|LabModifier|false|false||morenull|Episode of|Time|false|false||episodesnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Minute of time|Time|false|false||minutesnull|Minute Unit of Plane Angle|LabModifier|false|false||minutes
null|Minute (diminutive)|LabModifier|false|false||minutes
null|Small|LabModifier|false|false||minutesnull|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Morning|Time|false|false||morningnull|Much|Finding|false|false||muchnull|Smaller|Modifier|false|false||lessnull|Less Than|LabModifier|false|false||lessnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Episode of|Time|false|false||episode ofnull|Episode of|Time|false|false||episodenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Palpitations|Finding|true|false||palpitationsnull|Lightheadedness|Finding|true|false||lightheadednessnull|Dizziness|Finding|true|false||dizziness
null|Vertigo|Finding|true|false||dizzinessnull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|Vomiting|Finding|false|false||vomitingnull|Increased sweating|Finding|false|false||diaphoresisnull|Initial (abbreviation)|Finding|false|false||initialnull|Initially|Time|false|false||initialnull|Firstly|Modifier|false|false||initialnull|Laboratory test finding|Lab|false|false||Labsnull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|carbon dioxide|Drug|false|false||CO2
null|carbon dioxide|Drug|false|false||CO2null|MT-CO2 gene|Finding|false|false||CO2
null|null|Finding|false|false||CO2
null|C2 wt Allele|Finding|false|false||CO2null|Blood Urea Nitrogen|Drug|false|false||BUN
null|Blood Urea Nitrogen|Drug|false|false||BUNnull|Blood urea nitrogen measurement|Procedure|false|false||BUNnull|Leukocytes|Anatomy|false|false|C1424337;C0201617;C0472699;C0018935;C0019046|WBCnull|Hemoglobin|Drug|false|false|C0023516|Hgb
null|Hemoglobin|Drug|false|false|C0023516|Hgbnull|CYGB gene|Finding|false|false|C0023516|Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false|C0023516|Hct
null|Hematocrit Measurement|Procedure|false|false|C0023516|Hctnull|Primed lymphocyte test|Procedure|false|false|C0023516|Pltnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Integrated Neuromusculoskeletal Release|Procedure|false|false||INR
null|International Normalized Ratio|Procedure|false|false||INRnull|Coagulation tissue factor induced.INR|Attribute|false|false||INRnull|lactate|Drug|false|false||Lactate
null|lactate|Drug|false|false||Lactate
null|Lactates|Drug|false|false||Lactatenull|Lactic acid measurement|Procedure|false|false||Lactatenull|Imaging problem|Finding|false|false||Imagingnull|Diagnostic Imaging|Procedure|false|false||Imaging
null|Imaging Techniques|Procedure|false|false||Imagingnull|Imaging Technology|Title|false|false||Imagingnull|Plain chest X-ray|Procedure|false|false||CXRnull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Cardiovascular disease+Pulmonary disease|Disorder|false|false|C1184743;C0553534|cardiopulmonarynull|Cardiopulmonary|Anatomy|false|false|C4072686;C1522240;C4521054|cardiopulmonarynull|Process Pharmacologic Substance|Drug|true|false|C1184743|processnull|Process (qualifier value)|Finding|true|false|C0553534;C1184743|processnull|bony process|Anatomy|false|false|C1951340;C4072686;C1522240;C4521054|processnull|Process|Phenomenon|true|false|C1184743;C0553534|processnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|aspirin|Drug|false|false||Aspirin
null|aspirin|Drug|false|false||Aspirinnull|albuterol|Drug|false|false||Albuterol
null|albuterol|Drug|false|false||Albuterolnull|NEB protein, human|Drug|false|false||Neb
null|NEB protein, human|Drug|false|false||Neb
null|Nebulizer solution|Drug|false|false||Nebnull|NEB gene|Finding|false|false||Neb
null|mitotic nuclear membrane disassembly|Finding|false|false||Nebnull|ipratropium bromide|Drug|false|false||Ipratropium Bromide
null|ipratropium bromide|Drug|false|false||Ipratropium Bromidenull|ipratropium|Drug|false|false||Ipratropium
null|ipratropium|Drug|false|false||Ipratropiumnull|Bromides|Drug|false|false||Bromidenull|Bromides measurement|Procedure|false|false||Bromidenull|NEB protein, human|Drug|false|false||Neb
null|NEB protein, human|Drug|false|false||Neb
null|Nebulizer solution|Drug|false|false||Nebnull|NEB gene|Finding|false|false||Neb
null|mitotic nuclear membrane disassembly|Finding|false|false||Nebnull|potassium chloride|Drug|false|false||Potassium Chloride
null|potassium chloride|Drug|false|false||Potassium Chloridenull|Potassium Drug Class|Drug|false|false||Potassium
null|Dietary Potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassiumnull|Potassium metabolic function|Finding|false|false||Potassiumnull|Potassium measurement|Procedure|false|false||Potassiumnull|chloride ion|Drug|false|false||Chloride
null|Chlorides|Drug|false|false||Chloridenull|Chloride metabolic function|Finding|false|false||Chloridenull|Chloride measurement|Procedure|false|false||Chloridenull|mEq|LabModifier|false|false||mEqnull|mEq|LabModifier|false|false||mEqnull|potassium chloride|Drug|false|false||Potassium Chloride
null|potassium chloride|Drug|false|false||Potassium Chloridenull|Potassium Drug Class|Drug|false|false||Potassium
null|Dietary Potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassiumnull|Potassium metabolic function|Finding|false|false||Potassiumnull|Potassium measurement|Procedure|false|false||Potassiumnull|chloride ion|Drug|false|false||Chloride
null|Chlorides|Drug|false|false||Chloridenull|Chloride metabolic function|Finding|false|false||Chloridenull|Chloride measurement|Procedure|false|false||Chloridenull|null|Time|false|false||prior tonull|null|Time|false|false||priornull|Transfer - product ownership|Finding|false|false||transfer
null|Transfer Technique|Finding|false|false||transfer
null|ActClass - transfer|Finding|false|false||transfer
null|null|Finding|false|false||transfernull|Transfer (immobility management)|Procedure|false|false||transfernull|arrival - ActRelationshipType|Finding|false|false||arrivalnull|null|Event|false|false||arrivalnull|Floor (anatomic)|Anatomy|false|false||floornull|floor (object)|Device|false|false||floornull|Floor - story of building|Entity|false|false||floornull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Chest Pain|Finding|true|false|C1527391;C0817096|chest painnull|null|Attribute|true|false|C1527391;C0817096|chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0008031;C0741025;C2926613|chest
null|Anterior thoracic region|Anatomy|false|false|C0008031;C0741025;C2926613|chestnull|Administration Method - Pain|Finding|true|false||pain
null|Pain|Finding|true|false||painnull|null|Attribute|true|false||painnull|Breath|Finding|false|false||breathnull|Palpitations|Finding|false|false||palpitationsnull|Lightheadedness|Finding|false|false||lightheadednessnull|Dizziness|Finding|false|false||dizziness
null|Vertigo|Finding|false|false||dizzinessnull|Review of systems (procedure)|Procedure|false|false||REVIEW OF SYSTEMSnull|null|Attribute|false|false||REVIEW OF SYSTEMS
null|null|Attribute|false|false||REVIEW OF SYSTEMSnull|Review of|Finding|false|false||REVIEW OFnull|Review (Publication Type)|Finding|false|false||REVIEW
null|Act Class - review|Finding|false|false||REVIEWnull|System|Finding|false|false||SYSTEMSnull|Proline dehydrogenase deficiency|Disorder|false|false||HPInull|History of present illness (finding)|Finding|false|false||HPI
null|allene oxide synthase activity|Finding|false|false||HPInull|Asthma|Disorder|false|false||ASTHMAnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|Encounter due to tobacco use|Finding|false|false||Tobacco use
null|Tobacco user|Finding|false|false||Tobacco use
null|History of tobacco use|Finding|false|false||Tobacco use
null|Tobacco use|Finding|false|false||Tobacco usenull|null|Attribute|false|false||Tobacco usenull|tobacco leaf allergenic extract|Drug|false|false||Tobacco
null|Tobacco|Drug|false|false||Tobacco
null|Tobacco|Drug|false|false||Tobacco
null|tobacco leaf allergenic extract|Drug|false|false||Tobacconull|Nicotiana tabacum|Entity|false|false||Tobacconull|Use - dosing instruction imperative|Finding|false|false||use
null|utilization qualifier|Finding|false|false||use
null|Usage|Finding|false|false||usenull|Peripheral Arterial Diseases|Disorder|false|false|C0003842|Peripheral Arterial disease
null|Peripheral Vascular Diseases|Disorder|false|false|C0003842|Peripheral Arterial diseasenull|Peripheral|Modifier|false|false||Peripheralnull|Arteriopathic disease|Disorder|false|false|C0003842|Arterial diseasenull|Arteries|Anatomy|false|false|C1704436;C0085096;C0852949|Arterialnull|Arterial|Modifier|false|false||Arterialnull|Disease|Disorder|false|false||diseasenull|Recent|Time|false|false||recentnull|Common Specifications in HL7 V3 Publishing|Finding|false|false|C0020889|common
null|shared attribute|Finding|false|false|C0020889|commonnull|Common (qualifier value)|LabModifier|false|false||commonnull|iliac stents|Procedure|false|false|C0020889|iliac stentingnull|Bone structure of ilium|Anatomy|false|false|C3245511;C1522138;C0850459;C2348535|iliacnull|Stenting|Procedure|false|false|C0020889|stentingnull|null|Device|false|false||stentingnull|Atrial tachycardia|Disorder|false|false|C0018792|ATRIAL TACHYCARDIAnull|continuous electrocardiogram atrial tachycardia|Finding|false|false|C0018792|ATRIAL TACHYCARDIAnull|Heart Atrium|Anatomy|false|false|C2059391;C0546959|ATRIALnull|Tachycardia by ECG Finding|Finding|false|false||TACHYCARDIA
null|Tachycardia|Finding|false|false||TACHYCARDIAnull|Atypical chest pain|Finding|false|false|C1527391;C0817096|ATYPICAL CHEST PAINnull|atypia morphology|Finding|false|false||ATYPICALnull|Atypical|Modifier|false|false||ATYPICALnull|Chest Pain|Finding|false|false|C1527391;C0817096|CHEST PAINnull|null|Attribute|false|false|C1527391;C0817096|CHEST PAINnull|Chest problem|Finding|false|false|C1527391;C0817096|CHESTnull|Chest|Anatomy|false|false|C0262384;C0008031;C0741025;C2926613|CHEST
null|Anterior thoracic region|Anatomy|false|false|C0262384;C0008031;C0741025;C2926613|CHESTnull|Administration Method - Pain|Finding|false|false||PAIN
null|Pain|Finding|false|false||PAINnull|null|Attribute|false|false||PAINnull|Cervical radiculitis|Disorder|false|false|C0027530|CERVICAL RADICULITISnull|Neck|Anatomy|false|false|C0034544;C0263884|CERVICALnull|Cervical|Modifier|false|false||CERVICALnull|Radiculitis|Disorder|false|false|C0027530|RADICULITISnull|Cervical spondylosis without myelopathy|Disorder|false|false|C0027530|CERVICAL SPONDYLOSIS
null|Cervical spondylosis|Disorder|false|false|C0027530|CERVICAL SPONDYLOSISnull|Neck|Anatomy|false|false|C0158241;C1384641;C0038019|CERVICALnull|Cervical|Modifier|false|false||CERVICALnull|Spondylosis|Disorder|false|false|C0027530|SPONDYLOSISnull|Coronary artery|Anatomy|false|false||CORONARY ARTERYnull|Heart|Anatomy|false|false||CORONARYnull|Coronary|Modifier|false|false||CORONARYnull|Arterial system|Anatomy|false|false||ARTERY
null|Arteries|Anatomy|false|false||ARTERYnull|Disease|Disorder|false|false||DISEASEnull|Headache|Finding|false|false||HEADACHEnull|Prosthetic arthroplasty of hip (procedure)|Procedure|false|false|C0022122;C0228391;C0019552;C4299095|HIP REPLACEMENTnull|heme iron polypeptide|Drug|false|false|C0022122;C0228391;C0019552;C4299095|HIP
null|ST13 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|HIP
null|ST13 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|HIP
null|RPL29 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|HIP
null|RPL29 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|HIP
null|HHIP protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|HIP
null|HHIP protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|HIP
null|heme iron polypeptide|Drug|false|false|C0022122;C0228391;C0019552;C4299095|HIPnull|RPL29 wt Allele|Finding|false|false|C0022122;C0228391;C0019552;C4299095|HIP
null|REG3A gene|Finding|false|false|C0022122;C0228391;C0019552;C4299095|HIP
null|RPL29 gene|Finding|false|false|C0022122;C0228391;C0019552;C4299095|HIP
null|ST13 wt Allele|Finding|false|false|C0022122;C0228391;C0019552;C4299095|HIP
null|ST13 gene|Finding|false|false|C0022122;C0228391;C0019552;C4299095|HIP
null|HHIP gene|Finding|false|false|C0022122;C0228391;C0019552;C4299095|HIP
null|HHIP wt Allele|Finding|false|false|C0022122;C0228391;C0019552;C4299095|HIP
null|REG3A wt Allele|Finding|false|false|C0022122;C0228391;C0019552;C4299095|HIPnull|Procedure on hip|Procedure|false|false|C0022122;C0228391;C0019552;C4299095|HIPnull|Lower extremity>Hip|Anatomy|false|false|C0559956;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C1430701;C0529134;C1505163;C1654726;C0392806;C1292890;C1555302;C0035139|HIP
null|Hip structure|Anatomy|false|false|C0559956;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C1430701;C0529134;C1505163;C1654726;C0392806;C1292890;C1555302;C0035139|HIP
null|Structure of habenulopeduncular tract|Anatomy|false|false|C0559956;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C1430701;C0529134;C1505163;C1654726;C0392806;C1292890;C1555302;C0035139|HIP
null|Bone structure of ischium|Anatomy|false|false|C0559956;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C1430701;C0529134;C1505163;C1654726;C0392806;C1292890;C1555302;C0035139|HIPnull|Replacement|Finding|false|false|C0022122;C0228391;C0019552;C4299095|REPLACEMENTnull|Replacement - supply|Procedure|false|false|C0022122;C0228391;C0019552;C4299095|REPLACEMENT
null|Surgical Replantation|Procedure|false|false|C0022122;C0228391;C0019552;C4299095|REPLACEMENTnull|Hyperlipidemia|Disorder|false|false||HYPERLIPIDEMIA
null|Hyperlipoproteinemias|Disorder|false|false||HYPERLIPIDEMIAnull|Serum lipids high (finding)|Finding|false|false||HYPERLIPIDEMIAnull|Hypertensive disease|Disorder|false|false||HYPERTENSIONnull|Degenerative polyarthritis|Disorder|false|false||OSTEOARTHRITISnull|Herpes zoster (disorder)|Disorder|false|false||HERPES ZOSTER
null|herpesvirus 3, human|Disorder|false|false||HERPES ZOSTERnull|Herpes simplex dermatitis|Disorder|false|false||HERPES
null|null|Disorder|false|false||HERPESnull|Herpes <Hyperinae>|Entity|false|false||HERPESnull|Herpes zoster (disorder)|Disorder|false|false||ZOSTERnull|Tobacco Use Disorder|Disorder|false|false||TOBACCO ABUSEnull|tobacco leaf allergenic extract|Drug|false|false||TOBACCO
null|Tobacco|Drug|false|false||TOBACCO
null|Tobacco|Drug|false|false||TOBACCO
null|tobacco leaf allergenic extract|Drug|false|false||TOBACCOnull|Nicotiana tabacum|Entity|false|false||TOBACCOnull|Drug abuse|Disorder|false|false||ABUSEnull|Victim of abuse (finding)|Finding|false|false||ABUSEnull|Abuse|Event|false|false||ABUSEnull|Heart Atrium|Anatomy|false|false||ATRIALnull|Fibrillation|Disorder|false|false||FIBRILLATIONnull|Anxiety Disorders|Disorder|false|false||ANXIETY
null|Anxiety|Disorder|false|false||ANXIETYnull|Anxiety symptoms|Finding|false|false||ANXIETYnull|Gastrointestinal Hemorrhage|Finding|false|false||GASTROINTESTINAL BLEEDINGnull|Gastrointestinal attachment|Finding|false|false||GASTROINTESTINALnull|gastrointestinal|Modifier|false|false||GASTROINTESTINALnull|Hemorrhage|Finding|false|false||BLEEDINGnull|Degenerative polyarthritis|Disorder|false|false||OSTEOARTHRITISnull|Atherosclerosis|Disorder|false|false|C0007226;C3887460|ATHEROSCLEROTIC CARDIOVASCULAR DISEASEnull|atherosclerotic|Finding|false|false||ATHEROSCLEROTICnull|Cardiovascular Diseases|Disorder|false|false|C0007226;C3887460|CARDIOVASCULAR DISEASEnull|Cardiovascular system|Anatomy|false|false|C0085096;C0004153;C0012634;C0007222|CARDIOVASCULAR
null|Cardiovascular|Anatomy|false|false|C0085096;C0004153;C0012634;C0007222|CARDIOVASCULARnull|Peripheral Vascular Diseases|Disorder|false|false|C0005847;C0007226;C3887460|DISEASE, PERIPHERAL VASCULARnull|Disease|Disorder|false|false|C0007226;C3887460|DISEASEnull|Peripheral|Modifier|false|false||PERIPHERALnull|Blood Vessel|Anatomy|false|false|C0085096|VASCULARnull|Vascular|Modifier|false|false||VASCULARnull|Disease|Disorder|false|false||DISEASEnull|reported history of cataract surgery|Finding|false|false||CATARACT SURGERY
null|Consent Type - Cataract Surgery|Finding|false|false||CATARACT SURGERYnull|Cataract surgery|Procedure|false|false||CATARACT SURGERY
null|Cataract Extraction|Procedure|false|false||CATARACT SURGERYnull|Cataract surgery specialty (qualifier value)|Title|false|false||CATARACT SURGERYnull|Cataract|Disorder|false|false||CATARACTnull|cataract on exam (physical finding)|Finding|false|false||CATARACTnull|Level of Care - Surgery|Finding|false|false||SURGERY
null|Surgical procedure finding|Finding|false|false||SURGERY
null|Surgical aspects|Finding|false|false||SURGERYnull|Operative Surgical Procedures|Procedure|false|false||SURGERYnull|General surgery specialty|Title|false|false||SURGERY
null|Surgery specialty|Title|false|false||SURGERYnull|Level of Care - Surgery|Finding|false|false||Surgery
null|Surgical procedure finding|Finding|false|false||Surgery
null|Surgical aspects|Finding|false|false||Surgerynull|Operative Surgical Procedures|Procedure|false|false||Surgerynull|General surgery specialty|Title|false|false||Surgery
null|Surgery specialty|Title|false|false||Surgerynull|Bilateral|Modifier|false|false||BILATERALnull|Common iliac artery structure|Anatomy|false|false|C2348535;C3245511;C1522138|COMMON ILIAC ARTERYnull|Common Specifications in HL7 V3 Publishing|Finding|false|false|C1261084;C0020887|COMMON
null|shared attribute|Finding|false|false|C1261084;C0020887|COMMONnull|Common (qualifier value)|LabModifier|false|false||COMMONnull|Structure of iliac artery|Anatomy|false|false|C2348535;C3245511;C1522138|ILIAC ARTERYnull|Bone structure of ilium|Anatomy|false|false||ILIACnull|Arterial system|Anatomy|false|false|C2348535|ARTERY
null|Arteries|Anatomy|false|false|C2348535|ARTERYnull|Stenting|Procedure|false|false|C1261084;C0226004;C0003842;C0020887|STENTINGnull|null|Device|false|false||STENTINGnull|Silver bunionectomy|Procedure|false|false||BUNIONECTOMYnull|Prosthetic arthroplasty of hip (procedure)|Procedure|false|false|C0022122;C0228391;C0019552;C4299095|HIP REPLACEMENTnull|heme iron polypeptide|Drug|false|false|C0022122;C0228391;C0019552;C4299095|HIP
null|ST13 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|HIP
null|ST13 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|HIP
null|RPL29 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|HIP
null|RPL29 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|HIP
null|HHIP protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|HIP
null|HHIP protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|HIP
null|heme iron polypeptide|Drug|false|false|C0022122;C0228391;C0019552;C4299095|HIPnull|RPL29 wt Allele|Finding|false|false|C0022122;C0228391;C0019552;C4299095|HIP
null|REG3A gene|Finding|false|false|C0022122;C0228391;C0019552;C4299095|HIP
null|RPL29 gene|Finding|false|false|C0022122;C0228391;C0019552;C4299095|HIP
null|ST13 wt Allele|Finding|false|false|C0022122;C0228391;C0019552;C4299095|HIP
null|ST13 gene|Finding|false|false|C0022122;C0228391;C0019552;C4299095|HIP
null|HHIP gene|Finding|false|false|C0022122;C0228391;C0019552;C4299095|HIP
null|HHIP wt Allele|Finding|false|false|C0022122;C0228391;C0019552;C4299095|HIP
null|REG3A wt Allele|Finding|false|false|C0022122;C0228391;C0019552;C4299095|HIPnull|Procedure on hip|Procedure|false|false|C0022122;C0228391;C0019552;C4299095|HIPnull|Lower extremity>Hip|Anatomy|false|false|C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C1430701;C0529134;C1505163;C1654726;C0392806;C1555302;C0035139;C0559956;C1292890|HIP
null|Hip structure|Anatomy|false|false|C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C1430701;C0529134;C1505163;C1654726;C0392806;C1555302;C0035139;C0559956;C1292890|HIP
null|Structure of habenulopeduncular tract|Anatomy|false|false|C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C1430701;C0529134;C1505163;C1654726;C0392806;C1555302;C0035139;C0559956;C1292890|HIP
null|Bone structure of ischium|Anatomy|false|false|C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C1430701;C0529134;C1505163;C1654726;C0392806;C1555302;C0035139;C0559956;C1292890|HIPnull|Replacement|Finding|false|false|C0022122;C0228391;C0019552;C4299095|REPLACEMENTnull|Replacement - supply|Procedure|false|false|C0022122;C0228391;C0019552;C4299095|REPLACEMENT
null|Surgical Replantation|Procedure|false|false|C0022122;C0228391;C0019552;C4299095|REPLACEMENTnull|null|Time|false|false||PRIORnull|Cesarean section|Procedure|false|false||CESAREAN SECTIONnull|Cesarean|Procedure|false|false||CESAREANnull|section sample|Drug|false|false||SECTIONnull|Html Link Type - section|Finding|false|false||SECTION
null|Act Class - Section|Finding|false|false||SECTIONnull|Sectioning technique|Procedure|false|false||SECTIONnull|Section - Geographic Area|Entity|false|false||SECTION
null|Section (object)|Entity|false|false||SECTIONnull|Square Mile|LabModifier|false|false||SECTIONnull|Synovial Cyst|Disorder|false|false|C0017067|GANGLION CYST
null|Myxoid cyst|Disorder|false|false|C0017067|GANGLION CYSTnull|Synovial Cyst|Disorder|false|false|C0017067|GANGLION
null|Myxoid cyst|Disorder|false|false|C0017067|GANGLIONnull|Ganglia|Anatomy|false|false|C1258666;C0085648;C1258666;C0085648;C0010709;C1546594;C1550626|GANGLIONnull|Cyst|Disorder|false|false|C0017067|CYSTnull|SpecimenType - Cyst|Finding|false|false|C0017067|CYST
null|null|Finding|false|false|C0017067|CYSTnull|Cyst form of protozoa|Entity|false|false||CYSTnull|Relationship - Mother|Finding|false|false||Mothernull|Mother (person)|Subject|false|false||Mothernull|Hypertensive disease|Disorder|false|false||HTNnull|Indirect exposure mechanism - Father|Finding|false|false||Father
null|Relationship - Father|Finding|false|false||Father
null|Father - courtesy title|Finding|false|false||Fathernull|Father (person)|Subject|false|false||Fathernull|Brother - courtesy title|Finding|false|false||Brother
null|Relationship - Brother|Finding|false|false||Brothernull|Brothers|Subject|false|false||Brothernull|Brother - courtesy title|Finding|false|false||Brother
null|Relationship - Brother|Finding|false|false||Brothernull|Brothers|Subject|false|false||Brothernull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||Generalnull|General medical service|Procedure|false|false||Generalnull|Generalized|Modifier|false|false||Generalnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Admission Level of Care Code - Acute|Finding|true|false||acute
null|Acute - Triage Code|Finding|true|false||acutenull|acute|Time|false|false||acutenull|Emotional distress|Finding|true|false||distress
null|Distress|Finding|true|false||distressnull|HEENT|Anatomy|false|false||HEENTnull|Scleral Diseases|Disorder|false|false|C0036410|Scleranull|examination of sclera|Procedure|false|false|C0036410|Scleranull|Sclera|Anatomy|false|false|C2228481;C0205180;C0026987;C0036412|Scleranull|Anicteric|Finding|false|false|C0036410|anictericnull|Myelofibrosis|Disorder|false|false|C0694605;C0036410|MMMnull|Medial part of medial mammillary nucleus|Anatomy|false|false|C0026987|MMMnull|Oropharyngeal|Anatomy|false|false|C1550016|oropharynxnull|Remote control command - Clear|Finding|false|false|C0521367|clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|Pupil equal round and reacting to light|Finding|false|false||PERRLnull|Passive joint movement of neck (finding)|Finding|false|false|C0027530;C3159206|Neck
null|Neck problem|Finding|false|false|C0027530;C3159206|Necknull|dendritic spine neck|Anatomy|false|false|C0812434;C0684335|Neck
null|Neck|Anatomy|false|false|C0812434;C0684335|Necknull|Supple|Finding|false|false||Supplenull|Jugular venous pressure|Finding|false|false||JVPnull|Elevated|Modifier|false|false||elevated
null|High|Modifier|false|false||elevatednull|Leukocyte adhesion deficiency type 1|Disorder|true|false|C0226032|LAD
null|Leukocyte adhesion deficiency|Disorder|true|false|C0226032|LADnull|ITGB2 wt Allele|Finding|true|false|C0226032|LAD
null|DLD gene|Finding|true|false|C0226032|LADnull|Anterior descending branch of left coronary artery|Anatomy|true|false|C1414063;C1706333;C5550999;C0398738|LADnull|Ladino Language|Entity|true|false||LADnull|Regular|Modifier|false|false||Regularnull|Amount type - Rate|Finding|false|false||ratenull|Rating (action)|Event|false|false||ratenull|Rate|LabModifier|false|false||ratenull|Rhythm|Finding|false|false||rhythm
null|rhythmic process (biological)|Finding|false|false||rhythmnull|Systolic Murmurs|Finding|false|false||systolic murmurnull|Systole|Finding|false|false||systolicnull|Heart murmur|Finding|false|false||murmurnull|Pericardial friction rub|Finding|true|false||rubsnull|Lung|Anatomy|false|false||Lungsnull|Inspiration (function)|Finding|false|false||inspiratorynull|Expiratory wheezing|Finding|false|false||expiratory wheezesnull|Expiration, Respiratory|Finding|false|false||expiratorynull|Wheezing|Finding|false|false||wheezesnull|Basilar Rales|Finding|true|false||rales
null|Rales|Finding|true|false||ralesnull|Rhonchi|Finding|true|false||rhonchinull|Malignant neoplasm of abdomen|Disorder|false|false|C0230168;C0000726|Abdomennull|Abdomen problem|Finding|false|false|C0230168;C0000726|Abdomennull|Abdomen|Anatomy|false|false|C0153662;C0941288|Abdomen
null|Abdominal Cavity|Anatomy|false|false|C0153662;C0941288|Abdomennull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||Softnull|Soft|Modifier|false|false||Softnull|Bowel sounds|Finding|false|false|C0021853|bowel soundsnull|Intestines|Anatomy|false|false|C0232693|bowelnull|null|Device|false|false||soundsnull|null|Phenomenon|false|false||soundsnull|Present|Finding|false|false||present
null|Presentation|Finding|false|false||presentnull|Organomegaly|Finding|true|false||organomegalynull|Protective muscle spasm|Finding|true|false||guardingnull|Hereditary Multiple Exostoses|Disorder|false|false||Extnull|EXT1 wt Allele|Finding|false|false||Ext
null|EXT1 gene|Finding|false|false||Extnull|Feels warm|Finding|false|false||Warmnull|warming process|Phenomenon|false|false||Warmnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false||pulsesnull|Clubbing|Disorder|true|false||clubbingnull|Cyanosis|Finding|true|false||cyanosisnull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|infant weight for previous delivery (history)|Finding|false|false||Weight
null|Weight symptom (finding)|Finding|false|false||Weightnull|Weighing patient|Procedure|false|false||Weightnull|null|Attribute|false|false||Weightnull|Body Weight|Subject|false|false||Weightnull|Importance Weight|Modifier|false|false||Weightnull|Weight|LabModifier|false|false||Weightnull|infant weight for previous delivery (history)|Finding|false|false||Weight
null|Weight symptom (finding)|Finding|false|false||Weightnull|Weighing patient|Procedure|false|false||Weightnull|null|Attribute|false|false||Weightnull|Body Weight|Subject|false|false||Weightnull|Importance Weight|Modifier|false|false||Weightnull|Weight|LabModifier|false|false||Weightnull|On admission|Time|false|false||on admissionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||Generalnull|General medical service|Procedure|false|false||Generalnull|Generalized|Modifier|false|false||Generalnull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|HEENT|Anatomy|false|false||HEENTnull|Scleral Diseases|Disorder|false|false|C0036410|Scleranull|examination of sclera|Procedure|false|false|C0036410|Scleranull|Sclera|Anatomy|false|false|C2228481;C0036412;C0205180|Scleranull|Anicteric|Finding|false|false|C0036410|anictericnull|Passive joint movement of neck (finding)|Finding|false|false|C0027530;C3159206|Neck
null|Neck problem|Finding|false|false|C0027530;C3159206|Necknull|dendritic spine neck|Anatomy|false|false|C0812434;C0684335|Neck
null|Neck|Anatomy|false|false|C0812434;C0684335|Necknull|Jugular venous pressure|Finding|false|false||JVPnull|Elevated|Modifier|false|false||elevated
null|High|Modifier|false|false||elevatednull|Regular|Modifier|false|false||Regularnull|Rhythm|Finding|false|false||rhythm
null|rhythmic process (biological)|Finding|false|false||rhythmnull|Frequently|Time|false|false||frequentnull|Systolic Murmurs|Finding|false|false||systolic murmurnull|Systole|Finding|false|false||systolicnull|Heart murmur|Finding|false|false||murmurnull|Pericardial friction rub|Finding|true|false||rubsnull|Lung|Anatomy|false|false||Lungsnull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Expiratory wheezing|Finding|false|false||expiratory wheezesnull|Expiration, Respiratory|Finding|false|false||expiratorynull|Wheezing|Finding|false|false||wheezesnull|Diffuse|Modifier|false|false||diffusenull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Rhonchi|Finding|false|false||rhonchinull|Malignant neoplasm of abdomen|Disorder|false|false|C0230168;C0000726|Abdomennull|Abdomen problem|Finding|false|false|C0230168;C0000726|Abdomennull|Abdomen|Anatomy|false|false|C0153662;C0941288|Abdomen
null|Abdominal Cavity|Anatomy|false|false|C0153662;C0941288|Abdomennull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||Softnull|Soft|Modifier|false|false||Softnull|Bowel sounds|Finding|false|false|C0021853|bowel soundsnull|Intestines|Anatomy|false|false|C0232693|bowelnull|null|Device|false|false||soundsnull|null|Phenomenon|false|false||soundsnull|Present|Finding|false|false||present
null|Presentation|Finding|false|false||presentnull|Organomegaly|Finding|true|false||organomegalynull|Protective muscle spasm|Finding|true|false||guardingnull|Hereditary Multiple Exostoses|Disorder|false|false||Extnull|EXT1 wt Allele|Finding|false|false||Ext
null|EXT1 gene|Finding|false|false||Extnull|Feels warm|Finding|false|false||Warmnull|warming process|Phenomenon|false|false||Warmnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Edema|Finding|true|false||edemanull|null|Attribute|true|false||edemanull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|Laboratory test finding|Lab|false|false||Labsnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|lactate|Drug|false|false||LACTATE
null|lactate|Drug|false|false||LACTATE
null|Lactates|Drug|false|false||LACTATEnull|Lactic acid measurement|Procedure|false|false||LACTATEnull|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSEnull|Glucose measurement|Procedure|false|false||GLUCOSEnull|Glucose^1.5H post dose glucagon|Lab|false|false||GLUCOSEnull|urea|Drug|false|false||UREA
null|urea|Drug|false|false||UREA
null|urea|Drug|false|false||UREAnull|Urea measurement|Procedure|false|false||UREAnull|Sodium supplements|Drug|false|false||SODIUM
null|sodium|Drug|false|false||SODIUM
null|sodium|Drug|false|false||SODIUM
null|Sodium Drug Class|Drug|false|false||SODIUMnull|Sodium metabolic function|Finding|false|false||SODIUMnull|Sodium measurement|Procedure|false|false||SODIUMnull|Potassium Drug Class|Drug|false|false||POTASSIUM
null|Dietary Potassium|Drug|false|false||POTASSIUM
null|potassium|Drug|false|false||POTASSIUM
null|potassium|Drug|false|false||POTASSIUM
null|potassium|Drug|false|false||POTASSIUM
null|Potassium supplement|Drug|false|false||POTASSIUM
null|Potassium supplement|Drug|false|false||POTASSIUMnull|Potassium metabolic function|Finding|false|false||POTASSIUMnull|Potassium measurement|Procedure|false|false||POTASSIUMnull|chloride ion|Drug|false|false||CHLORIDE
null|Chlorides|Drug|false|false||CHLORIDEnull|Chloride metabolic function|Finding|false|false||CHLORIDEnull|Chloride measurement|Procedure|false|false||CHLORIDEnull|Total|Modifier|false|false||TOTALnull|carbon dioxide|Drug|false|false||CO2
null|carbon dioxide|Drug|false|false||CO2null|MT-CO2 gene|Finding|false|false||CO2
null|null|Finding|false|false||CO2
null|C2 wt Allele|Finding|false|false||CO2null|blood anion gap (lab test)|Procedure|false|false||ANION GAP
null|Anion gap measurement|Procedure|false|false||ANION GAPnull|Anion Gap|Attribute|false|false||ANION GAPnull|Anion gap result|Lab|false|false||ANION GAPnull|Anions|Drug|false|false||ANIONnull|Ras GTPase-Activating Protein 1, Human|Drug|false|false||GAP
null|Ras GTPase-Activating Protein 1, Human|Drug|false|false||GAP
null|GTPase-Activating Proteins|Drug|false|false||GAP
null|GTPase-Activating Proteins|Drug|false|false||GAPnull|RASA1 wt Allele|Finding|false|false||GAP
null|RASA1 gene|Finding|false|false||GAPnull|Gap (space)|Modifier|false|false||GAPnull|CALCIUM SUPPLEMENTS|Drug|false|false||CALCIUM
null|calcium|Drug|false|false||CALCIUM
null|calcium|Drug|false|false||CALCIUM
null|calcium|Drug|false|false||CALCIUM
null|CALCIUM SUPPLEMENTS|Drug|false|false||CALCIUM
null|Calcium, Dietary|Drug|false|false||CALCIUM
null|Calcium [EPC]|Drug|false|false||CALCIUM
null|Calcium Drug Class|Drug|false|false||CALCIUMnull|Calcium metabolic function|Finding|false|false||CALCIUMnull|Calcium measurement|Procedure|false|false||CALCIUMnull|phosphate ion|Drug|false|false||PHOSPHATE
null|Phosphates|Drug|false|false||PHOSPHATE
null|phosphate ion|Drug|false|false||PHOSPHATEnull|Phosphate measurement|Procedure|false|false||PHOSPHATEnull|Magnesium supplements, alimentary tract and metabolism|Drug|false|false||MAGNESIUM
null|magnesium|Drug|false|false||MAGNESIUM
null|magnesium|Drug|false|false||MAGNESIUM
null|Magnesium Drug Class|Drug|false|false||MAGNESIUM
null|Magnesium supplements, alimentary tract and metabolism|Drug|false|false||MAGNESIUMnull|Magnesium measurement|Procedure|false|false||MAGNESIUMnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C0014792;C1114281|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||HGB
null|Hemoglobin|Drug|false|false||HGBnull|CYGB gene|Finding|false|false||HGBnull|Hemoglobin concentration|Lab|false|false||HGBnull|Hemopoietic stem cell transplant|Procedure|false|false||HCT
null|Hematocrit Measurement|Procedure|false|false||HCTnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Monos|Drug|false|false||MONOS
null|Mono-S|Drug|false|false||MONOS
null|Monos|Drug|false|false||MONOSnull|SARCOIDOSIS, EARLY-ONSET|Disorder|false|false||EOS
null|Familial eosinophilia|Disorder|false|false||EOSnull|PRSS33 gene|Finding|false|false||EOS
null|IKZF4 gene|Finding|false|false||EOSnull|Eos <Loriini>|Entity|false|false||EOSnull|Primed lymphocyte test|Procedure|false|false||PLTnull|Count Dosing Unit|LabModifier|false|false||COUNT
null|Count|LabModifier|false|false||COUNTnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Laboratory test finding|Lab|false|false||Labsnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0851353;C0005768;C0229664;C0005767|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C0014792;C1114281|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Alanine Transaminase|Drug|false|false||ALT
null|Alanine Transaminase|Drug|false|false||ALTnull|Liposarcoma, well differentiated|Disorder|false|false|C1185650|ALT
null|Atypical Lipoma|Disorder|false|false|C1185650|ALTnull|null|Finding|false|false|C1185650|ALT
null|Alternative Billing Concepts|Finding|false|false|C1185650|ALT
null|GPT gene|Finding|false|false|C1185650|ALTnull|Antibiotic Lock Therapy|Procedure|false|false|C1185650|ALTnull|Southern Altai Language|Entity|false|false||ALTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false|C1185650|AST
null|Aspartate Transaminase|Drug|false|false|C1185650|AST
null|Aspartate Transaminase|Drug|false|false|C1185650|AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false|C1185650|AST
null|SLC17A5 protein, human|Drug|false|false|C1185650|AST
null|SLC17A5 protein, human|Drug|false|false|C1185650|ASTnull|Atypical Spitz Nevus|Disorder|false|false|C1185650|ASTnull|SLC17A5 wt Allele|Finding|false|false|C1185650|AST
null|SLC17A5 gene|Finding|false|false|C1185650|AST
null|GOT1 gene|Finding|false|false|C1185650|ASTnull|Asterion|Anatomy|false|false|C2257651;C1415274;C1140170;C4553172;C1266129;C1370889;C4522245;C0004002;C0242192;C1121182;C1415181;C1420113;C5960784;C0202113;C0851148|ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|Lactate Dehydrogenase|Drug|false|false||LDH
null|Lactate Dehydrogenase|Drug|false|false||LDHnull|Lifetime Drinking History|Finding|false|false|C1185650|LDHnull|Lactate dehydrogenase measurement|Procedure|false|false|C1185650|LDHnull|Alkaline Phosphatase|Drug|false|false||AlkPhos
null|Alkaline Phosphatase|Drug|false|false||AlkPhosnull|Blood calcium measurement|Procedure|false|false||BLOOD Calciumnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Scientific Study|Procedure|false|false||Studiesnull|Plain chest X-ray|Procedure|false|false||CXRnull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Cardiovascular disease+Pulmonary disease|Disorder|false|false|C1184743;C0553534|cardiopulmonarynull|Cardiopulmonary|Anatomy|false|false|C4521054;C4072686;C1522240|cardiopulmonarynull|Process Pharmacologic Substance|Drug|true|false|C1184743|processnull|Process (qualifier value)|Finding|true|false|C0553534;C1184743|processnull|bony process|Anatomy|false|false|C4072686;C1522240;C4521054;C1951340|processnull|Process|Phenomenon|true|false|C1184743;C0553534|processnull|Exercise stress test - endocrine|Procedure|false|false|C4318744|Exercise stress test
null|Exercise stress test|Procedure|false|false|C4318744|Exercise stress testnull|Exercise|Finding|false|false|C4318744|Exercisenull|Exercise Pain Management|Procedure|false|false|C4318744|Exercisenull|Exercise stress test|Procedure|false|false|C4318744|stress test
null|Stress Test|Procedure|false|false|C4318744|stress testnull|Stress bismuth subsalicylate|Drug|false|false||stress
null|Stress bismuth subsalicylate|Drug|false|false||stressnull|Stress|Finding|false|false|C4318744|stressnull|W stress|Attribute|false|false||stressnull|Tests (qualifier value)|Finding|false|false|C4318744|test
null|Testing|Finding|false|false|C4318744|testnull|Laboratory Procedures|Procedure|false|false|C4318744|testnull|Test - temporal region|Anatomy|false|false|C0039593;C0392366;C0015259;C0015260;C3494508;C0456984;C0038435;C1522704;C0430120;C0015260;C0022885|testnull|Test Result|Lab|false|false|C4318744|testnull|Test Dosing Unit|LabModifier|false|false||testnull|Interpretation Process|Finding|false|false||INTERPRETATIONnull|null|Attribute|false|false||INTERPRETATIONnull|Transaction counts and value totals - year|Finding|false|false||year
null|Precision - year|Finding|false|false||yearnull|year|Time|false|false||yearnull|Old|Time|false|false||oldnull|Woman|Subject|false|false||woman
null|Human, Female adult|Subject|false|false||womannull|Medical History|Finding|false|false|C3669270|history ofnull|History of present illness (finding)|Finding|false|false|C3669270|history
null|History of previous events|Finding|false|false|C3669270|history
null|Historical aspects qualifier|Finding|false|false|C3669270|history
null|Medical History|Finding|false|false|C3669270|history
null|Concept History|Finding|false|false|C3669270|historynull|History|Subject|false|false||historynull|Pad Dosage Form|Drug|false|false|C3669270|PADnull|Pad Mass|Disorder|false|false|C3669270|PAD
null|Peripheral Arterial Diseases|Disorder|false|false|C3669270|PADnull|PADI4 wt Allele|Finding|false|false|C3669270|PAD
null|PADI4 gene|Finding|false|false|C3669270|PAD
null|DHX40 gene|Finding|false|false|C3669270|PADnull|PAD Regimen|Procedure|false|false|C3669270|PADnull|Strucure of thick cushion of skin|Anatomy|false|false|C2347441;C0332568;C1704436;C0262926;C0262926;C1705255;C0019665;C0262512;C2004062;C3540603;C1425478;C1425244;C3814046|PADnull|Pad Device|Device|false|false||PAD
null|Pads|Device|false|false||PADnull|Pad (unit of presentation)|LabModifier|false|false||PAD
null|Pad Dosing Unit|LabModifier|false|false||PADnull|Left Bundle-Branch Block|Disorder|false|false||LBBBnull|null|Lab|false|false||LBBBnull|AML Lab Table|Finding|true|false||lab
null|LAT2 gene|Finding|true|false||lab
null|EWS Lab Table|Finding|true|false||labnull|Laboratory|Device|true|false||labnull|Labrador retriever|Entity|true|false||lab
null|Laboratory|Entity|true|false||labnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Periodicals|Finding|false|false||serialnull|Serial|Time|false|false||serialnull|Cardiac markers|Procedure|false|false|C0018787|cardiac markersnull|Cardiac attachment|Finding|false|false|C0018787|cardiacnull|Heart|Anatomy|false|false|C1271630;C0741025;C1314974;C2364135;C0235710|cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||cardiacnull|Marker Device|Device|false|false||markersnull|Processing type - Evaluation|Finding|false|false||evaluationnull|Evaluation procedure|Procedure|false|false||evaluation
null|Evaluation|Procedure|false|false||evaluationnull|Chest discomfort|Finding|false|false|C1527391;C0817096;C0018787|chest discomfortnull|Chest problem|Finding|false|false|C0018787;C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0235710;C2364135;C0741025|chest
null|Anterior thoracic region|Anatomy|false|false|C0235710;C2364135;C0741025|chestnull|Discomfort|Finding|false|false|C1527391;C0817096;C0018787|discomfortnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|dipyridamole|Drug|false|false||dipyridamole
null|dipyridamole|Drug|false|false||dipyridamolenull|Exercise stress test|Procedure|false|false|C4318744|stress test
null|Stress Test|Procedure|false|false|C4318744|stress testnull|Stress bismuth subsalicylate|Drug|false|false||stress
null|Stress bismuth subsalicylate|Drug|false|false||stressnull|Stress|Finding|false|false|C4318744|stressnull|W stress|Attribute|false|false||stressnull|Tests (qualifier value)|Finding|false|false|C4318744|test
null|Testing|Finding|false|false|C4318744|testnull|Laboratory Procedures|Procedure|false|false|C4318744|testnull|Test - temporal region|Anatomy|false|false|C0022885;C0456984;C0039593;C0392366;C0015260;C3494508;C0038435|testnull|Test Result|Lab|false|false|C4318744|testnull|Test Dosing Unit|LabModifier|false|false||testnull|theophylline|Drug|false|false||theophylline
null|theophylline|Drug|false|false||theophyllinenull|Assay of theophylline|Procedure|false|false||theophyllinenull|Therapy Object (animal model)|Finding|false|false||therapy
null|therapeutic aspects|Finding|false|false||therapynull|Therapeutic procedure|Procedure|false|false||therapynull|Able (qualifier value)|Finding|false|false||ablenull|Ability|Subject|false|false||ablenull|Frequently|Time|false|false||frequentnull|Heart Atrium|Anatomy|false|false||atrialnull|dobutamine|Drug|false|false||dobutamine
null|dobutamine|Drug|false|false||dobutaminenull|Walking (function)|Finding|false|false||walknull|Treadmill (physical activity)|Finding|false|false||treadmillnull|treadmill conditioning training|Procedure|false|false||treadmillnull|null|Device|false|false||treadmillnull|Minute of time|Time|false|false||minutesnull|Minute Unit of Plane Angle|LabModifier|false|false||minutes
null|Minute (diminutive)|LabModifier|false|false||minutes
null|Small|LabModifier|false|false||minutesnull|Changing|Finding|false|false||modifiednull|Protocol - answer to question|Finding|false|false||protocol
null|Study Protocol|Finding|false|false||protocol
null|Protocols documentation|Finding|false|false||protocol
null|Clinical trial protocol document|Finding|false|false||protocol
null|Library Protocol|Finding|false|false||protocolnull|Leg|Anatomy|false|false|C0021775;C1456822;C0311395|leg
null|Lower Extremity|Anatomy|false|false|C0021775;C1456822;C0311395|legnull|Intermittent Claudication|Disorder|false|false|C1140621;C0023216|claudicationnull|Claudication (finding)|Finding|false|false|C1140621;C0023216|claudication
null|Lameness|Finding|false|false|C1140621;C0023216|claudicationnull|Peak level|Modifier|false|false||peaknull|Capacity|LabModifier|false|false||capacitynull|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group|Finding|false|false||poor
null|Patient Condition Code - Poor|Finding|false|false||poornull|Poverty|Subject|false|false||poornull|Language Proficiency - Poor|Modifier|false|false||poor
null|Specimen Quality - Poor|Modifier|false|false||poor
null|Poor - grade|Modifier|false|false||poor
null|Poor - qualifier|Modifier|false|false||poornull|Functional capacity|Finding|false|false||functional capacitynull|Functional Relationship|Finding|false|false||functional
null|Function (attribute)|Finding|false|false||functional
null|Functional|Finding|false|false||functionalnull|Capacity|LabModifier|false|false||capacitynull|Glycation End Products, Advanced|Drug|false|false||age
null|Glycation End Products, Advanced|Drug|false|false||agenull|null|Attribute|false|false||agenull|Age|Subject|false|false||agenull|Anorectal Malformations|Disorder|true|false|C0446516;C1140618;C1269078|armnull|AKR1A1 wt Allele|Finding|true|false|C0446516;C1140618;C1269078|arm
null|ARMC9 gene|Finding|true|false|C0446516;C1140618;C1269078|armnull|Protocol Treatment Arm|Procedure|true|false|C0446516;C1140618;C1269078|arm
null|Axillary Reverse Mapping|Procedure|true|false|C0446516;C1140618;C1269078|arm
null|Study Arm|Procedure|true|false|C0446516;C1140618;C1269078|armnull|Upper arm|Anatomy|false|false|C1824218;C3715044;C1522541;C5400986;C4761640;C3495676;C0812434;C0684335|arm
null|null|Anatomy|false|false|C1824218;C3715044;C1522541;C5400986;C4761640;C3495676;C0812434;C0684335|arm
null|Upper Extremity|Anatomy|false|false|C1824218;C3715044;C1522541;C5400986;C4761640;C3495676;C0812434;C0684335|armnull|Passive joint movement of neck (finding)|Finding|true|false|C0446516;C1140618;C1269078;C0027530;C3159206|neck
null|Neck problem|Finding|true|false|C0446516;C1140618;C1269078;C0027530;C3159206|necknull|dendritic spine neck|Anatomy|false|false|C0741025;C0812434;C0684335|neck
null|Neck|Anatomy|false|false|C0741025;C0812434;C0684335|necknull|Chest problem|Finding|true|false|C0027530;C3159206;C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0741025|chest
null|Anterior thoracic region|Anatomy|false|false|C0741025|chestnull|Discomfort|Finding|false|false||discomfortnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Study Object|Finding|false|false||studynull|Scientific Study|Procedure|false|false||study
null|Study|Procedure|false|false||study
null|Clinical Research|Procedure|false|false||studynull|Room of building - Study|Device|false|false||studynull|Uninterpretable|Modifier|false|false||uninterpretablenull|Ischemia|Finding|false|false||ischemianull|Ischemia Procedure|Procedure|false|false||ischemianull|contextual factors|Finding|false|false||settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|BaseLine dental cement|Drug|false|false||baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|Left Bundle-Branch Block|Disorder|false|false||LBBBnull|null|Lab|false|false||LBBBnull|Rhythm|Finding|false|false||rhythm
null|rhythmic process (biological)|Finding|false|false||rhythmnull|Sinus brand of acetaminophen-pseudoephedrine|Drug|false|false|C1305231;C0030471|sinus
null|Sinus brand of acetaminophen-pseudoephedrine|Drug|false|false|C1305231;C0030471|sinusnull|pathologic fistula|Disorder|false|false|C1305231;C0030471|sinusnull|Sinus - general anatomical term|Anatomy|false|false|C0723346;C0016169|sinus
null|Nasal sinus|Anatomy|false|false|C0723346;C0016169|sinusnull|Frequently|Time|false|false||frequentnull|Bed Status - Isolated|Finding|false|false||isolated
null|Isolated|Finding|false|false||isolatednull|Infrequent|Time|false|false||occasionalnull|Heart Atrium|Anatomy|false|false||atrialnull|Paired ventricular premature complexes|Finding|false|false||coupletsnull|Does run (finding)|Finding|false|false||run
null|Running (physical activity)|Finding|false|false||run
null|Go Jogging or Running Question|Finding|false|false||run
null|Run action|Finding|false|false||runnull|Rundi language|Entity|false|false||runnull|Paroxysmal supraventricular tachycardia|Disorder|false|false||PSVTnull|Paroxysmal Supraventricular Tachycardia by ECG Finding|Finding|false|false||PSVTnull|Retinoic Acid Response Element|Finding|false|false||Rarenull|Infrequent|Time|false|false||Rarenull|Rare|Modifier|false|false||Rarenull|Bed Status - Isolated|Finding|false|false||isolated
null|Isolated|Finding|false|false||isolatednull|Premature ventricular contractions|Disorder|false|false||vpbsnull|Rest|Finding|false|false||Restingnull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Systole|Finding|false|false||systolicnull|Hypertensive disease|Disorder|false|false||hypertensionnull|Increase|Finding|false|false||increasenull|Exercise|Finding|false|false||exercisenull|Exercise Pain Management|Procedure|false|false||exercisenull|Recovery - healing process|Finding|false|false||recoverynull|null|Event|false|false||recoverynull|recovery - adjustment|LabModifier|false|false||recoverynull|impression (attitude)|Finding|false|false||IMPRESSION
null|EKG impression|Finding|false|false||IMPRESSIONnull|Type - ParameterizedDataType|Finding|false|false||type
null|SGCG gene|Finding|false|false||typenull|null|Modifier|false|false||typenull|Symptoms aspect|Finding|true|false||symptoms
null|Symptoms|Finding|true|false||symptomsnull|Message Waiting Priority - High|Finding|false|false||high
null|high - ActExposureLevelCode|Finding|false|false||high
null|IPSS Risk Category High|Finding|false|false||high
null|IPSS-R Risk Category High|Finding|false|false||high
null|High (finding)|Finding|false|false||highnull|Observation Value - High|Modifier|false|false||high
null|High|Modifier|false|false||high
null|Abnormally high|Modifier|false|false||highnull|Cardiac attachment|Finding|false|false|C0018787|cardiacnull|Heart|Anatomy|false|false|C1314974|cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||cardiacnull|Economic demand|Finding|false|false||demandnull|Demand (clinical)|Procedure|false|false||demandnull|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group|Finding|false|false||poor
null|Patient Condition Code - Poor|Finding|false|false||poornull|Poverty|Subject|false|false||poornull|Language Proficiency - Poor|Modifier|false|false||poor
null|Specimen Quality - Poor|Modifier|false|false||poor
null|Poor - grade|Modifier|false|false||poor
null|Poor - qualifier|Modifier|false|false||poornull|Functional capacity|Finding|false|false||functional capacitynull|Functional Relationship|Finding|false|false||functional
null|Function (attribute)|Finding|false|false||functional
null|Functional|Finding|false|false||functionalnull|Capacity|LabModifier|false|false||capacitynull|Nuclear (incident type)|Modifier|false|false||Nuclear
null|Nuclear (nucleus)|Modifier|false|false||Nuclearnull|Report (document)|Finding|false|false||reportnull|Reporting|Procedure|false|false||reportnull|null|Attribute|false|false||reportnull|Catheterization|Procedure|false|false||CATHnull|levomefolate calcium|Drug|false|false||LMCA
null|levomefolate calcium|Drug|false|false||LMCA
null|levomefolate calcium|Drug|false|false||LMCAnull|Shortened|Modifier|false|false||shortnull|Short Value|LabModifier|false|false||short
null|Short|LabModifier|false|false||shortnull|DFFB protein, human|Drug|true|false||CAD
null|DFFB protein, human|Drug|true|false||CADnull|Cold Hemagglutinin Disease|Disorder|true|false||CAD
null|Coronary heart disease|Disorder|true|false||CAD
null|Coronary Artery Disease|Disorder|true|false||CADnull|CAD gene|Finding|true|false||CAD
null|CALD1 wt Allele|Finding|true|false||CAD
null|B4GALNT2 gene|Finding|true|false||CAD
null|DFFB wt Allele|Finding|true|false||CAD
null|ACOD1 gene|Finding|true|false||CAD
null|DFFB gene|Finding|true|false||CADnull|cytarabine/daunorubicin protocol|Procedure|true|false||CAD
null|Computer Assisted Diagnosis|Procedure|true|false||CAD
null|Collision-Induced Dissociation|Procedure|true|false||CAD
null|CyADIC regimen|Procedure|true|false||CADnull|Caddo language|Entity|true|false||CADnull|Leukocyte adhesion deficiency type 1|Disorder|false|false|C0226032|LAD
null|Leukocyte adhesion deficiency|Disorder|false|false|C0226032|LADnull|ITGB2 wt Allele|Finding|false|false|C0226032|LAD
null|DLD gene|Finding|false|false|C0226032|LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false|C5550999;C0398738;C1414063;C1706333|LADnull|Ladino Language|Entity|false|false||LADnull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Focal origin|Finding|false|false||focal originnull|Focal|Modifier|false|false||focalnull|Participation Type - origin|Finding|false|false||origin
null|National origin|Finding|false|false||originnull|Beginning|Time|false|false||originnull|Disease|Disorder|false|false||diseasenull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Proximal Resection Margin|Attribute|false|false||proximalnull|Proximal|Modifier|false|false||proximalnull|Disease|Disorder|false|false||diseasenull|Methylcytosine Dioxygenase TET1|Drug|false|false||LCX
null|Methylcytosine Dioxygenase TET1|Drug|false|false||LCXnull|TET1 wt Allele|Finding|false|false||LCX
null|TET1 gene|Finding|false|false||LCXnull|Minimal|Modifier|false|false||minimal
null|Mild (qualifier value)|Modifier|false|false||minimal
null|Minimum|Modifier|false|false||minimalnull|Luminal|Drug|false|false||luminal
null|Luminal|Drug|false|false||luminalnull|Luminal region|Modifier|false|false||luminalnull|Equine Gonadotropins|Drug|false|false||ECG
null|Equine Gonadotropins|Drug|false|false||ECG
null|Equine Gonadotropins|Drug|false|false||ECGnull|Electrocardiogram image|Finding|false|false||ECG
null|Electrocardiogram|Finding|false|false||ECGnull|Electrocardiography|Procedure|false|false||ECGnull|Sinus rhythm|Finding|false|false|C1305231;C0030471|sinus rhythm
null|null|Finding|false|false|C1305231;C0030471|sinus rhythmnull|Sinus brand of acetaminophen-pseudoephedrine|Drug|false|false|C1305231;C0030471|sinus
null|Sinus brand of acetaminophen-pseudoephedrine|Drug|false|false|C1305231;C0030471|sinusnull|pathologic fistula|Disorder|false|false|C1305231;C0030471|sinusnull|Sinus - general anatomical term|Anatomy|false|false|C2041122;C0232201;C0016169;C0723346;C1523018;C0871269|sinus
null|Nasal sinus|Anatomy|false|false|C2041122;C0232201;C0016169;C0723346;C1523018;C0871269|sinusnull|Rhythm|Finding|false|false|C1305231;C0030471|rhythm
null|rhythmic process (biological)|Finding|false|false|C1305231;C0030471|rhythmnull|Numerous|LabModifier|false|false||multiplenull|Atrial Premature Complexes|Disorder|false|false||PACsnull|Picture Archiving and Communication Systems|Finding|false|false||PACsnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Fracture of second cervical vertebra|Disorder|false|false|C0004457|axisnull|Axis vertebra|Anatomy|false|false|C0349013|axisnull|Genus Axis|Entity|false|false||axisnull|Axis|Modifier|false|false||axisnull|Protocol Deviation|Finding|false|false||deviationnull|Spatial Displacement|Modifier|false|false||deviation
null|Variant|Modifier|false|false||deviationnull|Old|Time|false|false||oldnull|Left Bundle-Branch Block|Disorder|false|false||LBBBnull|null|Lab|false|false||LBBBnull|Equine Gonadotropins|Drug|true|false||ECG
null|Equine Gonadotropins|Drug|true|false||ECG
null|Equine Gonadotropins|Drug|true|false||ECGnull|Electrocardiogram image|Finding|true|false||ECG
null|Electrocardiogram|Finding|true|false||ECGnull|Electrocardiography|Procedure|true|false||ECGnull|Probable diagnosis|Finding|false|false||Likely
null|Probably|Finding|false|false||Likelynull|Atrial tachycardia|Disorder|false|false|C0018792|atrial tachycardianull|continuous electrocardiogram atrial tachycardia|Finding|false|false|C0018792|atrial tachycardianull|Heart Atrium|Anatomy|false|false|C2059391;C0546959;C3827868;C0039231|atrialnull|Tachycardia by ECG Finding|Finding|false|false|C0018792|tachycardia
null|Tachycardia|Finding|false|false|C0018792|tachycardianull|Table Cell Horizontal Align - left|Finding|false|false||Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|Macromolecular Branch|Drug|false|false||branchnull|Branch of|Modifier|false|false||branchnull|Block Dosage Form|Drug|false|false||blocknull|Fixed Block|Finding|false|false||block
null|Obstruction|Finding|false|false||block
null|Blocking|Finding|false|false||blocknull|Geographic Block|Entity|false|false||blocknull|Block (unit of presentation)|LabModifier|false|false||block
null|Block Dosing Unit|LabModifier|false|false||block
null|Block (unit of measure)|LabModifier|false|false||blocknull|Act Relationship Subset - previous|Time|false|false||previous
null|Previous|Time|false|false||previousnull|Atrial tachycardia|Disorder|false|false|C0018792|atrial tachycardianull|continuous electrocardiogram atrial tachycardia|Finding|false|false|C0018792|atrial tachycardianull|Heart Atrium|Anatomy|false|false|C0546959;C2059391|atrialnull|Tachycardia by ECG Finding|Finding|false|false||tachycardia
null|Tachycardia|Finding|false|false||tachycardianull|Sinus rhythm|Finding|false|false|C1305231;C0030471|sinus rhythm
null|null|Finding|false|false|C1305231;C0030471|sinus rhythmnull|Sinus brand of acetaminophen-pseudoephedrine|Drug|false|false|C1305231;C0030471|sinus
null|Sinus brand of acetaminophen-pseudoephedrine|Drug|false|false|C1305231;C0030471|sinusnull|pathologic fistula|Disorder|false|false|C1305231;C0030471|sinusnull|Sinus - general anatomical term|Anatomy|false|false|C0016169;C2041122;C0232201;C1523018;C0871269;C0033036;C0723346|sinus
null|Nasal sinus|Anatomy|false|false|C0016169;C2041122;C0232201;C1523018;C0871269;C0033036;C0723346|sinusnull|Rhythm|Finding|false|false|C1305231;C0030471|rhythm
null|rhythmic process (biological)|Finding|false|false|C1305231;C0030471|rhythmnull|Atrial Premature Complexes|Disorder|false|false|C0018792;C1305231;C0030471|premature atrial contractionsnull|null|Attribute|false|false|C0018792|premature atrial contractionsnull|Premature Birth|Finding|false|false||premature
null|Too early|Finding|false|false||prematurenull|Immature|Modifier|false|false||prematurenull|Heart Atrium|Anatomy|false|false|C0033036;C0488348;C1140999|atrialnull|Contraction (finding)|Finding|false|false|C0018792|contractionsnull|Table Cell Horizontal Align - left|Finding|false|false||Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|Bundle-Branch Block|Disorder|false|false||bundle-branch blocknull|Macromolecular Branch|Drug|false|false||branchnull|Branch of|Modifier|false|false||branchnull|Block Dosage Form|Drug|false|false||blocknull|Fixed Block|Finding|false|false||block
null|Obstruction|Finding|false|false||block
null|Blocking|Finding|false|false||blocknull|Geographic Block|Entity|false|false||blocknull|Block (unit of presentation)|LabModifier|false|false||block
null|Block Dosing Unit|LabModifier|false|false||block
null|Block (unit of measure)|LabModifier|false|false||blocknull|ECHO protocol|Procedure|false|false||ECHO
null|Extension for Community Healthcare Outcomes|Procedure|false|false||ECHOnull|Echo <Calopterygidae>|Entity|false|false||ECHOnull|Conclusion|Finding|false|false||Conclusionsnull|Left atrial structure|Anatomy|false|false|C1552822|left atriumnull|Table Cell Horizontal Align - left|Finding|false|false|C0018792;C0225860|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Heart Atrium|Anatomy|false|false|C1552822|atriumnull|size|Modifier|false|false||sizenull|size - solid dosage form|LabModifier|false|false||sizenull|Atrial Septal Defects|Disorder|true|false|C0018792|atrial septal defectnull|Heart Atrium|Anatomy|false|false|C0018816;C5779791;C1457869;C0018817;C1861101|atrialnull|Congenital septal defect of heart|Disorder|true|false|C0018792|septal defect
null|Heart Septal Defects|Disorder|true|false|C0018792|septal defectnull|Septal|Modifier|false|false||septalnull|THYROID HORMONE PLASMA MEMBRANE TRANSPORT DEFECT|Disorder|true|false|C0018792|defectnull|Defect|Finding|true|false|C0018792|defectnull|Color doppler ultrasound|Procedure|false|false||color Dopplernull|color additive|Drug|false|false||color
null|Coloring Excipient|Drug|false|false||colornull|color - solid dosage form|Modifier|false|false||color
null|Color|Modifier|false|false||colornull|Color quantity|LabModifier|false|false||colornull|Doppler studies|Procedure|false|false||Dopplernull|Right atrial pressure|Attribute|false|false|C0018792|right atrial pressure
null|null|Attribute|false|false|C0018792|right atrial pressurenull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Atrial Pressure|Finding|false|false|C0018792|atrial pressurenull|Heart Atrium|Anatomy|false|false|C0460139;C1306345;C0234222;C0456165;C4050168;C0033095;C0428877|atrialnull|Pressure (finding)|Finding|false|false|C0018792|pressure
null|null|Finding|false|false|C0018792|pressure
null|Baresthesia|Finding|false|false|C0018792|pressurenull|null|Phenomenon|false|false|C0018792|pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|mmHg|LabModifier|false|false||mmHgnull|Wall of left ventricle|Anatomy|false|false|C2024242;C1552822;C1510420;C0011334|Left ventricular wallnull|Table Cell Horizontal Align - left|Finding|false|false|C0504053|Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|cardiac evaluation of ventricular wall thickness|Finding|false|false|C0018827;C0504053;C0507618|ventricular wall thicknessnull|Wall of ventricle|Anatomy|false|false|C2024242|ventricular wallnull|Heart Ventricle|Anatomy|false|false|C2024242|ventricularnull|Ventricular|Modifier|false|false||ventricularnull|Walls of a building|Device|false|false||wallnull|Thick|Modifier|false|false||thicknessnull|Dental caries|Disorder|false|false|C0504053;C0333343|cavity
null|Cavitation|Disorder|false|false|C0504053;C0333343|cavitynull|Body cavities|Anatomy|false|false|C1510420;C0011334|cavitynull|size|Modifier|false|false||sizenull|size - solid dosage form|LabModifier|false|false||sizenull|regional|Modifier|false|false||regional
null|Local|Modifier|false|false||regionalnull|Global|Modifier|false|false||global
null|Generalized|Modifier|false|false||globalnull|Systole|Finding|false|false||systolicnull|Function (attribute)|Finding|false|false||function
null|physiological aspects|Finding|false|false||function
null|Mathematical Operator|Finding|false|false||function
null|Functional Status|Finding|false|false||functionnull|Function Axis|Subject|false|false||functionnull|LVEF (procedure)|Procedure|false|false||LVEFnull|Left ventricular ejection fraction|Attribute|false|false||LVEFnull|Variability|Finding|false|false|C0018827|variabilitynull|Table Cell Horizontal Align - left|Finding|false|false|C0018827|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Heart Ventricle|Anatomy|false|false|C1552822;C2827666|ventricularnull|Ventricular|Modifier|false|false||ventricularnull|stress echo measurements ejection fraction|Finding|false|false||ejection fraction
null|Ejection fraction|Finding|false|false||ejection fractionnull|Ejection fraction (procedure)|Procedure|false|false||ejection fractionnull|Ejection as a Sports activity|Finding|false|false||ejectionnull|Ejection time|Attribute|false|false||ejectionnull|Ejection as a Circumstance of Injury|Phenomenon|false|false||ejectionnull|MDFAttributeType - Fraction|Finding|false|false||fractionnull|Fraction of|LabModifier|false|false||fractionnull|Irregular|Modifier|false|false||irregularnull|Rhythm|Finding|false|false||rhythm
null|rhythmic process (biological)|Finding|false|false||rhythmnull|Premature Cardiac Complex|Disorder|false|false||premature beatsnull|Premature Birth|Finding|false|false||premature
null|Too early|Finding|false|false||prematurenull|Immature|Modifier|false|false||prematurenull|Tissue Specimen Code|Finding|false|false|C0040300|Tissuenull|Body tissue|Anatomy|false|false|C0554756;C1547928;C0079595;C0011923;C0740845|Tissuenull|Doppler studies|Procedure|false|false|C0040300|Dopplernull|Imaging problem|Finding|false|false|C0040300|imagingnull|Diagnostic Imaging|Procedure|false|false|C0040300|imaging
null|Imaging Techniques|Procedure|false|false|C0040300|imagingnull|Imaging Technology|Title|false|false||imagingnull|Table Cell Horizontal Align - left|Finding|false|false|C0018827|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Heart Ventricle|Anatomy|false|false|C1552822|ventricularnull|Ventricular|Modifier|false|false||ventricularnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|Pulmonary Wedge Pressure|Attribute|false|false||PCWPnull|Table Cell Horizontal Align - right|Finding|false|false||Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|Heart Ventricle|Anatomy|false|false||ventricularnull|Ventricular|Modifier|false|false||ventricularnull|chamber [body part]|Anatomy|false|false||chambernull|Chamber (physical object)|Device|false|false||chambernull|size|Modifier|false|false||sizenull|size - solid dosage form|LabModifier|false|false||sizenull|Free of (attribute)|Finding|false|false||freenull|Empty (qualifier)|Modifier|false|false||freenull|Wall motion|Attribute|false|false||wall motionnull|Walls of a building|Device|false|false||wallnull|Motion|Phenomenon|false|false||motionnull|Aortic valve structure|Anatomy|false|false||aortic valve
null|Chest>Aortic valve|Anatomy|false|false||aortic valvenull|Aorta|Anatomy|false|false||aorticnull|Anatomical valve|Anatomy|false|false||valvenull|Valve (physical object)|Device|false|false||valve
null|Valve Device|Device|false|false||valve
null|medical valve|Device|false|false||valvenull|MILDLY|Modifier|false|false||mildly
null|Mild (qualifier value)|Modifier|false|false||mildlynull|AORTIC VALVE DISEASE 3|Disorder|true|false|C0003483;C1186983;C4533215;C0003501|aortic valve stenosis
null|Stenosis of aorta|Disorder|true|false|C0003483;C1186983;C4533215;C0003501|aortic valve stenosisnull|Aortic Valve Stenosis|Finding|true|false|C1186983;C4533215;C0003501;C0003483|aortic valve stenosisnull|Aortic valve structure|Anatomy|false|false|C0003507;C1261287;C5700069;C5193127|aortic valve
null|Chest>Aortic valve|Anatomy|false|false|C0003507;C1261287;C5700069;C5193127|aortic valvenull|Aorta|Anatomy|false|false|C5700069;C5193127;C0003507|aorticnull|Anatomical valve|Anatomy|false|false|C0003507;C5700069;C5193127|valvenull|Valve (physical object)|Device|false|false||valve
null|Valve Device|Device|false|false||valve
null|medical valve|Device|false|false||valvenull|Stenosis|Finding|true|false|C4533215;C0003501|stenosisnull|Stenosis <Pimeliinae>|Entity|true|false||stenosisnull|Stenosis Morphology|Modifier|false|false||stenosisnull|Aortic Valve Insufficiency|Disorder|false|false|C0003483|aortic regurgitationnull|Aorta|Anatomy|false|false|C0003504;C0232605;C2004489|aorticnull|Regurgitation|Finding|false|false|C0003483|regurgitation
null|Regurgitates after swallowing|Finding|false|false|C0003483|regurgitationnull|Regurgitation - mechanism|Phenomenon|false|false||regurgitationnull|Mitral Valve|Anatomy|false|false||mitral valvenull|mitral|Modifier|false|false||mitralnull|Anatomical valve|Anatomy|false|false||valvenull|Valve (physical object)|Device|false|false||valve
null|Valve Device|Device|false|false||valve
null|medical valve|Device|false|false||valvenull|MILDLY|Modifier|false|false||mildly
null|Mild (qualifier value)|Modifier|false|false||mildlynull|Mitral Valve Prolapse Syndrome|Disorder|true|false|C0026264;C1186983|mitral valve prolapsenull|Mitral Valve|Anatomy|false|false|C0026267;C0033377|mitral valvenull|mitral|Modifier|false|false||mitralnull|Anatomical valve|Anatomy|false|false|C0026267;C0033377|valvenull|Valve (physical object)|Device|false|false||valve
null|Valve Device|Device|false|false||valve
null|medical valve|Device|false|false||valvenull|Ptosis|Disorder|true|false|C1186983;C0026264|prolapsenull|Physiological|Finding|false|false||Physiologicnull|Mitral Valve Insufficiency|Disorder|false|false||mitral regurgitationnull|mitral|Modifier|false|false||mitralnull|Regurgitation|Finding|false|false||regurgitation
null|Regurgitates after swallowing|Finding|false|false||regurgitationnull|Regurgitation - mechanism|Phenomenon|false|false||regurgitationnull|null|Finding|false|false||within normal limitsnull|Limited (extensiveness)|Finding|false|false||limitsnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Heart Ventricle|Anatomy|false|false||ventricularnull|Ventricular|Modifier|false|false||ventricularnull|Patterns|Modifier|false|false||patternnull|Relaxation|Event|false|false||relaxationnull|Pulmonary artery systolic pressure|Finding|false|false|C0034052;C0226004;C0003842;C0024109|pulmonary artery systolic pressurenull|Pulmonary artery structure|Anatomy|false|false|C0039155;C0460139;C1306345;C0234222;C0428643;C4522268;C0871470;C0033095|pulmonary arterynull|Pulmonary (intended site)|Finding|false|false|C0034052;C0226004;C0003842;C0024109|pulmonarynull|Lung|Anatomy|false|false|C4522268;C0428643;C2707265|pulmonarynull|null|Attribute|false|false|C0024109|pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Arterial system|Anatomy|false|false|C0428643;C4522268;C0033095;C0039155;C0460139;C1306345;C0234222|artery
null|Arteries|Anatomy|false|false|C0428643;C4522268;C0033095;C0039155;C0460139;C1306345;C0234222|arterynull|Systolic Pressure|Attribute|false|false|C0034052|systolic pressurenull|Systole|Finding|false|false|C0034052;C0226004;C0003842|systolicnull|Pressure (finding)|Finding|false|false|C0034052;C0226004;C0003842|pressure
null|null|Finding|false|false|C0034052;C0226004;C0003842|pressure
null|Baresthesia|Finding|false|false|C0034052;C0226004;C0003842|pressurenull|null|Phenomenon|false|false|C0226004;C0003842;C0034052|pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|Pericardial effusion|Disorder|true|false|C0031050;C0442031|pericardial effusionnull|Pericardial effusion body substance|Finding|true|false|C0031050;C0442031|pericardial effusionnull|Pericardial (qualifier value)|Anatomy|false|false|C1253937;C0031039;C2317432;C1546613;C0013687|pericardial
null|Pericardial sac structure|Anatomy|false|false|C1253937;C0031039;C2317432;C1546613;C0013687|pericardialnull|Effusion (substance)|Finding|true|false|C0031050;C0442031|effusion
null|null|Finding|true|false|C0031050;C0442031|effusion
null|effusion|Finding|true|false|C0031050;C0442031|effusionnull|null|Time|false|false||priornull|Study Object|Finding|false|false||studynull|Scientific Study|Procedure|false|false||study
null|Study|Procedure|false|false||study
null|Clinical Research|Procedure|false|false||studynull|Room of building - Study|Device|false|false||studynull|Frequently|Time|false|false||frequentnull|Atrial arrhythmia|Finding|false|false|C0018792|atrial ectopynull|Heart Atrium|Anatomy|false|false|C0085611|atrialnull|biventricular|Modifier|false|false||biventricularnull|Function (attribute)|Finding|false|false||function
null|physiological aspects|Finding|false|false||function
null|Mathematical Operator|Finding|false|false||function
null|Functional Status|Finding|false|false||functionnull|Function Axis|Subject|false|false||functionnull|Similarity|Modifier|false|false||similarnull|Micro (prefix)|Finding|false|false||Micro
null|Microbiology - Laboratory Class|Finding|false|false||Micronull|Microbiology procedure|Procedure|false|false||Micronull|Unit Of Measure Prefix - micro|LabModifier|false|false||Micronull|Pending - Allergy Clinical Status|Finding|false|false||pending
null|Pending - referral status|Finding|false|false||pendingnull|Pending - status|Time|false|false||pendingnull|pending - ManagedParticipationStatus|Modifier|false|false||pending
null|pending - RoleStatus|Modifier|false|false||pending
null|Pending - Day type|Modifier|false|false||pendingnull|PMH - past medical history|Finding|false|false||PMH
null|Medical History|Finding|false|false||PMHnull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Peripheral Vascular Diseases|Disorder|false|false||PVDnull|Pomalidomide/Bortezomib/Dexamethasone Regimen|Procedure|false|false||PVDnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|Recurrent|Time|false|false||recurrent
null|Episodic|Time|false|false||recurrentnull|Retrosternal pain|Finding|false|false|C1527391;C0817096|substernal chest painnull|Chest Pain|Finding|false|false|C1527391;C0817096|chest painnull|null|Attribute|false|false|C1527391;C0817096|chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0741025;C1549543;C0030193;C0151826;C0008031;C2926613|chest
null|Anterior thoracic region|Anatomy|false|false|C0741025;C1549543;C0030193;C0151826;C0008031;C2926613|chestnull|Administration Method - Pain|Finding|false|false|C1527391;C0817096|pain
null|Pain|Finding|false|false|C1527391;C0817096|painnull|null|Attribute|false|false||painnull|Has patient|Finding|false|false||patient hasnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Laboratory test finding|Lab|false|false||labsnull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|Negative|Finding|false|false||for negativenull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Troponin|Drug|false|false||troponins
null|Troponin|Drug|false|false||troponinsnull|Electrocardiogram image|Finding|false|false||EKG
null|Electrocardiogram|Finding|false|false||EKGnull|Electrocardiography|Procedure|false|false||EKGnull|Ischemic|Finding|false|false||ischemicnull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Numerous|LabModifier|false|false||multiplenull|Episode of|Time|false|false||episodesnull|Atrial tachycardia|Disorder|false|false|C0018792|atrial tachycardianull|continuous electrocardiogram atrial tachycardia|Finding|false|false|C0018792|atrial tachycardianull|Heart Atrium|Anatomy|false|false|C0546959;C2059391;C0004238;C3827868;C0039231|atrialnull|Tachycardia by ECG Finding|Finding|false|false|C0018792|tachycardia
null|Tachycardia|Finding|false|false|C0018792|tachycardianull|Atrial Fibrillation|Disorder|false|false|C0018792|AFibnull|Atrial Fibrillation by ECG Finding|Lab|false|false||AFibnull|amiodarone|Drug|false|false||Amiodarone
null|amiodarone|Drug|false|false||Amiodaronenull|Drug assay amiodarone|Procedure|false|false||Amiodaronenull|Amount type - Rate|Finding|false|false||ratenull|Rating (action)|Event|false|false||ratenull|Rate|LabModifier|false|false||ratenull|Rhythm|Finding|false|false||rhythm
null|rhythmic process (biological)|Finding|false|false||rhythmnull|Control brand of phenylpropanolamine|Drug|false|false||control
null|CONTROL veterinary product|Drug|false|false||control
null|control substance|Drug|false|false||control
null|Control brand of phenylpropanolamine|Drug|false|false||controlnull|Control - Relationship modifier|Finding|false|false||control
null|Control function|Finding|false|false||control
null|Scientific Control|Finding|false|false||controlnull|Control Groups|Subject|false|false||controlnull|True Control Status|Modifier|false|false||control
null|control aspects|Modifier|false|false||controlnull|rivaroxaban|Drug|false|false||Rivaroxaban
null|rivaroxaban|Drug|false|false||Rivaroxabannull|ANTICOAGULATION (finding)|Finding|false|false||anticoagulation
null|Anticoagulation function|Finding|false|false||anticoagulation
null|Decreased Coagulation Activity [PE]|Finding|false|false||anticoagulationnull|Anticoagulation Therapy|Procedure|false|false||anticoagulationnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|diltiazem|Drug|false|false||Diltiazem
null|diltiazem|Drug|false|false||Diltiazemnull|rate control|Finding|false|false||rate controlnull|Amount type - Rate|Finding|false|false||ratenull|Rating (action)|Event|false|false||ratenull|Rate|LabModifier|false|false||ratenull|Control brand of phenylpropanolamine|Drug|false|false||control
null|CONTROL veterinary product|Drug|false|false||control
null|control substance|Drug|false|false||control
null|Control brand of phenylpropanolamine|Drug|false|false||controlnull|Control - Relationship modifier|Finding|false|false||control
null|Control function|Finding|false|false||control
null|Scientific Control|Finding|false|false||controlnull|Control Groups|Subject|false|false||controlnull|True Control Status|Modifier|false|false||control
null|control aspects|Modifier|false|false||controlnull|Episode of|Time|false|false||episodesnull|Chest Pain|Finding|false|false|C1527391;C0817096|chest painnull|null|Attribute|false|false|C1527391;C0817096|chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C2926613;C1549543;C0030193;C0008031;C0741025|chest
null|Anterior thoracic region|Anatomy|false|false|C2926613;C1549543;C0030193;C0008031;C0741025|chestnull|Administration Method - Pain|Finding|false|false|C1527391;C0817096|pain
null|Pain|Finding|false|false|C1527391;C0817096|painnull|null|Attribute|false|false||painnull|during hospitalization|Time|false|false||during hospitalizationnull|Hospitalization|Procedure|false|false||hospitalizationnull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Atrial fibrillation and flutter|Finding|false|false|C0018792|atrial fibrillation/flutternull|Atrial Fibrillation|Disorder|false|false|C0018792|atrial fibrillationnull|null|Attribute|false|false|C0018792|atrial fibrillationnull|Atrial Fibrillation by ECG Finding|Lab|false|false|C0018792|atrial fibrillationnull|Heart Atrium|Anatomy|false|false|C0016385;C0232197;C2926591;C0155709;C0344434;C0004238|atrialnull|Fibrillation|Disorder|false|false|C0018792|fibrillationnull|Cardiac Flutter|Finding|false|false|C0018792|flutternull|Flutter (respiratory device)|Device|false|false||flutternull|Primary care provider|Subject|false|false||primary care doctornull|Location Service Code - Primary Care|Finding|false|false||primary carenull|Primary Health Care|Procedure|false|false||primary carenull|True primary (qualifier value)|Time|false|false||primarynull|Primary|Modifier|false|false||primarynull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Doctor - Title|Finding|false|false||doctornull|Physicians|Subject|false|false||doctornull|Vague|Modifier|false|false||vaguenull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0741025|chest
null|Anterior thoracic region|Anatomy|false|false|C0741025|chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Admission Level of Care Code - Acute|Finding|false|false||Acute
null|Acute - Triage Code|Finding|false|false||Acutenull|acute|Time|false|false||Acutenull|Atrial tachycardia|Disorder|false|false|C0018792|Atrial Tachycardianull|continuous electrocardiogram atrial tachycardia|Finding|false|false|C0018792|Atrial Tachycardianull|Heart Atrium|Anatomy|false|false|C0546959;C2059391;C3827868;C0039231|Atrialnull|Tachycardia by ECG Finding|Finding|false|false|C0018792|Tachycardia
null|Tachycardia|Finding|false|false|C0018792|Tachycardianull|During admission|Time|false|false||During admissionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Does run (finding)|Finding|false|false||runsnull|Widening|Modifier|false|false||widenull|complex (molecular entity)|Drug|false|false||complexnull|Complex|Modifier|false|false||complexnull|Thought|Finding|false|false||thought
null|null|Finding|false|false||thoughtnull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Participation Type - origin|Finding|false|false||origin
null|National origin|Finding|false|false||originnull|Beginning|Time|false|false||originnull|Rapid atrial fibrillation|Disorder|false|false|C0018792|rapid Atrial Fibrillationnull|Rapid|Modifier|false|false||rapidnull|Atrial fibrillation and flutter|Finding|false|false|C0018792|Atrial Fibrillation/ Flutternull|Atrial Fibrillation|Disorder|false|false|C0018792|Atrial Fibrillationnull|null|Attribute|false|false|C0018792|Atrial Fibrillationnull|Atrial Fibrillation by ECG Finding|Lab|false|false|C0018792|Atrial Fibrillationnull|Heart Atrium|Anatomy|false|false|C0155709;C2926591;C0016385;C0004238;C1281999;C0344434;C0232197|Atrialnull|Fibrillation|Disorder|false|false|C0018792|Fibrillationnull|Cardiac Flutter|Finding|false|false|C0018792|Flutternull|Flutter (respiratory device)|Device|false|false||Flutternull|Heart Atrium|Anatomy|false|false||atrialnull|Tachycardia by ECG Finding|Finding|false|false||tachycardia
null|Tachycardia|Finding|false|false||tachycardianull|complex (molecular entity)|Drug|false|false||complexesnull|Similarity|Modifier|false|false||similarnull|Physical shape|Finding|false|false||morphologynull|Science of Morphology|Title|false|false||morphologynull|Morphology (property)|Modifier|false|false||morphology
null|Morphology|Modifier|false|false||morphology
null|morphological|Modifier|false|false||morphologynull|Kind of quantity - Morphology|LabModifier|false|false||morphologynull|Native (qualifier value)|Finding|false|false||nativenull|Left Bundle-Branch Block|Disorder|false|false||LBBBnull|null|Lab|false|false||LBBBnull|diltiazem|Drug|false|false||Diltiazem
null|diltiazem|Drug|false|false||Diltiazemnull|amiodarone|Drug|false|false||Amiodarone
null|amiodarone|Drug|false|false||Amiodaronenull|Drug assay amiodarone|Procedure|false|false||Amiodaronenull|Episode of|Time|false|false||episodesnull|Tachycardia by ECG Finding|Finding|false|false||tachycardia
null|Tachycardia|Finding|false|false||tachycardianull|Team|Subject|false|false||teamnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|ANTICOAGULATION (finding)|Finding|false|false||anticoagulation
null|Anticoagulation function|Finding|false|false||anticoagulation
null|Decreased Coagulation Activity [PE]|Finding|false|false||anticoagulationnull|Anticoagulation Therapy|Procedure|false|false||anticoagulationnull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|Follow-up status|Finding|false|false||follow upnull|follow-up|Procedure|false|false||follow upnull|Follow - dosing instruction imperative|Finding|false|false||follow
null|Follow|Finding|false|false||follownull|Followed by|Time|false|false||follownull|Cardiac electrophysiology study|Procedure|false|false||EP studynull|Study Object|Finding|false|false||studynull|Scientific Study|Procedure|false|false||study
null|Study|Procedure|false|false||study
null|Clinical Research|Procedure|false|false||studynull|Room of building - Study|Device|false|false||studynull|Possible|Finding|false|false||possiblenull|Possible diagnosis|Modifier|false|false||possible
null|Possibly Related to Intervention|Modifier|false|false||possiblenull|Ablation|Procedure|false|false|C0018792|ablation
null|Destructive procedure (surgical)|Procedure|false|false|C0018792|ablationnull|Atrial Flutter|Finding|false|false|C0018792|Atrial Flutternull|Atrial Flutter by ECG Finding|Lab|false|false|C0018792|Atrial Flutternull|Heart Atrium|Anatomy|false|false|C0016385;C0344423;C0004239;C0547070;C1261381|Atrialnull|Cardiac Flutter|Finding|false|false|C0018792|Flutternull|Flutter (respiratory device)|Device|false|false||Flutternull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Heart|Anatomy|false|false||Heartsnull|Monitor brand of insecticide|Drug|false|false||monitor
null|Monitor brand of insecticide|Drug|false|false||monitornull|Monitor Device|Device|false|false||monitor
null|Monitoring Device|Device|false|false||monitornull|Monitor, occupation|Subject|false|false||monitornull|amiodarone|Drug|false|false||Amiodarone
null|amiodarone|Drug|false|false||Amiodaronenull|Drug assay amiodarone|Procedure|false|false||Amiodaronenull|Twice a day|Time|false|false||twice dailynull|Daily|Time|false|false||dailynull|1 Week|Time|false|false||1 weeknull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|Daily|Time|false|false||dailynull|diltiazem|Drug|false|false||Diltiazem
null|diltiazem|Drug|false|false||Diltiazemnull|At home|Finding|false|false||at homenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|rivaroxaban|Drug|false|false||Rivaroxaban
null|rivaroxaban|Drug|false|false||Rivaroxabannull|ANTICOAGULATION (finding)|Finding|false|false||anticoagulation
null|Anticoagulation function|Finding|false|false||anticoagulation
null|Decreased Coagulation Activity [PE]|Finding|false|false||anticoagulationnull|Anticoagulation Therapy|Procedure|false|false||anticoagulationnull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|Cardiologists|Subject|false|false||cardiologistnull|Plavix|Drug|false|false||plavix
null|Plavix|Drug|false|false||plavixnull|TNFSF14 protein, human|Drug|false|false||light
null|TNFSF14 protein, human|Drug|false|false||lightnull|Light - subjective measurement|Finding|false|false||light
null|TNFSF14 wt Allele|Finding|false|false||light
null|TNFSF14 gene|Finding|false|false||light
null|Light color|Finding|false|false||lightnull|Phototherapy|Procedure|false|false||lightnull|Light|Phenomenon|false|false||lightnull|Light (qualifier)|Modifier|false|false||lightnull|In addition to|Finding|false|false||addition
null|Add - instruction imperative|Finding|false|false||additionnull|rivaroxaban|Drug|false|false||Rivaroxaban
null|rivaroxaban|Drug|false|false||Rivaroxabannull|Interested|Finding|false|false||interestnull|Triplicate|LabModifier|false|false||triplenull|Therapy Object (animal model)|Finding|false|false||therapy
null|therapeutic aspects|Finding|false|false||therapynull|Therapeutic procedure|Procedure|false|false||therapynull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Appointments|Event|false|false||appointmentsnull|Processing type - Evaluation|Finding|false|false||evaluationnull|Evaluation procedure|Procedure|false|false||evaluation
null|Evaluation|Procedure|false|false||evaluationnull|2 Months|Time|false|false||2 monthsnull|month|Time|false|false||monthsnull|Chest Pain|Finding|false|false|C1527391;C0817096|Chest painnull|null|Attribute|false|false|C1527391;C0817096|Chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|Chestnull|Chest|Anatomy|false|false|C0008031;C0741025;C1549543;C0030193;C2926613|Chest
null|Anterior thoracic region|Anatomy|false|false|C0008031;C0741025;C1549543;C0030193;C2926613|Chestnull|Administration Method - Pain|Finding|false|false|C1527391;C0817096|pain
null|Pain|Finding|false|false|C1527391;C0817096|painnull|null|Attribute|false|false||painnull|Retrosternal pain|Finding|false|false|C1527391;C0817096|substernal chest painnull|Chest Pain|Finding|false|false|C1527391;C0817096|chest painnull|null|Attribute|false|false||chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0741025;C0008031;C0151826|chest
null|Anterior thoracic region|Anatomy|false|false|C0741025;C0008031;C0151826|chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|At rest (qualifier value)|Finding|false|false||at restnull|REST protein, human|Drug|false|false||rest
null|REST protein, human|Drug|false|false||restnull|REST gene|Finding|false|false||rest
null|site-specific telomere resolvase activity|Finding|false|false||rest
null|Rest|Finding|false|false||restnull|Troponin|Drug|true|false||troponin
null|Troponin|Drug|true|false||troponinnull|Troponin measurement|Procedure|true|false||troponinnull|Elevation procedure|Procedure|false|false||elevationnull|Elevation|Modifier|false|false||elevationnull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|Equine Gonadotropins|Drug|false|false||ECG
null|Equine Gonadotropins|Drug|false|false||ECG
null|Equine Gonadotropins|Drug|false|false||ECGnull|Electrocardiogram image|Finding|false|false||ECG
null|Electrocardiogram|Finding|false|false||ECGnull|Electrocardiography|Procedure|false|false||ECGnull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|Chest Pain|Finding|false|false|C1527391;C0817096|chest painnull|null|Attribute|false|false|C1527391;C0817096|chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0741025;C0008031;C2926613|chest
null|Anterior thoracic region|Anatomy|false|false|C0741025;C0008031;C2926613|chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Menstruation|Finding|false|false||periodsnull|Tachycardia by ECG Finding|Finding|false|false||tachycardia
null|Tachycardia|Finding|false|false||tachycardianull|Organization unit type - Hospital|Finding|false|false|C0018792;C1527391;C0817096|hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Diarrhea|Finding|false|false||the runsnull|Does run (finding)|Finding|false|false|C0018792|runsnull|Atrial tachycardia|Disorder|false|false|C0018792|atrial tachycardianull|continuous electrocardiogram atrial tachycardia|Finding|false|false|C0018792|atrial tachycardianull|Heart Atrium|Anatomy|false|false|C1547192;C0546959;C2059391;C3827868;C0039231;C0600140|atrialnull|Tachycardia by ECG Finding|Finding|false|false|C0018792|tachycardia
null|Tachycardia|Finding|false|false|C0018792|tachycardianull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C1547192;C0741025|chest
null|Anterior thoracic region|Anatomy|false|false|C1547192;C0741025|chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Episode of|Time|false|false||episodesnull|Chest Pain|Finding|false|false|C1527391;C0817096|chest painnull|null|Attribute|false|false|C1527391;C0817096|chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0741025;C2926613;C0008031|chest
null|Anterior thoracic region|Anatomy|false|false|C0741025;C2926613;C0008031|chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Hospitalization|Procedure|false|false||hospitalizationnull|Heart Atrium|Anatomy|false|false||atrialnull|Fibrillation|Disorder|false|false||fibrillationnull|Cardiac Flutter|Finding|false|false||flutternull|Flutter (respiratory device)|Device|false|false||flutternull|Primary care provider|Subject|false|false||primary care doctornull|Location Service Code - Primary Care|Finding|false|false||primary carenull|Primary Health Care|Procedure|false|false||primary carenull|True primary (qualifier value)|Time|false|false||primarynull|Primary|Modifier|false|false||primarynull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Doctor - Title|Finding|false|false||doctornull|Physicians|Subject|false|false||doctornull|Vague|Modifier|false|false||vaguenull|Chest Pain|Finding|false|false|C1527391;C0817096|chest painnull|null|Attribute|false|false|C1527391;C0817096|chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0741025;C2926613;C0008031|chest
null|Anterior thoracic region|Anatomy|false|false|C0741025;C2926613;C0008031|chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Dry Eyes brand of ocular lubricant|Drug|false|false|C0015392|Dry eyesnull|Dry Eye Syndromes|Disorder|false|false|C0015392|Dry eyes
null|Keratoconjunctivitis Sicca|Disorder|false|false|C0015392|Dry eyesnull|Dryness of eye|Finding|false|false|C0015392|Dry eyesnull|Eye|Anatomy|false|false|C0720056;C0022575;C0013238;C0314719;C5848506|eyesnull|null|Attribute|false|false|C0015392|eyesnull|Erythema|Disorder|false|false|C4266572;C0015392;C0700042|erythemanull|Administration Method - Pain|Finding|false|false|C4266572;C0015392;C0700042|pain
null|Pain|Finding|false|false|C4266572;C0015392;C0700042|painnull|null|Attribute|false|false||painnull|null|Attribute|false|false|C4266572;C0015392;C0700042|R eyenull|Carcinoma in situ of eye|Disorder|false|false|C4266572;C0015392;C0700042|eye
null|Disorder of eye|Disorder|false|false|C4266572;C0015392;C0700042|eyenull|Eye - Specimen Source Code|Finding|false|false|C4266572;C0015392;C0700042|eye
null|Eye problem|Finding|false|false|C4266572;C0015392;C0700042|eye
null|Eye Specimen|Finding|false|false|C4266572;C0015392;C0700042|eyenull|Head>Eye|Anatomy|false|false|C0041834;C1549543;C0030193;C0154094;C0015397;C1550636;C1546630;C0262477;C5886197|eye
null|Eye|Anatomy|false|false|C0041834;C1549543;C0030193;C0154094;C0015397;C1550636;C1546630;C0262477;C5886197|eye
null|Orbital region|Anatomy|false|false|C0041834;C1549543;C0030193;C0154094;C0015397;C1550636;C1546630;C0262477;C5886197|eyenull|Eye|Anatomy|false|false|C5848506|eyesnull|null|Attribute|false|false|C0015392|eyesnull|artificial tears (medication)|Drug|false|false||Artificial tears
null|Lubricant Eye Drops|Drug|false|false||Artificial tears
null|Artificial Tears|Drug|false|false||Artificial tearsnull|Artificial (qualifier value)|Modifier|false|false||Artificialnull|Tears (substance)|Finding|false|false||tears
null|null|Finding|false|false||tears
null|Tears specimen|Finding|false|false||tearsnull|erythromycin|Drug|false|false|C4266572;C0015392;C0700042|erythromycin
null|erythromycin|Drug|false|false|C4266572;C0015392;C0700042|erythromycinnull|Eye drops brand of Tetrahydrozoline|Drug|false|false|C4266572;C0015392;C0700042|eye drops
null|Eye Drops|Drug|false|false|C4266572;C0015392;C0700042|eye drops
null|Eye drops brand of Tetrahydrozoline|Drug|false|false|C4266572;C0015392;C0700042|eye dropsnull|Carcinoma in situ of eye|Disorder|false|false|C4266572;C0015392;C0700042|eye
null|Disorder of eye|Disorder|false|false|C4266572;C0015392;C0700042|eyenull|Eye - Specimen Source Code|Finding|false|false|C4266572;C0015392;C0700042|eye
null|Eye problem|Finding|false|false|C4266572;C0015392;C0700042|eye
null|Eye Specimen|Finding|false|false|C4266572;C0015392;C0700042|eyenull|Head>Eye|Anatomy|false|false|C0015399;C1154269;C1550636;C1546630;C0262477;C0154094;C0015397;C0014806|eye
null|Eye|Anatomy|false|false|C0015399;C1154269;C1550636;C1546630;C0262477;C0154094;C0015397;C0014806|eye
null|Orbital region|Anatomy|false|false|C0015399;C1154269;C1550636;C1546630;C0262477;C0154094;C0015397;C0014806|eyenull|Drops - Drug Form|Drug|false|false||dropsnull|Drop Dosing Unit|LabModifier|false|false||dropsnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Appointments|Event|false|false||appointmentnull|Attending (action)|Finding|false|false||attendnull|Appointments|Event|false|false||appointmentnull|Chronic - Admission Level of Care Code|Finding|false|false||Chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||Chronicnull|chronic|Time|false|false||Chronicnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|BaseLine dental cement|Drug|false|false||baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|Respiratory Status|Finding|false|false||respiratory statusnull|null|Attribute|false|false||respiratory statusnull|Respiratory attachment|Finding|false|false||respiratory
null|respiratory|Finding|false|false||respiratory
null|null|Finding|false|false||respiratory
null|Respiratory specimen|Finding|false|false||respiratorynull|Respiratory rate|Attribute|false|false||respiratorynull|What subject filter - Status|Finding|false|false||statusnull|null|Attribute|false|false||statusnull|Social status|Modifier|false|false||status
null|Status|Modifier|false|false||statusnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|albuterol|Drug|false|false||albuterol
null|albuterol|Drug|false|false||albuterolnull|NEB protein, human|Drug|false|false||neb
null|NEB protein, human|Drug|false|false||neb
null|Nebulizer solution|Drug|false|false||nebnull|NEB gene|Finding|false|false||neb
null|mitotic nuclear membrane disassembly|Finding|false|false||nebnull|albuterol|Drug|false|false||albuterol
null|albuterol|Drug|false|false||albuterolnull|Inhaler (unit of presentation)|Finding|false|false||inhalernull|Inhaler|Device|false|false||inhalernull|Inhaler Dosing Unit|LabModifier|false|false||inhalernull|null|Drug|false|false|C0028429|Fluticasone nasalnull|fluticasone|Drug|false|false||Fluticasone
null|fluticasone|Drug|false|false||Fluticasonenull|Nasal Spray brand of phenylephrine|Drug|false|false|C0028429|nasal spraynull|Nasal spray (device)|Device|false|false||nasal spray
null|Nasal Sprays|Device|false|false||nasal spray
null|Nasal Spray|Device|false|false||nasal spraynull|Nasal brand of oxymetazoline|Drug|false|false|C0028429|nasal
null|Nasal brand of oxymetazoline|Drug|false|false|C0028429|nasal
null|Nasal dosage form|Drug|false|false|C0028429|nasalnull|Nasal Route of Administration|Finding|false|false|C0028429|nasal
null|Nasal (intended site)|Finding|false|false|C0028429|nasalnull|null|Anatomy|false|false|C4520890;C1522019;C1272939;C0721966;C0360577;C4521772;C2608294;C2003858|nasalnull|Spray Dosage Form|Drug|false|false||spraynull|Spray (administration method)|Finding|false|false|C0028429|spraynull|Spray (action)|Event|false|false|C0028429|spraynull|Spray Dosing Unit|LabModifier|false|false||spraynull|Fluticasone-Salmeterol Diskus|Drug|false|false||fluticasone-salmeterol diskus
null|Fluticasone-Salmeterol Diskus|Drug|false|false||fluticasone-salmeterol diskusnull|fluticasone / salmeterol|Drug|false|false||fluticasone-salmeterolnull|fluticasone|Drug|false|false||fluticasone
null|fluticasone|Drug|false|false||fluticasonenull|salmeterol|Drug|false|false||salmeterol
null|salmeterol|Drug|false|false||salmeterolnull|Diskus|Device|false|false||diskusnull|tiotropium bromide|Drug|false|false||tiotropium bromide
null|tiotropium bromide|Drug|false|false||tiotropium bromidenull|tiotropium|Drug|false|false||tiotropium
null|tiotropium|Drug|false|false||tiotropiumnull|Bromides|Drug|false|false||bromidenull|Bromides measurement|Procedure|false|false||bromidenull|Nebulizer solution|Drug|false|false||nebsnull|theophylline|Drug|false|false||theophylline
null|theophylline|Drug|false|false||theophyllinenull|Assay of theophylline|Procedure|false|false||theophyllinenull|Pad Dosage Form|Drug|false|false|C3669270|PADnull|Pad Mass|Disorder|false|false|C3669270|PAD
null|Peripheral Arterial Diseases|Disorder|false|false|C3669270|PADnull|PADI4 wt Allele|Finding|false|false|C3669270|PAD
null|PADI4 gene|Finding|false|false|C3669270|PAD
null|DHX40 gene|Finding|false|false|C3669270|PADnull|PAD Regimen|Procedure|false|false|C3669270|PADnull|Strucure of thick cushion of skin|Anatomy|false|false|C3814046;C2347441;C3540603;C1425478;C1425244;C0332568;C1704436|PADnull|Pad Device|Device|false|false||PAD
null|Pads|Device|false|false||PADnull|Pad (unit of presentation)|LabModifier|false|false||PAD
null|Pad Dosing Unit|LabModifier|false|false||PADnull|Table Frame - above|Finding|false|false||abovenull|Upper|Modifier|false|false||abovenull|clopidogrel|Drug|false|false||Clopidogrel
null|clopidogrel|Drug|false|false||Clopidogrelnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|rivaroxaban|Drug|false|false||Rivaroxaban
null|rivaroxaban|Drug|false|false||Rivaroxabannull|Triplicate|LabModifier|false|false||triplenull|Therapy Object (animal model)|Finding|false|false||therapy
null|therapeutic aspects|Finding|false|false||therapynull|Therapeutic procedure|Procedure|false|false||therapynull|Cardiologists|Subject|false|false||cardiologistnull|Marketing basis - Transitional|Finding|false|false||Transitionalnull|Transitional cell morphology|Modifier|false|false||Transitionalnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|amiodarone|Drug|false|false||Amiodarone
null|amiodarone|Drug|false|false||Amiodaronenull|Drug assay amiodarone|Procedure|false|false||Amiodaronenull|Twice a day|Time|false|false||twice dailynull|Daily|Time|false|false||dailynull|1 Week|Time|false|false||one weeknull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|Daily|Time|false|false||dailynull|Appointments|Event|false|false||appointmentnull|Approximate|Modifier|false|false||approximatelynull|2 Months|Time|false|false||2 monthsnull|month|Time|false|false||monthsnull|rivaroxaban|Drug|false|false||Rivaroxaban
null|rivaroxaban|Drug|false|false||Rivaroxabannull|QPM|Time|false|false||qpm
null|Once a day, in the evening|Time|false|false||qpmnull|With dinner|Time|false|false||with dinnernull|Dinner|Finding|false|false||dinnernull|With dinner|Time|false|false||dinnernull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|Heart|Anatomy|false|false||Heartsnull|Monitor brand of insecticide|Drug|false|false||monitor
null|Monitor brand of insecticide|Drug|false|false||monitornull|Monitor Device|Device|false|false||monitor
null|Monitoring Device|Device|false|false||monitornull|Monitor, occupation|Subject|false|false||monitornull|Cardiologists|Subject|false|false||Cardiologistnull|Chest Pain|Finding|false|false|C1527391;C0817096|chest painnull|null|Attribute|false|false|C1527391;C0817096|chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0008031;C2926613;C0741025|chest
null|Anterior thoracic region|Anatomy|false|false|C0008031;C2926613;C0741025|chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Biological Markers|Attribute|false|false||biomarkersnull|Electrocardiogram image|Finding|false|false||EKG
null|Electrocardiogram|Finding|false|false||EKGnull|Electrocardiography|Procedure|false|false||EKGnull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|Myocardium|Anatomy|false|false|C2681922;C1883709;C0010957|myocardialnull|Myocardial|Modifier|false|false||myocardialnull|Tissue damage|Disorder|false|false|C0027061|damagenull|Damage|Finding|false|false|C0027061|damage
null|MAGEE1 gene|Finding|false|false|C0027061|damagenull|Asymptomatic diagnosis of|Finding|false|false||asymptomatic
null|Asymptomatic (finding)|Finding|false|false||asymptomaticnull|Menstruation|Finding|false|false||periodsnull|Supraventricular tachycardia|Disorder|false|false||supraventricular tachycardianull|Supraventricular Tachycardia by ECG Finding|Finding|false|false||supraventricular tachycardianull|Tachycardia by ECG Finding|Finding|false|false||tachycardia
null|Tachycardia|Finding|false|false||tachycardianull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|Exercise stress test|Procedure|false|false|C4318744|stress test
null|Stress Test|Procedure|false|false|C4318744|stress testnull|Stress bismuth subsalicylate|Drug|false|false||stress
null|Stress bismuth subsalicylate|Drug|false|false||stressnull|Stress|Finding|false|false|C4318744|stressnull|W stress|Attribute|false|false||stressnull|Tests (qualifier value)|Finding|false|false|C4318744|test
null|Testing|Finding|false|false|C4318744|testnull|Laboratory Procedures|Procedure|false|false|C4318744|testnull|Test - temporal region|Anatomy|false|false|C0015260;C3494508;C0456984;C0039593;C0392366;C0038435;C0022885|testnull|Test Result|Lab|false|false|C4318744|testnull|Test Dosing Unit|LabModifier|false|false||testnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|null|Attribute|false|false|C4266572;C0015392;C0700042|R eyenull|Eye pain|Finding|false|false|C4266572;C0015392;C0700042|eye painnull|Carcinoma in situ of eye|Disorder|false|false|C4266572;C0015392;C0700042|eye
null|Disorder of eye|Disorder|false|false|C4266572;C0015392;C0700042|eyenull|Eye - Specimen Source Code|Finding|false|false|C4266572;C0015392;C0700042|eye
null|Eye problem|Finding|false|false|C4266572;C0015392;C0700042|eye
null|Eye Specimen|Finding|false|false|C4266572;C0015392;C0700042|eyenull|Head>Eye|Anatomy|false|false|C1550636;C1546630;C0262477;C0154094;C0015397;C0151827;C5886197|eye
null|Eye|Anatomy|false|false|C1550636;C1546630;C0262477;C0154094;C0015397;C0151827;C5886197|eye
null|Orbital region|Anatomy|false|false|C1550636;C1546630;C0262477;C0154094;C0015397;C0151827;C5886197|eyenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Erythema|Disorder|false|false||rednessnull|Redness|Finding|false|false||rednessnull|Red color|Modifier|false|false||rednessnull|Dry Eyes brand of ocular lubricant|Drug|false|false|C0015392|dry eyesnull|Dry Eye Syndromes|Disorder|false|false|C0015392|dry eyes
null|Keratoconjunctivitis Sicca|Disorder|false|false|C0015392|dry eyesnull|Dryness of eye|Finding|false|false|C0015392|dry eyesnull|Eye|Anatomy|false|false|C0314719;C0720056;C5848506;C0022575;C0013238|eyesnull|null|Attribute|false|false|C0015392|eyesnull|erythromycin|Drug|false|false||erythromycin
null|erythromycin|Drug|false|false||erythromycinnull|Drops - Drug Form|Drug|false|false||dropsnull|Drop Dosing Unit|LabModifier|false|false||dropsnull|Tears (substance)|Finding|false|false||tears
null|null|Finding|false|false||tears
null|Tears specimen|Finding|false|false||tearsnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|4-azido-7-phenylpyrazolo-(1,5a)-1,3,5-triazine|Drug|false|false||appt
null|4-azido-7-phenylpyrazolo-(1,5a)-1,3,5-triazine|Drug|false|false||apptnull|5 Days|Time|false|false||5 daysnull|day|Time|false|false||daysnull|Full|Modifier|false|false||Fullnull|MDF Attribute Type - Code|Finding|false|false||Code
null|A Codes|Finding|false|false||Code
null|Code|Finding|false|false||Codenull|Coding|Event|false|false||Codenull|Contact - HL7 Attribution|Finding|false|false||Contact
null|Contact with|Finding|false|false||Contact
null|Communication Contact|Finding|false|false||Contactnull|contact person|Subject|false|false||Contactnull|Physical contact|Phenomenon|false|false||Contactnull|Personal Contact|Event|false|false||Contactnull|Contact - HL7 Attribution|Finding|false|false||CONTACT
null|Contact with|Finding|false|false||CONTACT
null|Communication Contact|Finding|false|false||CONTACTnull|contact person|Subject|false|false||CONTACTnull|Physical contact|Phenomenon|false|false||CONTACTnull|Personal Contact|Event|false|false||CONTACTnull|husband|Subject|false|false||husbandnull|Daughter|Subject|false|false||daughternull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|MEDICATION LIST|Finding|false|false||Medication listnull|Pharmaceutical Preparations|Drug|false|false||Medicationnull|medication - HL7 publishing domain|Finding|false|false||Medication
null|Medications|Finding|false|false||Medicationnull|List|Finding|false|false||list
null|Sequence Data Type|Finding|false|false||listnull|Accurate (qualifier value)|Modifier|false|false||accuratenull|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||completenull|Completion Status for valid values - Complete|Finding|false|false||complete
null|Data operation - complete|Finding|false|false||complete
null|Finish - dosing instruction imperative|Finding|false|false||completenull|Complete|Modifier|false|false||completenull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Every four hours|Time|false|false||Q4Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|albuterol|Drug|false|false||Albuterol
null|albuterol|Drug|false|false||Albuterolnull|NEB protein, human|Drug|false|false||Neb
null|NEB protein, human|Drug|false|false||Neb
null|Nebulizer solution|Drug|false|false||Nebnull|NEB gene|Finding|false|false||Neb
null|mitotic nuclear membrane disassembly|Finding|false|false||Nebnull|NEB protein, human|Drug|false|false||NEB
null|NEB protein, human|Drug|false|false||NEB
null|Nebulizer solution|Drug|false|false||NEBnull|NEB gene|Finding|false|false||NEB
null|mitotic nuclear membrane disassembly|Finding|false|false||NEBnull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Breath|Finding|false|false||breathnull|aspirin|Drug|false|false||Aspirin
null|aspirin|Drug|false|false||Aspirinnull|Daily|Time|false|false||DAILYnull|atorvastatin|Drug|false|false||Atorvastatin
null|atorvastatin|Drug|false|false||Atorvastatinnull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|clopidogrel|Drug|false|false||Clopidogrel
null|clopidogrel|Drug|false|false||Clopidogrelnull|Daily|Time|false|false||DAILYnull|diltiazem|Drug|false|false||Diltiazem
null|diltiazem|Drug|false|false||Diltiazemnull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Daily|Time|false|false||DAILYnull|fluticasone propionate|Drug|false|false||Fluticasone Propionate
null|fluticasone propionate|Drug|false|false||Fluticasone Propionatenull|fluticasone|Drug|false|false||Fluticasone
null|fluticasone|Drug|false|false||Fluticasonenull|propionate|Drug|false|false||Propionate
null|Propionates|Drug|false|false||Propionatenull|Nasal brand of oxymetazoline|Drug|false|false|C0028429|NASAL
null|Nasal brand of oxymetazoline|Drug|false|false|C0028429|NASAL
null|Nasal dosage form|Drug|false|false|C0028429|NASALnull|Nasal Route of Administration|Finding|false|false|C0028429|NASAL
null|Nasal (intended site)|Finding|false|false|C0028429|NASALnull|null|Anatomy|false|false|C1272939;C0721966;C4520890;C1522019|NASALnull|Daily|Time|false|false||DAILYnull|CIAO3 gene|Finding|false|false|C0028429|PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Nasal brand of oxymetazoline|Drug|false|false|C0028429|nasal
null|Nasal brand of oxymetazoline|Drug|false|false|C0028429|nasal
null|Nasal dosage form|Drug|false|false|C0028429|nasalnull|Nasal Route of Administration|Finding|false|false|C0028429|nasal
null|Nasal (intended site)|Finding|false|false|C0028429|nasalnull|null|Anatomy|false|false|C1422467;C4520890;C1522019;C1272939;C0721966|nasalnull|Congestion|Finding|false|false||congestionnull|Fluticasone-Salmeterol Diskus|Drug|false|false||Fluticasone-Salmeterol Diskus
null|Fluticasone-Salmeterol Diskus|Drug|false|false||Fluticasone-Salmeterol Diskusnull|fluticasone / salmeterol|Drug|false|false||Fluticasone-Salmeterolnull|fluticasone|Drug|false|false||Fluticasone
null|fluticasone|Drug|false|false||Fluticasonenull|salmeterol|Drug|false|false||Salmeterol
null|salmeterol|Drug|false|false||Salmeterolnull|Diskus|Device|false|false||Diskusnull|Inhalant dose form|Drug|false|false||INH
null|isoniazid|Drug|false|false||INH
null|isoniazid|Drug|false|false||INHnull|Inhalation Route of Administration|Finding|false|false||INHnull|Ingush language|Entity|false|false||INHnull|Inhalation Dosing Unit|LabModifier|false|false||INHnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|hydrochlorothiazide|Drug|false|false||Hydrochlorothiazide
null|hydrochlorothiazide|Drug|false|false||Hydrochlorothiazidenull|Daily|Time|false|false||DAILYnull|isosorbide mononitrate|Drug|false|false||Isosorbide Mononitrate
null|isosorbide mononitrate|Drug|false|false||Isosorbide Mononitratenull|isosorbide|Drug|false|false||Isosorbide
null|isosorbide|Drug|false|false||Isosorbidenull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Daily|Time|false|false||DAILYnull|latanoprost|Drug|false|false||Latanoprost
null|latanoprost|Drug|false|false||Latanoprostnull|Ophthalmic Route of Administration|Finding|false|false||Ophthnull|Drops - Drug Form|Drug|false|false|C0229090|DROPnull|Dropping|Event|false|false|C0229090|DROPnull|Drop (unit of presentation)|LabModifier|false|false||DROP
null|Drop British|LabModifier|false|false||DROP
null|Drop Dosing Unit|LabModifier|false|false||DROP
null|Medical Drop|LabModifier|false|false||DROP
null|Drop Unit of Volume|LabModifier|false|false||DROPnull|examination of left eye|Procedure|false|false|C4266572;C0015392;C0700042;C0229090|LEFT EYEnull|Left eye structure|Anatomy|false|false|C1705648;C1550636;C1546630;C0262477;C0991568;C2141124;C1552822;C0154094;C0015397|LEFT EYEnull|Table Cell Horizontal Align - left|Finding|false|false|C4266572;C0015392;C0700042;C0229090|LEFTnull|Left sided|Modifier|false|false||LEFT
null|Left|Modifier|false|false||LEFTnull|Carcinoma in situ of eye|Disorder|false|false|C4266572;C0015392;C0700042;C0229090|EYE
null|Disorder of eye|Disorder|false|false|C4266572;C0015392;C0700042;C0229090|EYEnull|Eye - Specimen Source Code|Finding|false|false|C0229090;C4266572;C0015392;C0700042|EYE
null|Eye problem|Finding|false|false|C0229090;C4266572;C0015392;C0700042|EYE
null|Eye Specimen|Finding|false|false|C0229090;C4266572;C0015392;C0700042|EYEnull|Head>Eye|Anatomy|false|false|C2141124;C1550636;C1546630;C0262477;C0154094;C0015397;C1552822|EYE
null|Eye|Anatomy|false|false|C2141124;C1550636;C1546630;C0262477;C0154094;C0015397;C1552822|EYE
null|Orbital region|Anatomy|false|false|C2141124;C1550636;C1546630;C0262477;C0154094;C0015397;C1552822|EYEnull|lorazepam|Drug|false|false||Lorazepam
null|lorazepam|Drug|false|false||Lorazepamnull|Once a day, at bedtime|Time|false|false||QHSnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Insomnia homeopathic medication|Drug|false|false||insomnianull|Sleeplessness|Finding|false|false||insomnianull|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin Drug Class|Drug|false|false||Multivitamins
null|Multivitamin Drug Class|Drug|false|false||Multivitaminsnull|Minerals|Drug|false|false||mineralsnull|Tablet Dosage Form|Drug|false|false||TABnull|Tablet Dosing Unit|LabModifier|false|false||TABnull|Daily|Time|false|false||DAILYnull|ranitidine|Drug|false|false||Ranitidine
null|ranitidine|Drug|false|false||Ranitidinenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|tramadol|Drug|false|false||TraMADOL
null|tramadol|Drug|false|false||TraMADOLnull|Tramadol measurement (procedure)|Procedure|false|false||TraMADOLnull|Ultram|Drug|false|false||Ultram
null|Ultram|Drug|false|false||Ultramnull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Theophylline ER|Drug|false|false||Theophylline ER
null|Theophylline ER|Drug|false|false||Theophylline ERnull|theophylline|Drug|false|false||Theophylline
null|theophylline|Drug|false|false||Theophyllinenull|Assay of theophylline|Procedure|false|false||Theophyllinenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|tiotropium bromide|Drug|false|false||Tiotropium Bromide
null|tiotropium bromide|Drug|false|false||Tiotropium Bromidenull|tiotropium|Drug|false|false||Tiotropium
null|tiotropium|Drug|false|false||Tiotropiumnull|Bromides|Drug|false|false||Bromidenull|Bromides measurement|Procedure|false|false||Bromidenull|capsule (pharmacologic)|Drug|false|false||CAPnull|CATARACT, ANTERIOR POLAR|Disorder|false|false||CAPnull|BRD4 wt Allele|Finding|false|false||CAP
null|HACD1 gene|Finding|false|false||CAP
null|SERPINB6 gene|Finding|false|false||CAP
null|BRD4 gene|Finding|false|false||CAP
null|CAP1 gene|Finding|false|false||CAP
null|SORBS1 gene|Finding|false|false||CAP
null|LNPEP gene|Finding|false|false||CAPnull|CAP Regimen|Procedure|false|false||CAP
null|cisplatin/cyclophosphamide/doxorubicin protocol|Procedure|false|false||CAP
null|cyclophosphamide/doxorubicin/prednisone protocol|Procedure|false|false||CAPnull|Cap (physical object)|Device|false|false||CAP
null|Syringe Caps|Device|false|false||CAP
null|Cap device|Device|false|false||CAPnull|College of American Pathologists|Subject|false|false||CAPnull|Controlled Attenuation Parameter|Modifier|false|false||CAPnull|Capsule Dosing Unit|LabModifier|false|false||CAPnull|Daily|Time|false|false||DAILYnull|guaifenesin|Drug|false|false||Guaifenesin
null|guaifenesin|Drug|false|false||Guaifenesinnull|codeine phosphate|Drug|false|false||CODEINE Phosphate
null|codeine phosphate|Drug|false|false||CODEINE Phosphatenull|codeine|Drug|false|false||CODEINE
null|codeine|Drug|false|false||CODEINEnull|phosphate ion|Drug|false|false||Phosphate
null|Phosphates|Drug|false|false||Phosphate
null|phosphate ion|Drug|false|false||Phosphatenull|Phosphate measurement|Procedure|false|false||Phosphatenull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|cod liver oil|Drug|false|false|C4037986;C1278929;C0023884|cod liver oil
null|cod liver oil|Drug|false|false|C4037986;C1278929;C0023884|cod liver oil
null|cod liver oil|Drug|false|false|C4037986;C1278929;C0023884|cod liver oilnull|cod, unspecified preparation|Drug|false|false||cod
null|null|Drug|false|false||cod
null|Cyclophosphamide/Dacarbazine/Vincristine|Drug|false|false||cod
null|cod, unspecified preparation|Drug|false|false||cod
null|codfish allergenic extract|Drug|false|false||cod
null|codfish allergenic extract|Drug|false|false||codnull|Cancerization of Pancreatic Ducts|Finding|false|false|C4037986;C1278929;C0023884|cod
null|Cemento-osseous dysplasia|Finding|false|false|C4037986;C1278929;C0023884|cod
null|SNRPB gene|Finding|false|false|C4037986;C1278929;C0023884|cod
null|Cause of Death|Finding|false|false|C4037986;C1278929;C0023884|codnull|Cod|Entity|false|false||codnull|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|liver
null|liver extract|Drug|false|false|C4037986;C1278929;C0023884|liver
null|liver extract|Drug|false|false|C4037986;C1278929;C0023884|liver
null|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|liver
null|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|livernull|Benign neoplasm of liver|Disorder|false|false|C4037986;C1278929;C0023884|liver
null|Liver diseases|Disorder|false|false|C4037986;C1278929;C0023884|livernull|Liver problem|Finding|false|false|C4037986;C1278929;C0023884|livernull|Procedures on liver|Procedure|false|false|C4037986;C1278929;C0023884|livernull|Abdomen>Liver|Anatomy|false|false|C0721399;C0023899;C0009213;C0023895;C0496870;C0577060;C0872387;C5444130;C0457523;C1420285;C0007465|liver
null|null|Anatomy|false|false|C0721399;C0023899;C0009213;C0023895;C0496870;C0577060;C0872387;C5444130;C0457523;C1420285;C0007465|liver
null|Liver|Anatomy|false|false|C0721399;C0023899;C0009213;C0023895;C0496870;C0577060;C0872387;C5444130;C0457523;C1420285;C0007465|livernull|oil ingredients|Drug|false|false||oil
null|oil ingredients|Drug|false|false||oil
null|Oil Dosage Form|Drug|false|false||oil
null|Oils|Drug|false|false||oil
null|Food Oil|Drug|false|false||oilnull|Storage Unit|Device|false|false||unit
null|Unit device|Device|false|false||unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||unit
null|Unit of Measure|LabModifier|false|false||unit
null|Unit|LabModifier|false|false||unit
null|Enzyme Unit|LabModifier|false|false||unitnull|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C4546282;C1527415;C4521986;C1332410;C1272919|oralnull|Oral|Modifier|false|false||oralnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false|C0226896|BIDnull|BID gene|Finding|false|false|C0226896|BIDnull|Twice a day|Time|false|false||BIDnull|CalCarb|Drug|false|false||Calcarbnull|Vitamin D Drug Class|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|D Vitamin|Drug|false|false||Vitamin D
null|Vitamin D [EPC]|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|Vitamin D Drug Class|Drug|false|false||Vitamin Dnull|Vitamin D measurement|Procedure|false|false||Vitamin Dnull|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitaminnull|calcium carbonate|Drug|false|false||calcium carbonate
null|calcium carbonate|Drug|false|false||calcium carbonatenull|CALCIUM SUPPLEMENTS|Drug|false|false||calcium
null|calcium|Drug|false|false||calcium
null|calcium|Drug|false|false||calcium
null|calcium|Drug|false|false||calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||calcium
null|Calcium, Dietary|Drug|false|false||calcium
null|Calcium [EPC]|Drug|false|false||calcium
null|Calcium Drug Class|Drug|false|false||calciumnull|Calcium metabolic function|Finding|false|false||calciumnull|Calcium measurement|Procedure|false|false||calciumnull|carbonate ion|Drug|false|false||carbonate
null|Carbonates|Drug|false|false||carbonate
null|Carbonates|Drug|false|false||carbonatenull|vitamin D3|Drug|false|false||vitamin D3
null|vitamin D3|Drug|false|false||vitamin D3
null|cholecalciferol|Drug|false|false||vitamin D3
null|cholecalciferol|Drug|false|false||vitamin D3
null|cholecalciferol|Drug|false|false||vitamin D3null|Vitamins|Drug|false|false||vitamin
null|Vitamins|Drug|false|false||vitamin
null|Vitamins|Drug|false|false||vitaminnull|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C1527415;C4521986;C1272919|oralnull|Oral|Modifier|false|false||oralnull|Daily|Time|false|false||dailynull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|amiodarone|Drug|false|false||Amiodarone
null|amiodarone|Drug|false|false||Amiodaronenull|Drug assay amiodarone|Procedure|false|false||Amiodaronenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|amiodarone|Drug|false|false||amiodarone
null|amiodarone|Drug|false|false||amiodaronenull|Drug assay amiodarone|Procedure|false|false||amiodaronenull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false|C0230028;C0226896|by mouthnull|Oral cavity|Anatomy|false|false|C1527415;C1561538;C1561539|mouth
null|Oral region|Anatomy|false|false|C1527415;C1561538;C1561539|mouthnull|Twice a day|Time|false|false||twice a daynull|Transaction counts and value totals - day|Finding|false|false|C0230028;C0226896|day
null|Precision - day|Finding|false|false|C0230028;C0226896|daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|rivaroxaban|Drug|false|false||Rivaroxaban
null|rivaroxaban|Drug|false|false||Rivaroxabannull|Dinner|Finding|false|false||DINNERnull|With dinner|Time|false|false||DINNERnull|rivaroxaban|Drug|false|false||rivaroxaban
null|rivaroxaban|Drug|false|false||rivaroxabannull|Xarelto|Drug|false|false||Xarelto
null|Xarelto|Drug|false|false||Xareltonull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false|C0230028;C0226896|by mouthnull|Oral cavity|Anatomy|false|false|C1527415|mouth
null|Oral region|Anatomy|false|false|C1527415|mouthnull|QPM|Time|false|false||qpm
null|Once a day, in the evening|Time|false|false||qpmnull|PRSS30P gene|Finding|false|false||Dispnull|Dispense (activity)|Event|false|false||Dispnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Every four hours|Time|false|false||Q4Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|albuterol|Drug|false|false||Albuterol
null|albuterol|Drug|false|false||Albuterolnull|NEB protein, human|Drug|false|false||Neb
null|NEB protein, human|Drug|false|false||Neb
null|Nebulizer solution|Drug|false|false||Nebnull|NEB gene|Finding|false|false||Neb
null|mitotic nuclear membrane disassembly|Finding|false|false||Nebnull|NEB protein, human|Drug|false|false||NEB
null|NEB protein, human|Drug|false|false||NEB
null|Nebulizer solution|Drug|false|false||NEBnull|NEB gene|Finding|false|false||NEB
null|mitotic nuclear membrane disassembly|Finding|false|false||NEBnull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Breath|Finding|false|false||breathnull|aspirin|Drug|false|false||Aspirin
null|aspirin|Drug|false|false||Aspirinnull|Daily|Time|false|false||DAILYnull|atorvastatin|Drug|false|false||Atorvastatin
null|atorvastatin|Drug|false|false||Atorvastatinnull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|diltiazem|Drug|false|false||Diltiazem
null|diltiazem|Drug|false|false||Diltiazemnull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Daily|Time|false|false||DAILYnull|fluticasone propionate|Drug|false|false||Fluticasone Propionate
null|fluticasone propionate|Drug|false|false||Fluticasone Propionatenull|fluticasone|Drug|false|false||Fluticasone
null|fluticasone|Drug|false|false||Fluticasonenull|propionate|Drug|false|false||Propionate
null|Propionates|Drug|false|false||Propionatenull|Nasal brand of oxymetazoline|Drug|false|false|C0028429|NASAL
null|Nasal brand of oxymetazoline|Drug|false|false|C0028429|NASAL
null|Nasal dosage form|Drug|false|false|C0028429|NASALnull|Nasal Route of Administration|Finding|false|false|C0028429|NASAL
null|Nasal (intended site)|Finding|false|false|C0028429|NASALnull|null|Anatomy|false|false|C1272939;C0721966;C4520890;C1522019|NASALnull|Daily|Time|false|false||DAILYnull|CIAO3 gene|Finding|false|false|C0028429|PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Nasal brand of oxymetazoline|Drug|false|false|C0028429|nasal
null|Nasal brand of oxymetazoline|Drug|false|false|C0028429|nasal
null|Nasal dosage form|Drug|false|false|C0028429|nasalnull|Nasal Route of Administration|Finding|false|false|C0028429|nasal
null|Nasal (intended site)|Finding|false|false|C0028429|nasalnull|null|Anatomy|false|false|C1272939;C0721966;C4520890;C1522019;C1422467|nasalnull|Congestion|Finding|false|false||congestionnull|Fluticasone-Salmeterol Diskus|Drug|false|false||Fluticasone-Salmeterol Diskus
null|Fluticasone-Salmeterol Diskus|Drug|false|false||Fluticasone-Salmeterol Diskusnull|fluticasone / salmeterol|Drug|false|false||Fluticasone-Salmeterolnull|fluticasone|Drug|false|false||Fluticasone
null|fluticasone|Drug|false|false||Fluticasonenull|salmeterol|Drug|false|false||Salmeterol
null|salmeterol|Drug|false|false||Salmeterolnull|Diskus|Device|false|false||Diskusnull|Inhalant dose form|Drug|false|false||INH
null|isoniazid|Drug|false|false||INH
null|isoniazid|Drug|false|false||INHnull|Inhalation Route of Administration|Finding|false|false||INHnull|Ingush language|Entity|false|false||INHnull|Inhalation Dosing Unit|LabModifier|false|false||INHnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|guaifenesin|Drug|false|false||Guaifenesin
null|guaifenesin|Drug|false|false||Guaifenesinnull|codeine phosphate|Drug|false|false||CODEINE Phosphate
null|codeine phosphate|Drug|false|false||CODEINE Phosphatenull|codeine|Drug|false|false||CODEINE
null|codeine|Drug|false|false||CODEINEnull|phosphate ion|Drug|false|false||Phosphate
null|Phosphates|Drug|false|false||Phosphate
null|phosphate ion|Drug|false|false||Phosphatenull|Phosphate measurement|Procedure|false|false||Phosphatenull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|hydrochlorothiazide|Drug|false|false||Hydrochlorothiazide
null|hydrochlorothiazide|Drug|false|false||Hydrochlorothiazidenull|Daily|Time|false|false||DAILYnull|isosorbide mononitrate|Drug|false|false||Isosorbide Mononitrate
null|isosorbide mononitrate|Drug|false|false||Isosorbide Mononitratenull|isosorbide|Drug|false|false||Isosorbide
null|isosorbide|Drug|false|false||Isosorbidenull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Daily|Time|false|false||DAILYnull|latanoprost|Drug|false|false||Latanoprost
null|latanoprost|Drug|false|false||Latanoprostnull|Ophthalmic Route of Administration|Finding|false|false||Ophthnull|Drops - Drug Form|Drug|false|false|C0229090|DROPnull|Dropping|Event|false|false|C0229090|DROPnull|Drop (unit of presentation)|LabModifier|false|false||DROP
null|Drop British|LabModifier|false|false||DROP
null|Drop Dosing Unit|LabModifier|false|false||DROP
null|Medical Drop|LabModifier|false|false||DROP
null|Drop Unit of Volume|LabModifier|false|false||DROPnull|examination of left eye|Procedure|false|false|C0229090;C4266572;C0015392;C0700042|LEFT EYEnull|Left eye structure|Anatomy|false|false|C0154094;C0015397;C1550636;C1546630;C0262477;C2141124;C1705648;C0991568;C1552822|LEFT EYEnull|Table Cell Horizontal Align - left|Finding|false|false|C4266572;C0015392;C0700042;C0229090|LEFTnull|Left sided|Modifier|false|false||LEFT
null|Left|Modifier|false|false||LEFTnull|Carcinoma in situ of eye|Disorder|false|false|C0229090;C4266572;C0015392;C0700042|EYE
null|Disorder of eye|Disorder|false|false|C0229090;C4266572;C0015392;C0700042|EYEnull|Eye - Specimen Source Code|Finding|false|false|C0229090;C4266572;C0015392;C0700042|EYE
null|Eye problem|Finding|false|false|C0229090;C4266572;C0015392;C0700042|EYE
null|Eye Specimen|Finding|false|false|C0229090;C4266572;C0015392;C0700042|EYEnull|Head>Eye|Anatomy|false|false|C0154094;C0015397;C1552822;C1550636;C1546630;C0262477;C2141124|EYE
null|Eye|Anatomy|false|false|C0154094;C0015397;C1552822;C1550636;C1546630;C0262477;C2141124|EYE
null|Orbital region|Anatomy|false|false|C0154094;C0015397;C1552822;C1550636;C1546630;C0262477;C2141124|EYEnull|lorazepam|Drug|false|false||Lorazepam
null|lorazepam|Drug|false|false||Lorazepamnull|Once a day, at bedtime|Time|false|false||QHSnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Insomnia homeopathic medication|Drug|false|false||insomnianull|Sleeplessness|Finding|false|false||insomnianull|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin Drug Class|Drug|false|false||Multivitamins
null|Multivitamin Drug Class|Drug|false|false||Multivitaminsnull|Minerals|Drug|false|false||mineralsnull|Tablet Dosage Form|Drug|false|false||TABnull|Tablet Dosing Unit|LabModifier|false|false||TABnull|Daily|Time|false|false||DAILYnull|ranitidine|Drug|false|false||Ranitidine
null|ranitidine|Drug|false|false||Ranitidinenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Theophylline ER|Drug|false|false||Theophylline ER
null|Theophylline ER|Drug|false|false||Theophylline ERnull|theophylline|Drug|false|false||Theophylline
null|theophylline|Drug|false|false||Theophyllinenull|Assay of theophylline|Procedure|false|false||Theophyllinenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|tiotropium bromide|Drug|false|false||Tiotropium Bromide
null|tiotropium bromide|Drug|false|false||Tiotropium Bromidenull|tiotropium|Drug|false|false||Tiotropium
null|tiotropium|Drug|false|false||Tiotropiumnull|Bromides|Drug|false|false||Bromidenull|Bromides measurement|Procedure|false|false||Bromidenull|capsule (pharmacologic)|Drug|false|false||CAPnull|CATARACT, ANTERIOR POLAR|Disorder|false|false||CAPnull|BRD4 wt Allele|Finding|false|false||CAP
null|HACD1 gene|Finding|false|false||CAP
null|SERPINB6 gene|Finding|false|false||CAP
null|BRD4 gene|Finding|false|false||CAP
null|CAP1 gene|Finding|false|false||CAP
null|SORBS1 gene|Finding|false|false||CAP
null|LNPEP gene|Finding|false|false||CAPnull|CAP Regimen|Procedure|false|false||CAP
null|cisplatin/cyclophosphamide/doxorubicin protocol|Procedure|false|false||CAP
null|cyclophosphamide/doxorubicin/prednisone protocol|Procedure|false|false||CAPnull|Cap (physical object)|Device|false|false||CAP
null|Syringe Caps|Device|false|false||CAP
null|Cap device|Device|false|false||CAPnull|College of American Pathologists|Subject|false|false||CAPnull|Controlled Attenuation Parameter|Modifier|false|false||CAPnull|Capsule Dosing Unit|LabModifier|false|false||CAPnull|Daily|Time|false|false||DAILYnull|tramadol|Drug|false|false||TraMADOL
null|tramadol|Drug|false|false||TraMADOLnull|Tramadol measurement (procedure)|Procedure|false|false||TraMADOLnull|Ultram|Drug|false|false||Ultram
null|Ultram|Drug|false|false||Ultramnull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|artificial tears (medication)|Drug|false|false||Artificial Tears
null|Lubricant Eye Drops|Drug|false|false||Artificial Tears
null|Artificial Tears|Drug|false|false||Artificial Tearsnull|Artificial (qualifier value)|Modifier|false|false||Artificialnull|Tears (substance)|Finding|false|false||Tears
null|null|Finding|false|false||Tears
null|Tears specimen|Finding|false|false||Tearsnull|Preserving|Finding|false|false||Preservnull|Biologic Preservation|Procedure|false|false||Preservnull|Free of (attribute)|Finding|false|false||Freenull|Empty (qualifier)|Modifier|false|false||Freenull|Drops - Drug Form|Drug|false|false||DROPnull|Dropping|Event|false|false||DROPnull|Drop (unit of presentation)|LabModifier|false|false||DROP
null|Drop British|LabModifier|false|false||DROP
null|Drop Dosing Unit|LabModifier|false|false||DROP
null|Medical Drop|LabModifier|false|false||DROP
null|Drop Unit of Volume|LabModifier|false|false||DROPnull|Structure of both eyes|Anatomy|false|false||BOTH EYESnull|Eye|Anatomy|false|false|C5848506|EYESnull|null|Attribute|false|false|C0015392|EYESnull|CIAO3 gene|Finding|false|false|C4266572;C0015392;C0700042|PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Carcinoma in situ of eye|Disorder|false|false|C4266572;C0015392;C0700042|eye
null|Disorder of eye|Disorder|false|false|C4266572;C0015392;C0700042|eyenull|Eye - Specimen Source Code|Finding|false|false|C4266572;C0015392;C0700042|eye
null|Eye problem|Finding|false|false|C4266572;C0015392;C0700042|eye
null|Eye Specimen|Finding|false|false|C4266572;C0015392;C0700042|eyenull|Head>Eye|Anatomy|false|false|C1550636;C1546630;C0262477;C1422467;C0154094;C0015397|eye
null|Eye|Anatomy|false|false|C1550636;C1546630;C0262477;C1422467;C0154094;C0015397|eye
null|Orbital region|Anatomy|false|false|C1550636;C1546630;C0262477;C1422467;C0154094;C0015397|eyenull|Have Vulvar Irritation question|Finding|false|false||irritation
null|Irritability - emotion|Finding|false|false||irritation
null|Irritation (finding)|Finding|false|false||irritationnull|Irritation|Phenomenon|false|false||irritationnull|dextran 70|Drug|false|false||dextran 70
null|dextran 70|Drug|false|false||dextran 70null|dextran|Drug|false|false||dextran
null|dextran|Drug|false|false||dextran
null|Dextrans|Drug|false|false||dextran
null|Dextrans|Drug|false|false||dextrannull|hypromellose|Drug|false|false||hypromellose
null|hypromellose|Drug|false|false||hypromellosenull|artificial tears (medication)|Drug|false|false||Artificial Tears
null|Lubricant Eye Drops|Drug|false|false||Artificial Tears
null|Artificial Tears|Drug|false|false||Artificial Tearsnull|Artificial (qualifier value)|Modifier|false|false||Artificialnull|Tears (substance)|Finding|false|false||Tears
null|null|Finding|false|false||Tears
null|Tears specimen|Finding|false|false||Tearsnull|Drops - Drug Form|Drug|false|false||dropnull|Dropping|Event|false|false||dropnull|Drop (unit of presentation)|LabModifier|false|false||drop
null|Drop British|LabModifier|false|false||drop
null|Drop Dosing Unit|LabModifier|false|false||drop
null|Medical Drop|LabModifier|false|false||drop
null|Drop Unit of Volume|LabModifier|false|false||dropnull|Four times daily|Time|false|false||QIDnull|CIAO3 gene|Finding|false|false||prnnull|As required|Time|false|false||prn
null|Pro Re Nata|Time|false|false||prnnull|refill|Finding|false|false||Refillsnull|dextran 70|Drug|false|false||dextran 70
null|dextran 70|Drug|false|false||dextran 70null|dextran|Drug|false|false||dextran
null|dextran|Drug|false|false||dextran
null|Dextrans|Drug|false|false||dextran
null|Dextrans|Drug|false|false||dextrannull|hypromellose|Drug|false|false||hypromellose
null|hypromellose|Drug|false|false||hypromellosenull|artificial tears (medication)|Drug|false|false||Artificial Tears
null|Lubricant Eye Drops|Drug|false|false||Artificial Tears
null|Artificial Tears|Drug|false|false||Artificial Tearsnull|Artificial (qualifier value)|Modifier|false|false||Artificialnull|Tears (substance)|Finding|false|false||Tears
null|null|Finding|false|false||Tears
null|Tears specimen|Finding|false|false||Tearsnull|Drops - Drug Form|Drug|false|false||dropsnull|Drop Dosing Unit|LabModifier|false|false||dropsnull|Carcinoma in situ of eye|Disorder|false|false|C4266572;C0015392;C0700042|eye
null|Disorder of eye|Disorder|false|false|C4266572;C0015392;C0700042|eyenull|Eye - Specimen Source Code|Finding|false|false|C4266572;C0015392;C0700042|eye
null|Eye problem|Finding|false|false|C4266572;C0015392;C0700042|eye
null|Eye Specimen|Finding|false|false|C4266572;C0015392;C0700042|eyenull|Head>Eye|Anatomy|false|false|C1550636;C1546630;C0262477;C1704709;C0154094;C0015397|eye
null|Eye|Anatomy|false|false|C1550636;C1546630;C0262477;C1704709;C0154094;C0015397|eye
null|Orbital region|Anatomy|false|false|C1550636;C1546630;C0262477;C1704709;C0154094;C0015397|eyenull|Computer program package|Finding|false|false|C4266572;C0015392;C0700042|Packagenull|medical supply, miscellaneous MISCELL PACKAGE|Device|false|false||Package
null|Package|Device|false|false||Packagenull|Package Dosing Unit|LabModifier|false|false||Packagenull|refill|Finding|false|false||Refillsnull|erythromycin|Drug|false|false|C0229089|Erythromycin
null|erythromycin|Drug|false|false|C0229089|Erythromycinnull|Ophthalmic Route of Administration|Finding|false|false|C4266572;C0015392;C0700042;C0229089|Ophthnull|Ointments|Drug|false|false|C0229089|Ointnull|examination of right eye|Procedure|false|false|C4266572;C0015392;C0700042;C0229089|RIGHT EYEnull|Right eye|Anatomy|false|false|C0154094;C0015397;C1550636;C1546630;C0262477;C1522230;C0014806;C2177784;C0028912;C1552823|RIGHT EYEnull|Table Cell Horizontal Align - right|Finding|false|false|C4266572;C0015392;C0700042;C0229089|RIGHTnull|Right sided|Modifier|false|false||RIGHT
null|Right|Modifier|false|false||RIGHTnull|Carcinoma in situ of eye|Disorder|false|false|C0229089;C4266572;C0015392;C0700042|EYE
null|Disorder of eye|Disorder|false|false|C0229089;C4266572;C0015392;C0700042|EYEnull|Eye - Specimen Source Code|Finding|false|false|C4266572;C0015392;C0700042;C0229089|EYE
null|Eye problem|Finding|false|false|C4266572;C0015392;C0700042;C0229089|EYE
null|Eye Specimen|Finding|false|false|C4266572;C0015392;C0700042;C0229089|EYEnull|Head>Eye|Anatomy|false|false|C1550636;C1546630;C0262477;C2177784;C1522230;C0154094;C0015397;C1552823|EYE
null|Eye|Anatomy|false|false|C1550636;C1546630;C0262477;C2177784;C1522230;C0154094;C0015397;C1552823|EYE
null|Orbital region|Anatomy|false|false|C1550636;C1546630;C0262477;C2177784;C1522230;C0154094;C0015397;C1552823|EYEnull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|erythromycin|Drug|false|false||erythromycin
null|erythromycin|Drug|false|false||erythromycinnull|gram|LabModifier|false|false||gramnull|Inch Unit of Length|LabModifier|false|false||inchnull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|CIAO3 gene|Finding|false|false||prnnull|As required|Time|false|false||prn
null|Pro Re Nata|Time|false|false||prnnull|refill|Finding|false|false||Refillsnull|CalCarb|Drug|false|false||Calcarbnull|Vitamin D Drug Class|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|D Vitamin|Drug|false|false||Vitamin D
null|Vitamin D [EPC]|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|Vitamin D Drug Class|Drug|false|false||Vitamin Dnull|Vitamin D measurement|Procedure|false|false||Vitamin Dnull|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitaminnull|calcium carbonate|Drug|false|false||calcium carbonate
null|calcium carbonate|Drug|false|false||calcium carbonatenull|CALCIUM SUPPLEMENTS|Drug|false|false||calcium
null|calcium|Drug|false|false||calcium
null|calcium|Drug|false|false||calcium
null|calcium|Drug|false|false||calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||calcium
null|Calcium, Dietary|Drug|false|false||calcium
null|Calcium [EPC]|Drug|false|false||calcium
null|Calcium Drug Class|Drug|false|false||calciumnull|Calcium metabolic function|Finding|false|false||calciumnull|Calcium measurement|Procedure|false|false||calciumnull|carbonate ion|Drug|false|false||carbonate
null|Carbonates|Drug|false|false||carbonate
null|Carbonates|Drug|false|false||carbonatenull|vitamin D3|Drug|false|false||vitamin D3
null|vitamin D3|Drug|false|false||vitamin D3
null|cholecalciferol|Drug|false|false||vitamin D3
null|cholecalciferol|Drug|false|false||vitamin D3
null|cholecalciferol|Drug|false|false||vitamin D3null|Vitamins|Drug|false|false||vitamin
null|Vitamins|Drug|false|false||vitamin
null|Vitamins|Drug|false|false||vitaminnull|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C1272919;C1527415;C4521986|oralnull|Oral|Modifier|false|false||oralnull|Daily|Time|false|false||dailynull|cod liver oil|Drug|false|false|C4037986;C1278929;C0023884|cod liver oil
null|cod liver oil|Drug|false|false|C4037986;C1278929;C0023884|cod liver oil
null|cod liver oil|Drug|false|false|C4037986;C1278929;C0023884|cod liver oilnull|cod, unspecified preparation|Drug|false|false||cod
null|null|Drug|false|false||cod
null|Cyclophosphamide/Dacarbazine/Vincristine|Drug|false|false||cod
null|cod, unspecified preparation|Drug|false|false||cod
null|codfish allergenic extract|Drug|false|false||cod
null|codfish allergenic extract|Drug|false|false||codnull|Cancerization of Pancreatic Ducts|Finding|false|false|C4037986;C1278929;C0023884|cod
null|Cemento-osseous dysplasia|Finding|false|false|C4037986;C1278929;C0023884|cod
null|SNRPB gene|Finding|false|false|C4037986;C1278929;C0023884|cod
null|Cause of Death|Finding|false|false|C4037986;C1278929;C0023884|codnull|Cod|Entity|false|false||codnull|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|liver
null|liver extract|Drug|false|false|C4037986;C1278929;C0023884|liver
null|liver extract|Drug|false|false|C4037986;C1278929;C0023884|liver
null|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|liver
null|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|livernull|Benign neoplasm of liver|Disorder|false|false|C4037986;C1278929;C0023884|liver
null|Liver diseases|Disorder|false|false|C4037986;C1278929;C0023884|livernull|Liver problem|Finding|false|false|C4037986;C1278929;C0023884|livernull|Procedures on liver|Procedure|false|false|C4037986;C1278929;C0023884|livernull|Abdomen>Liver|Anatomy|false|false|C0872387;C0577060;C0721399;C0023899;C0009213;C5444130;C0457523;C1420285;C0007465;C0023895;C0496870|liver
null|null|Anatomy|false|false|C0872387;C0577060;C0721399;C0023899;C0009213;C5444130;C0457523;C1420285;C0007465;C0023895;C0496870|liver
null|Liver|Anatomy|false|false|C0872387;C0577060;C0721399;C0023899;C0009213;C5444130;C0457523;C1420285;C0007465;C0023895;C0496870|livernull|oil ingredients|Drug|false|false||oil
null|oil ingredients|Drug|false|false||oil
null|Oil Dosage Form|Drug|false|false||oil
null|Oils|Drug|false|false||oil
null|Food Oil|Drug|false|false||oilnull|Storage Unit|Device|false|false||unit
null|Unit device|Device|false|false||unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||unit
null|Unit of Measure|LabModifier|false|false||unit
null|Unit|LabModifier|false|false||unit
null|Enzyme Unit|LabModifier|false|false||unitnull|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C1272919;C1527415;C4521986|oralnull|Oral|Modifier|false|false||oralnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Rapid atrial fibrillation|Disorder|false|false|C0018792|Rapid Atrial Fibrillationnull|Rapid|Modifier|false|false||Rapidnull|Atrial fibrillation and flutter|Finding|false|false|C0018792|Atrial Fibrillation/Flutternull|Atrial Fibrillation|Disorder|false|false|C0018792|Atrial Fibrillationnull|null|Attribute|false|false|C0018792|Atrial Fibrillationnull|Atrial Fibrillation by ECG Finding|Lab|false|false|C0018792|Atrial Fibrillationnull|Heart Atrium|Anatomy|false|false|C0016385;C2926591;C0155709;C1281999;C0004238;C0344434;C0232197|Atrialnull|Fibrillation|Disorder|false|false|C0018792|Fibrillationnull|Cardiac Flutter|Finding|false|false|C0018792|Flutternull|Flutter (respiratory device)|Device|false|false||Flutternull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Coordination of Benefits - Independent|Finding|false|false||Independent
null|Religious Affiliation - Independent|Finding|false|false||Independent
null|Independence|Finding|false|false||Independent
null|Independently able|Finding|false|false||Independentnull|FBXW7-AS1 gene|Finding|false|false||Dearnull|Chest Pain|Finding|false|false|C1527391;C0817096|chest painnull|null|Attribute|false|false|C1527391;C0817096|chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0008031;C0741025;C2926613|chest
null|Anterior thoracic region|Anatomy|false|false|C0008031;C0741025;C2926613|chestnull|Pain|Finding|false|false||pain symptomsnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Infrequent|Time|false|false||infrequentnull|Bursting sensation quality|Modifier|false|false||burstsnull|Rapid|Modifier|false|false||rapidnull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787|heart
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787|heartnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|heartnull|Chest>Heart|Anatomy|false|false|C0153957;C0153500;C0795691|heart
null|Heart|Anatomy|false|false|C0153957;C0153500;C0795691|heartnull|Amount type - Rate|Finding|false|false||ratenull|Rating (action)|Event|false|false||ratenull|Rate|LabModifier|false|false||ratenull|Rapid|Modifier|false|false||rapidnull|Amount type - Rate|Finding|false|false||ratenull|Rating (action)|Event|false|false||ratenull|Rate|LabModifier|false|false||ratenull|Increased risk|Finding|false|false||increased risknull|Risk|Finding|false|false||risknull|Cerebrovascular accident|Disorder|false|false||strokenull|Stroke (heart beat)|Finding|false|false||strokenull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Thinning Weight Loss|Finding|false|false||thinningnull|Decreased thickness|Modifier|false|false||thinningnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|rivaroxaban|Drug|false|false||Rivaroxaban
null|rivaroxaban|Drug|false|false||Rivaroxabannull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Specialized|Finding|false|false||specializednull|Special|Modifier|false|false||specializednull|Cardiologists|Subject|false|false||cardiologistsnull|Electrical (qualifier value)|Finding|false|false|C4037974;C0018787|electricalnull|Electricity|Phenomenon|false|false||electricalnull|Rhythm|Finding|false|false|C4037974;C0018787|rhythm
null|rhythmic process (biological)|Finding|false|false|C4037974;C0018787|rhythmnull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787|heart
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787|heartnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|heartnull|Chest>Heart|Anatomy|false|false|C0442828;C0153957;C0153500;C0795691;C1523018;C0871269|heart
null|Heart|Anatomy|false|false|C0442828;C0153957;C0153500;C0795691;C1523018;C0871269|heartnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|amiodarone|Drug|false|false||amiodarone
null|amiodarone|Drug|false|false||amiodaronenull|Drug assay amiodarone|Procedure|false|false||amiodaronenull|Clinic|Device|false|false||clinic
null|Ambulatory Care Facilities|Device|false|false||clinicnull|Clinic|Entity|false|false||clinic
null|Ambulatory Care Facilities|Entity|false|false||clinicnull|Patient location type - Clinic|Modifier|false|false||clinic
null|Person location type - Clinic|Modifier|false|false||clinicnull|Observation Interpretation - Abnormal|Finding|false|false||abnormal
null|Abnormal|Finding|false|false||abnormalnull|Rhythm|Finding|false|false||rhythm
null|rhythmic process (biological)|Finding|false|false||rhythmnull|Holter Electrocardiography|Procedure|false|false||Holter monitornull|Holter Monitors|Device|false|false||Holter monitornull|Monitor brand of insecticide|Drug|false|false||monitor
null|Monitor brand of insecticide|Drug|false|false||monitornull|Monitor Device|Device|false|false||monitor
null|Monitoring Device|Device|false|false||monitornull|Monitor, occupation|Subject|false|false||monitornull|null|Finding|false|false|C4037974;C0018787|heart ratenull|examination of heart rate|Procedure|false|false|C4037974;C0018787|heart ratenull|heart rate|Attribute|false|false|C4037974;C0018787|heart rate
null|null|Attribute|false|false|C4037974;C0018787|heart ratenull|Mean Heart Rate|LabModifier|false|false||heart ratenull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787|heart
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787|heartnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|heartnull|Chest>Heart|Anatomy|false|false|C2041121;C0795691;C0018810;C0488794;C0153957;C0153500;C2197023|heart
null|Heart|Anatomy|false|false|C2041121;C0795691;C0018810;C0488794;C0153957;C0153500;C2197023|heartnull|Amount type - Rate|Finding|false|false||ratenull|Rating (action)|Event|false|false||ratenull|Rate|LabModifier|false|false||ratenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Very Important|Finding|false|false||very importantnull|Very|Modifier|false|false||verynull|Important|Modifier|false|false||importantnull|Cardiologists|Subject|false|false||cardiologistnull|Vitelliform Macular Dystrophy|Disorder|false|false||bestnull|BEST1 wt Allele|Finding|false|false||best
null|BEST1 gene|Finding|false|false||bestnull|best (quality)|Modifier|false|false||bestnull|Care team|Finding|false|false||care teamnull|null|Attribute|false|false||care teamnull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Team|Subject|false|false||teamnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions