CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Level of Care - Surgery|Finding|false|false||SURGERY
null|Surgical procedure finding|Finding|false|false||SURGERY
null|Surgical aspects|Finding|false|false||SURGERYnull|Operative Surgical Procedures|Procedure|false|false||SURGERYnull|General surgery specialty|Title|false|false||SURGERY
null|Surgery specialty|Title|false|false||SURGERYnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Known|Modifier|false|false||Knownnull|Hypersensitivity|Finding|true|false||Allergiesnull|null|Attribute|true|false||Allergiesnull|Pharmaceutical Preparations|Drug|false|false||Drugsnull|Drugs - dental services|Procedure|false|false||Drugsnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Diverticulitis|Disorder|false|false||diverticulitisnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Laparoscopic-assisted sigmoid colectomy|Procedure|false|false|C0227391|laparoscopic sigmoid colectomy
null|Laparoscopic sigmoid colectomy|Procedure|false|false|C0227391|laparoscopic sigmoid colectomynull|Laparoscopy|Procedure|false|false||laparoscopicnull|Laparoscopic approach|Modifier|false|false||laparoscopicnull|Sigmoid colectomy|Procedure|false|false|C0227391|sigmoid colectomynull|Sigmoid colon|Anatomy|false|false|C0585462;C5890124;C0192866|sigmoidnull|Colectomy|Procedure|false|false||colectomynull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Recurrent|Time|false|false||recurrent
null|Episodic|Time|false|false||recurrentnull|Diverticulitis|Disorder|false|false||diverticulitisnull|One month|Time|false|false||one monthnull|Transaction counts and value totals - month|Finding|false|false||month
null|Precision - month|Finding|false|false||monthnull|month|Time|false|false||month
null|Monthly (qualifier value)|Time|false|false||monthnull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Structure of left lower quadrant of abdomen|Anatomy|false|false||LLQnull|Left lower quadrant|Modifier|false|false||LLQnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|With intensity|Modifier|false|false||intensitynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Course|Time|false|false||coursenull|Cipro|Drug|false|false||Cipro
null|Cipro|Drug|false|false||Cipronull|Flagyl|Drug|false|false||Flagyl
null|Flagyl|Drug|false|false||Flagylnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Abdominal Pain|Finding|false|false|C0000726|abdominal painnull|Abdomen|Anatomy|false|false|C0000737;C1549543;C0030193|abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Administration Method - Pain|Finding|false|false|C0000726|pain
null|Pain|Finding|false|false|C0000726|painnull|null|Attribute|false|false||painnull|1 Week|Time|false|false||one weeknull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|Antibiotics|Drug|false|false||antibioticnull|Course|Time|false|false||coursenull|Nausea or vomiting|Finding|true|false||nausea or vomitingnull|Nausea|Finding|true|false||nauseanull|null|Attribute|true|false||nauseanull|Vomiting|Finding|true|false||vomitingnull|Able (qualifier value)|Finding|false|false||ablenull|Ability|Subject|false|false||ablenull|Hydration status|Finding|false|false||hydration
null|Hydration|Finding|false|false||hydrationnull|Regular|Modifier|false|false||regularnull|Intake|Finding|false|false||intakenull|Measurement of fluid intake|Procedure|false|false||intake
null|Intake (treatment)|Procedure|false|false||intakenull|Desire for food|Finding|false|false||appetitenull|Somewhat|Finding|false|false||somewhatnull|Decreasing|Finding|false|false||decreased
null|Reduced|Finding|false|false||decreasednull|Decreased|LabModifier|false|false||decreasednull|Regular|Modifier|false|false||regularnull|Defecation|Finding|false|false|C0021853|bowel movementsnull|Intestines|Anatomy|false|false|C0011135|bowelnull|Movement|Finding|false|false||movementsnull|Several|LabModifier|false|false||severalnull|Small|LabModifier|false|false||smallnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||softnull|Soft|Modifier|false|false||softnull|Brown Tendon Sheath Syndrome|Disorder|false|false||brownnull|Brown color|Modifier|false|false||brownnull|Defecation|Finding|false|false|C0021853|bowel movementsnull|Intestines|Anatomy|false|false|C0011135|bowelnull|Movement|Finding|false|false||movementsnull|rectal discharge diarrhea (physical finding)|Finding|true|false||diarrhea
null|Diarrhea|Finding|true|false||diarrheanull|Direct - PostalAddressUse|Finding|false|false||direct
null|direct address|Finding|false|false||directnull|Direct type of relationship|Modifier|false|false||direct
null|Direct (qualifier)|Modifier|false|false||directnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Unresponsive to Treatment|Finding|false|false||refractorynull|Left lower quadrant pain|Finding|false|false|C0230180|LLQ painnull|Structure of left lower quadrant of abdomen|Anatomy|false|false|C1549543;C0030193;C0238551|LLQnull|Left lower quadrant|Modifier|false|false||LLQnull|Administration Method - Pain|Finding|false|false|C0230180|pain
null|Pain|Finding|false|false|C0230180|painnull|null|Attribute|false|false||painnull|Diverticulitis|Disorder|false|false||diverticulitisnull|Migraine Disorders|Disorder|false|false||Migrainesnull|Table Cell Horizontal Align - left|Finding|false|false|C4299059;C0851278;C0016129|Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|Upper extremity>Finger|Anatomy|false|false|C0007642;C1552822;C2025995|finger
null|Fingers|Anatomy|false|false|C0007642;C1552822;C2025995|finger
null|Fingers not including thumb|Anatomy|false|false|C0007642;C1552822;C2025995|fingernull|Cellulitis|Disorder|false|false|C4299059;C0851278;C0016129|cellulitisnull|cellulitis on exam (physical finding)|Finding|false|false|C4299059;C0851278;C0016129|cellulitisnull|Indirect exposure mechanism - Father|Finding|false|false||father
null|Relationship - Father|Finding|false|false||father
null|Father - courtesy title|Finding|false|false||fathernull|Father (person)|Subject|false|false||fathernull|Colitis|Disorder|false|false||colitisnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|C1orf210 gene|Finding|false|false||Tempnull|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Procedure|false|false||Tempnull|Temperature|LabModifier|false|false||Tempnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||Gen
null|GEN1 wt Allele|Finding|false|false||Gen
null|GEN1 gene|Finding|false|false||Gennull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|Respiratory, thoracic and mediastinal disorders|Disorder|false|false||RESPnull|Respiratory rate|Attribute|false|false||RESPnull|cetrimonium bromide|Drug|false|false||CTABnull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false|C0449202;C0000726|ABDnull|ABD (body structure)|Anatomy|false|false|C3811055|ABD
null|Abdomen|Anatomy|false|false|C3811055|ABDnull|Focal|Modifier|false|false||Focalnull|Emotional tenderness|Finding|false|false|C0230180|tenderness
null|Sore to touch|Finding|false|false|C0230180|tendernessnull|Structure of left lower quadrant of abdomen|Anatomy|false|false|C0684239;C0234233|LLQnull|Left lower quadrant|Modifier|false|false||LLQnull|Inferolateral|Modifier|false|false||inferolateralnull|Umbilical structure|Anatomy|false|false||umbilicusnull|Umbilicus <Crassulaceae>|Entity|false|false||umbilicusnull|Protective muscle spasm|Finding|true|false||guardingnull|Hereditary Multiple Exostoses|Disorder|false|false||EXTnull|EXT1 wt Allele|Finding|false|false||EXT
null|EXT1 gene|Finding|false|false||EXTnull|Edema|Finding|true|false||edemanull|null|Attribute|true|false||edemanull|radiology referral type|Finding|false|false||RADIOLOGY
null|Radiology Section ID|Finding|false|false||RADIOLOGY
null|Encounter due to radiological examination|Finding|false|false||RADIOLOGYnull|Radiology studies|Procedure|false|false||RADIOLOGY
null|Diagnostic radiologic examination|Procedure|false|false||RADIOLOGY
null|Radiographic imaging procedure|Procedure|false|false||RADIOLOGYnull|Radiology Specialty|Title|false|false||RADIOLOGYnull|Final report|Finding|false|false||Final Reportnull|Diagnosis Type - Final|Finding|false|false||Finalnull|Final|Time|false|false||Finalnull|End-stage|Modifier|false|false||Finalnull|Report (document)|Finding|false|false||Reportnull|Reporting|Procedure|false|false||Reportnull|null|Attribute|false|false||Reportnull|Computed tomography of pelvis|Procedure|false|false|C4266535;C0030797;C0559769|CT PELVISnull|null|Attribute|false|false|C4266535;C0030797;C0559769|CT PELVISnull|Malignant neoplasm of pelvis|Disorder|false|false|C4266535;C0030797;C0559769|PELVISnull|Pelvis problem|Finding|false|false|C4266535;C0030797;C0559769|PELVISnull|Pelvis+|Anatomy|false|false|C0412628;C0153663;C0882057;C0812455|PELVIS
null|Pelvic cavity structure|Anatomy|false|false|C0412628;C0153663;C0882057;C0812455|PELVIS
null|Pelvis|Anatomy|false|false|C0412628;C0153663;C0882057;C0812455|PELVISnull|Contrast Media|Drug|false|false||CONTRASTnull|Contrast|Modifier|false|false||CONTRASTnull|Medical Condition|Finding|false|false||MEDICAL CONDITIONnull|Medical referral type|Finding|false|false||MEDICAL
null|Medical|Finding|false|false||MEDICAL
null|Medical school type|Finding|false|false||MEDICALnull|Medical service|Procedure|false|false||MEDICALnull|Disease|Disorder|false|false||CONDITIONnull|Logical Condition|Finding|false|false||CONDITIONnull|null|Attribute|false|false||CONDITIONnull|Condition|Modifier|false|false||CONDITIONnull|Transaction counts and value totals - year|Finding|false|false||year
null|Precision - year|Finding|false|false||yearnull|year|Time|false|false||yearnull|Old|Time|false|false||oldnull|Woman|Subject|false|false||woman
null|Human, Female adult|Subject|false|false||womannull|Diverticulitis|Disorder|false|false||diverticulitisnull|Right lower quadrant pain|Finding|false|false|C0230178|RLQ painnull|Structure of right lower quadrant of abdomen|Anatomy|false|false|C0694551;C1549543;C0030193|RLQnull|Right lower quadrant|Modifier|false|false||RLQnull|Administration Method - Pain|Finding|false|false|C0230178|pain
null|Pain|Finding|false|false|C0230178|painnull|null|Attribute|false|false||painnull|impression (attitude)|Finding|false|false||IMPRESSION
null|EKG impression|Finding|false|false||IMPRESSIONnull|Moderate - Severity of Illness Code|Finding|false|false||Moderate
null|Moderate|Finding|false|false||Moderatenull|Moderate (severity modifier)|Modifier|false|false||Moderate
null|Moderate - Allergy Severity|Modifier|false|false||Moderate
null|Moderation|Modifier|false|false||Moderatenull|Uncomplicated|Modifier|false|false||uncomplicatednull|Diverticulitis|Disorder|false|false||diverticulitisnull|Junction Device|Device|false|false||junctionnull|Junctional|Modifier|false|false||junctionnull|Descending colon and sigmoid colon|Anatomy|false|false|C0009373;C0154061;C0496907;C0750873;C0750873;C1547177;C0009373;C0154061;C0496907;C0496863;C0153435;C0496864;C0153436|descending colon and sigmoid colonnull|Malignant neoplasm of descending colon|Disorder|false|false|C0391910;C0227391;C0009368;C4071907;C0545860;C0227389|descending colon
null|Benign neoplasm of descending colon|Disorder|false|false|C0391910;C0227391;C0009368;C4071907;C0545860;C0227389|descending colonnull|Descending colon|Anatomy|false|false|C0750873;C0750873;C0009373;C0154061;C0496907;C0496864;C0153436;C0009373;C0154061;C0496907;C0496863;C0153435|descending colonnull|Sequencing - Descending|Finding|false|false|C0545860;C0391910|descendingnull|Descending|Modifier|false|false||descendingnull|colon and sigmoid colon|Anatomy|false|false|C1547177;C0009373;C0154061;C0496907;C0750873;C0496864;C0153436;C0009373;C0154061;C0496907;C0496863;C0153435;C0750873|colon and sigmoid colonnull|Neoplasm of uncertain or unknown behavior of colon|Disorder|false|false|C0009368;C4071907;C0545860;C0391910;C0227389;C0227391;C0227391|colon
null|Colonic Diseases|Disorder|false|false|C0009368;C4071907;C0545860;C0391910;C0227389;C0227391;C0227391|colon
null|Carcinoma in situ of colon|Disorder|false|false|C0009368;C4071907;C0545860;C0391910;C0227389;C0227391;C0227391|colonnull|COLON PROBLEM|Finding|false|false|C0391910;C0227391;C0227389;C0009368;C4071907;C0545860|colonnull|Colon structure (body structure)|Anatomy|false|false|C0496864;C0153436;C0009373;C0154061;C0496907;C0009373;C0154061;C0496907;C0750873;C0750873;C0496863;C0153435|colon
null|Abdomen+Pelvis>Colon|Anatomy|false|false|C0496864;C0153436;C0009373;C0154061;C0496907;C0009373;C0154061;C0496907;C0750873;C0750873;C0496863;C0153435|colonnull|TUBE,COLON,22FR,RADIOPAQUE RUBBER B#7370|Device|false|false||colonnull|Colon <Coloninae>|Entity|false|false||colonnull|Malignant neoplasm of sigmoid colon|Disorder|false|false|C0009368;C4071907;C0009368;C4071907;C0227391;C0227391;C0545860;C0227389;C0391910|sigmoid colon
null|Benign neoplasm of sigmoid colon|Disorder|false|false|C0009368;C4071907;C0009368;C4071907;C0227391;C0227391;C0545860;C0227389;C0391910|sigmoid colonnull|Sigmoid colon|Anatomy|false|false|C0750873;C0009373;C0154061;C0496907;C0496863;C0153435;C0496864;C0153436;C0009373;C0154061;C0496907;C0750873|sigmoid colonnull|Sigmoid colon|Anatomy|false|false|C0496864;C0153436;C0009373;C0154061;C0496907;C0750873;C0009373;C0154061;C0496907|sigmoidnull|Neoplasm of uncertain or unknown behavior of colon|Disorder|false|false|C0391910;C0009368;C4071907;C0227391;C0227391;C0009368;C4071907;C0545860;C0227389|colon
null|Colonic Diseases|Disorder|false|false|C0391910;C0009368;C4071907;C0227391;C0227391;C0009368;C4071907;C0545860;C0227389|colon
null|Carcinoma in situ of colon|Disorder|false|false|C0391910;C0009368;C4071907;C0227391;C0227391;C0009368;C4071907;C0545860;C0227389|colonnull|COLON PROBLEM|Finding|false|false|C0391910;C0227389;C0227391;C0009368;C4071907;C0009368;C4071907;C0227391;C0545860|colonnull|Colon structure (body structure)|Anatomy|false|false|C0496864;C0153436;C0750873;C0009373;C0154061;C0496907|colon
null|Abdomen+Pelvis>Colon|Anatomy|false|false|C0496864;C0153436;C0750873;C0009373;C0154061;C0496907|colonnull|TUBE,COLON,22FR,RADIOPAQUE RUBBER B#7370|Device|false|false||colonnull|Colon <Coloninae>|Entity|false|false||colonnull|Patient Condition Code - Stable|Finding|false|false||Stablenull|Stable status|Modifier|false|false||Stablenull|Mildly enlarged|Finding|false|false|C0035359;C0024204|mildly enlargednull|MILDLY|Modifier|false|false||mildly
null|Mild (qualifier value)|Modifier|false|false||mildlynull|Enlargement procedure|Procedure|false|false|C0035359;C0024204|enlargednull|Enlarged|Modifier|false|false||enlargednull|Retroperitoneal Space|Anatomy|false|false|C0024202;C0154054;C1293134;C5425894|retroperitonealnull|benign neoplasm of lymph nodes|Disorder|false|false|C0035359;C0024204|lymph nodesnull|lymph nodes|Anatomy|false|false|C4722408;C0024202;C1293134;C0154054;C5425894|lymph nodesnull|Lymph|Finding|false|false|C0024204;C0035359|lymphnull|Reactive Therapy|Procedure|false|false|C0024204|reactivenull|Reactive|Modifier|false|false||reactivenull|Nature|Finding|false|false||nature
null|Natures|Finding|false|false||naturenull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|follow-up|Procedure|false|false||followupnull|week|Time|false|false||weeksnull|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||completenull|Completion Status for valid values - Complete|Finding|false|false||complete
null|Data operation - complete|Finding|false|false||complete
null|Finish - dosing instruction imperative|Finding|false|false||completenull|Complete|Modifier|false|false||completenull|physiologic resolution|Finding|false|false||resolution
null|Resolution|Finding|false|false||resolutionnull|Resolution Property|LabModifier|false|false||resolutionnull|findings aspects|Finding|false|false||findingsnull|null|Attribute|false|false||findingsnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0851353;C0005768;C0229664;C0005767|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C0014792;C1114281|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0851353;C0005768;C0229664;C0005767|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C0014792;C1114281|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0005768;C0229664;C0005767;C0851353|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C1114281;C0014792|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Alanine Transaminase|Drug|false|false||ALT
null|Alanine Transaminase|Drug|false|false||ALTnull|Liposarcoma, well differentiated|Disorder|false|false||ALT
null|Atypical Lipoma|Disorder|false|false||ALTnull|null|Finding|false|false||ALT
null|Alternative Billing Concepts|Finding|false|false||ALT
null|GPT gene|Finding|false|false||ALTnull|Antibiotic Lock Therapy|Procedure|false|false||ALTnull|Southern Altai Language|Entity|false|false||ALTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false|C1185650|AST
null|Aspartate Transaminase|Drug|false|false|C1185650|AST
null|Aspartate Transaminase|Drug|false|false|C1185650|AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false|C1185650|AST
null|SLC17A5 protein, human|Drug|false|false|C1185650|AST
null|SLC17A5 protein, human|Drug|false|false|C1185650|ASTnull|Atypical Spitz Nevus|Disorder|false|false|C1185650|ASTnull|SLC17A5 wt Allele|Finding|false|false|C1185650|AST
null|SLC17A5 gene|Finding|false|false|C1185650|AST
null|GOT1 gene|Finding|false|false|C1185650|ASTnull|Asterion|Anatomy|false|false|C1415181;C1420113;C5960784;C0004002;C0242192;C1121182;C4522245|ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|Lactate Dehydrogenase|Drug|false|false||LDH
null|Lactate Dehydrogenase|Drug|false|false||LDHnull|Lifetime Drinking History|Finding|false|false||LDHnull|Lactate dehydrogenase measurement|Procedure|false|false||LDHnull|Alkaline Phosphatase|Drug|false|false||AlkPhos
null|Alkaline Phosphatase|Drug|false|false||AlkPhosnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Alanine Transaminase|Drug|false|false||ALT
null|Alanine Transaminase|Drug|false|false||ALTnull|Liposarcoma, well differentiated|Disorder|false|false|C1185650|ALT
null|Atypical Lipoma|Disorder|false|false|C1185650|ALTnull|null|Finding|false|false|C1185650|ALT
null|Alternative Billing Concepts|Finding|false|false|C1185650|ALT
null|GPT gene|Finding|false|false|C1185650|ALTnull|Antibiotic Lock Therapy|Procedure|false|false|C1185650|ALTnull|Southern Altai Language|Entity|false|false||ALTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false|C1185650|AST
null|Aspartate Transaminase|Drug|false|false|C1185650|AST
null|Aspartate Transaminase|Drug|false|false|C1185650|AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false|C1185650|AST
null|SLC17A5 protein, human|Drug|false|false|C1185650|AST
null|SLC17A5 protein, human|Drug|false|false|C1185650|ASTnull|Atypical Spitz Nevus|Disorder|false|false|C1185650|ASTnull|SLC17A5 wt Allele|Finding|false|false|C1185650|AST
null|SLC17A5 gene|Finding|false|false|C1185650|AST
null|GOT1 gene|Finding|false|false|C1185650|ASTnull|Asterion|Anatomy|false|false|C1266129;C1370889;C4522245;C0202113;C4553172;C0851148;C0004002;C0242192;C1121182;C1415181;C1420113;C5960784;C2257651;C1415274;C1140170|ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|Lactate Dehydrogenase|Drug|false|false||LDH
null|Lactate Dehydrogenase|Drug|false|false||LDHnull|Lifetime Drinking History|Finding|false|false|C1185650|LDHnull|Lactate dehydrogenase measurement|Procedure|false|false|C1185650|LDHnull|Alkaline Phosphatase|Drug|false|false||AlkPhos
null|Alkaline Phosphatase|Drug|false|false||AlkPhosnull|amylase|Drug|false|false||Amylase
null|amylase|Drug|false|false||Amylase
null|amylase|Drug|false|false||Amylasenull|Amylase measurement|Procedure|false|false||Amylasenull|Blood albumin|Procedure|false|false||BLOOD Albuminnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Albumin|Drug|false|false||Albumin
null|Albumins|Drug|false|false||Albumin
null|Albumins|Drug|false|false||Albumin
null|Albumin|Drug|false|false||Albuminnull|Albumin metabolic function|Finding|false|false||Albumin
null|ALB gene|Finding|false|false||Albuminnull|Albumin measurement|Procedure|false|false||Albuminnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Blood albumin|Procedure|false|false||BLOOD Albuminnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Albumin|Drug|false|false||Albumin
null|Albumins|Drug|false|false||Albumin
null|Albumins|Drug|false|false||Albumin
null|Albumin|Drug|false|false||Albuminnull|Albumin metabolic function|Finding|false|false||Albumin
null|ALB gene|Finding|false|false||Albuminnull|Albumin measurement|Procedure|false|false||Albuminnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|vancomycin|Drug|false|false||Vanco
null|vancomycin|Drug|false|false||Vanconull|Swab Dosage Form|Drug|false|false||SWAB
null|Swab specimen|Drug|false|false||SWABnull|Taking of swab|Procedure|false|false|C1515974|SWABnull|Swab|Device|false|false||SWABnull|Swab Dosing Unit|LabModifier|false|false||SWABnull|null|Finding|false|false|C1515974|Sitenull|Anatomic Site|Anatomy|false|false|C0563454;C1546778|Sitenull|Study Site|Modifier|false|false||Site
null|Site|Modifier|false|false||Sitenull|Malignant neoplasm of abdomen|Disorder|false|false|C0230168;C0000726|ABDOMENnull|Abdomen problem|Finding|false|false|C0230168;C0000726|ABDOMENnull|Abdomen|Anatomy|false|false|C0941288;C0153662|ABDOMEN
null|Abdominal Cavity|Anatomy|false|false|C0941288;C0153662|ABDOMENnull|fluid - substance|Drug|false|false||Fluid
null|Liquid substance|Drug|false|false||Fluidnull|Fluid Specimen Code|Finding|false|false||Fluidnull|Fluid behavior|Modifier|false|false||Fluidnull|Swab Dosage Form|Drug|false|false||swab
null|Swab specimen|Drug|false|false||swabnull|Taking of swab|Procedure|false|false|C1254021;C0162867|swabnull|Swab|Device|false|false||swabnull|Swab Dosing Unit|LabModifier|false|false||swabnull|Transport Media,|Procedure|false|false|C1254021;C0162867|transport medianull|Biological Transport|Finding|false|false|C1254021;C0162867|transport
null|Transfer Technique|Finding|false|false|C1254021;C0162867|transport
null|Molecular Transport|Finding|false|false|C1254021;C0162867|transportnull|Transport Device|Device|false|false||transport
null|Mobility aid|Device|false|false||transportnull|Communications Media|Finding|false|false|C1254021;C0162867|media
null|PAMS Media|Finding|false|false|C1254021;C0162867|medianull|Tunica Media|Anatomy|false|false|C1519628;C0005528;C1705822;C1548752;C0563454;C0677540;C0009458|media
null|Media layer|Anatomy|false|false|C1519628;C0005528;C1705822;C1548752;C0563454;C0677540;C0009458|medianull|Liquid substance|Drug|false|false||fluidsnull|Mouse Body Fluid or Substance|Finding|false|false||fluidsnull|Fluid Therapy|Procedure|false|false||fluidsnull|Syringes|Device|false|false||syringenull|Syringe (unit of presentation)|LabModifier|false|false||syringe
null|Syringe Dosing Unit|LabModifier|false|false||syringenull|null|Finding|true|false||needlenull|Needle device|Device|true|false||needlenull|Needle Shape|Modifier|false|false||needlenull|Serum Collection Tube|Device|false|false||red top tubenull|DYRK3 gene|Finding|false|false||red
null|Redness|Finding|false|false||red
null|IK gene|Finding|false|false||rednull|Radiological Exposure Device|Device|false|false||rednull|Red color|Modifier|false|false||rednull|Unspecified tube|Finding|false|false||tube
null|TUBE1 gene|Finding|false|false||tubenull|biomedical tube device|Device|false|false||tube
null|Packaging Tube|Device|false|false||tubenull|tube|Modifier|false|false||tubenull|Tube (unit of presentation)|LabModifier|false|false||tube
null|Tube Dosing Unit|LabModifier|false|false||tubenull|Sterility, Reproductive|Finding|false|false||sterile
null|Infertility|Finding|false|false||sterilenull|Sterile (qualifier value)|Modifier|false|false||sterilenull|Carcinoma of unknown primary|Disorder|false|false||cupnull|Cup (physical object)|Device|false|false||cup
null|Cup Device|Device|false|false||cupnull|Cup (unit of presentation)|LabModifier|false|false||cup
null|Cup Dosing Unit|LabModifier|false|false||cupnull|Gram's stain|Drug|false|false||GRAM STAIN
null|Gram's stain|Drug|false|false||GRAM STAINnull|Bacterial stain, routine|Procedure|false|false||GRAM STAINnull|gram|LabModifier|false|false||GRAMnull|Stains|Drug|false|false||STAINnull|Staining method|Procedure|false|false||STAINnull|Diagnosis Type - Final|Finding|false|false||Finalnull|Final|Time|false|false||Finalnull|End-stage|Modifier|false|false||Finalnull|Knowledge Field|Finding|false|false||FIELD
null|Force Field|Finding|false|false||FIELD
null|Field|Finding|false|false||FIELDnull|field - patient encounter|Procedure|false|false||FIELDnull|Specimen Type - Leukocytes|Finding|false|false|C0023516|LEUKOCYTES
null|null|Finding|false|false|C0023516|LEUKOCYTESnull|Leukocytes|Anatomy|false|false|C1550647;C1547962|LEUKOCYTESnull|Knowledge Field|Finding|false|false||FIELD
null|Force Field|Finding|false|false||FIELD
null|Field|Finding|false|false||FIELDnull|field - patient encounter|Procedure|false|false||FIELDnull|Gram-Positive Cocci|Entity|false|false||GRAM POSITIVE COCCInull|gram|LabModifier|false|false||GRAMnull|BRAF Gene Rearrangement|Disorder|false|false||POSITIVEnull|Rh Positive Blood Group|Finding|false|false||POSITIVE
null|Positive Finding|Finding|false|false||POSITIVE
null|Positive|Finding|false|false||POSITIVEnull|Positive Charge|Modifier|false|false||POSITIVEnull|Positive Number|LabModifier|false|false||POSITIVEnull|Cocci bacteria|Entity|false|false||COCCInull|Chain device|Device|false|false||CHAINSnull|fluid - substance|Drug|false|false||FLUID
null|Liquid substance|Drug|false|false||FLUIDnull|Fluid Specimen Code|Finding|false|false||FLUIDnull|Fluid behavior|Modifier|false|false||FLUIDnull|Culture Dose Form|Drug|false|false||CULTUREnull|Culture (Anthropological)|Finding|false|false||CULTURE
null|Cultural aspects|Finding|false|false||CULTUREnull|Microbial culture (procedure)|Procedure|false|false||CULTURE
null|Laboratory culture|Procedure|false|false||CULTUREnull|Diagnosis Type - Final|Finding|false|false||Finalnull|Final|Time|false|false||Finalnull|End-stage|Modifier|false|false||Finalnull|Staphylococcus aureus|Entity|false|false||STAPH AUREUSnull|Staphylococcal Infections|Disorder|false|false||STAPHnull|Genus staphylococcus|Entity|false|false||STAPHnull|Blood coagulation tests|Procedure|false|false||COAGnull|Moderate growth|Modifier|false|false||MODERATE GROWTHnull|Moderate - Severity of Illness Code|Finding|false|false||MODERATE
null|Moderate|Finding|false|false||MODERATEnull|Moderate (severity modifier)|Modifier|false|false||MODERATE
null|Moderate - Allergy Severity|Modifier|false|false||MODERATE
null|Moderation|Modifier|false|false||MODERATEnull|Growth & development aspects|Finding|false|false||GROWTH
null|Tissue Growth|Finding|false|false||GROWTH
null|Growth|Finding|false|false||GROWTH
null|growth aspects|Finding|false|false||GROWTHnull|Growth action|Phenomenon|false|false||GROWTHnull|clindamycin|Drug|false|false|C0449201|CLINDAMYCIN
null|clindamycin|Drug|false|false|C0449201|CLINDAMYCINnull|PROGRESSIVE ENCEPHALOMYELITIS WITH RIGIDITY|Disorder|false|false|C0449201|PERnull|Per - dosing instruction fragment|Finding|false|false|C0449201|PER
null|PER1 gene|Finding|false|false|C0449201|PER
null|Follow|Finding|false|false|C0449201|PER
null|PER1 wt Allele|Finding|false|false|C0449201|PERnull|PER (body structure)|Anatomy|false|false|C0008947;C1861457;C3273590;C4281991;C1418464;C1704764|PERnull|Per (qualifier)|Modifier|false|false||PERnull|Isolate - microorganism|Drug|false|false||isolate
null|ISOLATE COMPOUND|Drug|false|false||isolatenull|Resistant (qualifier value)|Finding|false|false||resistant tonull|resistant - Observation Interpretation Susceptibility|Finding|false|false||resistant
null|Resistant (qualifier value)|Finding|false|false||resistantnull|Antimicrobial Resistance Result|Lab|false|false||resistantnull|clindamycin|Drug|false|false||clindamycin
null|clindamycin|Drug|false|false||clindamycinnull|Detection|Procedure|false|false||detectionnull|Induce (action)|Finding|false|false||induciblenull|Resistance (Psychotherapeutic)|Finding|false|false||resistance
null|social resistance|Finding|false|false||resistance
null|Resistance Process|Finding|false|false||resistancenull|Resistance|Attribute|false|false||resistancenull|Anaerobic microbial culture|Procedure|false|false||ANAEROBIC CULTUREnull|Anaerobic|Modifier|false|false||ANAEROBICnull|Culture Dose Form|Drug|false|false||CULTUREnull|Culture (Anthropological)|Finding|false|false||CULTURE
null|Cultural aspects|Finding|false|false||CULTUREnull|Microbial culture (procedure)|Procedure|false|false||CULTURE
null|Laboratory culture|Procedure|false|false||CULTUREnull|Preliminary|Time|false|false||Preliminarynull|Bacteria, Anaerobic|Entity|true|false||ANAEROBESnull|Acid fast stain|Drug|false|false||ACID FASTnull|Fas-activated serine/threonine kinase activity|Finding|false|false||FAST
null|FASTK Gene|Finding|false|false||FAST
null|FOXD3-AS1 gene|Finding|false|false||FAST
null|FASTK wt Allele|Finding|false|false||FAST
null|Fasting|Finding|false|false||FASTnull|Rapid|Modifier|false|false||FASTnull|Smearing technique|Finding|false|false||SMEARnull|Smear test|Procedure|false|false||SMEARnull|Smear - instruction imperative|Event|false|false||SMEARnull|Diagnosis Type - Final|Finding|false|false||Finalnull|Final|Time|false|false||Finalnull|End-stage|Modifier|false|false||Finalnull|Acid fast stain|Drug|true|false||ACID FASTnull|Fas-activated serine/threonine kinase activity|Finding|true|false||FAST
null|FASTK Gene|Finding|true|false||FAST
null|FOXD3-AS1 gene|Finding|true|false||FAST
null|FASTK wt Allele|Finding|true|false||FAST
null|Fasting|Finding|true|false||FASTnull|Rapid|Modifier|false|false||FASTnull|Bacilli <Bacillota>|Entity|true|false||BACILLI
null|Genus Bacillus|Entity|true|false||BACILLInull|Direct - PostalAddressUse|Finding|false|false||DIRECT
null|direct address|Finding|false|false||DIRECTnull|Direct type of relationship|Modifier|false|false||DIRECT
null|Direct (qualifier)|Modifier|false|false||DIRECTnull|Smearing technique|Finding|false|false||SMEARnull|Smear test|Procedure|false|false||SMEARnull|Smear - instruction imperative|Event|false|false||SMEARnull|Acid fast stain|Drug|false|false||ACID FASTnull|Fas-activated serine/threonine kinase activity|Finding|false|false||FAST
null|FASTK Gene|Finding|false|false||FAST
null|FOXD3-AS1 gene|Finding|false|false||FAST
null|FASTK wt Allele|Finding|false|false||FAST
null|Fasting|Finding|false|false||FASTnull|Rapid|Modifier|false|false||FASTnull|Culture Dose Form|Drug|false|false||CULTUREnull|Culture (Anthropological)|Finding|false|false||CULTURE
null|Cultural aspects|Finding|false|false||CULTUREnull|Microbial culture (procedure)|Procedure|false|false||CULTURE
null|Laboratory culture|Procedure|false|false||CULTUREnull|Preliminary|Time|false|false||Preliminarynull|Swab specimen|Drug|false|false||swab
null|Swab Dosage Form|Drug|false|false||swabnull|Taking of swab|Procedure|false|false||swabnull|Swab|Device|false|false||swabnull|Swab Dosing Unit|LabModifier|false|false||swabnull|Outpatient Physical Therapy Improvement in Movement and Assessment Log (OPTIMAL) Survey|Finding|false|false||optimalnull|Optimum|Modifier|false|false||optimalnull|Specimen|Drug|false|false||specimennull|Role Class - specimen|Finding|false|false||specimen
null|Biospecimen|Finding|false|false||specimennull|Recovery - healing process|Finding|false|false||recoverynull|null|Event|false|false||recoverynull|recovery - adjustment|LabModifier|false|false||recoverynull|Genus Mycobacterium|Entity|false|false||mycobacterianull|Filamentous fungus|Entity|false|false||filamentous funginull|Fungal|Finding|false|false||funginull|Fungi|Entity|false|false||funginull|Negative Results|Finding|false|false||negative resultnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|What subject filter - Result|Finding|false|false||result
null|Result|Finding|false|false||result
null|Experimental Result|Finding|false|false||resultnull|Possible|Finding|false|false||possiblenull|Possible diagnosis|Modifier|false|false||possible
null|Possibly Related to Intervention|Modifier|false|false||possiblenull|Tissue Specimen Code|Finding|false|false|C0040300|tissuenull|Body tissue|Anatomy|false|false|C1547928|tissuenull|biopsy characteristics|Finding|false|false||biopsy
null|null|Finding|false|false||biopsynull|Biopsy Procedures on the Pharynx, Adenoids, and Tonsils|Procedure|false|false||biopsy
null|Biopsy|Procedure|false|false||biopsy
null|Consent Type - biopsy|Procedure|false|false||biopsynull|Respiratory Aspiration|Disorder|false|false||aspiratednull|Pulmonary aspiration|Finding|false|false||aspiratednull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Mycology culture|Procedure|false|false||FUNGAL CULTUREnull|Fungal|Finding|false|false||FUNGALnull|Fungi|Entity|false|false||FUNGALnull|Culture Dose Form|Drug|false|false||CULTUREnull|Culture (Anthropological)|Finding|false|false||CULTURE
null|Cultural aspects|Finding|false|false||CULTUREnull|Microbial culture (procedure)|Procedure|false|false||CULTURE
null|Laboratory culture|Procedure|false|false||CULTUREnull|Preliminary|Time|false|false||Preliminarynull|Specimen fungus isolated|Lab|false|false||FUNGUS ISOLATEDnull|Fungus Present|Lab|true|false||FUNGUSnull|Fungi|Entity|true|false||FUNGUSnull|Swab specimen|Drug|false|false||swab
null|Swab Dosage Form|Drug|false|false||swabnull|Taking of swab|Procedure|false|false||swabnull|Swab|Device|false|false||swabnull|Swab Dosing Unit|LabModifier|false|false||swabnull|Outpatient Physical Therapy Improvement in Movement and Assessment Log (OPTIMAL) Survey|Finding|false|false||optimalnull|Optimum|Modifier|false|false||optimalnull|Specimen|Drug|false|false||specimennull|Role Class - specimen|Finding|false|false||specimen
null|Biospecimen|Finding|false|false||specimennull|Recovery - healing process|Finding|false|false||recoverynull|null|Event|false|false||recoverynull|recovery - adjustment|LabModifier|false|false||recoverynull|Genus Mycobacterium|Entity|false|false||mycobacterianull|Filamentous fungus|Entity|false|false||filamentous funginull|Fungal|Finding|false|false||funginull|Fungi|Entity|false|false||funginull|Negative Results|Finding|false|false||negative resultnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|What subject filter - Result|Finding|false|false||result
null|Result|Finding|false|false||result
null|Experimental Result|Finding|false|false||resultnull|Possible|Finding|false|false||possiblenull|Possible diagnosis|Modifier|false|false||possible
null|Possibly Related to Intervention|Modifier|false|false||possiblenull|Tissue Specimen Code|Finding|false|false|C0040300|tissuenull|Body tissue|Anatomy|false|false|C1547928|tissuenull|biopsy characteristics|Finding|false|false||biopsy
null|null|Finding|false|false||biopsynull|Biopsy Procedures on the Pharynx, Adenoids, and Tonsils|Procedure|false|false||biopsy
null|Biopsy|Procedure|false|false||biopsy
null|Consent Type - biopsy|Procedure|false|false||biopsynull|Respiratory Aspiration|Disorder|false|false||aspiratednull|Pulmonary aspiration|Finding|false|false||aspiratednull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Pathologic Examination|Procedure|false|false||Pathology Examinationnull|Pathology processes|Finding|false|false||Pathology
null|Pathological aspects|Finding|false|false||Pathologynull|Pathology procedure|Procedure|false|false||Pathologynull|Pathology|Title|false|false||Pathologynull|Physical Examination|Procedure|false|false||Examination
null|Medical Examination|Procedure|false|false||Examinationnull|Examination|Event|false|false||Examinationnull|Specimen|Drug|false|false||SPECIMENnull|Role Class - specimen|Finding|false|false||SPECIMEN
null|Biospecimen|Finding|false|false||SPECIMENnull|Malignant neoplasm of sigmoid colon|Disorder|false|false|C0227391;C0009368;C4071907;C0227391|sigmoid colon
null|Benign neoplasm of sigmoid colon|Disorder|false|false|C0227391;C0009368;C4071907;C0227391|sigmoid colonnull|Sigmoid colon|Anatomy|false|false|C0496864;C0153436;C0009373;C0154061;C0496907;C0750873|sigmoid colonnull|Sigmoid colon|Anatomy|false|false|C0009373;C0154061;C0496907;C0496864;C0153436|sigmoidnull|Neoplasm of uncertain or unknown behavior of colon|Disorder|false|false|C0009368;C4071907;C0227391;C0227391|colon
null|Colonic Diseases|Disorder|false|false|C0009368;C4071907;C0227391;C0227391|colon
null|Carcinoma in situ of colon|Disorder|false|false|C0009368;C4071907;C0227391;C0227391|colonnull|COLON PROBLEM|Finding|false|false|C0227391;C0009368;C4071907|colonnull|Colon structure (body structure)|Anatomy|false|false|C0009373;C0154061;C0496907;C0496864;C0153436;C0750873|colon
null|Abdomen+Pelvis>Colon|Anatomy|false|false|C0009373;C0154061;C0496907;C0496864;C0153436;C0750873|colonnull|TUBE,COLON,22FR,RADIOPAQUE RUBBER B#7370|Device|false|false||colonnull|Colon <Coloninae>|Entity|false|false||colonnull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Malignant neoplasm of sigmoid colon|Disorder|false|false|C0227391;C0009368;C4071907;C0227391|Sigmoid colon
null|Benign neoplasm of sigmoid colon|Disorder|false|false|C0227391;C0009368;C4071907;C0227391|Sigmoid colonnull|Sigmoid colon|Anatomy|false|false|C0750873;C0009373;C0154061;C0496907;C0496864;C0153436;C0015252;C0728940|Sigmoid colonnull|Sigmoid colon|Anatomy|false|false|C0009373;C0154061;C0496907;C0750873;C0496864;C0153436|Sigmoidnull|Neoplasm of uncertain or unknown behavior of colon|Disorder|false|false|C0227391;C0227391;C0009368;C4071907|colon
null|Colonic Diseases|Disorder|false|false|C0227391;C0227391;C0009368;C4071907|colon
null|Carcinoma in situ of colon|Disorder|false|false|C0227391;C0227391;C0009368;C4071907|colonnull|COLON PROBLEM|Finding|false|false|C0227391;C0009368;C4071907;C0227391|colonnull|Colon structure (body structure)|Anatomy|false|false|C0750873;C0496864;C0153436;C0009373;C0154061;C0496907|colon
null|Abdomen+Pelvis>Colon|Anatomy|false|false|C0750873;C0496864;C0153436;C0009373;C0154061;C0496907|colonnull|TUBE,COLON,22FR,RADIOPAQUE RUBBER B#7370|Device|false|false||colonnull|Colon <Coloninae>|Entity|false|false||colonnull|Segmental|Modifier|false|false||segmentalnull|removal technique|Procedure|false|false|C0227391|resection
null|Excision|Procedure|false|false|C0227391|resectionnull|Colon structure (body structure)|Anatomy|false|false|C1300196;C0000833|Colonicnull|Anatomical segmentation|Modifier|false|false||segmentnull|Organized|Finding|false|false|C0009368|organizingnull|Paracolic abscess|Disorder|false|false||pericolic abscessnull|Paracolic|Modifier|false|false||pericolicnull|Abscess|Disorder|false|false|C0009368|abscessnull|null|Finding|false|false||abscessnull|Consistent with|Finding|false|false||consistentnull|Perforated diverticulum|Disorder|false|false||ruptured diverticulumnull|Diverticulum|Disorder|false|false||diverticulumnull|null|Finding|false|false||diverticulumnull|null|Modifier|false|false||Unremarkablenull|Set of regional lymph nodes|Anatomy|false|false|C0154054;C0024202|regional lymph nodesnull|regional|Modifier|false|false||regional
null|Local|Modifier|false|false||regionalnull|benign neoplasm of lymph nodes|Disorder|false|false|C1184738;C0024204|lymph nodesnull|lymph nodes|Anatomy|false|false|C0024202;C0154054|lymph nodesnull|Lymph|Finding|false|false|C0024204;C1184738|lymphnull|Intrinsic origin|Finding|true|false|C0026724|intrinsicnull|Internal|Modifier|false|false||intrinsicnull|Mucous Membrane|Anatomy|false|false|C0000769;C0000768;C0439674|mucosalnull|Congenital Abnormality|Disorder|true|false|C0026724|abnormalitiesnull|teratologic|Finding|true|false|C0026724|abnormalitiesnull|Clinical NEC (not elsewhere classified in LNC)|Finding|false|false||Clinicalnull|Clinical|Modifier|false|false||Clinicalnull|Diverticulitis|Disorder|false|false||Diverticulitisnull|radiology referral type|Finding|false|false||RADIOLOGY
null|Radiology Section ID|Finding|false|false||RADIOLOGY
null|Encounter due to radiological examination|Finding|false|false||RADIOLOGYnull|Radiology studies|Procedure|false|false||RADIOLOGY
null|Diagnostic radiologic examination|Procedure|false|false||RADIOLOGY
null|Radiographic imaging procedure|Procedure|false|false||RADIOLOGYnull|Radiology Specialty|Title|false|false||RADIOLOGYnull|Final report|Finding|false|false||Final Reportnull|Diagnosis Type - Final|Finding|false|false||Finalnull|Final|Time|false|false||Finalnull|End-stage|Modifier|false|false||Finalnull|Report (document)|Finding|false|false||Reportnull|Reporting|Procedure|false|false||Reportnull|null|Attribute|false|false||Reportnull|CT of abdomen with contrast|Procedure|false|false|C0230168;C0000726|CT ABDOMEN W/CONTRASTnull|CT of abdomen|Procedure|false|false|C0230168;C0000726|CT ABDOMENnull|null|Attribute|false|false|C0230168;C0000726|CT ABDOMENnull|Malignant neoplasm of abdomen|Disorder|false|false|C0230168;C0000726|ABDOMENnull|Abdomen problem|Finding|false|false|C0230168;C0000726|ABDOMENnull|Abdomen|Anatomy|false|false|C0412620;C0153662;C0202840;C1644645;C0941288|ABDOMEN
null|Abdominal Cavity|Anatomy|false|false|C0412620;C0153662;C0202840;C1644645;C0941288|ABDOMENnull|Contrast Media|Drug|false|false||CONTRASTnull|Contrast|Modifier|false|false||CONTRASTnull|Indication of (contextual qualifier)|Finding|false|false||Reasonnull|Subcutaneous air|Finding|false|false||subcutaneous airnull|Subcutaneous Route of Administration|Finding|false|false||subcutaneousnull|subcutaneous|Modifier|false|false||subcutaneousnull|Air (substance)|Drug|false|false||air
null|air|Drug|false|false||air
null|air|Drug|false|false||airnull|ACUTE INSULIN RESPONSE|Finding|false|false||air
null|AIRN gene|Finding|false|false||air
null|AI/RHEUM|Finding|false|false||airnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|IV contrast|Drug|false|false||IV contrastnull|Contrast Media|Drug|false|false||contrastnull|Contrast|Modifier|false|false||contrastnull|History of present illness (finding)|Finding|false|false||HISTORY
null|History of previous events|Finding|false|false||HISTORY
null|Historical aspects qualifier|Finding|false|false||HISTORY
null|Medical History|Finding|false|false||HISTORY
null|Concept History|Finding|false|false||HISTORYnull|History|Subject|false|false||HISTORYnull|Females|Subject|false|false||female
null|Woman|Subject|false|false||femalenull|Female, Self-Report|Modifier|false|false||female
null|Female Phenotype|Modifier|false|false||femalenull|Recurrent|Time|false|false||recurrent
null|Episodic|Time|false|false||recurrentnull|Diverticulitis|Disorder|false|false||diverticulitisnull|Status post|Time|false|false||status post
null|Post|Time|false|false||status postnull|What subject filter - Status|Finding|false|false||statusnull|null|Attribute|false|false||statusnull|Social status|Modifier|false|false||status
null|Status|Modifier|false|false||statusnull|Laparoscopic-assisted sigmoid colectomy|Procedure|false|false|C0227391|laparoscopic sigmoid colectomy
null|Laparoscopic sigmoid colectomy|Procedure|false|false|C0227391|laparoscopic sigmoid colectomynull|Laparoscopy|Procedure|false|false||laparoscopicnull|Laparoscopic approach|Modifier|false|false||laparoscopicnull|Sigmoid colectomy|Procedure|false|false|C0227391|sigmoid colectomynull|Sigmoid colon|Anatomy|false|false|C0192866;C0585462;C5890124|sigmoidnull|Colectomy|Procedure|false|false||colectomynull|Surgical incisions|Procedure|false|false||incisionalnull|Erythema|Disorder|false|false||erythemanull|Subcutaneous air|Finding|false|false||subcutaneous airnull|Subcutaneous Route of Administration|Finding|false|false||subcutaneousnull|subcutaneous|Modifier|false|false||subcutaneousnull|Air (substance)|Drug|false|false||air
null|air|Drug|false|false||air
null|air|Drug|false|false||airnull|ACUTE INSULIN RESPONSE|Finding|false|false||air
null|AIRN gene|Finding|false|false||air
null|AI/RHEUM|Finding|false|false||airnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Status post|Time|false|false||Status post
null|Post|Time|false|false||Status postnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Sigmoid colectomy|Procedure|false|false|C0227391|sigmoid colectomynull|Sigmoid colon|Anatomy|false|false|C0192866|sigmoidnull|Colectomy|Procedure|false|false||colectomynull|Small amount|LabModifier|false|false||small amountnull|Small|LabModifier|false|false||smallnull|Amount class - Amount|Finding|false|false||amountnull|Quantity|LabModifier|false|false||amountnull|Postoperative Period|Time|false|false||post-operativenull|Free of (attribute)|Finding|false|false||freenull|Empty (qualifier)|Modifier|false|false||freenull|Intraperitoneal Route of Administration|Finding|false|false||intraperitoneal
null|Intraperitoneal (intended site)|Finding|false|false||intraperitonealnull|Intraperitoneal|Modifier|false|false||intraperitonealnull|Air (substance)|Drug|false|false||air
null|air|Drug|false|false||air
null|air|Drug|false|false||airnull|ACUTE INSULIN RESPONSE|Finding|false|false||air
null|AIRN gene|Finding|false|false||air
null|AI/RHEUM|Finding|false|false||airnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Malignant neoplasm of pelvis|Disorder|false|false|C4266535;C0030797;C0559769|pelvisnull|Pelvis problem|Finding|false|false|C4266535;C0030797;C0559769|pelvisnull|Pelvis+|Anatomy|false|false|C0812455;C0153663|pelvis
null|Pelvic cavity structure|Anatomy|false|false|C0812455;C0153663|pelvis
null|Pelvis|Anatomy|false|false|C0812455;C0153663|pelvisnull|Small amount|LabModifier|false|false||Small amountnull|Small|LabModifier|false|false||Smallnull|Amount class - Amount|Finding|false|false||amountnull|Quantity|LabModifier|false|false||amountnull|Scattered|Modifier|false|false||scatterednull|Subcutaneous air|Finding|false|false||subcutaneous airnull|Subcutaneous Route of Administration|Finding|false|false||subcutaneousnull|subcutaneous|Modifier|false|false||subcutaneousnull|Air (substance)|Drug|false|false||air
null|air|Drug|false|false||air
null|air|Drug|false|false||airnull|ACUTE INSULIN RESPONSE|Finding|false|false||air
null|AIRN gene|Finding|false|false||air
null|AI/RHEUM|Finding|false|false||airnull|Middle|Modifier|false|false||midnull|Lower anterior abdominal wall|Anatomy|false|false|C2003888;C0332290;C0751437;C0332290|lower anterior abdominal wallnull|Lower anterior|Modifier|false|false||lower anteriornull|Body Site Modifier - Lower|Anatomy|false|false|C2003888|lowernull|Lower (action)|Event|false|false|C2332167;C0230193;C1548802|lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Anterior abdominal wall|Anatomy|false|false|C0332290;C0332290;C2003888;C0751437|anterior abdominal wallnull|Adenohypophyseal Diseases|Disorder|false|false|C2332167;C0836916;C0230193|anteriornull|Anterior|Modifier|false|false||anteriornull|Abdominal wall structure|Anatomy|false|false|C0751437;C0332290|abdominal wallnull|Abdomen|Anatomy|false|false||abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Walls of a building|Device|false|false||wallnull|Consistent with|Finding|false|false|C2332167;C0230193|consistent withnull|Compatible|Modifier|false|false||consistent withnull|Consistent with|Finding|false|false|C0230193;C2332167;C0836916|consistentnull|Changing|Finding|false|false||changenull|Change - procedure|Procedure|false|false||changenull|Delta (difference)|LabModifier|false|false||change
null|Changed status|LabModifier|false|false||changenull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Separate|Modifier|false|false||discretenull|fluid - substance|Drug|true|false||fluid
null|Liquid substance|Drug|true|false||fluidnull|Fluid Specimen Code|Finding|true|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Collection Object - UML Entity|Finding|false|false||collection
null|Item Collection|Finding|false|false||collection
null|Collections (publication)|Finding|false|false||collection
null|Collection (action)|Finding|false|false||collectionnull|Direct (qualifier)|Modifier|false|false||directlynull|Address type - Office|Finding|false|false||officenull|Office|Device|false|false||officenull|Organization unit type - Office|Entity|false|false||officenull|Persistent|Time|false|false||persistentnull|Abdominal Pain|Finding|false|false|C0000726|abdominal painnull|Abdomen|Anatomy|false|false|C1549543;C0030193;C0000737|abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Administration Method - Pain|Finding|false|false|C0000726|pain
null|Pain|Finding|false|false|C0000726|painnull|null|Attribute|false|false||painnull|Adverse Event Probably Related to Intervention|Modifier|false|false||likely relatednull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Relate - vinyl resin|Drug|false|false||relatednull|Role Link Type - related|Finding|false|false||related
null|Related (finding)|Finding|false|false||relatednull|Definitely Related to Intervention|Modifier|false|false||related
null|Relationships|Modifier|false|false||relatednull|Diverticulitis|Disorder|false|false||diverticulitisnull|Flare|Finding|false|false||flare
null|Exacerbation of cGVHD|Finding|false|false||flarenull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Slightly (qualifier value)|Modifier|false|false||slightly
null|Slight (qualifier value)|Modifier|false|false||slightlynull|Hematocrit decreased|Finding|false|false||decreased hematocritnull|Hematocrit level|Finding|false|false||hematocritnull|Hematocrit Measurement|Procedure|false|false||hematocritnull|hematocrit attribute|Attribute|false|false||hematocritnull|On IV|Finding|false|false||on IVnull|Cipro|Drug|false|false||Cipro
null|Cipro|Drug|false|false||Cipronull|Flagyl|Drug|false|false||Flagyl
null|Flagyl|Drug|false|false||Flagylnull|NPO - Nothing by mouth|Procedure|false|false||NPOnull|null|Entity|false|false||NPOnull|Ventricular Fibrillation, Paroxysmal Familial, 1|Disorder|false|false|C0016520|IVFnull|SCN5A wt Allele|Finding|false|false|C0016520|IVF
null|SCN5A gene|Finding|false|false|C0016520|IVFnull|Assisted Reproductive Technologies|Procedure|false|false|C0016520|IVF
null|Fertilization in Vitro|Procedure|false|false|C0016520|IVFnull|Structure of interventricular foramen|Anatomy|false|false|C1419864;C4321334;C2751898;C0872104;C0015915|IVFnull|Hydration status|Finding|false|false||hydration
null|Hydration|Finding|false|false||hydrationnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Periodicals|Finding|false|false||serialnull|Serial|Time|false|false||serialnull|Abdomen|Anatomy|false|false||abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|HDAC2 protein, human|Drug|false|false||HD2
null|HDAC2 protein, human|Drug|false|false||HD2null|HDAC2 wt Allele|Finding|false|false||HD2null|HDAC7 protein, human|Drug|false|false||HD7
null|HDAC7 protein, human|Drug|false|false||HD7
null|HDAC9 protein, human|Drug|false|false||HD7
null|HDAC9 protein, human|Drug|false|false||HD7null|HDAC9 wt Allele|Finding|false|false||HD7
null|HDAC9 gene|Finding|false|false||HD7null|Absence of Biallelic TCRgamma Deletion|Disorder|false|false|C0449202;C0000726|abdnull|ABD (body structure)|Anatomy|false|false|C0040405;C3811055|abd
null|Abdomen|Anatomy|false|false|C0040405;C3811055|abdnull|X-Ray Computed Tomography|Procedure|false|false|C0449202;C0000726|CT scannull|Radionuclide Imaging|Procedure|false|false||scan
null|Scanning|Procedure|false|false||scannull|Uncomplicated|Modifier|false|false||uncomplicatednull|Diverticulitis|Disorder|false|false||diverticulitisnull|Table Frame - above|Finding|false|false||abovenull|Upper|Modifier|false|false||abovenull|Biomaterial Treatment|Finding|false|false||treatment
null|Treating|Finding|false|false||treatment
null|therapeutic aspects|Finding|false|false||treatmentnull|treatment - ActInformationManagementReason|Procedure|false|false||treatment
null|Administration (procedure)|Procedure|false|false||treatment
null|Therapeutic procedure|Procedure|false|false||treatmentnull|GDC Regimen Terminology|Finding|false|false||regimennull|Treatment Protocols|Procedure|false|false||regimennull|Abdominal Pain|Finding|false|false|C0000726|abdominal painnull|Abdomen|Anatomy|false|false|C1549543;C0030193;C0000737|abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Administration Method - Pain|Finding|false|false|C0000726|pain
null|Pain|Finding|false|false|C0000726|painnull|null|Attribute|false|false||painnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Dilaudid|Drug|false|false||Dilaudid
null|Dilaudid|Drug|false|false||Dilaudidnull|Numerous|LabModifier|false|false||multiplenull|Feces|Finding|false|false||stoolsnull|null|Attribute|false|false||stoolsnull|Stool seat|Device|false|false||stoolsnull|Ambulate|Finding|false|false||ambulatenull|Has difficulty doing (qualifier value)|Finding|false|false||difficultynull|Refused - Completion Status for valid values|Finding|false|false||refusednull|Refused|Event|false|false||refusednull|Injection Route of Administration|Finding|false|false||injectionsnull|Injection of therapeutic agent|Procedure|false|false||injections
null|Injection procedure|Procedure|false|false||injectionsnull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|treatment options|Finding|false|false||options
null|Options|Finding|false|false||optionsnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Level of Care - Surgery|Finding|false|false||Surgery
null|Surgical procedure finding|Finding|false|false||Surgery
null|Surgical aspects|Finding|false|false||Surgerynull|Operative Surgical Procedures|Procedure|false|false||Surgerynull|General surgery specialty|Title|false|false||Surgery
null|Surgery specialty|Title|false|false||Surgerynull|TAPBP protein, human|Drug|false|false||TPN
null|NADP|Drug|false|false||TPN
null|NADP|Drug|false|false||TPN
null|TAPBP protein, human|Drug|false|false||TPNnull|TAPBP wt Allele|Finding|false|false||TPN
null|TAPBP gene|Finding|false|false||TPNnull|Parenteral Nutrition, Total|Procedure|false|false||TPNnull|Peripherally Inserted Central Catheter Line Insertion|Procedure|false|false||PICCnull|Peripherally inserted central catheter (physical object)|Device|false|false||PICCnull|Ensure (product)|Drug|false|false||Ensurenull|null|Attribute|false|false||Operative consentnull|Operative|Time|false|false||Operativenull|Consent (record artifact)|Finding|false|false||consent
null|ActClass - consent|Finding|false|false||consent
null|Consent|Finding|false|false||consentnull|null|Attribute|false|false||consentnull|Plain chest X-ray|Procedure|false|false||CXRnull|Electrocardiogram image|Finding|false|false||EKG
null|Electrocardiogram|Finding|false|false||EKGnull|Electrocardiography|Procedure|false|false||EKGnull|HDAC8 protein, human|Drug|false|false||HD8
null|HDAC8 protein, human|Drug|false|false||HD8null|HDAC8 wt Allele|Finding|false|false||HD8null|NPO - Nothing by mouth|Procedure|false|false||NPOnull|null|Entity|false|false||NPOnull|Overnight|Time|false|false||overnightnull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Ventricular Fibrillation, Paroxysmal Familial, 1|Disorder|false|false|C0016520|IVFnull|SCN5A wt Allele|Finding|false|false|C0016520|IVF
null|SCN5A gene|Finding|false|false|C0016520|IVFnull|Assisted Reproductive Technologies|Procedure|false|false|C0016520|IVF
null|Fertilization in Vitro|Procedure|false|false|C0016520|IVFnull|Structure of interventricular foramen|Anatomy|false|false|C2751898;C0872104;C0015915;C1419864;C4321334|IVFnull|Level of Care - Surgery|Finding|false|false||Surgery
null|Surgical procedure finding|Finding|false|false||Surgery
null|Surgical aspects|Finding|false|false||Surgerynull|Operative Surgical Procedures|Procedure|false|false||Surgerynull|General surgery specialty|Title|false|false||Surgery
null|Surgery specialty|Title|false|false||Surgerynull|Operative|Time|false|false||operativenull|Course|Time|false|false||coursenull|Uncomplicated|Modifier|false|false||uncomplicatednull|Recovery Room|Device|false|false||PACUnull|Recovery Room|Entity|false|false||PACUnull|TCF21 wt Allele|Finding|false|false||POD1
null|CORO7 gene|Finding|false|false||POD1
null|TCF21 gene|Finding|false|false||POD1null|Ventricular Fibrillation, Paroxysmal Familial, 1|Disorder|false|false|C0016520|IVFnull|SCN5A wt Allele|Finding|false|false|C0016520|IVF
null|SCN5A gene|Finding|false|false|C0016520|IVFnull|Assisted Reproductive Technologies|Procedure|false|false|C0016520|IVF
null|Fertilization in Vitro|Procedure|false|false|C0016520|IVFnull|Structure of interventricular foramen|Anatomy|false|false|C2751898;C0872104;C0015915;C1419864;C4321334;C0419179|IVFnull|NPO - Nothing by mouth|Procedure|false|false|C0016520|NPOnull|null|Entity|false|false||NPOnull|pyrrolidonecarboxylic acid|Drug|false|false|C0149576|PCA
null|p-Chloroamphetamine|Drug|false|false|C0149576|PCA
null|p-Chloroamphetamine|Drug|false|false|C0149576|PCA
null|pyrrolidonecarboxylic acid|Drug|false|false|C0149576|PCA
null|pyrrolidonecarboxylic acid|Drug|false|false|C0149576|PCAnull|Posterior cortical atrophy syndrome|Disorder|false|false|C0149576|PCA
null|Familial lichen amyloidosis|Disorder|false|false|C0149576|PCAnull|PCA Message Structure|Finding|false|false|C0149576|PCA
null|CHOANAL ATRESIA, POSTERIOR|Finding|false|false|C0149576|PCA
null|FLVCR1 gene|Finding|false|false|C0149576|PCAnull|Patient controlled intravenous analgesia|Procedure|false|false|C0149576|PCA
null|Passive Cutaneous Anaphylaxis|Procedure|false|false|C0149576|PCA
null|Patient-Controlled Analgesia|Procedure|false|false|C0149576|PCAnull|Structure of posterior cerebral artery|Anatomy|false|false|C0034330;C0030131;C0002766;C0268398;C4275079;C0078944;C5968782;C0030625;C0376636;C1549543;C0030193;C1273870;C0001554;C0220723;C1836722;C1549860|PCAnull|Principal Component Analysis|LabModifier|false|false||PCAnull|Pain management (procedure)|Procedure|false|false|C0149576|pain managementnull|Pain Management (specialty)|Title|false|false||pain managementnull|Administration Method - Pain|Finding|false|false|C0149576|pain
null|Pain|Finding|false|false|C0149576|painnull|null|Attribute|false|false||painnull|Disease Management|Procedure|false|false|C0149576|managementnull|Management Occupations|Subject|false|false||managementnull|Management procedure|Event|false|false|C0149576|management
null|Administration occupational activities|Event|false|false|C0149576|managementnull|Adequate|Modifier|false|false||adequate
null|Sufficient|Modifier|false|false||adequatenull|Relief brand of phenylephrine|Drug|false|false||relief
null|Relief brand of phenylephrine|Drug|false|false||reliefnull|Feeling relief|Finding|false|false||reliefnull|Reported Information|Finding|false|false||Reported
null|Reported|Finding|false|false||Reported
null|Report (document)|Finding|false|false||Reportednull|Reporting|Procedure|false|false||Reportednull|null|Attribute|false|false||Reported
null|null|Attribute|false|false||Reported
null|null|Attribute|false|false||Reported
null|null|Attribute|false|false||Reported
null|null|Attribute|false|false||Reportednull|Flatulence|Finding|false|false||flatusnull|Small|LabModifier|false|false||smallnull|Malignant neoplasm of abdomen|Disorder|false|false|C0230168;C0000726|Abdomennull|Abdomen problem|Finding|false|false|C0230168;C0000726|Abdomennull|Abdomen|Anatomy|false|false|C0153662;C0941288|Abdomen
null|Abdominal Cavity|Anatomy|false|false|C0153662;C0941288|Abdomennull|thiamine triphosphorate|Drug|false|false||TTP
null|ZFP36 protein, human|Drug|false|false||TTP
null|ZFP36 protein, human|Drug|false|false||TTP
null|thiamine triphosphorate|Drug|false|false||TTPnull|Congenital Thrombotic Thrombocytopenic Purpura|Disorder|false|false||TTP
null|Purpura, Thrombotic Thrombocytopenic|Disorder|false|false||TTPnull|ZFP36 wt Allele|Finding|false|false||TTP
null|ZFP36 gene|Finding|false|false||TTP
null|ADAMTS13 gene|Finding|false|false||TTPnull|Time to Progression|Time|false|false||TTPnull|Bowel sounds|Finding|false|false|C0021853|bowel soundsnull|Intestines|Anatomy|false|false|C0232693|bowelnull|null|Device|false|false||soundsnull|null|Phenomenon|false|false||soundsnull|Surgical wound|Disorder|false|false|C2338258|incisionnull|Surgical incisions|Procedure|false|false|C2338258|incisionnull|Cranial incision point|Anatomy|false|false|C0184898;C0332803|incisionnull|Erythema|Disorder|false|false||erythemanull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|vancomycin|Drug|false|false||Vancomycin
null|vancomycin|Drug|false|false||Vancomycinnull|Vancomycin measurement|Procedure|false|false||Vancomycinnull|Improvement|Finding|false|false||improvementnull|Traumatic Wound|Disorder|false|false||wound
null|Wounds and Injuries|Disorder|false|false||wound
null|Traumatic injury|Disorder|false|false||woundnull|Route of Administration - Wound|Finding|false|false||wound
null|null|Finding|false|false||wound
null|Specimen Type - Wound|Finding|false|false||woundnull|HGS protein, human|Drug|false|false||hrs
null|HGS protein, human|Drug|false|false||hrsnull|Dentatorubral-Pallidoluysian Atrophy|Disorder|false|false||hrsnull|HARS1 wt Allele|Finding|false|false||hrs
null|HARS1 gene|Finding|false|false||hrs
null|HGS wt Allele|Finding|false|false||hrs
null|HGS gene|Finding|false|false||hrs
null|ATN1 wt Allele|Finding|false|false||hrs
null|SRSF5 gene|Finding|false|false||hrsnull|Hour|Time|false|false||hrsnull|Zosyn|Drug|false|false||Zosyn
null|Zosyn|Drug|false|false||Zosynnull|GDC Regimen Terminology|Finding|false|false||regimennull|Treatment Protocols|Procedure|false|false||regimennull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|matrix metalloproteinase 7 activity|Finding|false|false||pumpnull|null|Device|false|false||pumpnull|Pump Dosing Unit|LabModifier|false|false||pumpnull|C1orf210 gene|Finding|false|false||Tempnull|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Procedure|false|false||Tempnull|Temperature|LabModifier|false|false||Tempnull|Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE|Drug|false|false||antibiotics
null|Antibiotics|Drug|false|false||antibiotics
null|Antibiotics, ophthalmologic|Drug|false|false||antibiotics
null|Antibiotics, Gynecological|Drug|false|false||antibiotics
null|antibiotics, intestinal|Drug|false|false||antibiotics
null|Antibiotic throat preparations|Drug|false|false||antibiotics
null|Antibiotics, Antitubercular|Drug|false|false||antibiotics
null|Antibiotics for systemic use|Drug|false|false||antibiotics
null|Antifungal Antibiotics, Topical|Drug|false|false||antibioticsnull|Leukocytes|Anatomy|false|false||WBCnull|Bands|Device|false|false||bandsnull|Report (document)|Finding|false|false||Reportsnull|Reporting|Procedure|false|false||Reportsnull|Persistent|Time|false|false||persistentnull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|Zofran|Drug|false|false||zofran
null|Zofran|Drug|false|false||zofrannull|MILDLY|Modifier|false|false||mildly
null|Mild (qualifier value)|Modifier|false|false||mildlynull|Effective|Modifier|false|false||effective
null|Effectiveness|Modifier|false|false||effectivenull|Compazine|Drug|false|false||Compazine
null|Compazine|Drug|false|false||Compazinenull|GDC Regimen Terminology|Finding|false|false||regimennull|Treatment Protocols|Procedure|false|false||regimennull|Improved - answer to question|Finding|false|false||improved
null|Admission Level of Care Code - Improved|Finding|false|false||improved
null|Improved|Finding|false|false||improvednull|Better|Modifier|false|false||improvednull|Effect|Modifier|false|false||effectsnull|Ventricular Fibrillation, Paroxysmal Familial, 1|Disorder|false|false|C0016520|IVFnull|SCN5A wt Allele|Finding|false|false|C0016520|IVF
null|SCN5A gene|Finding|false|false|C0016520|IVFnull|Assisted Reproductive Technologies|Procedure|false|false|C0016520|IVF
null|Fertilization in Vitro|Procedure|false|false|C0016520|IVFnull|Structure of interventricular foramen|Anatomy|false|false|C2751898;C1419864;C4321334;C0872104;C0015915|IVFnull|Team|Subject|false|false||teamnull|Antibiotics|Drug|false|false||antibioticnull|GDC Regimen Terminology|Finding|false|false||regimennull|Treatment Protocols|Procedure|false|false||regimennull|X-Ray Computed Tomography|Procedure|false|false|C0449202;C0000726|CT scannull|Radionuclide Imaging|Procedure|false|false|C0449202;C0000726|scan
null|Scanning|Procedure|false|false|C0449202;C0000726|scannull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false|C0449202;C0000726|abdnull|ABD (body structure)|Anatomy|false|false|C0034606;C0441633;C3811055;C0040405|abd
null|Abdomen|Anatomy|false|false|C0034606;C0441633;C3811055;C0040405|abdnull|Traumatic Wound|Disorder|false|false||Wound
null|Wounds and Injuries|Disorder|false|false||Wound
null|Traumatic injury|Disorder|false|false||Woundnull|Route of Administration - Wound|Finding|false|false||Wound
null|null|Finding|false|false||Wound
null|Specimen Type - Wound|Finding|false|false||Woundnull|Open|Modifier|false|false||openednull|Culture (Anthropological)|Finding|false|false||Culturesnull|Serous|Modifier|false|false||serousnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|null|Finding|false|false|C1515974|Sitenull|Anatomic Site|Anatomy|false|false|C0152053;C0278286;C1546778|Sitenull|Study Site|Modifier|false|false||Site
null|Site|Modifier|false|false||Sitenull|Dressing Dosage Form|Drug|false|false||dressingnull|null|Finding|false|false||dressing
null|Ability to dress|Finding|false|false||dressingnull|Dressing patient (procedure)|Procedure|false|false|C1515974|dressing
null|Dressing of skin or wound|Procedure|false|false|C1515974|dressingnull|Medical dressing|Device|false|false||dressing
null|Dress (garment)|Device|false|false||dressing
null|Wound Dressings (device)|Device|false|false||dressingnull|Dressing (unit of presentation)|LabModifier|false|false||dressingnull|Communicable Diseases|Disorder|false|false||Infectiousnull|infectious - Entity Risk|Modifier|false|false||Infectiousnull|Reaction|Finding|false|false||reactionnull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Gas - SpecimenType|Drug|false|false||GAS
null|Gases|Drug|false|false||GAS
null|Gas Dosage Form|Drug|false|false||GASnull|Gas - Specimen Source Codes|Finding|false|false||GAS
null|gastrointestinal gas|Finding|false|false||GAS
null|PAGR1 wt Allele|Finding|false|false||GAS
null|GALNS wt Allele|Finding|false|false||GAS
null|GALNS gene|Finding|false|false||GAS
null|GAST wt Allele|Finding|false|false||GAS
null|GAST gene|Finding|false|false||GAS
null|germacrene-A synthase activity|Finding|false|false||GAS
null|PAGR1 gene|Finding|false|false||GASnull|Staphylococcus aureus infection|Disorder|false|false||staphylococcus aureusnull|Staphylococcus aureus|Entity|false|false||staphylococcus aureusnull|Unspecified Staphylococcus infection in conditions classified elsewhere and of unspecified site|Disorder|false|false||staphylococcusnull|Genus staphylococcus|Entity|false|false||staphylococcusnull|Nasal swab (specimen)|Finding|false|false|C0028429|Nasal swabnull|Nasal Swab Test|Procedure|false|false|C0028429|Nasal swabnull|Nasal Swabs|Device|false|false||Nasal swabnull|Nasal brand of oxymetazoline|Drug|false|false|C0028429|Nasal
null|Nasal brand of oxymetazoline|Drug|false|false|C0028429|Nasal
null|Nasal dosage form|Drug|false|false|C0028429|Nasalnull|Nasal Route of Administration|Finding|false|false|C0028429|Nasal
null|Nasal (intended site)|Finding|false|false|C0028429|Nasalnull|null|Anatomy|false|false|C1272939;C0721966;C4520890;C1522019;C0563454;C3669207;C4318939|Nasalnull|Swab Dosage Form|Drug|false|false||swab
null|Swab specimen|Drug|false|false||swabnull|Taking of swab|Procedure|false|false|C0028429|swabnull|Swab|Device|false|false||swabnull|Swab Dosing Unit|LabModifier|false|false||swabnull|Micro (prefix)|Finding|false|false||Micro
null|Microbiology - Laboratory Class|Finding|false|false||Micronull|Microbiology procedure|Procedure|false|false||Micronull|Unit Of Measure Prefix - micro|LabModifier|false|false||Micronull|clindamycin|Drug|false|false||Clindamycin
null|clindamycin|Drug|false|false||Clindamycinnull|GDC Regimen Terminology|Finding|false|false||regimennull|Treatment Protocols|Procedure|false|false||regimennull|Culture (Anthropological)|Finding|false|false||Culturesnull|Wounds and Injuries|Disorder|false|false||wound
null|Traumatic Wound|Disorder|false|false||wound
null|Traumatic injury|Disorder|false|false||woundnull|Route of Administration - Wound|Finding|false|false||wound
null|null|Finding|false|false||wound
null|Specimen Type - Wound|Finding|false|false||woundnull|MAX protein, human|Drug|false|false||max
null|MAX protein, human|Drug|false|false||maxnull|Max (cigarettes)|Finding|false|false||max
null|Oncogene MAX|Finding|false|false||max
null|MAX gene|Finding|false|false||maxnull|Maximum|LabModifier|false|false||maxnull|creatinine|Drug|false|false||creatinine
null|creatinine|Drug|false|false||creatininenull|Creatinine metabolic function|Finding|false|false||creatininenull|Creatinine measurement|Procedure|false|false||creatininenull|Wound Culture|Procedure|false|false||wound culturenull|Traumatic Wound|Disorder|false|false||wound
null|Wounds and Injuries|Disorder|false|false||wound
null|Traumatic injury|Disorder|false|false||woundnull|Route of Administration - Wound|Finding|false|false||wound
null|null|Finding|false|false||wound
null|Specimen Type - Wound|Finding|false|false||woundnull|Culture positive|Finding|false|false||culture positivenull|Culture Dose Form|Drug|false|false||culturenull|Culture (Anthropological)|Finding|false|false||culture
null|Cultural aspects|Finding|false|false||culturenull|Microbial culture (procedure)|Procedure|false|false||culture
null|Laboratory culture|Procedure|false|false||culturenull|Positive|Finding|false|false||positive fornull|BRAF Gene Rearrangement|Disorder|false|false||positivenull|Rh Positive Blood Group|Finding|false|false||positive
null|Positive Finding|Finding|false|false||positive
null|Positive|Finding|false|false||positivenull|Positive Charge|Modifier|false|false||positivenull|Positive Number|LabModifier|false|false||positivenull|Encounter due to being carrier or suspected carrier of Methicillin susceptible Staphylococcus aureus|Finding|false|false||MSSAnull|Methicillin susceptible Staphylococcus aureus|Entity|false|false||MSSAnull|nafcillin|Drug|false|false||Nafcillin
null|nafcillin|Drug|false|false||Nafcillinnull|vancomycin|Drug|false|false||Vanco
null|vancomycin|Drug|false|false||Vanconull|Zosyn|Drug|false|false||Zosyn
null|Zosyn|Drug|false|false||Zosynnull|Culture (Anthropological)|Finding|false|false||culturesnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Nasal swab (specimen)|Finding|false|false|C0028429|Nasal swabnull|Nasal Swab Test|Procedure|false|false|C0028429|Nasal swabnull|Nasal Swabs|Device|false|false||Nasal swabnull|Nasal brand of oxymetazoline|Drug|false|false|C0028429|Nasal
null|Nasal brand of oxymetazoline|Drug|false|false|C0028429|Nasal
null|Nasal dosage form|Drug|false|false|C0028429|Nasalnull|Nasal Route of Administration|Finding|false|false|C0028429|Nasal
null|Nasal (intended site)|Finding|false|false|C0028429|Nasalnull|null|Anatomy|false|false|C4520890;C1522019;C0563454;C1272939;C0721966;C0038160;C3669207;C4318939|Nasalnull|Swab Dosage Form|Drug|false|false||swab
null|Swab specimen|Drug|false|false||swabnull|Taking of swab|Procedure|false|false|C0028429|swabnull|Swab|Device|false|false||swabnull|Swab Dosing Unit|LabModifier|false|false||swabnull|Staphylococcal Infections|Disorder|false|false|C0028429|Staphnull|Genus staphylococcus|Entity|false|false||Staphnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Report (document)|Finding|false|false||reportsnull|Reporting|Procedure|false|false||reportsnull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|Still|Disorder|false|false||stillnull|Present|Finding|false|false||present
null|Presentation|Finding|false|false||presentnull|Observation Interpretation - better|Finding|false|false||betternull|Better|Modifier|false|false||betternull|Small|LabModifier|false|false||smallnull|Amount class - Amount|Finding|false|false||amountnull|Quantity|LabModifier|false|false||amountnull|Regular|Modifier|false|false||regularnull|Food allergenic extracts|Drug|false|false||food
null|Food|Drug|false|false||food
null|Food allergenic extracts|Drug|false|false||foodnull|Continuous|Finding|false|false||continuednull|Flatulence|Finding|false|false||flatusnull|Liquid Stool substance|Finding|false|false||liquid stool
null|Loose stool|Finding|false|false||liquid stoolnull|Liquid Dosage Form|Drug|false|false||liquid
null|Liquid substance|Drug|false|false||liquidnull|Liquid (finding)|Finding|false|false||liquidnull|Liquid diet|Procedure|false|false||liquidnull|Liquid (state of matter)|Modifier|false|false||liquidnull|Feces|Finding|false|false||stoolnull|Stool seat|Device|false|false||stoolnull|Production Processing ID|Finding|false|false||productionnull|production|Event|false|false||productionnull|Ventricular Fibrillation, Paroxysmal Familial, 1|Disorder|false|false|C0016520|IVFnull|SCN5A wt Allele|Finding|false|false|C0016520|IVF
null|SCN5A gene|Finding|false|false|C0016520|IVFnull|Assisted Reproductive Technologies|Procedure|false|false|C0016520|IVF
null|Fertilization in Vitro|Procedure|false|false|C0016520|IVFnull|Structure of interventricular foramen|Anatomy|false|false|C1419864;C4321334;C0872104;C0015915;C2751898|IVFnull|creatinine|Drug|false|false||Creatinine
null|creatinine|Drug|false|false||Creatininenull|Creatinine metabolic function|Finding|false|false||Creatininenull|Creatinine measurement|Procedure|false|false||Creatininenull|Adequate|Modifier|false|false||Adequate
null|Sufficient|Modifier|false|false||Adequatenull|monitoring of urine output for fluid balance|Procedure|false|false||urine outputnull|null|Attribute|false|false||urine output
null|null|Attribute|false|false||urine outputnull|Urine volume finding|LabModifier|false|false||urine outputnull|Portion of urine|Finding|false|false||urine
null|null|Finding|false|false||urine
null|Urine|Finding|false|false||urine
null|In Urine|Finding|false|false||urine
null|Urine specimen|Finding|false|false||urinenull|system output|Finding|false|false||outputnull|Measurement of fluid output|Procedure|false|false||outputnull|Liver Function Tests|Procedure|false|false||LFT'snull|Isolated lipoma of filum terminale|Disorder|false|false||LFTnull|LIX1 gene|Finding|false|false||LFTnull|Liver Function Tests|Procedure|false|false||LFTnull|Slightly (qualifier value)|Modifier|false|false||slightly
null|Slight (qualifier value)|Modifier|false|false||slightlynull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|clindamycin|Drug|false|false||Clindamycin
null|clindamycin|Drug|false|false||Clindamycinnull|Culture Dose Form|Drug|false|false||culturenull|Culture (Anthropological)|Finding|false|false||culture
null|Cultural aspects|Finding|false|false||culturenull|Microbial culture (procedure)|Procedure|false|false||culture
null|Laboratory culture|Procedure|false|false||culturenull|Resistance (Psychotherapeutic)|Finding|false|false||resistance
null|social resistance|Finding|false|false||resistance
null|Resistance Process|Finding|false|false||resistancenull|Resistance|Attribute|false|false||resistancenull|nafcillin|Drug|false|false||Nafcillin
null|nafcillin|Drug|false|false||Nafcillinnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|What subject filter - Status|Finding|false|false||statusnull|null|Attribute|false|false||statusnull|Social status|Modifier|false|false||status
null|Status|Modifier|false|false||statusnull|Apyrexial|Finding|false|false||afebrilenull|White blood cell count decreased|Finding|false|false|C0023516|decreased WBCnull|Leukocytes|Anatomy|false|false|C0750394|WBCnull|Admission Level of Care Code - Improved|Finding|false|false||improved
null|Improved - answer to question|Finding|false|false||improved
null|Improved|Finding|false|false||improvednull|Better|Modifier|false|false||improvednull|patient appearance regarding mental status exam|Procedure|false|false||appearancenull|null|Attribute|false|false||appearancenull|Personal appearance|Subject|false|false||appearancenull|Appearance|Modifier|false|false||appearancenull|Kind of quantity - Appearance|LabModifier|false|false||appearancenull|Traumatic Wound|Disorder|false|false||wound
null|Wounds and Injuries|Disorder|false|false||wound
null|Traumatic injury|Disorder|false|false||woundnull|Route of Administration - Wound|Finding|false|false||wound
null|null|Finding|false|false||wound
null|Specimen Type - Wound|Finding|false|false||woundnull|Erythema|Disorder|false|false||erythemanull|Ventricular Fibrillation, Paroxysmal Familial, 1|Disorder|false|false|C0016520|IVFnull|SCN5A wt Allele|Finding|false|false|C0016520|IVF
null|SCN5A gene|Finding|false|false|C0016520|IVFnull|Assisted Reproductive Technologies|Procedure|false|false|C0016520|IVF
null|Fertilization in Vitro|Procedure|false|false|C0016520|IVFnull|Structure of interventricular foramen|Anatomy|false|false|C0872104;C0015915;C1419864;C4321334;C2751898|IVFnull|Maintenance|Event|false|false||maintenancenull|Nasal swab (specimen)|Finding|false|false|C0028429|Nasal swabnull|Nasal Swab Test|Procedure|false|false|C0028429|Nasal swabnull|Nasal Swabs|Device|false|false||Nasal swabnull|Nasal brand of oxymetazoline|Drug|false|false|C0028429|Nasal
null|Nasal brand of oxymetazoline|Drug|false|false|C0028429|Nasal
null|Nasal dosage form|Drug|false|false|C0028429|Nasalnull|Nasal Route of Administration|Finding|false|false|C0028429|Nasal
null|Nasal (intended site)|Finding|false|false|C0028429|Nasalnull|null|Anatomy|false|false|C4318939;C1272939;C0721966;C0220844;C0018270;C1457898;C1621966;C3669207;C4520890;C1522019;C0563454|Nasalnull|Swab Dosage Form|Drug|false|false||swab
null|Swab specimen|Drug|false|false||swabnull|Taking of swab|Procedure|false|false|C0028429|swabnull|Swab|Device|false|false||swabnull|Swab Dosing Unit|LabModifier|false|false||swabnull|Growth & development aspects|Finding|true|false|C0028429|growth
null|Tissue Growth|Finding|true|false|C0028429|growth
null|Growth|Finding|true|false|C0028429|growth
null|growth aspects|Finding|true|false|C0028429|growthnull|Growth action|Phenomenon|true|false||growthnull|Ventricular Fibrillation, Paroxysmal Familial, 1|Disorder|false|false|C0016520|IVFnull|SCN5A wt Allele|Finding|false|false|C0016520|IVF
null|SCN5A gene|Finding|false|false|C0016520|IVFnull|Assisted Reproductive Technologies|Procedure|false|false|C0016520|IVF
null|Fertilization in Vitro|Procedure|false|false|C0016520|IVFnull|Structure of interventricular foramen|Anatomy|false|false|C0872104;C0015915;C2751898;C1419864;C4321334;C0027324|IVFnull|nafcillin|Drug|false|false|C0016520|Nafcillin
null|nafcillin|Drug|false|false|C0016520|Nafcillinnull|Intake|Finding|false|false||intakenull|Measurement of fluid intake|Procedure|false|false||intake
null|Intake (treatment)|Procedure|false|false||intakenull|Complaint (finding)|Finding|false|false||complaintsnull|Intermittent|Time|false|false||intermittentnull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|Slow|Modifier|false|false||slowlynull|Responsive|Finding|false|false||responsivenull|Compazine|Drug|false|false||Compazine
null|Compazine|Drug|false|false||Compazinenull|Apyrexial|Finding|false|false||afebrilenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|creatinine|Drug|false|false||Creatinine
null|creatinine|Drug|false|false||Creatininenull|Creatinine metabolic function|Finding|false|false||Creatininenull|Creatinine measurement|Procedure|false|false||Creatininenull|Current (present time)|Time|false|false||Currentlynull|Finding of creatinine level|Finding|false|false||Creatinine levelnull|creatinine|Drug|false|false||Creatinine
null|creatinine|Drug|false|false||Creatininenull|Creatinine metabolic function|Finding|false|false||Creatininenull|Creatinine measurement|Procedure|false|false||Creatininenull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|Food allergenic extracts|Drug|false|false||food
null|Food|Drug|false|false||food
null|Food allergenic extracts|Drug|false|false||foodnull|Intermittent|Time|false|false||intermittentnull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|Eating|Finding|false|false||eatingnull|Narcotics|Drug|false|false||narcotics
null|Narcotics|Drug|false|false||narcoticsnull|Keflex|Drug|false|false||Keflex
null|Keflex|Drug|false|false||Keflexnull|Suspension substance|Drug|false|false||suspension
null|Suspensions|Drug|false|false||suspensionnull|Suspension (action)|Finding|false|false||suspensionnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Observation Interpretation - better|Finding|false|false||betternull|Better|Modifier|false|false||betternull|Able (qualifier value)|Finding|false|false||ablenull|Ability|Subject|false|false||ablenull|Wound care management|Procedure|false|false||wound care
null|wound care|Procedure|false|false||wound carenull|Wound Care kit|Device|false|false||wound carenull|Traumatic Wound|Disorder|false|false||wound
null|Wounds and Injuries|Disorder|false|false||wound
null|Traumatic injury|Disorder|false|false||woundnull|Route of Administration - Wound|Finding|false|false||wound
null|null|Finding|false|false||wound
null|Specimen Type - Wound|Finding|false|false||woundnull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|Lexapro|Drug|false|false||Lexapro
null|Lexapro|Drug|false|false||Lexapronull|Nasonex|Drug|false|false||nasonex
null|Nasonex|Drug|false|false||nasonexnull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|escitalopram|Drug|false|false||Escitalopram
null|escitalopram|Drug|false|false||Escitalopramnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|fluticasone|Drug|false|false||Fluticasone
null|fluticasone|Drug|false|false||Fluticasonenull|mcg/actuation|LabModifier|false|false||mcg/Actuationnull|microgram|LabModifier|false|false||mcgnull|Actuation (unit of presentation)|LabModifier|false|false||Actuationnull|SPRAY, SUSPENSION|Drug|false|false||Spray, Suspensionnull|Spray Dosage Form|Drug|false|false||Spraynull|Spray (administration method)|Finding|false|false||Spraynull|Spray (action)|Event|false|false||Spraynull|Spray Dosing Unit|LabModifier|false|false||Spraynull|Suspension substance|Drug|false|false||Suspension
null|Suspensions|Drug|false|false||Suspensionnull|Suspension (action)|Finding|false|false||Suspensionnull|Spray Dosage Form|Drug|false|false||Spraynull|Spray (administration method)|Finding|false|false|C0028429|Spraynull|Spray (action)|Event|false|false|C0028429|Spraynull|Spray Dosing Unit|LabModifier|false|false||Spraynull|Nasal brand of oxymetazoline|Drug|false|false|C0028429|Nasal
null|Nasal brand of oxymetazoline|Drug|false|false|C0028429|Nasal
null|Nasal dosage form|Drug|false|false|C0028429|Nasalnull|Nasal Route of Administration|Finding|false|false|C0028429|Nasal
null|Nasal (intended site)|Finding|false|false|C0028429|Nasalnull|null|Anatomy|false|false|C2003858;C4520890;C1522019;C1272939;C0721966;C4521772|Nasalnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|Colace|Drug|false|false||Colace
null|Colace|Drug|false|false||Colacenull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0006935|Capsule
null|Structure of organ capsule|Anatomy|false|false|C0006935|Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0006935;C1561538;C1561539|Capsule
null|Structure of organ capsule|Anatomy|false|false|C0006935;C1561538;C1561539|Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Twice a day|Time|false|false||twice a daynull|Transaction counts and value totals - day|Finding|false|false|C0524463;C1325531|day
null|Precision - day|Finding|false|false|C0524463;C1325531|daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Constipation|Finding|false|false||constipationnull|month|Time|false|false||monthsnull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0006935|Capsule
null|Structure of organ capsule|Anatomy|false|false|C0006935|Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|refill|Finding|false|false||Refillsnull|lorazepam|Drug|false|false||Lorazepam
null|lorazepam|Drug|false|false||Lorazepamnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Every eight hours|Time|false|false||Q8Hnull|Hour|Time|false|false||hoursnull|Anxiety Disorders|Disorder|false|false||anxiety
null|Anxiety|Disorder|false|false||anxietynull|Anxiety symptoms|Finding|false|false||anxietynull|hydrocortisone|Drug|false|false||Hydrocortisone
null|hydrocortisone|Drug|false|false||Hydrocortisone
null|hydrocortisone|Drug|false|false||Hydrocortisonenull|Cortisol Measurement|Procedure|false|false||Hydrocortisonenull|Emollient Cream|Drug|false|false||Cream
null|Cream|Drug|false|false||Cream
null|Dairy Cream|Drug|false|false||Creamnull|APPL1 gene|Finding|false|false||Applnull|Rectal Dosage Form|Drug|false|false||Rectalnull|Rectal Route of Administration|Finding|false|false||Rectal
null|Rectal (intended site)|Finding|false|false||Rectalnull|TUBE,RECTAL,24FR,PLASTIC B#6510|Device|false|false||Rectalnull|rectal|Modifier|false|false||Rectalnull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Hemorrhoids|Disorder|false|false||hemorrhoidsnull|cephalexin|Drug|false|false||Cephalexin
null|cephalexin|Drug|false|false||Cephalexinnull|Suspension for Reconstitution Dosage Form|Drug|false|false||Suspension for Reconstitutionnull|Suspension substance|Drug|false|false||Suspension
null|Suspensions|Drug|false|false||Suspensionnull|Suspension (action)|Finding|false|false||Suspensionnull|5 Days|Time|false|false||5 daysnull|day|Time|false|false||daysnull|refill|Finding|false|false||Refillsnull|Tylenol|Drug|false|false||Tylenol
null|Tylenol|Drug|false|false||Tylenolnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Hour|Time|false|false||hoursnull|Fever symptoms (finding)|Finding|false|false||fever
null|Fever|Finding|false|false||fevernull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Referral category - Outpatient|Finding|false|false||Outpatient
null|Patient Class - Outpatient|Finding|false|false||Outpatientnull|Outpatients|Subject|false|false||Outpatientnull|AML Lab Table|Finding|false|false||Lab
null|LAT2 gene|Finding|false|false||Lab
null|EWS Lab Table|Finding|false|false||Labnull|Laboratory|Device|false|false||Labnull|Labrador retriever|Entity|false|false||Lab
null|Laboratory|Entity|false|false||Labnull|Work|Event|false|false||Worknull|Serum creatinine level|Finding|false|false||serum Creatininenull|Creatinine measurement, serum (procedure)|Procedure|false|false||serum Creatininenull|Cell Culture Serum|Drug|false|false||serumnull|Serum specimen|Finding|false|false||serum
null|null|Finding|false|false||serum
null|Serum|Finding|false|false||serumnull|creatinine|Drug|false|false||Creatinine
null|creatinine|Drug|false|false||Creatininenull|Creatinine metabolic function|Finding|false|false||Creatininenull|Creatinine measurement|Procedure|false|false||Creatininenull|What subject filter - Result|Finding|false|false||result
null|Result|Finding|false|false||result
null|Experimental Result|Finding|false|false||resultnull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|ADMIN.FACILITY|Finding|false|false||Facilitynull|Facility (object)|Device|false|false||Facilitynull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|True primary (qualifier value)|Time|false|false||Primarynull|Primary|Modifier|false|false||Primarynull|Recurrent|Time|false|false||Recurrent
null|Episodic|Time|false|false||Recurrentnull|Diverticulitis|Disorder|false|false||Diverticulitisnull|Wound cellulitis|Disorder|false|false||wound cellulitisnull|Traumatic Wound|Disorder|false|false||wound
null|Wounds and Injuries|Disorder|false|false||wound
null|Traumatic injury|Disorder|false|false||woundnull|Route of Administration - Wound|Finding|false|false||wound
null|null|Finding|false|false||wound
null|Specimen Type - Wound|Finding|false|false||woundnull|Cellulitis|Disorder|false|false||cellulitisnull|cellulitis on exam (physical finding)|Finding|false|false||cellulitisnull|Hypovolemia|Finding|false|false||hypovolemianull|Fever symptoms (finding)|Finding|false|false||fever
null|Fever|Finding|false|false||fevernull|Neoplasm Metastasis|Disorder|false|false||Secondarynull|metastatic qualifier|Finding|false|false||Secondarynull|Secondary to|Modifier|false|false||Secondarynull|second (number)|LabModifier|false|false||Secondarynull|Anxiety Disorders|Disorder|false|false||Anxiety
null|Anxiety|Disorder|false|false||Anxietynull|Anxiety symptoms|Finding|false|false||Anxietynull|Diverticulosis|Disorder|false|false||diverticulosisnull|Patient Condition Code - Stable|Finding|false|false||Stablenull|Stable status|Modifier|false|false||Stablenull|Regular|Modifier|false|false||regularnull|IPSS-R Risk Category Low|Finding|false|false||low
null|IPSS Risk Category Low|Finding|false|false||low
null|low confidentiality|Finding|false|false||lownull|Low - MessageWaitingPriority|Modifier|false|false||low
null|low|Modifier|false|false||low
null|low exposure|Modifier|false|false||lownull|null|LabModifier|false|false||lownull|Residue|Finding|false|false||residuenull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Adequate|Modifier|false|false||Adequate
null|Sufficient|Modifier|false|false||Adequatenull|Demonstrates adequate pain control|Finding|false|false||pain controlnull|Pain control|Procedure|false|false||pain control
null|Pain management (procedure)|Procedure|false|false||pain controlnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Control brand of phenylpropanolamine|Drug|false|false||control
null|CONTROL veterinary product|Drug|false|false||control
null|control substance|Drug|false|false||control
null|Control brand of phenylpropanolamine|Drug|false|false||controlnull|Control - Relationship modifier|Finding|false|false||control
null|Control function|Finding|false|false||control
null|Scientific Control|Finding|false|false||controlnull|Control Groups|Subject|false|false||controlnull|True Control Status|Modifier|false|false||control
null|control aspects|Modifier|false|false||controlnull|Oral medication (substance)|Drug|false|false||oral medicationnull|Oral Medication|Procedure|false|false|C0226896|oral medicationnull|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C1272919;C0175795;C1527415;C4521986|oralnull|Oral|Modifier|false|false||oralnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Doctor - Title|Finding|false|false||doctornull|Physicians|Subject|false|false||doctornull|Return to (contextual qualifier) (qualifier value)|Modifier|false|false||return tonull|Return to (contextual qualifier) (qualifier value)|Modifier|false|false||returnnull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|Chest Pain|Finding|false|false|C1527391;C0817096|chest painnull|null|Attribute|false|false|C1527391;C0817096|chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0741025;C0008031;C2926613|chest
null|Anterior thoracic region|Anatomy|false|false|C0741025;C0008031;C2926613|chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|Tightness sensation quality|Modifier|false|false||tightnessnull|Query Status Code - new|Finding|false|false||New
null|Act Status - new|Finding|false|false||Newnull|Newar Language|Entity|false|false||Newnull|New|Modifier|false|false||Newnull|Patient Outcome - Worsening|Finding|false|false||worseningnull|Worsening (qualifier value)|Modifier|false|false||worseningnull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|Wheezing|Finding|false|false||wheezingnull|Vomiting|Finding|false|false||vomitingnull|Liquid substance|Drug|false|false||fluidsnull|Mouse Body Fluid or Substance|Finding|false|false||fluidsnull|Fluid Therapy|Procedure|false|false||fluidsnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Dehydration|Disorder|false|false||dehydratednull|Vomiting|Finding|false|false||vomitingnull|rectal discharge diarrhea (physical finding)|Finding|false|false||diarrhea
null|Diarrhea|Finding|false|false||diarrheanull|Indication of (contextual qualifier)|Finding|false|false||reasonsnull|Signs of dehydration|Finding|false|false||Signs of dehydrationnull|Aspects of signs|Finding|false|false||Signs
null|Physical findings|Finding|false|false||Signsnull|Manufactured sign|Device|false|false||Signsnull|dehydration (Na, H2O)|Disorder|false|false||dehydration
null|Dehydration|Disorder|false|false||dehydrationnull|Dehydration procedure|Procedure|false|false||dehydrationnull|Oral cavity|Anatomy|false|false|C0849959;C1527305;C0425583;C4554554;C0039070;C0039231|mouth
null|Oral region|Anatomy|false|false|C0849959;C1527305;C0425583;C4554554;C0039070;C0039231|mouthnull|Tachycardia|Finding|false|false|C0230028;C0226896|rapid heartbeatnull|Rapid|Modifier|false|false||rapidnull|Heart beat|Finding|false|false|C0230028;C0226896|heartbeatnull|Pulse Rate|Attribute|false|false||heartbeatnull|feeling dizzy|Finding|false|false|C0230028;C0226896|feeling dizzynull|Feelings|Finding|false|false|C0230028;C0226896|feelingnull|Dizziness|Finding|false|false||dizzynull|Faint - appearance|Finding|false|false|C0230028;C0226896|faint
null|Syncope|Finding|false|false|C0230028;C0226896|faintnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Dark color|Modifier|false|false||darknull|Black - ethnic group (ethnic group)|Subject|false|false||black
null|Black race|Subject|false|false||black
null|African|Subject|false|false||blacknull|Black - Structured Product Labeling Color|Modifier|false|false||black
null|Black color|Modifier|false|false||blacknull|Materials|Drug|false|false||materialnull|Defecation|Finding|false|false|C0021853|bowel movementnull|Intestines|Anatomy|false|false|C0011135|bowelnull|Movement|Finding|false|false||movementnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Hour|Time|false|false||hoursnull|Within 24 hours|Time|false|false||within 24 hoursnull|24 Hours|Time|false|false||24 hoursnull|Hour|Time|false|false||hoursnull|Call - dosing instruction fragment|Finding|false|false||Call
null|Call (Instruction)|Finding|false|false||Call
null|Decision|Finding|false|false||Call
null|CHL1 gene|Finding|false|false||Callnull|Return to (contextual qualifier) (qualifier value)|Modifier|false|false||returnnull|Stat (do immediately)|Time|false|false||immediatelynull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Observation Interpretation - worse|Finding|false|false||worse
null|Worse|Finding|false|false||worsenull|Worsening (qualifier value)|Modifier|false|false||worsenull|Changing|Finding|false|false|C1515974|changingnull|Changed status|LabModifier|false|false||changingnull|Transaction counts and value totals - location|Finding|false|false|C1515974|locationnull|Anatomic Site|Anatomy|false|false|C0741025;C1555588;C0392747|locationnull|location participation type|Device|false|false||locationnull|location participation type|Entity|false|false||locationnull|Location|Modifier|false|false||locationnull|Chest problem|Finding|false|false|C1527391;C0817096;C1515974|chestnull|Chest|Anatomy|false|false|C0741025|chest
null|Anterior thoracic region|Anatomy|false|false|C0741025|chestnull|heavy machinery|Device|false|false||heavy machinerynull|Heavy (weight) (qualifier value)|Modifier|false|false||heavy
null|Heavy (amount)|Modifier|false|false||heavynull|Contact with machinery|Disorder|false|false||machinerynull|Industrial machine|Device|false|false||machinerynull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Chills|Finding|false|false||chillsnull|Fever symptoms (finding)|Finding|false|false||fever
null|Fever|Finding|false|false||fevernull|Greater Than|LabModifier|false|false||greater thannull|Greater|LabModifier|false|false||greaternull|Academic degree|Finding|false|false||degreesnull|Degree or extent|LabModifier|false|false||degreesnull|Academic degree|Finding|false|false||degreesnull|Degree or extent|LabModifier|false|false||degreesnull|Equipment Alert Level - Serious|Finding|false|false||serious
null|Device Alert Level - Serious|Finding|false|false||serious
null|Alert level - Serious|Finding|false|false||seriousnull|Serious|Modifier|false|false||seriousnull|Changing|Finding|false|false||changenull|Change - procedure|Procedure|false|false||changenull|Delta (difference)|LabModifier|false|false||change
null|Changed status|LabModifier|false|false||changenull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Concern|Finding|false|false||concernnull|Regular|Modifier|false|false||regularnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|MICROCEPHALY, EPILEPSY, AND DIABETES SYNDROME 1|Disorder|false|false||medsnull|Medications|Finding|false|false||medsnull|Several times per day|Finding|false|false||several times per daynull|Several|LabModifier|false|false||severalnull|times/day|LabModifier|false|false||times per daynull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|per day|Time|false|false||per daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Wound care management|Procedure|false|false||WOUND CARE
null|wound care|Procedure|false|false||WOUND CAREnull|Wound Care kit|Device|false|false||WOUND CAREnull|Traumatic Wound|Disorder|false|false||WOUND
null|Wounds and Injuries|Disorder|false|false||WOUND
null|Traumatic injury|Disorder|false|false||WOUNDnull|Route of Administration - Wound|Finding|false|false||WOUND
null|null|Finding|false|false||WOUND
null|Specimen Type - Wound|Finding|false|false||WOUNDnull|In care (finding)|Finding|false|false||CARE
null|Continuity Assessment Record and Evaluation|Finding|false|false||CAREnull|care activity|Event|false|false||CAREnull|Surgical wound|Disorder|false|false|C1515974|surgical woundnull|Surgical wound finding|Finding|false|false|C1515974|surgical woundnull|Operative Surgical Procedures|Procedure|false|false||surgical
null|Surgical service|Procedure|false|false||surgicalnull|Traumatic Wound|Disorder|false|false|C1515974|wound
null|Wounds and Injuries|Disorder|false|false|C1515974|wound
null|Traumatic injury|Disorder|false|false|C1515974|woundnull|Route of Administration - Wound|Finding|false|false|C1515974|wound
null|null|Finding|false|false|C1515974|wound
null|Specimen Type - Wound|Finding|false|false|C1515974|woundnull|null|Finding|false|false|C1515974|sitenull|Anatomic Site|Anatomy|false|false|C1546778;C3263723;C0043251;C0043250;C1628502;C1549529;C1547965;C1550680;C0332803|sitenull|Study Site|Modifier|false|false||site
null|Site|Modifier|false|false||sitenull|Daily|Time|false|false||dailynull|Changing|Finding|false|false||Changenull|Change - procedure|Procedure|false|false||Changenull|Delta (difference)|LabModifier|false|false||Change
null|Changed status|LabModifier|false|false||Changenull|Packing Dosage Form|Drug|false|false||packingnull|Insertion of pack (procedure)|Procedure|false|false||packingnull|Packing material|Device|false|false||packingnull|Packing (action)|Event|false|false||packingnull|Once daily|Time|false|false||once per daynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|per day|Time|false|false||per daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Pack|Drug|false|false||Packnull|Pack (physical object)|Device|false|false||Pack
null|Pack unit|Device|false|false||Packnull|Packing (action)|Event|false|false||Packnull|Package Dosing Unit|LabModifier|false|false||Packnull|Gauzes|Device|false|false||gauzenull|Saline Solution|Drug|false|false||Saline
null|Saline Solution|Drug|false|false||Salinenull|Saline method|Procedure|false|false||Salinenull|Surgical incisions|Procedure|false|false||incisionalnull|Dental caries|Disorder|false|false|C0333343|cavity
null|Cavitation|Disorder|false|false|C0333343|cavitynull|Body cavities|Anatomy|false|false|C1510420;C0011334|cavitynull|Gauzes|Device|false|false||gauzenull|Fix|Phenomenon|false|false||adherenull|TAPE,PAPER|Device|false|false||paper tapenull|Paper Authorization|Finding|false|false||papernull|Paper|Device|false|false||papernull|Paper Dosing Unit|LabModifier|false|false||papernull|Tape Dosage Form|Drug|false|false||tapenull|CC2D1A gene|Finding|false|false||tapenull|Biomedical tape|Device|false|false||tape
null|Tape Device|Device|false|false||tapenull|Changing|Finding|false|false||Changednull|Changed status|LabModifier|false|false||Changednull|Gauzes|Device|false|false||gauzenull|Saturated|Phenomenon|false|false||saturatednull|Have Vulvar Irritation question|Finding|false|false||irritation
null|Irritability - emotion|Finding|false|false||irritation
null|Irritation (finding)|Finding|false|false||irritationnull|Irritation|Phenomenon|false|false||irritationnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false|C1123023;C4520765|skin
null|Skin and subcutaneous tissue disorders|Disorder|false|false|C1123023;C4520765|skinnull|Skin Specimen Source Code|Finding|false|false|C1123023;C4520765|skin
null|Skin Specimen|Finding|false|false|C1123023;C4520765|skinnull|Skin, Human|Anatomy|false|false|C1546781;C0444099;C0178298;C0496955|skin
null|Skin|Anatomy|false|false|C1546781;C0444099;C0178298;C0496955|skinnull|Traumatic Wound|Disorder|false|false||wound
null|Wounds and Injuries|Disorder|false|false||wound
null|Traumatic injury|Disorder|false|false||woundnull|Route of Administration - Wound|Finding|false|false||wound
null|null|Finding|false|false||wound
null|Specimen Type - Wound|Finding|false|false||woundnull|Pack|Drug|false|false||packnull|Pack (physical object)|Device|false|false||pack
null|Pack unit|Device|false|false||packnull|Packing (action)|Event|false|false||packnull|Package Dosing Unit|LabModifier|false|false||packnull|Aquacel|Drug|false|false||Aquacelnull|Disorders of Sex Development|Disorder|false|false||DSD
null|Diaphanospondylodysostosis|Disorder|false|false||DSDnull|Wash Dosage Form|Drug|false|false||washnull|Wash - dosing instruction imperative|Finding|false|false||wash
null|Wash - Specimen Source Codes|Finding|false|false||wash
null|WASHC1 gene|Finding|false|false||wash
null|Wash - Administration Method|Finding|false|false||washnull|Cell Wash|Procedure|false|false||washnull|Wash (cleansing action)|Event|false|false||washnull|Surgical wound|Disorder|false|false||surgical incisionsnull|Surgical incisions|Procedure|false|false||surgical incisionsnull|Operative Surgical Procedures|Procedure|false|false||surgical
null|Surgical service|Procedure|false|false||surgicalnull|Surgical incisions|Procedure|false|false||incisionsnull|swimming (history)|Finding|false|false||swimming
null|Swimming|Finding|false|false||swimmingnull|TUB gene|Finding|false|false||tubnull|Tub - container|Device|false|false||tubnull|Tub Dosing Unit|LabModifier|false|false||tubnull|Bathing|Procedure|false|false||bathsnull|Baths (medical device)|Device|false|false||bathsnull|Wounds and Injuries|Disorder|false|false||wound
null|Traumatic Wound|Disorder|false|false||wound
null|Traumatic injury|Disorder|false|false||woundnull|Route of Administration - Wound|Finding|false|false||wound
null|null|Finding|false|false||wound
null|Specimen Type - Wound|Finding|false|false||woundnull|Completely - dosing instruction fragment|Finding|false|false||completelynull|Complete|Modifier|false|false||completelynull|Doctor - Title|Finding|false|false||doctornull|Physicians|Subject|false|false||doctornull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|Erythema|Disorder|false|false||rednessnull|Redness|Finding|false|false||rednessnull|Red color|Modifier|false|false||rednessnull|Body Substance Discharge|Finding|false|false||drainage
null|Body Fluid Discharge|Finding|false|false||drainagenull|Drainage procedure|Procedure|false|false||drainagenull|Site of incision|Modifier|false|false||incision sitesnull|Surgical wound|Disorder|false|false|C2338258|incisionnull|Surgical incisions|Procedure|false|false|C2338258|incisionnull|Cranial incision point|Anatomy|false|false|C0332803;C0184898|incisionnull|Site|Modifier|false|false||sitesnull|creatinine|Drug|false|false||CREATININE
null|creatinine|Drug|false|false||CREATININEnull|Creatinine metabolic function|Finding|false|false||CREATININEnull|Creatinine measurement|Procedure|false|false||CREATININEnull|creatinine|Drug|false|false||creatinine
null|creatinine|Drug|false|false||creatininenull|Creatinine metabolic function|Finding|false|false||creatininenull|Creatinine measurement|Procedure|false|false||creatininenull|Call - dosing instruction fragment|Finding|false|false||call
null|Call (Instruction)|Finding|false|false||call
null|Decision|Finding|false|false||call
null|CHL1 gene|Finding|false|false||callnull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|Address type - Office|Finding|false|false||officenull|Office|Device|false|false||officenull|Organization unit type - Office|Entity|false|false||officenull|What subject filter - Result|Finding|false|false||result
null|Result|Finding|false|false||result
null|Experimental Result|Finding|false|false||resultnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions