 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|25,29
No|30,32
:|32,33
_|36,37
_|37,38
_|38,39
<EOL>|39,40
<EOL>|41,42
Admission|42,51
Date|52,56
:|56,57
_|59,60
_|60,61
_|61,62
Discharge|76,85
Date|86,90
:|90,91
_|94,95
_|95,96
_|96,97
<EOL>|97,98
<EOL>|99,100
Date|100,104
of|105,107
Birth|108,113
:|113,114
_|116,117
_|117,118
_|118,119
Sex|132,135
:|135,136
F|139,140
<EOL>|140,141
<EOL>|142,143
Service|143,150
:|150,151
MEDICINE|152,160
<EOL>|160,161
<EOL>|162,163
Allergies|163,172
:|172,173
<EOL>|174,175
IV|175,177
Dye|178,181
,|181,182
Iodine|183,189
Containing|190,200
Contrast|201,209
Media|210,215
/|216,217
Oxycodone|218,227
/|228,229
<EOL>|230,231
cilostazol|231,241
/|242,243
Varenicline|244,255
<EOL>|255,256
<EOL>|257,258
Attending|258,267
:|267,268
_|269,270
_|270,271
_|271,272
.|272,273
<EOL>|273,274
<EOL>|275,276
Chief|276,281
Complaint|282,291
:|291,292
<EOL>|292,293
Shortness|293,302
of|303,305
breath|306,312
<EOL>|312,313
<EOL>|314,315
Major|315,320
Surgical|321,329
or|330,332
Invasive|333,341
Procedure|342,351
:|351,352
<EOL>|352,353
None|353,357
<EOL>|357,358
<EOL>|358,359
<EOL>|360,361
History|361,368
of|369,371
Present|372,379
Illness|380,387
:|387,388
<EOL>|388,389
Ms.|389,392
_|393,394
_|394,395
_|395,396
is|397,399
a|400,401
_|402,403
_|403,404
_|404,405
yo|406,408
woman|409,414
with|415,419
a|420,421
PMH|422,425
notable|426,433
for|434,437
COPD|438,442
on|443,445
<EOL>|446,447
home|447,451
O2|452,454
(|454,455
hospitalized|455,467
_|468,469
_|469,470
_|470,471
,|471,472
multiple|473,481
recent|482,488
ED|489,491
visits|492,498
)|498,499
,|499,500
Afib|501,505
on|506,508
<EOL>|509,510
apixaban|510,518
,|518,519
HTN|520,523
,|523,524
CAD|525,528
,|528,529
and|530,533
HLD|534,537
who|538,541
presents|542,550
with|551,555
several|556,563
days|564,568
of|569,571
<EOL>|572,573
worsening|573,582
dyspnea|583,590
.|590,591
<EOL>|591,592
<EOL>|592,593
Patient|593,600
has|601,604
had|605,608
several|609,616
ED|617,619
visits|620,626
for|627,630
dyspnea|631,638
and|639,642
a|643,644
recent|645,651
<EOL>|652,653
hospitalization|653,668
for|669,672
a|673,674
COPD|675,679
exacerbation|680,692
in|693,695
_|696,697
_|697,698
_|698,699
.|699,700
She|701,704
has|705,708
<EOL>|709,710
been|710,714
on|715,717
steroid|718,725
therapy|726,733
with|734,738
several|739,746
attempts|747,755
to|756,758
taper|759,764
over|765,769
the|770,773
<EOL>|774,775
last|775,779
several|780,787
months|788,794
.|794,795
After|796,801
her|802,805
most|806,810
recent|811,817
ED|818,820
visit|821,826
on|827,829
_|830,831
_|831,832
_|832,833
<EOL>|834,835
she|835,838
was|839,842
on|843,845
placed|846,852
on|853,855
60|856,858
mg|859,861
PO|862,864
prednisone|865,875
with|876,880
a|881,882
taper|883,888
down|889,893
by|894,896
10|897,899
<EOL>|900,901
mg|901,903
each|904,908
day|909,912
.|912,913
Her|914,917
SOB|918,921
worsened|922,930
with|931,935
the|936,939
taper|940,945
and|946,949
she|950,953
was|954,957
seen|958,962
on|963,965
<EOL>|966,967
_|967,968
_|968,969
_|969,970
by|971,973
her|974,977
PCP|978,981
who|982,985
started|986,993
her|994,997
on|998,1000
a|1001,1002
course|1003,1009
of|1010,1012
prednisone|1013,1023
30|1024,1026
mg|1027,1029
<EOL>|1030,1031
PO|1031,1033
to|1034,1036
be|1037,1039
tapered|1040,1047
down|1048,1052
by|1053,1055
5|1056,1057
mg|1058,1060
every|1061,1066
3|1067,1068
days|1069,1073
.|1073,1074
With|1075,1079
the|1080,1083
taper|1084,1089
she|1090,1093
<EOL>|1094,1095
is|1095,1097
currently|1098,1107
on|1108,1110
prednisone|1111,1121
25|1122,1124
mg|1125,1127
QD|1128,1130
.|1130,1131
<EOL>|1131,1132
<EOL>|1132,1133
She|1133,1136
reports|1137,1144
that|1145,1149
her|1150,1153
SOB|1154,1157
improved|1158,1166
slightly|1167,1175
after|1176,1181
starting|1182,1190
the|1191,1194
<EOL>|1195,1196
steroids|1196,1204
on|1205,1207
_|1208,1209
_|1209,1210
_|1210,1211
.|1211,1212
However|1213,1220
,|1220,1221
last|1222,1226
night|1227,1232
it|1233,1235
acutely|1236,1243
worsened|1244,1252
and|1253,1256
she|1257,1260
<EOL>|1261,1262
was|1262,1265
unable|1266,1272
to|1273,1275
sleep|1276,1281
.|1281,1282
She|1283,1286
usually|1287,1294
uses|1295,1299
3|1300,1301
pillows|1302,1309
to|1310,1312
sleep|1313,1318
but|1319,1322
was|1323,1326
<EOL>|1327,1328
only|1328,1332
comfortable|1333,1344
seated|1345,1351
upright|1352,1359
last|1360,1364
night|1365,1370
.|1370,1371
This|1372,1376
morning|1377,1384
she|1385,1388
<EOL>|1389,1390
increased|1390,1399
her|1400,1403
oxygen|1404,1410
to|1411,1413
3L|1414,1416
and|1417,1420
felt|1421,1425
better|1426,1432
.|1432,1433
She|1434,1437
is|1438,1440
usually|1441,1448
on|1449,1451
2L|1452,1454
<EOL>|1455,1456
NC|1456,1458
at|1459,1461
home|1462,1466
.|1466,1467
She|1468,1471
reports|1472,1479
that|1480,1484
for|1485,1488
the|1489,1492
last|1493,1497
several|1498,1505
months|1506,1512
she|1513,1516
has|1517,1520
<EOL>|1521,1522
been|1522,1526
using|1527,1532
two|1533,1536
different|1537,1546
albuterol|1547,1556
inhalers|1557,1565
each|1566,1570
every|1571,1576
_|1577,1578
_|1578,1579
_|1579,1580
<EOL>|1581,1582
hours|1582,1587
.|1587,1588
She|1589,1592
knows|1593,1598
that|1599,1603
this|1604,1608
is|1609,1611
more|1612,1616
than|1617,1621
they|1622,1626
are|1627,1630
prescribed|1631,1641
for|1642,1645
<EOL>|1646,1647
but|1647,1650
it|1651,1653
makes|1654,1659
her|1660,1663
comfortable|1664,1675
.|1675,1676
She|1677,1680
mostly|1681,1687
stays|1688,1693
put|1694,1697
on|1698,1700
the|1701,1704
second|1705,1711
<EOL>|1712,1713
floor|1713,1718
of|1719,1721
her|1722,1725
home|1726,1730
.|1730,1731
She|1732,1735
states|1736,1742
that|1743,1747
she|1748,1751
can|1752,1755
walk|1756,1760
to|1761,1763
the|1764,1767
bathroom|1768,1776
<EOL>|1777,1778
without|1778,1785
being|1786,1791
short|1792,1797
of|1798,1800
breath|1801,1807
,|1807,1808
but|1809,1812
does|1813,1817
not|1818,1821
use|1822,1825
the|1826,1829
stairs|1830,1836
<EOL>|1837,1838
unless|1838,1844
she|1845,1848
has|1849,1852
to|1853,1855
leave|1856,1861
the|1862,1865
house|1866,1871
because|1872,1879
it|1880,1882
worsens|1883,1890
her|1891,1894
<EOL>|1895,1896
breathing|1896,1905
.|1905,1906
She|1907,1910
endorses|1911,1919
a|1920,1921
cough|1922,1927
occasionally|1928,1940
productive|1941,1951
of|1952,1954
_|1955,1956
_|1956,1957
_|1957,1958
<EOL>|1959,1960
sputum|1960,1966
.|1966,1967
This|1968,1972
is|1973,1975
consistent|1976,1986
with|1987,1991
her|1992,1995
baseline|1996,2004
.|2004,2005
She|2006,2009
endorses|2010,2018
one|2019,2022
<EOL>|2023,2024
episode|2024,2031
of|2032,2034
non-exertional|2035,2049
chest|2050,2055
pain|2056,2060
today|2061,2066
that|2067,2071
spontaneously|2072,2085
<EOL>|2086,2087
resolved|2087,2095
.|2095,2096
She|2097,2100
denies|2101,2107
fever|2108,2113
,|2113,2114
chills|2115,2121
,|2121,2122
recent|2123,2129
sick|2130,2134
contacts|2135,2143
,|2143,2144
and|2145,2148
<EOL>|2149,2150
lower|2150,2155
extremity|2156,2165
edema|2166,2171
.|2171,2172
<EOL>|2172,2173
<EOL>|2173,2174
In|2174,2176
the|2177,2180
ED|2181,2183
,|2183,2184
initial|2185,2192
vital|2193,2198
signs|2199,2204
were|2205,2209
:|2209,2210
T|2211,2212
98.5|2213,2217
P|2218,2219
80|2220,2222
BP|2223,2225
154|2226,2229
/|2229,2230
97|2230,2232
R|2233,2234
20|2235,2237
<EOL>|2238,2239
O2|2239,2241
sat|2242,2245
97|2246,2248
%|2248,2249
NC|2250,2252
.|2252,2253
<EOL>|2255,2256
-|2256,2257
Exam|2258,2262
notable|2263,2270
for|2271,2274
:|2274,2275
Diffuse|2276,2283
expiratory|2284,2294
wheezing|2295,2303
,|2303,2304
prolonged|2305,2314
<EOL>|2315,2316
expiratory|2316,2326
phase|2327,2332
,|2332,2333
left|2334,2338
inspiratory|2339,2350
crackles|2351,2359
,|2359,2360
irregularly|2361,2372
<EOL>|2373,2374
irregular|2374,2383
rhthym|2384,2390
,|2390,2391
minimal|2392,2399
pedal|2400,2405
edema|2406,2411
<EOL>|2413,2414
-|2414,2415
Labs|2416,2420
were|2421,2425
notable|2426,2433
for|2434,2437
CBC|2438,2441
wnl|2442,2445
,|2445,2446
proBNP|2447,2453
235|2454,2457
,|2457,2458
Trop|2459,2463
0.02|2464,2468
,|2468,2469
chem|2470,2474
<EOL>|2475,2476
notable|2476,2483
for|2484,2487
bicarb|2488,2494
31|2495,2497
,|2497,2498
AG|2499,2501
13|2502,2504
,|2504,2505
UA|2506,2508
notable|2509,2516
for|2517,2520
40|2521,2523
RBCs|2524,2528
<EOL>|2530,2531
-|2531,2532
Studies|2533,2540
performed|2541,2550
include|2551,2558
CXR|2559,2562
with|2563,2567
stable|2568,2574
mild|2575,2579
/|2579,2580
moderate|2580,2588
<EOL>|2589,2590
cardiomegaly|2590,2602
,|2602,2603
atelectasis|2604,2615
at|2616,2618
bases|2619,2624
,|2624,2625
otherwise|2626,2635
clear|2636,2641
lung|2642,2646
fields|2647,2653
<EOL>|2653,2654
-|2654,2655
Patient|2656,2663
was|2664,2667
given|2668,2673
Albuterol|2674,2683
neb|2684,2687
x|2688,2689
1|2690,2691
,|2691,2692
ipratropium|2693,2704
neb|2705,2708
x|2709,2710
1|2711,2712
,|2712,2713
<EOL>|2714,2715
Azithromycin|2715,2727
500|2728,2731
mg|2732,2734
PO|2735,2737
,|2737,2738
Prednisone|2739,2749
25|2750,2752
mg|2753,2755
PO|2756,2758
<EOL>|2758,2759
<EOL>|2759,2760
Upon|2760,2764
arrival|2765,2772
to|2773,2775
the|2776,2779
floor|2780,2785
,|2785,2786
the|2787,2790
patient|2791,2798
states|2799,2805
that|2806,2810
she|2811,2814
is|2815,2817
doing|2818,2823
<EOL>|2824,2825
well|2825,2829
.|2829,2830
She|2831,2834
says|2835,2839
that|2840,2844
her|2845,2848
SOB|2849,2852
has|2853,2856
improved|2857,2865
since|2866,2871
this|2872,2876
morning|2877,2884
and|2885,2888
<EOL>|2889,2890
is|2890,2892
better|2893,2899
than|2900,2904
last|2905,2909
night|2910,2915
when|2916,2920
she|2921,2924
could|2925,2930
not|2931,2934
sleep|2935,2940
.|2940,2941
<EOL>|2943,2944
<EOL>|2945,2946
Review|2946,2952
of|2953,2955
Systems|2956,2963
:|2963,2964
<EOL>|2966,2967
(|2968,2969
+|2969,2970
)|2970,2971
per|2972,2975
HPI|2976,2979
<EOL>|2981,2982
(|2983,2984
-|2984,2985
)|2985,2986
fever|2987,2992
,|2992,2993
chills|2994,3000
,|3000,3001
night|3002,3007
sweats|3008,3014
,|3014,3015
headache|3016,3024
,|3024,3025
vision|3026,3032
changes|3033,3040
,|3040,3041
<EOL>|3042,3043
rhinorrhea|3043,3053
,|3053,3054
congestion|3055,3065
,|3065,3066
sore|3067,3071
throat|3072,3078
,|3078,3079
abdominal|3080,3089
pain|3090,3094
,|3094,3095
nausea|3096,3102
,|3102,3103
<EOL>|3104,3105
vomiting|3105,3113
,|3113,3114
diarrhea|3115,3123
,|3123,3124
constipation|3125,3137
,|3137,3138
BRBPR|3139,3144
,|3144,3145
melena|3146,3152
,|3152,3153
hematochezia|3154,3166
,|3166,3167
<EOL>|3168,3169
dysuria|3169,3176
,|3176,3177
hematuria|3178,3187
.|3187,3188
<EOL>|3190,3191
<EOL>|3192,3193
Past|3193,3197
Medical|3198,3205
History|3206,3213
:|3213,3214
<EOL>|3214,3215
ASTHMA|3215,3221
/|3221,3222
COPD|3222,3226
<EOL>|3228,3229
ATYPICAL|3229,3237
CHEST|3238,3243
PAIN|3244,3248
<EOL>|3250,3251
CERVICAL|3251,3259
RADICULITIS|3260,3271
<EOL>|3273,3274
CERVICAL|3274,3282
SPONDYLOSIS|3283,3294
<EOL>|3296,3297
CORONARY|3297,3305
ARTERY|3306,3312
DISEASE|3313,3320
<EOL>|3322,3323
HEADACHE|3323,3331
<EOL>|3333,3334
HIP|3334,3337
REPLACEMENT|3338,3349
<EOL>|3351,3352
HYPERLIPIDEMIA|3352,3366
<EOL>|3368,3369
HYPERTENSION|3369,3381
<EOL>|3383,3384
OSTEOARTHRITIS|3384,3398
<EOL>|3400,3401
HERPES|3401,3407
ZOSTER|3408,3414
<EOL>|3416,3417
ATRIAL|3417,3423
FIBRILLATION|3424,3436
<EOL>|3438,3439
ANXIETY|3439,3446
<EOL>|3448,3449
GASTROINTESTINAL|3449,3465
BLEEDING|3466,3474
<EOL>|3476,3477
OSTEOARTHRITIS|3477,3491
<EOL>|3495,3496
PERIPHERAL|3496,3506
VASCULAR|3507,3515
DISEASE|3516,3523
(|3524,3525
s|3525,3526
/|3526,3527
p|3527,3528
bilateral|3529,3538
iliac|3539,3544
stents|3545,3551
)|3551,3552
<EOL>|3552,3553
<EOL>|3554,3555
Social|3555,3561
History|3562,3569
:|3569,3570
<EOL>|3570,3571
_|3571,3572
_|3572,3573
_|3573,3574
<EOL>|3574,3575
Family|3575,3581
History|3582,3589
:|3589,3590
<EOL>|3590,3591
Mother|3591,3597
:|3597,3598
_|3599,3600
_|3600,3601
_|3601,3602
,|3602,3603
HTN|3604,3607
<EOL>|3609,3610
Father|3610,3616
:|3616,3617
_|3618,3619
_|3619,3620
_|3620,3621
CA|3622,3624
<EOL>|3626,3627
Brother|3627,3634
:|3634,3635
CA|3636,3638
?|3638,3639
<EOL>|3641,3642
Brother|3642,3649
:|3649,3650
_|3651,3652
_|3652,3653
_|3653,3654
<EOL>|3655,3656
<EOL>|3657,3658
Physical|3658,3666
_|3667,3668
_|3668,3669
_|3669,3670
:|3670,3671
<EOL>|3671,3672
=|3672,3673
=|3673,3674
=|3674,3675
=|3675,3676
=|3676,3677
=|3677,3678
=|3678,3679
=|3679,3680
=|3680,3681
=|3681,3682
=|3682,3683
=|3683,3684
=|3684,3685
=|3685,3686
=|3686,3687
=|3687,3688
=|3688,3689
<EOL>|3689,3690
ADMISSION|3690,3699
EXAM|3700,3704
:|3704,3705
<EOL>|3705,3706
=|3706,3707
=|3707,3708
=|3708,3709
=|3709,3710
=|3710,3711
=|3711,3712
=|3712,3713
=|3713,3714
=|3714,3715
=|3715,3716
=|3716,3717
=|3717,3718
=|3718,3719
=|3719,3720
=|3720,3721
=|3721,3722
=|3722,3723
<EOL>|3723,3724
Vitals|3724,3730
-|3730,3731
T|3732,3733
98.0|3734,3738
BP|3739,3741
148|3742,3745
/|3745,3746
70|3746,3748
HR|3749,3751
70|3752,3754
RR|3755,3757
24|3758,3760
O2Sat|3761,3766
96|3767,3769
%|3769,3770
on|3771,3773
2L|3774,3776
NC|3777,3779
<EOL>|3781,3782
GENERAL|3782,3789
:|3789,3790
AOx3|3791,3795
,|3795,3796
NAD|3797,3800
,|3800,3801
sitting|3802,3809
up|3810,3812
in|3813,3815
bed|3816,3819
<EOL>|3819,3820
HEENT|3820,3825
:|3825,3826
Normocephalic|3827,3840
,|3840,3841
atraumatic|3842,3852
.|3852,3853
Pupils|3855,3861
equal|3862,3867
,|3867,3868
round|3869,3874
,|3874,3875
and|3876,3879
<EOL>|3880,3881
reactive|3881,3889
bilaterally|3890,3901
,|3901,3902
extraocular|3903,3914
muscles|3915,3922
intact|3923,3929
.|3929,3930
No|3932,3934
<EOL>|3935,3936
conjunctival|3936,3948
pallor|3949,3955
or|3956,3958
injection|3959,3968
,|3968,3969
sclera|3970,3976
anicteric|3977,3986
and|3987,3990
without|3991,3998
<EOL>|3999,4000
injection|4000,4009
.|4009,4010
Moist|4011,4016
mucous|4017,4023
membranes|4024,4033
,|4033,4034
good|4035,4039
dentition|4040,4049
.|4049,4050
Oropharynx|4052,4062
<EOL>|4063,4064
is|4064,4066
clear|4067,4072
.|4072,4073
<EOL>|4073,4074
NECK|4074,4078
:|4078,4079
Supple|4080,4086
.|4086,4087
JVD|4088,4091
not|4092,4095
visualized|4096,4106
.|4106,4107
<EOL>|4107,4108
CARDIAC|4108,4115
:|4115,4116
Irregularly|4117,4128
irregular|4129,4138
,|4138,4139
_|4140,4141
_|4141,4142
_|4142,4143
systolic|4144,4152
murmur|4153,4159
best|4160,4164
at|4165,4167
the|4168,4171
<EOL>|4172,4173
LSB|4173,4176
,|4176,4177
no|4178,4180
rubs|4181,4185
or|4186,4188
gallops|4189,4196
.|4196,4197
<EOL>|4197,4198
LUNGS|4198,4203
:|4203,4204
Poor|4205,4209
air|4210,4213
movement|4214,4222
throughout|4223,4233
.|4233,4234
Mild|4235,4239
diffuse|4240,4247
inspiratory|4248,4259
<EOL>|4260,4261
and|4261,4264
expiratory|4265,4275
wheezes|4276,4283
.|4283,4284
No|4285,4287
use|4288,4291
of|4292,4294
accessory|4295,4304
muscles|4305,4312
of|4313,4315
<EOL>|4316,4317
breathing|4317,4326
.|4326,4327
No|4328,4330
rhonchi|4331,4338
or|4339,4341
rales|4342,4347
.|4347,4348
<EOL>|4348,4349
BACK|4349,4353
:|4353,4354
No|4355,4357
CVA|4358,4361
tenderness|4362,4372
<EOL>|4373,4374
ABDOMEN|4374,4381
:|4381,4382
Normal|4384,4390
bowels|4391,4397
sounds|4398,4404
,|4404,4405
non|4406,4409
distended|4410,4419
,|4419,4420
non-tender|4421,4431
to|4432,4434
<EOL>|4435,4436
deep|4436,4440
palpation|4441,4450
in|4451,4453
all|4454,4457
four|4458,4462
quadrants|4463,4472
.|4472,4473
No|4474,4476
organomegaly|4477,4489
.|4489,4490
<EOL>|4490,4491
EXTREMITIES|4491,4502
:|4502,4503
No|4504,4506
clubbing|4507,4515
or|4516,4518
cyanosis|4519,4527
.|4527,4528
Bilateral|4529,4538
pitting|4539,4546
edema|4547,4552
to|4553,4555
<EOL>|4556,4557
the|4557,4560
mid|4561,4564
shin|4565,4569
.|4569,4570
Pulses|4571,4577
DP|4578,4580
/|4580,4581
Radial|4581,4587
2|4588,4589
+|4589,4590
bilaterally|4591,4602
.|4602,4603
<EOL>|4603,4604
SKIN|4604,4608
:|4608,4609
No|4610,4612
rash|4613,4617
or|4618,4620
ulcers|4621,4627
<EOL>|4627,4628
NEUROLOGIC|4628,4638
:|4638,4639
CN2|4640,4643
-|4643,4644
12|4644,4646
intact|4647,4653
.|4653,4654
Moves|4656,4661
all|4662,4665
extremities|4666,4677
spontaneously|4678,4691
.|4691,4692
<EOL>|4693,4694
Normal|4695,4701
sensation|4702,4711
.|4711,4712
<EOL>|4713,4714
=|4714,4715
=|4715,4716
=|4716,4717
=|4717,4718
=|4718,4719
=|4719,4720
=|4720,4721
=|4721,4722
=|4722,4723
=|4723,4724
=|4724,4725
=|4725,4726
=|4726,4727
=|4727,4728
=|4728,4729
=|4729,4730
=|4730,4731
<EOL>|4731,4732
DISCHARGE|4732,4741
EXAM|4742,4746
:|4746,4747
<EOL>|4747,4748
=|4748,4749
=|4749,4750
=|4750,4751
=|4751,4752
=|4752,4753
=|4753,4754
=|4754,4755
=|4755,4756
=|4756,4757
=|4757,4758
=|4758,4759
=|4759,4760
=|4760,4761
=|4761,4762
=|4762,4763
=|4763,4764
=|4764,4765
<EOL>|4765,4766
Vitals|4766,4772
-|4772,4773
T|4774,4775
98.7|4776,4780
BP|4781,4783
154|4784,4787
/|4787,4788
85|4788,4790
HR|4791,4793
77|4794,4796
RR|4797,4799
18|4800,4802
O2Sat|4803,4808
99|4809,4811
%|4811,4812
on|4813,4815
3L|4816,4818
NC|4819,4821
<EOL>|4823,4824
GENERAL|4824,4831
:|4831,4832
AOx3|4833,4837
,|4837,4838
NAD|4839,4842
,|4842,4843
sitting|4844,4851
up|4852,4854
in|4855,4857
bed|4858,4861
<EOL>|4861,4862
HEENT|4862,4867
:|4867,4868
NCAT|4869,4873
.|4873,4874
PERRL|4876,4881
.|4881,4882
EOMI|4883,4887
.|4887,4888
Sclera|4889,4895
anicteric|4896,4905
and|4906,4909
not|4910,4913
injected|4914,4922
.|4922,4923
<EOL>|4924,4925
MMM|4925,4928
.|4928,4929
Oropharynx|4932,4942
is|4943,4945
clear|4946,4951
.|4951,4952
<EOL>|4952,4953
NECK|4953,4957
:|4957,4958
Supple|4959,4965
.|4965,4966
No|4967,4969
LAD|4970,4973
.|4973,4974
JVP|4975,4978
not|4979,4982
appreciated|4983,4994
at|4995,4997
45|4998,5000
degrees|5001,5008
.|5008,5009
<EOL>|5009,5010
CARDIAC|5010,5017
:|5017,5018
Irregularly|5019,5030
irregular|5031,5040
,|5040,5041
normal|5042,5048
rate|5049,5053
.|5053,5054
_|5055,5056
_|5056,5057
_|5057,5058
systolic|5059,5067
murmur|5068,5074
<EOL>|5075,5076
at|5076,5078
the|5079,5082
RUSB|5083,5087
.|5087,5088
No|5089,5091
rubs|5092,5096
or|5097,5099
gallops|5100,5107
.|5107,5108
<EOL>|5108,5109
LUNGS|5109,5114
:|5114,5115
Poor|5116,5120
air|5121,5124
movement|5125,5133
throughout|5134,5144
all|5145,5148
zones|5149,5154
of|5155,5157
the|5158,5161
lungs|5162,5167
.|5167,5168
No|5169,5171
<EOL>|5172,5173
wheezes|5173,5180
.|5180,5181
No|5182,5184
prolonged|5185,5194
expiratory|5195,5205
phase|5206,5211
.|5211,5212
No|5213,5215
rhonchi|5216,5223
or|5224,5226
rales|5227,5232
.|5232,5233
<EOL>|5234,5235
Does|5235,5239
typically|5240,5249
sit|5250,5253
cross|5254,5259
legged|5260,5266
in|5267,5269
the|5270,5273
bed|5274,5277
with|5278,5282
forearms|5283,5291
on|5292,5294
her|5295,5298
<EOL>|5299,5300
legs|5300,5304
in|5305,5307
a|5308,5309
tripod|5310,5316
position|5317,5325
.|5325,5326
<EOL>|5326,5327
BACK|5327,5331
:|5331,5332
No|5333,5335
CVA|5336,5339
tenderness|5340,5350
.|5350,5351
<EOL>|5352,5353
ABDOMEN|5353,5360
:|5360,5361
+|5363,5364
BS|5364,5366
,|5366,5367
soft|5368,5372
,|5372,5373
nontender|5374,5383
,|5383,5384
nondistended|5385,5397
<EOL>|5397,5398
EXTREMITIES|5398,5409
:|5409,5410
Trace|5411,5416
pitting|5417,5424
edema|5425,5430
to|5431,5433
the|5434,5437
mid|5438,5441
shin|5442,5446
.|5446,5447
2|5448,5449
+|5449,5450
DP|5451,5453
pulses|5454,5460
<EOL>|5461,5462
bilaterally|5462,5473
.|5473,5474
No|5475,5477
TTP|5478,5481
.|5481,5482
<EOL>|5482,5483
SKIN|5483,5487
:|5487,5488
No|5489,5491
rash|5492,5496
or|5497,5499
ulcers|5500,5506
.|5506,5507
<EOL>|5507,5508
NEUROLOGIC|5508,5518
:|5518,5519
CN2|5520,5523
-|5523,5524
12|5524,5526
intact|5527,5533
.|5533,5534
Moves|5536,5541
all|5542,5545
extremities|5546,5557
spontaneously|5558,5571
.|5571,5572
<EOL>|5573,5574
Normal|5575,5581
sensation|5582,5591
.|5591,5592
<EOL>|5593,5594
<EOL>|5595,5596
Pertinent|5596,5605
Results|5606,5613
:|5613,5614
<EOL>|5614,5615
=|5615,5616
=|5616,5617
=|5617,5618
=|5618,5619
=|5619,5620
=|5620,5621
=|5621,5622
=|5622,5623
=|5623,5624
=|5624,5625
=|5625,5626
=|5626,5627
=|5627,5628
=|5628,5629
=|5629,5630
=|5630,5631
=|5631,5632
=|5632,5633
<EOL>|5633,5634
ADMISSION|5634,5643
LABS|5644,5648
:|5648,5649
<EOL>|5649,5650
=|5650,5651
=|5651,5652
=|5652,5653
=|5653,5654
=|5654,5655
=|5655,5656
=|5656,5657
=|5657,5658
=|5658,5659
=|5659,5660
=|5660,5661
=|5661,5662
=|5662,5663
=|5663,5664
=|5664,5665
=|5665,5666
=|5666,5667
=|5667,5668
<EOL>|5668,5669
_|5669,5670
_|5670,5671
_|5671,5672
02|5673,5675
:|5675,5676
27PM|5676,5680
BLOOD|5681,5686
WBC|5687,5690
-|5690,5691
7.4|5691,5694
RBC|5695,5698
-|5698,5699
4|5699,5700
.|5700,5701
57|5701,5703
Hgb|5704,5707
-|5707,5708
12.3|5708,5712
Hct|5713,5716
-|5716,5717
39.3|5717,5721
MCV|5722,5725
-|5725,5726
86|5726,5728
<EOL>|5729,5730
MCH|5730,5733
-|5733,5734
26.9|5734,5738
MCHC|5739,5743
-|5743,5744
31|5744,5746
.|5746,5747
3|5747,5748
*|5748,5749
RDW|5750,5753
-|5753,5754
23|5754,5756
.|5756,5757
6|5757,5758
*|5758,5759
RDWSD|5760,5765
-|5765,5766
70|5766,5768
.|5768,5769
9|5769,5770
*|5770,5771
Plt|5772,5775
_|5776,5777
_|5777,5778
_|5778,5779
<EOL>|5779,5780
_|5780,5781
_|5781,5782
_|5782,5783
02|5784,5786
:|5786,5787
27PM|5787,5791
BLOOD|5792,5797
Neuts|5798,5803
-|5803,5804
86|5804,5806
.|5806,5807
5|5807,5808
*|5808,5809
Lymphs|5810,5816
-|5816,5817
6|5817,5818
.|5818,5819
1|5819,5820
*|5820,5821
Monos|5822,5827
-|5827,5828
6.6|5828,5831
<EOL>|5832,5833
Eos|5833,5836
-|5836,5837
0|5837,5838
.|5838,5839
0|5839,5840
*|5840,5841
Baso|5842,5846
-|5846,5847
0.0|5847,5850
Im|5851,5853
_|5854,5855
_|5855,5856
_|5856,5857
AbsNeut|5858,5865
-|5865,5866
6|5866,5867
.|5867,5868
38|5868,5870
*|5870,5871
AbsLymp|5872,5879
-|5879,5880
0|5880,5881
.|5881,5882
45|5882,5884
*|5884,5885
<EOL>|5886,5887
AbsMono|5887,5894
-|5894,5895
0|5895,5896
.|5896,5897
49|5897,5899
AbsEos|5900,5906
-|5906,5907
0|5907,5908
.|5908,5909
00|5909,5911
*|5911,5912
AbsBaso|5913,5920
-|5920,5921
0|5921,5922
.|5922,5923
00|5923,5925
*|5925,5926
<EOL>|5926,5927
_|5927,5928
_|5928,5929
_|5929,5930
02|5931,5933
:|5933,5934
27PM|5934,5938
BLOOD|5939,5944
Glucose|5945,5952
-|5952,5953
132|5953,5956
*|5956,5957
UreaN|5958,5963
-|5963,5964
17|5964,5966
Creat|5967,5972
-|5972,5973
1.0|5973,5976
Na|5977,5979
-|5979,5980
137|5980,5983
<EOL>|5984,5985
K|5985,5986
-|5986,5987
3.7|5987,5990
Cl|5991,5993
-|5993,5994
93|5994,5996
*|5996,5997
HCO3|5998,6002
-|6002,6003
31|6003,6005
AnGap|6006,6011
-|6011,6012
17|6012,6014
<EOL>|6014,6015
=|6015,6016
=|6016,6017
=|6017,6018
=|6018,6019
=|6019,6020
=|6020,6021
=|6021,6022
=|6022,6023
=|6023,6024
=|6024,6025
=|6025,6026
=|6026,6027
=|6027,6028
=|6028,6029
=|6029,6030
=|6030,6031
=|6031,6032
=|6032,6033
<EOL>|6033,6034
PERTINENT|6034,6043
RESULTS|6044,6051
:|6051,6052
<EOL>|6052,6053
=|6053,6054
=|6054,6055
=|6055,6056
=|6056,6057
=|6057,6058
=|6058,6059
=|6059,6060
=|6060,6061
=|6061,6062
=|6062,6063
=|6063,6064
=|6064,6065
=|6065,6066
=|6066,6067
=|6067,6068
=|6068,6069
=|6069,6070
=|6070,6071
<EOL>|6071,6072
LABS|6072,6076
:|6076,6077
<EOL>|6077,6078
=|6078,6079
=|6079,6080
=|6080,6081
=|6081,6082
=|6082,6083
=|6083,6084
=|6084,6085
=|6085,6086
=|6086,6087
=|6087,6088
=|6088,6089
=|6089,6090
=|6090,6091
=|6091,6092
=|6092,6093
=|6093,6094
=|6094,6095
=|6095,6096
<EOL>|6096,6097
_|6097,6098
_|6098,6099
_|6099,6100
12|6101,6103
:|6103,6104
15AM|6104,6108
BLOOD|6109,6114
_|6115,6116
_|6116,6117
_|6117,6118
pO2|6119,6122
-|6122,6123
103|6123,6126
pCO2|6127,6131
-|6131,6132
49|6132,6134
*|6134,6135
pH|6136,6138
-|6138,6139
7.42|6139,6143
<EOL>|6144,6145
calTCO2|6145,6152
-|6152,6153
33|6153,6155
*|6155,6156
Base|6157,6161
XS|6162,6164
-|6164,6165
5|6165,6166
<EOL>|6166,6167
=|6167,6168
=|6168,6169
=|6169,6170
<EOL>|6170,6171
_|6171,6172
_|6172,6173
_|6173,6174
02|6175,6177
:|6177,6178
27PM|6178,6182
BLOOD|6183,6188
cTropnT|6189,6196
-|6196,6197
0|6197,6198
.|6198,6199
02|6199,6201
*|6201,6202
proBNP|6203,6209
-|6209,6210
235|6210,6213
<EOL>|6213,6214
_|6214,6215
_|6215,6216
_|6216,6217
09|6218,6220
:|6220,6221
05PM|6221,6225
BLOOD|6226,6231
CK|6232,6234
-|6234,6235
MB|6235,6237
-|6237,6238
6|6238,6239
cTropnT|6240,6247
-|6247,6248
<|6248,6249
0|6249,6250
.|6250,6251
01|6251,6253
<EOL>|6253,6254
_|6254,6255
_|6255,6256
_|6256,6257
07|6258,6260
:|6260,6261
45AM|6261,6265
BLOOD|6266,6271
CK|6272,6274
-|6274,6275
MB|6275,6277
-|6277,6278
6|6278,6279
cTropnT|6280,6287
-|6287,6288
0|6288,6289
.|6289,6290
02|6290,6292
*|6292,6293
<EOL>|6293,6294
=|6294,6295
=|6295,6296
=|6296,6297
<EOL>|6297,6298
_|6298,6299
_|6299,6300
_|6300,6301
07|6302,6304
:|6304,6305
45AM|6305,6309
BLOOD|6310,6315
THEOPHYLLINE|6316,6328
-|6328,6329
17.3|6329,6333
(|6334,6335
10.0|6335,6339
-|6339,6340
20.0|6340,6344
)|6344,6345
<EOL>|6345,6346
=|6346,6347
=|6347,6348
=|6348,6349
=|6349,6350
=|6350,6351
=|6351,6352
=|6352,6353
=|6353,6354
=|6354,6355
=|6355,6356
=|6356,6357
=|6357,6358
=|6358,6359
=|6359,6360
=|6360,6361
=|6361,6362
=|6362,6363
=|6363,6364
<EOL>|6364,6365
IMAGING|6365,6372
:|6372,6373
<EOL>|6373,6374
=|6374,6375
=|6375,6376
=|6376,6377
=|6377,6378
=|6378,6379
=|6379,6380
=|6380,6381
=|6381,6382
=|6382,6383
=|6383,6384
=|6384,6385
=|6385,6386
=|6386,6387
=|6387,6388
=|6388,6389
=|6389,6390
=|6390,6391
=|6391,6392
<EOL>|6392,6393
CXR|6393,6396
(|6397,6398
_|6398,6399
_|6399,6400
_|6400,6401
)|6401,6402
:|6402,6403
PA|6404,6406
and|6407,6410
lateral|6411,6418
views|6419,6424
the|6425,6428
chest|6429,6434
provided|6435,6443
.|6443,6444
Biapical|6445,6453
<EOL>|6454,6455
pleural|6455,6462
parenchymal|6463,6474
scarring|6475,6483
noted|6484,6489
.|6489,6490
No|6492,6494
focal|6495,6500
consolidation|6501,6514
<EOL>|6515,6516
concerning|6516,6526
for|6527,6530
pneumonia|6531,6540
.|6540,6541
No|6542,6544
effusion|6545,6553
or|6554,6556
pneumothorax|6557,6569
.|6569,6570
No|6572,6574
signs|6575,6580
<EOL>|6581,6582
of|6582,6584
congestion|6585,6595
or|6596,6598
edema|6599,6604
.|6604,6605
Cardiomediastinal|6606,6623
silhouette|6624,6634
is|6635,6637
stable|6638,6644
<EOL>|6645,6646
with|6646,6650
an|6651,6653
unfolded|6654,6662
thoracic|6663,6671
aorta|6672,6677
and|6678,6681
top|6682,6685
-|6685,6686
normal|6686,6692
heart|6693,6698
size|6699,6703
.|6703,6704
Bony|6705,6709
<EOL>|6710,6711
structures|6711,6721
are|6722,6725
intact|6726,6732
.|6732,6733
<EOL>|6733,6734
=|6734,6735
=|6735,6736
=|6736,6737
<EOL>|6737,6738
CT|6738,6740
Chest|6741,6746
(|6747,6748
_|6748,6749
_|6749,6750
_|6750,6751
)|6751,6752
:|6752,6753
<EOL>|6753,6754
1.|6754,6756
Moderate|6758,6766
upper|6767,6772
lobe|6773,6777
predominant|6778,6789
centrilobular|6790,6803
and|6804,6807
paraseptal|6808,6818
<EOL>|6819,6820
emphysema|6820,6829
.|6829,6830
<EOL>|6830,6831
2.|6831,6833
New|6835,6838
left|6839,6843
lower|6844,6849
lobe|6850,6854
nodule|6855,6861
,|6861,6862
potentially|6863,6874
measuring|6875,6884
as|6885,6887
large|6888,6893
<EOL>|6894,6895
as|6895,6897
6|6898,6899
x|6900,6901
8|6902,6903
mm|6904,6906
,|6906,6907
warrants|6908,6916
close|6917,6922
follow|6923,6929
-|6929,6930
up|6930,6932
.|6932,6933
Stable|6935,6941
to|6942,6944
slightly|6945,6953
<EOL>|6954,6955
smaller|6955,6962
4|6963,6964
mm|6965,6967
right|6968,6973
middle|6974,6980
lobe|6981,6985
nodule|6986,6992
.|6992,6993
<EOL>|6993,6994
3.|6994,6996
Severe|6998,7004
coronary|7005,7013
artery|7014,7020
calcifications|7021,7035
.|7035,7036
Aortic|7038,7044
valve|7045,7050
<EOL>|7051,7052
calcifications|7052,7066
.|7066,7067
<EOL>|7068,7069
4.|7069,7071
Enlargement|7073,7084
of|7085,7087
the|7088,7091
main|7092,7096
and|7097,7100
right|7101,7106
pulmonary|7107,7116
arteries|7117,7125
is|7126,7128
<EOL>|7129,7130
suggestive|7130,7140
of|7141,7143
chronic|7144,7151
pulmonary|7152,7161
arterial|7162,7170
hypertension|7171,7183
.|7183,7184
<EOL>|7185,7186
5.|7186,7188
Fusiform|7190,7198
aneurysmal|7199,7209
dilatation|7210,7220
of|7221,7223
the|7224,7227
abdominal|7228,7237
aorta|7238,7243
<EOL>|7244,7245
measuring|7245,7254
up|7255,7257
to|7258,7260
3.7|7261,7264
cm|7265,7267
has|7268,7271
progressed|7272,7282
compared|7283,7291
to|7292,7294
prior|7295,7300
<EOL>|7301,7302
examination|7302,7313
.|7313,7314
<EOL>|7314,7315
=|7315,7316
=|7316,7317
=|7317,7318
=|7318,7319
=|7319,7320
=|7320,7321
=|7321,7322
=|7322,7323
=|7323,7324
=|7324,7325
=|7325,7326
=|7326,7327
=|7327,7328
=|7328,7329
=|7329,7330
=|7330,7331
=|7331,7332
=|7332,7333
<EOL>|7333,7334
DISCHARGE|7334,7343
LABS|7344,7348
:|7348,7349
<EOL>|7349,7350
=|7350,7351
=|7351,7352
=|7352,7353
=|7353,7354
=|7354,7355
=|7355,7356
=|7356,7357
=|7357,7358
=|7358,7359
=|7359,7360
=|7360,7361
=|7361,7362
=|7362,7363
=|7363,7364
=|7364,7365
=|7365,7366
=|7366,7367
=|7367,7368
<EOL>|7368,7369
_|7369,7370
_|7370,7371
_|7371,7372
07|7373,7375
:|7375,7376
45AM|7376,7380
BLOOD|7381,7386
WBC|7387,7390
-|7390,7391
7.8|7391,7394
RBC|7395,7398
-|7398,7399
4|7399,7400
.|7400,7401
74|7401,7403
Hgb|7404,7407
-|7407,7408
12.7|7408,7412
Hct|7413,7416
-|7416,7417
41.0|7417,7421
MCV|7422,7425
-|7425,7426
87|7426,7428
<EOL>|7429,7430
MCH|7430,7433
-|7433,7434
26.8|7434,7438
MCHC|7439,7443
-|7443,7444
31|7444,7446
.|7446,7447
0|7447,7448
*|7448,7449
RDW|7450,7453
-|7453,7454
23|7454,7456
.|7456,7457
7|7457,7458
*|7458,7459
RDWSD|7460,7465
-|7465,7466
71|7466,7468
.|7468,7469
7|7469,7470
*|7470,7471
Plt|7472,7475
_|7476,7477
_|7477,7478
_|7478,7479
<EOL>|7479,7480
_|7480,7481
_|7481,7482
_|7482,7483
07|7484,7486
:|7486,7487
45AM|7487,7491
BLOOD|7492,7497
Glucose|7498,7505
-|7505,7506
94|7506,7508
UreaN|7509,7514
-|7514,7515
18|7515,7517
Creat|7518,7523
-|7523,7524
1.0|7524,7527
Na|7528,7530
-|7530,7531
135|7531,7534
<EOL>|7535,7536
K|7536,7537
-|7537,7538
3.3|7538,7541
Cl|7542,7544
-|7544,7545
93|7545,7547
*|7547,7548
HCO3|7549,7553
-|7553,7554
31|7554,7556
AnGap|7557,7562
-|7562,7563
14|7563,7565
<EOL>|7565,7566
_|7566,7567
_|7567,7568
_|7568,7569
07|7570,7572
:|7572,7573
45AM|7573,7577
BLOOD|7578,7583
Calcium|7584,7591
-|7591,7592
9.8|7592,7595
Phos|7596,7600
-|7600,7601
2.8|7601,7604
Mg|7605,7607
-|7607,7608
2.0|7608,7611
<EOL>|7611,7612
<EOL>|7613,7614
Brief|7614,7619
Hospital|7620,7628
Course|7629,7635
:|7635,7636
<EOL>|7636,7637
Ms.|7637,7640
_|7641,7642
_|7642,7643
_|7643,7644
is|7645,7647
a|7648,7649
_|7650,7651
_|7651,7652
_|7652,7653
y|7654,7655
/|7655,7656
o|7656,7657
woman|7658,7663
with|7664,7668
a|7669,7670
PMH|7671,7674
notable|7675,7682
for|7683,7686
COPD|7687,7691
on|7692,7694
<EOL>|7695,7696
home|7696,7700
O2|7701,7703
(|7704,7705
hospitalized|7705,7717
_|7718,7719
_|7719,7720
_|7720,7721
,|7721,7722
multiple|7723,7731
recent|7732,7738
ED|7739,7741
visits|7742,7748
)|7748,7749
,|7749,7750
Afib|7751,7755
<EOL>|7756,7757
on|7757,7759
apixaban|7760,7768
,|7768,7769
HTN|7770,7773
,|7773,7774
CAD|7775,7778
,|7778,7779
and|7780,7783
HLD|7784,7787
who|7788,7791
presented|7792,7801
with|7802,7806
dyspnea|7807,7814
and|7815,7818
<EOL>|7819,7820
orthopnea|7820,7829
in|7830,7832
the|7833,7836
setting|7837,7844
of|7845,7847
a|7848,7849
steroid|7850,7857
taper|7858,7863
for|7864,7867
recent|7868,7874
COPD|7875,7879
<EOL>|7880,7881
exacerbation|7881,7893
.|7893,7894
Her|7895,7898
dyspnea|7899,7906
was|7907,7910
thought|7911,7918
to|7919,7921
be|7922,7924
multifactorial|7925,7939
due|7940,7943
<EOL>|7944,7945
to|7945,7947
her|7948,7951
severe|7952,7958
COPD|7959,7963
and|7964,7967
with|7968,7972
a|7973,7974
component|7975,7984
of|7985,7987
anxiety|7988,7995
.|7995,7996
The|7997,8000
patient|8001,8008
<EOL>|8009,8010
was|8010,8013
not|8014,8017
thought|8018,8025
to|8026,8028
be|8029,8031
having|8032,8038
an|8039,8041
acute|8042,8047
COPD|8048,8052
exacerbation|8053,8065
.|8065,8066
<EOL>|8066,8067
<EOL>|8067,8068
=|8068,8069
=|8069,8070
=|8070,8071
=|8071,8072
=|8072,8073
=|8073,8074
=|8074,8075
=|8075,8076
=|8076,8077
=|8077,8078
=|8078,8079
=|8079,8080
=|8080,8081
=|8081,8082
=|8082,8083
=|8083,8084
<EOL>|8084,8085
ACTIVE|8085,8091
ISSUES|8092,8098
:|8098,8099
<EOL>|8099,8100
=|8100,8101
=|8101,8102
=|8102,8103
=|8103,8104
=|8104,8105
=|8105,8106
=|8106,8107
=|8107,8108
=|8108,8109
=|8109,8110
=|8110,8111
=|8111,8112
=|8112,8113
=|8113,8114
=|8114,8115
=|8115,8116
<EOL>|8116,8117
<EOL>|8117,8118
#|8118,8119
Dyspnea|8120,8127
:|8127,8128
Patient|8129,8136
was|8137,8140
admitted|8141,8149
after|8150,8155
one|8156,8159
night|8160,8165
of|8166,8168
worsened|8169,8177
<EOL>|8178,8179
orthopnea|8179,8188
and|8189,8192
dyspnea|8193,8200
in|8201,8203
the|8204,8207
setting|8208,8215
of|8216,8218
a|8219,8220
steroid|8221,8228
taper|8229,8234
from|8235,8239
30|8240,8242
<EOL>|8243,8244
mg|8244,8246
to|8247,8249
25|8250,8252
mg|8253,8255
.|8255,8256
Her|8257,8260
dyspnea|8261,8268
was|8269,8272
thought|8273,8280
to|8281,8283
be|8284,8286
multifactorial|8287,8301
due|8302,8305
to|8306,8308
<EOL>|8309,8310
her|8310,8313
severe|8314,8320
COPD|8321,8325
and|8326,8329
with|8330,8334
a|8335,8336
component|8337,8346
of|8347,8349
anxiety|8350,8357
.|8357,8358
The|8359,8362
patient|8363,8370
was|8371,8374
<EOL>|8375,8376
not|8376,8379
thought|8380,8387
to|8388,8390
be|8391,8393
having|8394,8400
an|8401,8403
acute|8404,8409
COPD|8410,8414
exacerbation|8415,8427
.|8427,8428
The|8429,8432
patient|8433,8440
<EOL>|8441,8442
was|8442,8445
treated|8446,8453
with|8454,8458
occasional|8459,8469
duonebs|8470,8477
and|8478,8481
lorazepam|8482,8491
0.5|8492,8495
mg|8496,8498
PRN|8499,8502
<EOL>|8503,8504
that|8504,8508
helped|8509,8515
relieve|8516,8523
her|8524,8527
dyspnea|8528,8535
.|8535,8536
Pulmonology|8537,8548
was|8549,8552
consulted|8553,8562
.|8562,8563
The|8564,8567
<EOL>|8568,8569
patient|8569,8576
underwent|8577,8586
CT|8587,8589
that|8590,8594
showed|8595,8601
emphysema|8602,8611
but|8612,8615
no|8616,8618
evidence|8619,8627
of|8628,8630
<EOL>|8631,8632
infection|8632,8641
such|8642,8646
as|8647,8649
_|8650,8651
_|8651,8652
_|8652,8653
.|8653,8654
The|8655,8658
patient|8659,8666
was|8667,8670
initiated|8671,8680
on|8681,8683
a|8684,8685
steroid|8686,8693
<EOL>|8694,8695
taper|8695,8700
on|8701,8703
_|8704,8705
_|8705,8706
_|8706,8707
of|8708,8710
prednisone|8711,8721
30|8722,8724
mg|8725,8727
for|8728,8731
3|8732,8733
days|8734,8738
,|8738,8739
then|8740,8744
20|8745,8747
mg|8748,8750
for|8751,8754
3|8755,8756
<EOL>|8757,8758
days|8758,8762
,|8762,8763
then|8764,8768
10|8769,8771
mg|8772,8774
until|8775,8780
outpatient|8781,8791
follow|8792,8798
-|8798,8799
up|8799,8801
.|8801,8802
Pulmonology|8803,8814
<EOL>|8815,8816
recommended|8816,8827
increasing|8828,8838
her|8839,8842
Advair|8843,8849
dose|8850,8854
to|8855,8857
500|8858,8861
/|8861,8862
50|8862,8864
,|8864,8865
which|8866,8871
was|8872,8875
<EOL>|8876,8877
done|8877,8881
.|8881,8882
They|8883,8887
also|8888,8892
recommended|8893,8904
switching|8905,8914
from|8915,8919
theophylline|8920,8932
to|8933,8935
<EOL>|8936,8937
roflumilast|8937,8948
and|8949,8952
initiation|8953,8963
of|8964,8966
long|8967,8971
-|8971,8972
term|8972,8976
azithromycin|8977,8989
therapy|8990,8997
<EOL>|8998,8999
provided|8999,9007
the|9008,9011
patient|9012,9019
's|9019,9021
QTc|9022,9025
was|9026,9029
not|9030,9033
prolonged|9034,9043
;|9043,9044
this|9045,9049
was|9050,9053
deferred|9054,9062
<EOL>|9063,9064
to|9064,9066
the|9067,9070
outpatient|9071,9081
setting|9082,9089
.|9089,9090
Throughout|9091,9101
her|9102,9105
admission|9106,9115
she|9116,9119
had|9120,9123
O2|9124,9126
<EOL>|9127,9128
sats|9128,9132
greater|9133,9140
than|9141,9145
95|9146,9148
%|9148,9149
on|9150,9152
2L|9153,9155
NC|9156,9158
.|9158,9159
She|9160,9163
did|9164,9167
not|9168,9171
desaturate|9172,9182
on|9183,9185
<EOL>|9186,9187
ambulation|9187,9197
.|9197,9198
<EOL>|9199,9200
<EOL>|9200,9201
#|9201,9202
Anxiety|9203,9210
/|9210,9211
Insomnia|9211,9219
:|9219,9220
Patient|9221,9228
with|9229,9233
a|9234,9235
history|9236,9243
of|9244,9246
anxiety|9247,9254
and|9255,9258
<EOL>|9259,9260
insomnia|9260,9268
,|9268,9269
thought|9270,9277
to|9278,9280
be|9281,9283
contributing|9284,9296
to|9297,9299
her|9300,9303
experience|9304,9314
of|9315,9317
<EOL>|9318,9319
dyspnea|9319,9326
.|9326,9327
The|9328,9331
patient|9332,9339
was|9340,9343
discharged|9344,9354
with|9355,9359
lorazepam|9360,9369
Q8H|9370,9373
as|9374,9376
needed|9377,9383
<EOL>|9384,9385
for|9385,9388
anxiety|9389,9396
.|9396,9397
The|9398,9401
patient|9402,9409
would|9410,9415
likely|9416,9422
benefit|9423,9430
from|9431,9435
therapy|9436,9443
with|9444,9448
<EOL>|9449,9450
an|9450,9452
SSRI|9453,9457
.|9457,9458
<EOL>|9458,9459
<EOL>|9459,9460
#|9460,9461
Demand|9462,9468
Ischemia|9469,9477
:|9477,9478
Patient|9479,9486
with|9487,9491
troponin|9492,9500
0.02|9501,9505
,|9505,9506
<|9507,9508
0.01|9508,9512
,|9512,9513
then|9514,9518
0.02|9519,9523
.|9523,9524
<EOL>|9525,9526
ECG|9526,9529
without|9530,9537
acute|9538,9543
ischemic|9544,9552
changes|9553,9560
.|9560,9561
<EOL>|9561,9562
<EOL>|9562,9563
#|9563,9564
Microscopic|9565,9576
hematuria|9577,9586
:|9586,9587
On|9588,9590
admission|9591,9600
the|9601,9604
patient|9605,9612
had|9613,9616
a|9617,9618
UA|9619,9621
with|9622,9626
<EOL>|9627,9628
40|9628,9630
RBCs|9631,9635
.|9635,9636
Occasional|9637,9647
UAs|9648,9651
over|9652,9656
the|9657,9660
last|9661,9665
year|9666,9670
in|9671,9673
OMR|9674,9677
with|9678,9682
<EOL>|9683,9684
microscopic|9684,9695
hematuria|9696,9705
.|9705,9706
Would|9707,9712
recommend|9713,9722
repeat|9723,9729
UA|9730,9732
as|9733,9735
an|9736,9738
<EOL>|9739,9740
outpatient|9740,9750
or|9751,9753
work|9754,9758
-|9758,9759
up|9759,9761
for|9762,9765
microscopic|9766,9777
hematuria|9778,9787
.|9787,9788
<EOL>|9788,9789
<EOL>|9789,9790
=|9790,9791
=|9791,9792
=|9792,9793
=|9793,9794
=|9794,9795
=|9795,9796
=|9796,9797
=|9797,9798
=|9798,9799
=|9799,9800
=|9800,9801
=|9801,9802
=|9802,9803
=|9803,9804
=|9804,9805
=|9805,9806
<EOL>|9806,9807
CHRONIC|9807,9814
ISSUES|9815,9821
:|9821,9822
<EOL>|9822,9823
=|9823,9824
=|9824,9825
=|9825,9826
=|9826,9827
=|9827,9828
=|9828,9829
=|9829,9830
=|9830,9831
=|9831,9832
=|9832,9833
=|9833,9834
=|9834,9835
=|9835,9836
=|9836,9837
=|9837,9838
=|9838,9839
<EOL>|9839,9840
<EOL>|9840,9841
#|9841,9842
Smoking|9843,9850
:|9850,9851
Patient|9852,9859
recently|9860,9868
quit|9869,9873
smoking|9874,9881
one|9882,9885
month|9886,9891
ago|9892,9895
.|9895,9896
Patient|9897,9904
<EOL>|9905,9906
was|9906,9909
provided|9910,9918
with|9919,9923
a|9924,9925
nicotine|9926,9934
patch|9935,9940
7|9941,9942
mg|9943,9945
while|9946,9951
in|9952,9954
house|9955,9960
;|9960,9961
could|9962,9967
<EOL>|9968,9969
consider|9969,9977
continuing|9978,9988
as|9989,9991
an|9992,9994
outpatient|9995,10005
if|10006,10008
patient|10009,10016
endorses|10017,10025
<EOL>|10026,10027
cravings|10027,10035
.|10035,10036
<EOL>|10036,10037
<EOL>|10037,10038
#|10038,10039
Atrial|10040,10046
fibrillation|10047,10059
:|10059,10060
Patient|10061,10068
continued|10069,10078
on|10079,10081
diltiazem|10082,10091
240|10092,10095
mg|10096,10098
PO|10099,10101
<EOL>|10102,10103
BID|10103,10106
and|10107,10110
apixaban|10111,10119
5|10120,10121
mg|10122,10124
BID|10125,10128
.|10128,10129
<EOL>|10129,10130
<EOL>|10130,10131
#|10131,10132
HTN|10133,10136
:|10136,10137
Patient|10138,10145
with|10146,10150
a|10151,10152
history|10153,10160
of|10161,10163
hypertension|10164,10176
.|10176,10177
Blood|10178,10183
pressure|10184,10192
<EOL>|10193,10194
well|10194,10198
-|10198,10199
controlled|10199,10209
.|10209,10210
Continued|10211,10220
on|10221,10223
isosorbide|10224,10234
mononitrate|10235,10246
ER|10247,10249
240|10250,10253
mg|10254,10256
<EOL>|10257,10258
PO|10258,10260
daily|10261,10266
and|10267,10270
hydrochlorothiazide|10271,10290
50|10291,10293
mg|10294,10296
PO|10297,10299
daily|10300,10305
.|10305,10306
<EOL>|10306,10307
<EOL>|10307,10308
#|10308,10309
CAD|10310,10313
:|10313,10314
Cardiac|10315,10322
catheterization|10323,10338
in|10339,10341
_|10342,10343
_|10343,10344
_|10344,10345
without|10346,10353
evidence|10354,10362
of|10363,10365
<EOL>|10366,10367
significant|10367,10378
stenosis|10379,10387
of|10388,10390
coronaries|10391,10401
.|10401,10402
ECHO|10403,10407
on|10408,10410
_|10411,10412
_|10412,10413
_|10413,10414
with|10415,10419
EF|10420,10422
>|10422,10423
55|10423,10425
%|10425,10426
<EOL>|10427,10428
and|10428,10431
no|10432,10434
regional|10435,10443
or|10444,10446
global|10447,10453
wall|10454,10458
motion|10459,10465
abnormalities|10466,10479
.|10479,10480
The|10481,10484
patient|10485,10492
<EOL>|10493,10494
was|10494,10497
continued|10498,10507
on|10508,10510
aspirin|10511,10518
81|10519,10521
mg|10522,10524
daily|10525,10530
and|10531,10534
atorvastatin|10535,10547
10|10548,10550
mg|10551,10553
QPM|10554,10557
.|10557,10558
<EOL>|10558,10559
<EOL>|10559,10560
=|10560,10561
=|10561,10562
=|10562,10563
=|10563,10564
=|10564,10565
=|10565,10566
=|10566,10567
=|10567,10568
=|10568,10569
=|10569,10570
=|10570,10571
=|10571,10572
=|10572,10573
=|10573,10574
=|10574,10575
=|10575,10576
=|10576,10577
=|10577,10578
=|10578,10579
<EOL>|10579,10580
TRANSITIONAL|10580,10592
ISSUES|10593,10599
:|10599,10600
<EOL>|10600,10601
=|10601,10602
=|10602,10603
=|10603,10604
=|10604,10605
=|10605,10606
=|10606,10607
=|10607,10608
=|10608,10609
=|10609,10610
=|10610,10611
=|10611,10612
=|10612,10613
=|10613,10614
=|10614,10615
=|10615,10616
=|10616,10617
=|10617,10618
=|10618,10619
=|10619,10620
<EOL>|10620,10621
#|10621,10622
New|10622,10625
Medications|10626,10637
:|10637,10638
<EOL>|10638,10639
-|10639,10640
Prednisone|10640,10650
30|10651,10653
mg|10654,10656
PO|10657,10659
QD|10660,10662
through|10663,10670
_|10671,10672
_|10672,10673
_|10673,10674
,|10674,10675
then|10676,10680
on|10681,10683
_|10684,10685
_|10685,10686
_|10686,10687
mg|10688,10690
for|10691,10694
3|10695,10696
<EOL>|10697,10698
days|10698,10702
,|10702,10703
then|10704,10708
on|10709,10711
_|10712,10713
_|10713,10714
_|10714,10715
mg|10716,10718
until|10719,10724
outpatient|10725,10735
follow|10736,10742
-|10742,10743
up|10743,10745
<EOL>|10745,10746
-|10746,10747
Increased|10747,10756
Advair|10757,10763
(|10764,10765
Fluticasone|10765,10776
-|10776,10777
Salmeterol|10777,10787
)|10787,10788
to|10789,10791
500|10792,10795
/|10795,10796
50|10796,10798
dose|10799,10803
<EOL>|10803,10804
-|10804,10805
Lorazepam|10805,10814
0.5|10815,10818
mg|10819,10821
PO|10822,10824
Q8H|10825,10828
PRN|10829,10832
for|10833,10836
anxiety|10837,10844
<EOL>|10844,10845
<EOL>|10845,10846
#|10846,10847
Follow|10847,10853
-|10853,10854
up|10854,10856
:|10856,10857
<EOL>|10857,10858
-|10858,10859
Appointment|10859,10870
arranged|10871,10879
with|10880,10884
PCP|10885,10888
,|10888,10889
_|10890,10891
_|10891,10892
_|10892,10893
_|10894,10895
_|10895,10896
_|10896,10897
<EOL>|10897,10898
-|10898,10899
Appointment|10899,10910
arranged|10911,10919
with|10920,10924
Pulmonologist|10925,10938
,|10938,10939
Dr.|10940,10943
_|10944,10945
_|10945,10946
_|10946,10947
,|10947,10948
_|10949,10950
_|10950,10951
_|10951,10952
<EOL>|10952,10953
<EOL>|10953,10954
#|10954,10955
COPD|10955,10959
:|10959,10960
Patient|10961,10968
was|10969,10972
seen|10973,10977
by|10978,10980
pulmonology|10981,10992
during|10993,10999
admission|11000,11009
who|11010,11013
had|11014,11017
<EOL>|11018,11019
the|11019,11022
following|11023,11032
recommendations|11033,11048
to|11049,11051
consider|11052,11060
as|11061,11063
an|11064,11066
outpatient|11067,11077
.|11077,11078
<EOL>|11078,11079
-|11079,11080
Switch|11080,11086
to|11087,11089
roflumilast|11090,11101
from|11102,11106
theophylline|11107,11119
<EOL>|11119,11120
-|11120,11121
Daily|11121,11126
azithromycin|11127,11139
for|11140,11143
treatment|11144,11153
of|11154,11156
chronic|11157,11164
inflammation|11165,11177
<EOL>|11178,11179
provided|11179,11187
QTc|11188,11191
within|11192,11198
normal|11199,11205
limits|11206,11212
.|11212,11213
<EOL>|11213,11214
-|11214,11215
Patient|11215,11222
may|11223,11226
benefit|11227,11234
from|11235,11239
treatment|11240,11249
of|11250,11252
anxiety|11253,11260
with|11261,11265
an|11266,11268
SSRI|11269,11273
,|11273,11274
as|11275,11277
<EOL>|11278,11279
her|11279,11282
anxiety|11283,11290
is|11291,11293
likely|11294,11300
contributing|11301,11313
to|11314,11316
her|11317,11320
experience|11321,11331
of|11332,11334
dyspnea|11335,11342
.|11342,11343
<EOL>|11343,11344
-|11344,11345
In|11345,11347
the|11348,11351
future|11352,11358
,|11358,11359
palliative|11360,11370
care|11371,11375
consult|11376,11383
for|11384,11387
consideration|11388,11401
of|11402,11404
<EOL>|11405,11406
opioid|11406,11412
treatment|11413,11422
of|11423,11425
dyspnea|11426,11433
<EOL>|11433,11434
<EOL>|11434,11435
#|11435,11436
Microscopic|11436,11447
hematuria|11448,11457
:|11457,11458
Patient|11459,11466
had|11467,11470
a|11471,11472
UA|11473,11475
with|11476,11480
40|11481,11483
RBCs|11484,11488
on|11489,11491
<EOL>|11492,11493
admission|11493,11502
<EOL>|11503,11504
-|11504,11505
Recommend|11505,11514
repeat|11515,11521
UA|11522,11524
as|11525,11527
an|11528,11530
outpatient|11531,11541
or|11542,11544
work|11545,11549
-|11549,11550
up|11550,11552
for|11553,11556
microscopic|11557,11568
<EOL>|11569,11570
hematuria|11570,11579
<EOL>|11579,11580
<EOL>|11580,11581
#|11581,11582
Lung|11582,11586
nodule|11587,11593
:|11593,11594
New|11595,11598
left|11599,11603
lower|11604,11609
lobe|11610,11614
nodule|11615,11621
,|11621,11622
potentially|11623,11634
measuring|11635,11644
<EOL>|11645,11646
as|11646,11648
large|11649,11654
as|11655,11657
6|11658,11659
x|11660,11661
8|11662,11663
mm|11664,11666
,|11666,11667
warrants|11668,11676
close|11677,11682
follow|11683,11689
-|11689,11690
up|11690,11692
.|11692,11693
Stable|11695,11701
to|11702,11704
<EOL>|11705,11706
slightly|11706,11714
smaller|11715,11722
4|11723,11724
mm|11725,11727
right|11728,11733
middle|11734,11740
lobe|11741,11745
nodule|11746,11752
.|11752,11753
Follow|11754,11760
-|11760,11761
up|11761,11763
CT|11764,11766
in|11767,11769
<EOL>|11770,11771
_|11771,11772
_|11772,11773
_|11773,11774
months|11775,11781
as|11782,11784
per|11785,11788
_|11789,11790
_|11790,11791
_|11791,11792
guidelines|11793,11803
for|11804,11807
evaluation|11808,11818
<EOL>|11819,11820
of|11820,11822
new|11823,11826
left|11827,11831
lower|11832,11837
lobe|11838,11842
pulmonary|11843,11852
nodule|11853,11859
.|11859,11860
<EOL>|11860,11861
<EOL>|11861,11862
#|11862,11863
Code|11863,11867
Status|11868,11874
:|11874,11875
Full|11876,11880
code|11881,11885
<EOL>|11885,11886
#|11886,11887
Emergency|11887,11896
Contact|11897,11904
/|11904,11905
HCP|11905,11908
:|11908,11909
_|11910,11911
_|11911,11912
_|11912,11913
(|11914,11915
HUSBAND|11915,11922
)|11922,11923
_|11924,11925
_|11925,11926
_|11926,11927
<EOL>|11927,11928
<EOL>|11929,11930
Medications|11930,11941
on|11942,11944
Admission|11945,11954
:|11954,11955
<EOL>|11955,11956
The|11956,11959
Preadmission|11960,11972
Medication|11973,11983
list|11984,11988
is|11989,11991
accurate|11992,12000
and|12001,12004
complete|12005,12013
.|12013,12014
<EOL>|12014,12015
1.|12015,12017
PredniSONE|12018,12028
5|12029,12030
mg|12031,12033
PO|12034,12036
DAILY|12037,12042
<EOL>|12043,12044
Tapered|12044,12051
dose|12052,12056
-|12057,12058
DOWN|12059,12063
<EOL>|12064,12065
2.|12065,12067
Acetaminophen|12068,12081
325|12082,12085
mg|12086,12088
PO|12089,12091
Q4H|12092,12095
:|12095,12096
PRN|12096,12099
Pain|12100,12104
<EOL>|12105,12106
3.|12106,12108
Ipratropium|12109,12120
Bromide|12121,12128
Neb|12129,12132
1|12133,12134
NEB|12135,12138
IH|12139,12141
Q6H|12142,12145
:|12145,12146
PRN|12146,12149
Wheezing|12150,12158
<EOL>|12159,12160
4.|12160,12162
Tiotropium|12163,12173
Bromide|12174,12181
1|12182,12183
CAP|12184,12187
IH|12188,12190
DAILY|12191,12196
<EOL>|12197,12198
5.|12198,12200
Guaifenesin|12201,12212
1|12213,12214
teaspoon|12215,12223
PO|12224,12226
Q3H|12227,12230
:|12230,12231
PRN|12231,12234
cough|12235,12240
<EOL>|12241,12242
6.|12242,12244
Lorazepam|12245,12254
0.5|12255,12258
mg|12259,12261
PO|12262,12264
QHS|12265,12268
vertigo|12269,12276
/|12276,12277
insomnia|12277,12285
<EOL>|12286,12287
7.|12287,12289
Diltiazem|12290,12299
Extended|12300,12308
-|12308,12309
Release|12309,12316
240|12317,12320
mg|12321,12323
PO|12324,12326
BID|12327,12330
<EOL>|12331,12332
8.|12332,12334
Dorzolamide|12335,12346
2|12347,12348
%|12348,12349
Ophth|12350,12355
.|12355,12356
Soln.|12357,12362
1|12363,12364
DROP|12365,12369
BOTH|12370,12374
EYES|12375,12379
BID|12380,12383
<EOL>|12384,12385
9.|12385,12387
Docusate|12388,12396
Sodium|12397,12403
100|12404,12407
mg|12408,12410
PO|12411,12413
BID|12414,12417
<EOL>|12418,12419
10.|12419,12422
Fluticasone|12423,12434
Propionate|12435,12445
NASAL|12446,12451
2|12452,12453
SPRY|12454,12458
NU|12459,12461
DAILY|12462,12467
:|12467,12468
PRN|12468,12471
allergies|12472,12481
<EOL>|12482,12483
11|12483,12485
.|12485,12486
Apixaban|12487,12495
5|12496,12497
mg|12498,12500
PO|12501,12503
BID|12504,12507
<EOL>|12508,12509
12.|12509,12512
Ranitidine|12513,12523
300|12524,12527
mg|12528,12530
PO|12531,12533
DAILY|12534,12539
<EOL>|12540,12541
13.|12541,12544
Atorvastatin|12545,12557
10|12558,12560
mg|12561,12563
PO|12564,12566
QPM|12567,12570
<EOL>|12571,12572
14.|12572,12575
Ferrous|12576,12583
Sulfate|12584,12591
325|12592,12595
mg|12596,12598
PO|12599,12601
DAILY|12602,12607
<EOL>|12608,12609
15.|12609,12612
Multivitamins|12613,12626
1|12627,12628
TAB|12629,12632
PO|12633,12635
DAILY|12636,12641
<EOL>|12642,12643
16|12643,12645
.|12645,12646
Isosorbide|12647,12657
Mononitrate|12658,12669
(|12670,12671
Extended|12671,12679
Release|12680,12687
)|12687,12688
240|12689,12692
mg|12693,12695
PO|12696,12698
DAILY|12699,12704
<EOL>|12705,12706
17.|12706,12709
Fluticasone|12710,12721
-|12721,12722
Salmeterol|12722,12732
Diskus|12733,12739
(|12740,12741
250|12741,12744
/|12744,12745
50|12745,12747
)|12747,12748
1|12750,12751
INH|12752,12755
IH|12756,12758
BID|12759,12762
<EOL>|12763,12764
18.|12764,12767
Latanoprost|12768,12779
0.005|12780,12785
%|12785,12786
Ophth|12787,12792
.|12792,12793
Soln.|12794,12799
1|12800,12801
DROP|12802,12806
BOTH|12807,12811
EYES|12812,12816
QHS|12817,12820
<EOL>|12821,12822
19|12822,12824
.|12824,12825
Calcitrate|12826,12836
-|12836,12837
Vitamin|12837,12844
D|12845,12846
(|12847,12848
calcium|12848,12855
citrate|12856,12863
-|12863,12864
vitamin|12864,12871
D3|12872,12874
)|12874,12875
315|12876,12879
mg|12880,12882
-|12883,12884
<EOL>|12885,12886
200|12886,12889
units|12890,12895
oral|12897,12901
DAILY|12902,12907
<EOL>|12908,12909
20|12909,12911
.|12911,12912
Theophylline|12913,12925
SR|12926,12928
300|12929,12932
mg|12933,12935
PO|12936,12938
BID|12939,12942
<EOL>|12943,12944
21|12944,12946
.|12946,12947
Aspirin|12948,12955
81|12956,12958
mg|12959,12961
PO|12962,12964
DAILY|12965,12970
<EOL>|12971,12972
22.|12972,12975
albuterol|12976,12985
sulfate|12986,12993
90|12994,12996
mcg|12997,13000
/|13000,13001
actuation|13001,13010
inhalation|13011,13021
Q4H|13022,13025
<EOL>|13026,13027
23|13027,13029
.|13029,13030
Hydrochlorothiazide|13031,13050
50|13051,13053
mg|13054,13056
PO|13057,13059
DAILY|13060,13065
<EOL>|13066,13067
24.|13067,13070
cod|13071,13074
liver|13075,13080
oil|13081,13084
1|13085,13086
capsule|13087,13094
oral|13096,13100
BID|13101,13104
<EOL>|13105,13106
<EOL>|13106,13107
<EOL>|13108,13109
Discharge|13109,13118
Medications|13119,13130
:|13130,13131
<EOL>|13131,13132
1.|13132,13134
Acetaminophen|13135,13148
325|13149,13152
mg|13153,13155
PO|13156,13158
Q4H|13159,13162
:|13162,13163
PRN|13163,13166
Pain|13167,13171
<EOL>|13172,13173
2.|13173,13175
Apixaban|13176,13184
5|13185,13186
mg|13187,13189
PO|13190,13192
BID|13193,13196
<EOL>|13197,13198
3.|13198,13200
Aspirin|13201,13208
81|13209,13211
mg|13212,13214
PO|13215,13217
DAILY|13218,13223
<EOL>|13224,13225
4.|13225,13227
Atorvastatin|13228,13240
10|13241,13243
mg|13244,13246
PO|13247,13249
QPM|13250,13253
<EOL>|13254,13255
5.|13255,13257
Diltiazem|13258,13267
Extended|13268,13276
-|13276,13277
Release|13277,13284
240|13285,13288
mg|13289,13291
PO|13292,13294
BID|13295,13298
<EOL>|13299,13300
6.|13300,13302
Docusate|13303,13311
Sodium|13312,13318
100|13319,13322
mg|13323,13325
PO|13326,13328
BID|13329,13332
<EOL>|13333,13334
7.|13334,13336
Dorzolamide|13337,13348
2|13349,13350
%|13350,13351
Ophth|13352,13357
.|13357,13358
Soln.|13359,13364
1|13365,13366
DROP|13367,13371
BOTH|13372,13376
EYES|13377,13381
BID|13382,13385
<EOL>|13386,13387
8.|13387,13389
Ferrous|13390,13397
Sulfate|13398,13405
325|13406,13409
mg|13410,13412
PO|13413,13415
DAILY|13416,13421
<EOL>|13422,13423
9.|13423,13425
Fluticasone|13426,13437
Propionate|13438,13448
NASAL|13449,13454
2|13455,13456
SPRY|13457,13461
NU|13462,13464
DAILY|13465,13470
:|13470,13471
PRN|13471,13474
allergies|13475,13484
<EOL>|13485,13486
10.|13486,13489
Hydrochlorothiazide|13490,13509
50|13510,13512
mg|13513,13515
PO|13516,13518
DAILY|13519,13524
<EOL>|13525,13526
11.|13526,13529
Isosorbide|13530,13540
Mononitrate|13541,13552
(|13553,13554
Extended|13554,13562
Release|13563,13570
)|13570,13571
240|13572,13575
mg|13576,13578
PO|13579,13581
DAILY|13582,13587
<EOL>|13588,13589
12.|13589,13592
Latanoprost|13593,13604
0.005|13605,13610
%|13610,13611
Ophth|13612,13617
.|13617,13618
Soln.|13619,13624
1|13625,13626
DROP|13627,13631
BOTH|13632,13636
EYES|13637,13641
QHS|13642,13645
<EOL>|13646,13647
13.|13647,13650
Multivitamins|13651,13664
1|13665,13666
TAB|13667,13670
PO|13671,13673
DAILY|13674,13679
<EOL>|13680,13681
14.|13681,13684
PredniSONE|13685,13695
30|13696,13698
mg|13699,13701
PO|13702,13704
DAILY|13705,13710
<EOL>|13711,13712
RX|13712,13714
*|13715,13716
prednisone|13716,13726
10|13727,13729
mg|13730,13732
3|13733,13734
tablet|13735,13741
(|13741,13742
s|13742,13743
)|13743,13744
by|13745,13747
mouth|13748,13753
Daily|13754,13759
Disp|13760,13764
#|13765,13766
*|13766,13767
30|13767,13769
Tablet|13770,13776
<EOL>|13777,13778
Refills|13778,13785
:|13785,13786
*|13786,13787
0|13787,13788
<EOL>|13788,13789
15.|13789,13792
Ranitidine|13793,13803
300|13804,13807
mg|13808,13810
PO|13811,13813
DAILY|13814,13819
<EOL>|13820,13821
16|13821,13823
.|13823,13824
Theophylline|13825,13837
SR|13838,13840
300|13841,13844
mg|13845,13847
PO|13848,13850
BID|13851,13854
<EOL>|13855,13856
17.|13856,13859
Tiotropium|13860,13870
Bromide|13871,13878
1|13879,13880
CAP|13881,13884
IH|13885,13887
DAILY|13888,13893
<EOL>|13894,13895
18.|13895,13898
Guaifenesin|13899,13910
1|13911,13912
teaspoon|13913,13921
PO|13922,13924
Q3H|13925,13928
:|13928,13929
PRN|13929,13932
cough|13933,13938
<EOL>|13939,13940
19|13940,13942
.|13942,13943
Ipratropium|13944,13955
Bromide|13956,13963
Neb|13964,13967
1|13968,13969
NEB|13970,13973
IH|13974,13976
Q6H|13977,13980
:|13980,13981
PRN|13981,13984
Wheezing|13985,13993
<EOL>|13994,13995
20.|13995,13998
cod|13999,14002
liver|14003,14008
oil|14009,14012
1|14013,14014
capsule|14015,14022
oral|14024,14028
BID|14029,14032
<EOL>|14033,14034
21|14034,14036
.|14036,14037
Calcitrate|14038,14048
-|14048,14049
Vitamin|14049,14056
D|14057,14058
(|14059,14060
calcium|14060,14067
citrate|14068,14075
-|14075,14076
vitamin|14076,14083
D3|14084,14086
)|14086,14087
315|14088,14091
mg|14092,14094
-|14095,14096
<EOL>|14097,14098
200|14098,14101
units|14102,14107
oral|14109,14113
DAILY|14114,14119
<EOL>|14120,14121
22.|14121,14124
albuterol|14125,14134
sulfate|14135,14142
90|14143,14145
mcg|14146,14149
/|14149,14150
actuation|14150,14159
inhalation|14160,14170
Q4H|14171,14174
<EOL>|14175,14176
23|14176,14178
.|14178,14179
Fluticasone|14180,14191
-|14191,14192
Salmeterol|14192,14202
Diskus|14203,14209
(|14210,14211
500|14211,14214
/|14214,14215
50|14215,14217
)|14217,14218
1|14220,14221
INH|14222,14225
IH|14226,14228
BID|14229,14232
<EOL>|14233,14234
RX|14234,14236
*|14237,14238
fluticasone|14238,14249
-|14249,14250
salmeterol|14250,14260
[|14261,14262
Advair|14262,14268
Diskus|14269,14275
]|14275,14276
500|14277,14280
mcg|14281,14284
-|14284,14285
50|14285,14287
mcg|14288,14291
/|14291,14292
dose|14292,14296
1|14297,14298
<EOL>|14299,14300
dose|14300,14304
Inhaled|14305,14312
Twice|14313,14318
a|14319,14320
day|14321,14324
Disp|14325,14329
#|14330,14331
*|14331,14332
1|14332,14333
Disk|14334,14338
Refills|14339,14346
:|14346,14347
*|14347,14348
1|14348,14349
<EOL>|14349,14350
24|14350,14352
.|14352,14353
Lorazepam|14354,14363
0.5|14364,14367
mg|14368,14370
PO|14371,14373
Q8H|14374,14377
:|14377,14378
PRN|14378,14381
Anxiety|14382,14389
<EOL>|14390,14391
RX|14391,14393
*|14394,14395
lorazepam|14395,14404
[|14405,14406
Ativan|14406,14412
]|14412,14413
0.5|14414,14417
mg|14418,14420
0.5|14421,14424
(|14425,14426
One|14426,14429
half|14430,14434
)|14434,14435
mg|14436,14438
by|14439,14441
mouth|14442,14447
Every|14448,14453
8|14454,14455
<EOL>|14456,14457
hours|14457,14462
Disp|14463,14467
#|14468,14469
*|14469,14470
30|14470,14472
Tablet|14473,14479
Refills|14480,14487
:|14487,14488
*|14488,14489
0|14489,14490
<EOL>|14490,14491
<EOL>|14491,14492
<EOL>|14493,14494
Discharge|14494,14503
Disposition|14504,14515
:|14515,14516
<EOL>|14516,14517
Home|14517,14521
With|14522,14526
Service|14527,14534
<EOL>|14534,14535
<EOL>|14536,14537
Facility|14537,14545
:|14545,14546
<EOL>|14546,14547
_|14547,14548
_|14548,14549
_|14549,14550
<EOL>|14550,14551
<EOL>|14552,14553
Discharge|14553,14562
Diagnosis|14563,14572
:|14572,14573
<EOL>|14573,14574
Primary|14574,14581
Diagnosis|14582,14591
:|14591,14592
<EOL>|14592,14593
Chronic|14593,14600
obstruction|14601,14612
pulmonary|14613,14622
disease|14623,14630
exacerbation|14631,14643
<EOL>|14643,14644
<EOL>|14644,14645
Secondary|14645,14654
Diagnoses|14655,14664
:|14664,14665
<EOL>|14665,14666
Tobacco|14666,14673
use|14674,14677
disorder|14678,14686
<EOL>|14686,14687
Atrial|14687,14693
fibrillation|14694,14706
<EOL>|14706,14707
Hypertension|14707,14719
<EOL>|14719,14720
Anxiety|14720,14727
<EOL>|14727,14728
Coronary|14728,14736
Artery|14737,14743
Disease|14744,14751
<EOL>|14751,14752
<EOL>|14752,14753
<EOL>|14754,14755
Discharge|14755,14764
Condition|14765,14774
:|14774,14775
<EOL>|14775,14776
Mental|14776,14782
Status|14783,14789
:|14789,14790
Clear|14791,14796
and|14797,14800
coherent|14801,14809
.|14809,14810
<EOL>|14810,14811
Level|14811,14816
of|14817,14819
Consciousness|14820,14833
:|14833,14834
Alert|14835,14840
and|14841,14844
interactive|14845,14856
.|14856,14857
<EOL>|14857,14858
Activity|14858,14866
Status|14867,14873
:|14873,14874
Ambulatory|14875,14885
-|14886,14887
Independent|14888,14899
.|14899,14900
<EOL>|14900,14901
<EOL>|14901,14902
<EOL>|14903,14904
Discharge|14904,14913
Instructions|14914,14926
:|14926,14927
<EOL>|14927,14928
Dear|14928,14932
Ms.|14933,14936
_|14937,14938
_|14938,14939
_|14939,14940
,|14940,14941
<EOL>|14941,14942
<EOL>|14942,14943
It|14943,14945
was|14946,14949
a|14950,14951
privilege|14952,14961
taking|14962,14968
care|14969,14973
of|14974,14976
you|14977,14980
during|14981,14987
your|14988,14992
admission|14993,15002
to|15003,15005
<EOL>|15006,15007
_|15007,15008
_|15008,15009
_|15009,15010
.|15010,15011
You|15012,15015
were|15016,15020
admitted|15021,15029
to|15030,15032
the|15033,15036
hospital|15037,15045
for|15046,15049
<EOL>|15050,15051
shortness|15051,15060
of|15061,15063
breath|15064,15070
and|15071,15074
concern|15075,15082
that|15083,15087
you|15088,15091
were|15092,15096
having|15097,15103
a|15104,15105
flare|15106,15111
of|15112,15114
<EOL>|15115,15116
your|15116,15120
COPD|15121,15125
.|15125,15126
<EOL>|15126,15127
<EOL>|15127,15128
While|15128,15133
in|15134,15136
the|15137,15140
hospital|15141,15149
we|15150,15152
increased|15153,15162
your|15163,15167
dose|15168,15172
of|15173,15175
steroids|15176,15184
to|15185,15187
help|15188,15192
<EOL>|15193,15194
your|15194,15198
breathing|15199,15208
.|15208,15209
You|15210,15213
also|15214,15218
received|15219,15227
several|15228,15235
nebulizer|15236,15245
treatments|15246,15256
<EOL>|15257,15258
that|15258,15262
helped|15263,15269
your|15270,15274
breathing|15275,15284
.|15284,15285
You|15286,15289
were|15290,15294
also|15295,15299
expressing|15300,15310
some|15311,15315
<EOL>|15316,15317
anxiety|15317,15324
that|15325,15329
may|15330,15333
have|15334,15338
been|15339,15343
contributing|15344,15356
to|15357,15359
your|15360,15364
shortness|15365,15374
of|15375,15377
<EOL>|15378,15379
breath|15379,15385
.|15385,15386
You|15387,15390
were|15391,15395
given|15396,15401
a|15402,15403
medication|15404,15414
called|15415,15421
Ativan|15422,15428
for|15429,15432
your|15433,15437
<EOL>|15438,15439
anxiety|15439,15446
that|15447,15451
also|15452,15456
seemed|15457,15463
to|15464,15466
help|15467,15471
your|15472,15476
breathing|15477,15486
.|15486,15487
<EOL>|15487,15488
<EOL>|15488,15489
During|15489,15495
your|15496,15500
admission|15501,15510
you|15511,15514
were|15515,15519
seen|15520,15524
by|15525,15527
the|15528,15531
pulmonary|15532,15541
<EOL>|15542,15543
specialists|15543,15554
.|15554,15555
They|15556,15560
recommended|15561,15572
a|15573,15574
CT|15575,15577
scan|15578,15582
that|15583,15587
showed|15588,15594
that|15595,15599
you|15600,15603
<EOL>|15604,15605
have|15605,15609
extensive|15610,15619
COPD|15620,15624
but|15625,15628
did|15629,15632
not|15633,15636
show|15637,15641
any|15642,15645
infection|15646,15655
.|15655,15656
They|15657,15661
also|15662,15666
<EOL>|15667,15668
suggested|15668,15677
increasing|15678,15688
the|15689,15692
dose|15693,15697
of|15698,15700
your|15701,15705
Advair|15706,15712
inhaler|15713,15720
,|15720,15721
which|15722,15727
we|15728,15730
<EOL>|15731,15732
did|15732,15735
.|15735,15736
<EOL>|15736,15737
<EOL>|15737,15738
If|15738,15740
you|15741,15744
feel|15745,15749
short|15750,15755
of|15756,15758
breath|15759,15765
,|15765,15766
first|15767,15772
please|15773,15779
check|15780,15785
your|15786,15790
oxygen|15791,15797
<EOL>|15798,15799
level|15799,15804
.|15804,15805
If|15806,15808
it|15809,15811
is|15812,15814
less|15815,15819
than|15820,15824
90|15825,15827
,|15827,15828
you|15829,15832
can|15833,15836
use|15837,15840
oxygen|15841,15847
and|15848,15851
your|15852,15856
<EOL>|15857,15858
inhaler|15858,15865
.|15865,15866
If|15867,15869
not|15870,15873
,|15873,15874
try|15875,15878
to|15879,15881
wait|15882,15886
a|15887,15888
few|15889,15892
minutes|15893,15900
,|15900,15901
take|15902,15906
a|15907,15908
few|15909,15912
deep|15913,15917
<EOL>|15918,15919
breaths|15919,15926
and|15927,15930
see|15931,15934
if|15935,15937
your|15938,15942
shortness|15943,15952
of|15953,15955
breath|15956,15962
improves|15963,15971
.|15971,15972
You|15973,15976
can|15977,15980
<EOL>|15981,15982
use|15982,15985
the|15986,15989
medication|15990,16000
called|16001,16007
Ativan|16008,16014
(|16014,16015
lorazepam|16015,16024
)|16024,16025
to|16026,16028
help|16029,16033
with|16034,16038
the|16039,16042
<EOL>|16043,16044
shortness|16044,16053
of|16054,16056
breath|16057,16063
(|16063,16064
no|16064,16066
more|16067,16071
than|16072,16076
three|16077,16082
times|16083,16088
a|16089,16090
day|16091,16094
)|16094,16095
.|16095,16096
If|16097,16099
still|16100,16105
<EOL>|16106,16107
not|16107,16110
improved|16111,16119
,|16119,16120
you|16121,16124
can|16125,16128
use|16129,16132
one|16133,16136
of|16137,16139
the|16140,16143
inhalers|16144,16152
/|16152,16153
oxygen|16153,16159
.|16159,16160
<EOL>|16161,16162
<EOL>|16162,16163
Please|16163,16169
follow|16170,16176
-|16176,16177
up|16177,16179
with|16180,16184
all|16185,16188
your|16189,16193
appointments|16194,16206
as|16207,16209
listed|16210,16216
below|16217,16222
and|16223,16226
<EOL>|16227,16228
continue|16228,16236
to|16237,16239
take|16240,16244
all|16245,16248
of|16249,16251
your|16252,16256
medications|16257,16268
as|16269,16271
prescribed|16272,16282
.|16282,16283
If|16284,16286
you|16287,16290
<EOL>|16291,16292
experience|16292,16302
any|16303,16306
of|16307,16309
the|16310,16313
danger|16314,16320
signs|16321,16326
listed|16327,16333
you|16334,16337
should|16338,16344
call|16345,16349
your|16350,16354
<EOL>|16355,16356
doctor|16356,16362
immediately|16363,16374
or|16375,16377
go|16378,16380
to|16381,16383
the|16384,16387
Emergency|16388,16397
Room|16398,16402
.|16402,16403
<EOL>|16403,16404
<EOL>|16404,16405
We|16405,16407
wish|16408,16412
you|16413,16416
the|16417,16420
best|16421,16425
!|16425,16426
<EOL>|16426,16427
<EOL>|16427,16428
Sincerely|16428,16437
,|16437,16438
<EOL>|16438,16439
Your|16439,16443
_|16444,16445
_|16445,16446
_|16446,16447
Care|16448,16452
Team|16453,16457
<EOL>|16457,16458
<EOL>|16459,16460
Followup|16460,16468
Instructions|16469,16481
:|16481,16482
<EOL>|16482,16483
_|16483,16484
_|16484,16485
_|16485,16486
<EOL>|16486,16487

