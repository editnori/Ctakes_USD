CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|true|false||Unit
null|Unit device|Device|true|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|true|false||Unit
null|Unit of Measure|LabModifier|true|false||Unit
null|Unit|LabModifier|true|false||Unit
null|Enzyme Unit|LabModifier|true|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Psychiatry Specialty|Title|false|false||PSYCHIATRYnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|Relationship modifier - Patient|Finding|true|false||Patient
null|Specimen Type - Patient|Finding|true|false||Patient
null|Mail Claim Party - Patient|Finding|true|false||Patient
null|Report source - Patient|Finding|true|false||Patient
null|null|Finding|true|false||Patient
null|Disabled Person Code - Patient|Finding|true|false||Patientnull|Patients|Subject|true|false||Patientnull|Veterinary Patient|Entity|true|false||Patientnull|Known|Modifier|true|false||Knownnull|Hypersensitivity|Finding|true|false||Allergiesnull|null|Attribute|true|false||Allergiesnull|Pharmaceutical Preparations|Drug|true|false||Drugsnull|Drugs - dental services|Procedure|true|false||Drugsnull|Attending (action)|Finding|true|false||Attendingnull|Attending (provider role)|Subject|true|false||Attendingnull|Chief complaint (finding)|Finding|false|false||Chief Complaintnull|Complaint (finding)|Finding|false|false||Complaintnull|null|Attribute|false|false||Complaintnull|Suicidal|Disorder|false|false||suicidalnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|History of present illness (finding)|Finding|true|false||History of Present Illnessnull|null|Attribute|true|false||History of Present Illnessnull|Medical History|Finding|true|false||History ofnull|History of present illness (finding)|Finding|true|false||History
null|History of previous events|Finding|true|false||History
null|Historical aspects qualifier|Finding|true|false||History
null|Medical History|Finding|true|false||History
null|Concept History|Finding|true|false||Historynull|History|Subject|true|false||Historynull|Present illness|Finding|true|false||Present Illnessnull|Present|Finding|true|false||Present
null|Presentation|Finding|true|false||Presentnull|Illness (finding)|Finding|true|false||Illnessnull|Proline dehydrogenase deficiency|Disorder|false|false||HPInull|History of present illness (finding)|Finding|false|false||HPI
null|allene oxide synthase activity|Finding|false|false||HPInull|Depressed mood|Disorder|false|false||depressed moodnull|Depressed mood|Disorder|false|false||depressednull|Mood (psychological function)|Finding|false|false||mood
null|mood (physical finding)|Finding|false|false||mood
null|Mood (attribute)|Finding|false|false||moodnull|null|Attribute|false|false||moodnull|Anxiety symptoms|Finding|false|false||anxiety symptomsnull|Anxiety Disorders|Disorder|false|false||anxiety
null|Anxiety|Disorder|false|false||anxietynull|Anxiety symptoms|Finding|false|false||anxietynull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Panic|Finding|false|false||panicnull|Recommendation|Finding|false|false||recommendationnull|therapist|Subject|false|false||therapistnull|month|Time|false|false||monthsnull|Processing type - Evaluation|Finding|false|false||evaluationnull|Evaluation procedure|Procedure|false|false||evaluation
null|Evaluation|Procedure|false|false||evaluationnull|3 Weeks|Time|false|false||3 weeksnull|week|Time|false|false||weeksnull|Cancer patients and suicide and depression|Disorder|false|false||depression
null|Mental Depression|Disorder|false|false||depression
null|Depressive disorder|Disorder|false|false||depression
null|Depressed mood|Disorder|false|false||depressionnull|Depression - motion|Finding|false|false||depression
null|null|Finding|false|false||depressionnull|Depression - recess|Modifier|false|false||depressionnull|Social Anhedonia|Disorder|false|false||anhedonia, socialnull|Anhedonia|Disorder|false|false||anhedonianull|Social isolation|Finding|false|false||social isolationnull|Social|Finding|false|false||socialnull|Social isolation|Finding|false|false||isolation
null|Isolated|Finding|false|false||isolation
null|Privacy Level - Isolation|Finding|false|false||isolation
null|Level of Care - Isolation|Finding|false|false||isolation
null|Need for isolation|Finding|false|false||isolationnull|Isolation procedure|Procedure|false|false||isolation
null|isolation aspects|Procedure|false|false||isolationnull|Accommodation - Isolation|Device|false|false||isolationnull|Specialty Type - Isolation|Title|false|false||isolationnull|Withdrawal (dysfunction)|Disorder|false|false||withdrawalnull|Withdrawal - birth control|Procedure|false|false||withdrawalnull|Withdraw (activity)|Event|false|false||withdrawalnull|Guilt|Finding|false|false||feelings of guiltnull|Subject's Feelings|Finding|false|false||feelings
null|Feelings|Finding|false|false||feelingsnull|Guilt|Finding|false|false||guiltnull|Difficulty sleeping|Finding|false|false||poor sleepnull|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group|Finding|false|false||poor
null|Patient Condition Code - Poor|Finding|false|false||poornull|Poverty|Subject|false|false||poornull|Language Proficiency - Poor|Modifier|false|false||poor
null|Specimen Quality - Poor|Modifier|false|false||poor
null|Poor - grade|Modifier|false|false||poor
null|Poor - qualifier|Modifier|false|false||poornull|Sleep brand of diphenhydramine hydrochloride|Drug|false|false||sleep
null|Sleep brand of diphenhydramine hydrochloride|Drug|false|false||sleepnull|Sleep|Finding|false|false||sleepnull|Neoplasm Metastasis|Disorder|false|false||secondarynull|metastatic qualifier|Finding|false|false||secondarynull|Secondary to|Modifier|false|false||secondarynull|second (number)|LabModifier|false|false||secondarynull|Rumination Disorders|Disorder|false|false||ruminationsnull|Rumination|Phenomenon|false|false||ruminationsnull|Guilt|Finding|false|false||guiltnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Class|Finding|false|false||classesnull|Classes - encounter|Procedure|false|false||classesnull|Cancer patients and suicide and depression|Disorder|false|false||depression
null|Mental Depression|Disorder|false|false||depression
null|Depressive disorder|Disorder|false|false||depression
null|Depressed mood|Disorder|false|false||depressionnull|Depression - motion|Finding|false|false||depression
null|null|Finding|false|false||depressionnull|Depression - recess|Modifier|false|false||depressionnull|Anxiety Disorders|Disorder|false|false||anxiety
null|Anxiety|Disorder|false|false||anxietynull|Anxiety symptoms|Finding|false|false||anxietynull|Legal fine|Entity|false|false||finenull|Fine (qualifier value)|Modifier|false|false||finenull|Continuity Assessment Record and Evaluation|Finding|false|false||care
null|In care (finding)|Finding|false|false||carenull|care activity|Event|false|false||carenull|Hygiene|Title|false|false||hygienenull|Recent|Time|false|false||recentnull|bout|Time|false|false||boutnull|Anxiety Disorders|Disorder|false|false||anxiety
null|Anxiety|Disorder|false|false||anxietynull|Anxiety symptoms|Finding|false|false||anxietynull|Stress bismuth subsalicylate|Drug|false|false||stress
null|Stress bismuth subsalicylate|Drug|false|false||stressnull|Stress|Finding|false|false||stressnull|W stress|Attribute|false|false||stressnull|Entity Name Part Qualifier - professional|Finding|false|false||professional
null|Charge type - professional|Finding|false|false||professionalnull|professional occupation status|Subject|false|false||professional
null|Professional Occupation|Subject|false|false||professionalnull|Concept Relationship|Finding|false|false||relationship
null|Object Relationship|Finding|false|false||relationshipnull|Relationships|Modifier|false|false||relationshipnull|Teacher|Subject|false|false||teachersnull|Program|Drug|false|false||program
null|Program|Drug|false|false||programnull|Program - framework of goals|Finding|false|false||program
null|Programs - Publication Format|Finding|false|false||program
null|Programs|Finding|false|false||programnull|Indication of (contextual qualifier)|Finding|true|false||reasonsnull|Completely - dosing instruction fragment|Finding|true|false||completelynull|Complete|Modifier|true|false||completelynull|Remote control command - Clear|Finding|true|false||clearnull|Clear|Modifier|true|false||clear
null|Transparent (qualitative concept)|Modifier|true|false||clearnull|Relationship modifier - Patient|Finding|true|false||patient
null|Specimen Type - Patient|Finding|true|false||patient
null|Mail Claim Party - Patient|Finding|true|false||patient
null|Report source - Patient|Finding|true|false||patient
null|null|Finding|true|false||patient
null|Disabled Person Code - Patient|Finding|true|false||patientnull|Patients|Subject|true|false||patientnull|Veterinary Patient|Entity|true|false||patientnull|LOINC class types|Finding|false|false||class
null|Class|Finding|false|false||class
null|Classification|Finding|false|false||class
null|Taxonomic|Finding|false|false||class
null|Taxonomic Class|Finding|false|false||classnull|Kind of quantity - Class|LabModifier|false|false||classnull|Instructor|Subject|false|false||instructor
null|Teacher|Subject|false|false||instructornull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Speak - language ability|Finding|false|false||speak
null|Speaking (function)|Finding|false|false||speak
null|Does speak|Finding|false|false||speaknull|Availability of|Finding|true|false||availablenull|Relationship modifier - Patient|Finding|true|false||patient
null|Specimen Type - Patient|Finding|true|false||patient
null|Mail Claim Party - Patient|Finding|true|false||patient
null|Report source - Patient|Finding|true|false||patient
null|null|Finding|true|false||patient
null|Disabled Person Code - Patient|Finding|true|false||patientnull|Patients|Subject|true|false||patientnull|Veterinary Patient|Entity|true|false||patientnull|Floor - story of building|Entity|false|false||storynull|detail - Response Level|Finding|false|false||detailnull|Details|Modifier|false|false||detailnull|FACT Complex|Drug|false|false||fact
null|FACT Complex|Drug|false|false||factnull|SSRP1 wt Allele|Finding|false|false||fact
null|SUPT16H gene|Finding|false|false||factnull|Foundation for the Accreditation of Cellular Therapy|Subject|false|false||factnull|Panic|Finding|false|false||panicnull|Attack (finding)|Finding|false|false||attack
null|Attack behavior|Finding|false|false||attacknull|Attack device|Device|false|false||attacknull|Does talk|Finding|false|false||talk
null|Speech|Finding|false|false||talk
null|Speaking (function)|Finding|false|false||talknull|week|Time|false|false||weeksnull|LOINC class types|Finding|false|false||class
null|Class|Finding|false|false||class
null|Classification|Finding|false|false||class
null|Taxonomic|Finding|false|false||class
null|Taxonomic Class|Finding|false|false||classnull|Kind of quantity - Class|LabModifier|false|false||classnull|null|Finding|true|false||lettersnull|Message|Finding|true|false||messagesnull|Instructor|Subject|true|false||instructor
null|Teacher|Subject|true|false||instructornull|Communication Response|Finding|true|false||response
null|Disease Response|Finding|true|false||response
null|Answer (statement)|Finding|true|false||responsenull|Response process|Subject|true|false||responsenull|Lacking|Modifier|false|false||lacknull|Communication Response|Finding|false|false||response
null|Disease Response|Finding|false|false||response
null|Answer (statement)|Finding|false|false||responsenull|Response process|Subject|false|false||responsenull|Patterns|Modifier|false|false||patternnull|Guilt|Finding|false|false||guiltnull|Cutting self|Disorder|false|false||cuttingnull|self-mutilation by cutting (history)|Finding|false|false||cuttingnull|Transection (procedure)|Procedure|false|false||cuttingnull|Cutting sensation quality|Modifier|false|false||cuttingnull|knife|Device|true|false||knifenull|Incised wound|Disorder|true|false||cutnull|reported cut of tissue (history)|Finding|true|false||cut
null|CUX1 gene|Finding|true|false||cutnull|Cuneate tubercle structure|Anatomy|true|false||cutnull|Structure of left wrist|Anatomy|true|false||left wristnull|Table Cell Horizontal Align - left|Finding|true|false||leftnull|Left sided|Modifier|true|false||left
null|Left|Modifier|true|false||leftnull|Upper extremity>Wrist|Anatomy|true|false||wrist
null|Wrist joint|Anatomy|true|false||wrist
null|Wrist|Anatomy|true|false||wristnull|Last|Modifier|false|false||Lastnull|Night time|Time|false|false||nightnull|Application Context|Finding|true|false||context
null|Context|Finding|true|false||context
null|contextual factors|Finding|true|false||contextnull|Guilt|Finding|true|false||guiltnull|More|LabModifier|true|false||morenull|Anxiety Disorders|Disorder|true|false||anxiety
null|Anxiety|Disorder|true|false||anxietynull|Anxiety symptoms|Finding|true|false||anxietynull|Feeling suicidal (finding)|Finding|false|false||feeling suicidalnull|Suicidal|Disorder|false|false||suicidalnull|Infantile Neuroaxonal Dystrophy|Disorder|false|false||plannull|Treatment Plan|Finding|false|false||plan
null|Planned|Finding|false|false||plan
null|null|Finding|false|false||plannull|knife|Device|false|false||knifenull|Subject's Feelings|Finding|false|false||feelings
null|Feelings|Finding|false|false||feelingsnull|Cancer patients and suicide and depression|Disorder|false|false||suicidenull|Suicide|Finding|false|false||suicidenull|counselor|Finding|false|false||counselornull|Counselors|Subject|false|false||counselornull|null|Finding|false|false||thoughts
null|Thought|Finding|false|false||thoughtsnull|counselor|Finding|false|false||counselornull|Counselors|Subject|false|false||counselornull|Never - AcknowledgementCondition|Time|false|false||never
null|Never (frequency)|Time|false|false||nevernull|Greater Than|LabModifier|true|false||more thannull|More|LabModifier|true|false||morenull|Transaction counts and value totals - day|Finding|true|false||day
null|Precision - day|Finding|true|false||daynull|Land Dayak Languages|Entity|true|false||daynull|day|Time|true|false||day
null|Daily|Time|true|false||daynull|Never - AcknowledgementCondition|Time|false|false||never
null|Never (frequency)|Time|false|false||nevernull|Sleep brand of diphenhydramine hydrochloride|Drug|true|false||sleep
null|Sleep brand of diphenhydramine hydrochloride|Drug|true|false||sleepnull|Sleep|Finding|true|false||sleepnull|Impaired decision-making|Finding|false|false||impaired decision-makingnull|Impaired|Finding|false|false||impairednull|Decision Making|Finding|false|false||decision-makingnull|Decision|Finding|false|false||decisionnull|spending|LabModifier|false|false||spendingnull|Too much|Finding|false|false||too muchnull|Much|Finding|false|false||muchnull|Indiscriminate|Modifier|false|false||indiscriminatenull|Sexual relationships|Finding|false|false||sexual relationshipsnull|Sex Behavior|Finding|false|false||sexualnull|Relationships|Modifier|false|false||relationshipsnull|Etc.|Finding|false|false||etcnull|Psychotic symptom|Finding|false|false||psychotic symptomsnull|Psychotic Disorders|Disorder|false|false||psychoticnull|Psychotic symptom present|Finding|false|false||psychoticnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Guilt|Finding|false|false||guiltnull|Psychotic Disorders|Disorder|false|false||psychoticnull|Psychotic symptom present|Finding|false|false||psychoticnull|Proportion|LabModifier|false|false||proportionnull|Instructor|Subject|true|false||instructor
null|Teacher|Subject|true|false||instructornull|Never - AcknowledgementCondition|Time|false|false||never
null|Never (frequency)|Time|false|false||nevernull|Instructor|Subject|true|false||instructor
null|Teacher|Subject|true|false||instructornull|Email|Finding|true|false||emailsnull|Instructor|Subject|true|false||instructor
null|Teacher|Subject|true|false||instructornull|null|Finding|true|false||thoughts
null|Thought|Finding|true|false||thoughtsnull|Instructor|Subject|false|false||instructor
null|Teacher|Subject|false|false||instructornull|Anxiety|Disorder|false|false||feeling anxiousnull|Anxious mood|Finding|false|false||feeling anxiousnull|Anxiety|Disorder|false|false||anxiousnull|RXFP2 gene|Finding|false|false||greatnull|Greater|LabModifier|false|false||great
null|Large|LabModifier|false|false||greatnull|Retinoic Acid Response Element|Finding|false|false||rarenull|Infrequent|Time|false|false||rarenull|Rare|Modifier|false|false||rarenull|Panic Attacks|Disorder|false|false||panic attacknull|Panic|Finding|false|false||panicnull|Attack (finding)|Finding|false|false||attack
null|Attack behavior|Finding|false|false||attacknull|Attack device|Device|false|false||attacknull|PMH - past medical history|Finding|false|false||Past Medical History
null|Medical History|Finding|false|false||Past Medical Historynull|Medical History|Finding|false|false||Medical Historynull|Medical referral type|Finding|false|false||Medical
null|Medical|Finding|false|false||Medical
null|Medical school type|Finding|false|false||Medicalnull|Medical service|Procedure|false|false||Medicalnull|Medical History|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|History of present illness (finding)|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Psychiatric problem|Disorder|false|false||PSYCH
null|Mental disorders|Disorder|false|false||PSYCHnull|Act Relationship Subset - previous|Time|true|false||previous
null|Previous|Time|true|false||previousnull|Pharmaceutical Preparations|Drug|true|false||medicationnull|medication - HL7 publishing domain|Finding|true|false||medication
null|Medications|Finding|true|false||medicationnull|Referral type - Psychiatric|Finding|true|false||psychiatric
null|Psychiatric|Finding|true|false||psychiatricnull|Psychiatric service|Procedure|true|false||psychiatricnull|Psychiatry Specialty|Title|true|false||psychiatricnull|Hospitalization|Procedure|true|false||hospitalizationsnull|Act Relationship Subset - previous|Time|false|false||previous
null|Previous|Time|false|false||previousnull|Episode of|Time|false|false||episode ofnull|Episode of|Time|false|false||episodenull|Referral type - Psychiatric|Finding|false|false||psychiatric
null|Psychiatric|Finding|false|false||psychiatricnull|Psychiatric service|Procedure|false|false||psychiatricnull|Psychiatry Specialty|Title|false|false||psychiatricnull|Application Context|Finding|false|false||context
null|Context|Finding|false|false||context
null|contextual factors|Finding|false|false||contextnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Panic Attacks|Disorder|false|false||panic attacknull|Panic|Finding|false|false||panicnull|Attack (finding)|Finding|false|false||attack
null|Attack behavior|Finding|false|false||attacknull|Attack device|Device|false|false||attacknull|Infrequent|Time|false|false||occasionalnull|Panic Attacks|Disorder|false|false||panic attacksnull|Panic|Finding|false|false||panicnull|Attack (finding)|Finding|false|false||attacks
null|Attack behavior|Finding|false|false||attacksnull|Frequently|Time|true|false||frequentlynull|Diagnosis Classification - Diagnosis|Finding|true|false||diagnosis
null|diagnosis aspects|Finding|true|false||diagnosisnull|Diagnosis|Procedure|true|false||diagnosisnull|null|Attribute|true|false||diagnosisnull|Panic|Finding|false|false||panicnull|counselor|Finding|false|false||counselornull|Counselors|Subject|false|false||counselornull|month|Time|false|false||monthsnull|null|Time|true|false||Prior tonull|null|Time|true|false||Priornull|3 Weeks|Time|true|false||3 weeksnull|week|Time|true|false||weeksnull|FBXW7 wt Allele|Finding|true|false||ago
null|FBXW7 gene|Finding|true|false||agonull|Self-Injurious Behavior|Finding|true|false||self-injurious behaviorsnull|subscriber - self|Finding|true|false||self
null|Self|Finding|true|false||selfnull|Behaviors and observations relating to behavior|Finding|true|false||behaviors
null|Behavior|Finding|true|false||behaviorsnull|Suicidal thoughts|Finding|false|false||suicidal ideationnull|null|Attribute|false|false||suicidal ideationnull|Suicidal|Disorder|false|false||suicidalnull|ideation|Finding|false|false||ideationnull|One to two times|Time|false|false||once or twicenull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|null|Time|false|false||prior tonull|null|Time|false|false||priornull|Last|Modifier|false|false||lastnull|Night time|Time|false|false||nightnull|Never - AcknowledgementCondition|Time|false|false||never
null|Never (frequency)|Time|false|false||nevernull|Act Mood - intent|Finding|true|false||intent
null|null|Finding|true|false||intentnull|intent|Modifier|true|false||intentnull|counselor|Finding|false|false||counselornull|Counselors|Subject|false|false||counselornull|high school level|Finding|false|false||high schoolnull|High Schools|Device|false|false||high schoolnull|High School Graduate|Subject|false|false||high schoolnull|High Schools|Entity|false|false||high schoolnull|Message Waiting Priority - High|Finding|false|false||high
null|high - ActExposureLevelCode|Finding|false|false||high
null|IPSS Risk Category High|Finding|false|false||high
null|IPSS-R Risk Category High|Finding|false|false||high
null|High (finding)|Finding|false|false||highnull|Observation Value - High|Modifier|false|false||high
null|High|Modifier|false|false||high
null|Abnormally high|Modifier|false|false||highnull|School|Device|false|false||schoolnull|School|Entity|false|false||schoolnull|Child coping with hospitalization|Finding|false|false||coping
null|Coping Behavior|Finding|false|false||copingnull|COPING - Dental Restorative Procedure|Procedure|false|false||coping
null|COPING - Fixed Prosthodontics|Procedure|false|false||copingnull|Feelings|Finding|false|false||feelingnull|Different|Modifier|false|false||differentnull|School|Device|false|false||schoolnull|School|Entity|false|false||schoolnull|null|Finding|false|false||thoughts
null|Thought|Finding|false|false||thoughtsnull|student|Subject|false|false||studentnull|month|Time|false|false||monthsnull|FBXW7 wt Allele|Finding|false|false||ago
null|FBXW7 gene|Finding|false|false||agonull|Encounter due to counseling|Finding|false|false||counseling
null|duration of counseling|Finding|false|false||counselingnull|Counseling|Procedure|false|false||counseling
null|Counselling service|Procedure|false|false||counselingnull|Details|Modifier|true|false||detailsnull|Able (qualifier value)|Finding|false|false||ablenull|Ability|Subject|false|false||ablenull|Person Info|Finding|false|false||personnull|null|Attribute|false|false||personnull|Persons|Subject|false|false||personnull|Violent|Disorder|true|false||violentnull|Behavior|Finding|true|false||behaviornull|null|Attribute|true|false||behaviornull|PMH - past medical history|Finding|false|false||PMH
null|Medical History|Finding|false|false||PMHnull|Healthy|Modifier|false|false||healthynull|Young|Time|false|false||youngnull|Male population group|Subject|false|false||man
null|Homo sapiens|Subject|false|false||man
null|Males|Subject|false|false||mannull|Mandinka Language|Entity|false|false||mannull|Repair of meniscus|Procedure|false|false||repair of meniscusnull|Repair|Finding|false|false||repair
null|Wound Healing|Finding|false|false||repairnull|Repair - Remedial Action|Procedure|false|false||repair
null|Surgical repair|Procedure|false|false||repairnull|Meniscus structure of joint|Anatomy|false|false||meniscusnull|Genus Meniscus|Entity|false|false||meniscusnull|Structure of left knee region|Anatomy|false|false||left knee
null|Structure of left knee|Anatomy|false|false||left kneenull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Examination of knee joint|Procedure|false|false||kneenull|Knee region structure|Anatomy|false|false||knee
null|Knee|Anatomy|false|false||knee
null|Lower extremity>Knee|Anatomy|false|false||knee
null|Knee joint|Anatomy|false|false||kneenull|Several|LabModifier|false|false||severalnull|month|Time|false|false||monthsnull|FBXW7 wt Allele|Finding|false|false||ago
null|FBXW7 gene|Finding|false|false||agonull|Secondary to|Modifier|false|false||secondary tonull|Neoplasm Metastasis|Disorder|false|false||secondarynull|metastatic qualifier|Finding|false|false||secondarynull|Secondary to|Modifier|false|false||secondarynull|second (number)|LabModifier|false|false||secondarynull|Traumatic AND/OR non-traumatic injury|Disorder|false|false||injury
null|Traumatic injury|Disorder|false|false||injurynull|Operative Surgical Procedures|Procedure|true|false||surgeriesnull|Social and personal history|Finding|false|false||Social History
null|Social History|Finding|false|false||Social Historynull|Social|Finding|false|false||Socialnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Social/family|Finding|false|false||SOCIAL/FAMILYnull|Social|Finding|false|false||SOCIALnull|Entity Name Part Type - family|Finding|false|false||FAMILY
null|Last Name|Finding|false|false||FAMILY
null|Living Arrangement - Family|Finding|false|false||FAMILY
null|Family (taxonomic)|Finding|false|false||FAMILY
null|Family Collection|Finding|false|false||FAMILYnull|Family|Subject|false|false||FAMILYnull|Is an only child|Subject|false|false||Only childnull|Relationship - Child|Finding|false|false||childnull|Child Individual|Subject|false|false||child
null|Offspring|Subject|false|false||child
null|Child|Subject|false|false||childnull|Divorced parents (family) (social concept)|Subject|false|false||divorced parentsnull|Divorced state|Finding|false|false||divorcednull|parent|Subject|false|false||parentsnull|parent|Subject|false|false||Parentsnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Relationship - Mother|Finding|false|false||mothernull|Mother (person)|Subject|false|false||mothernull|Concept Relationship|Finding|false|false||relationship
null|Object Relationship|Finding|false|false||relationshipnull|Relationships|Modifier|false|false||relationshipnull|Relationship - Father|Finding|false|false||father
null|Father - courtesy title|Finding|false|false||father
null|Indirect exposure mechanism - Father|Finding|false|false||fathernull|Father (person)|Subject|false|false||fathernull|Indirect exposure mechanism - Father|Finding|false|false||Father
null|Relationship - Father|Finding|false|false||Father
null|Father - courtesy title|Finding|false|false||Fathernull|Father (person)|Subject|false|false||Fathernull|Alcoholic Intoxication, Chronic|Disorder|false|false||alcohol dependencenull|Alcohols|Drug|false|false||alcohol
null|Alcohols|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcoholnull|Alcohol - Recreational Drug Use Code|Finding|false|false||alcoholnull|Dependence|Disorder|false|false||dependencenull|emotional dependency|Finding|false|false||dependencenull|year|Time|false|false||yearsnull|Relationship modifier - Patient|Finding|true|false||Patient
null|Specimen Type - Patient|Finding|true|false||Patient
null|Mail Claim Party - Patient|Finding|true|false||Patient
null|Report source - Patient|Finding|true|false||Patient
null|null|Finding|true|false||Patient
null|Disabled Person Code - Patient|Finding|true|false||Patientnull|Patients|Subject|true|false||Patientnull|Veterinary Patient|Entity|true|false||Patientnull|physical examination (physical finding)|Finding|true|false||physical
null|Physical|Finding|true|false||physicalnull|Physical Examination|Procedure|true|false||physicalnull|Sexual abuse|Disorder|true|false||sexual abusenull|Sex Behavior|Finding|true|false||sexualnull|Drug abuse|Disorder|true|false||abusenull|Victim of abuse (finding)|Finding|true|false||abusenull|Abuse|Event|true|false||abusenull|Different|Modifier|false|false||differentnull|Seizures|Finding|false|false||fittingnull|null|Procedure|false|false||fittingnull|More|LabModifier|true|false||morenull|Details|Modifier|true|false||detailsnull|Behavior|Finding|false|false||behavioralnull|School|Device|false|false||schoolnull|School|Entity|false|false||schoolnull|Relationship - Child|Finding|false|false||childnull|Child Individual|Subject|false|false||child
null|Offspring|Subject|false|false||child
null|Child|Subject|false|false||childnull|3 times|Finding|false|false||3 timesnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|high school level|Finding|false|false||high schoolnull|High Schools|Device|false|false||high schoolnull|High School Graduate|Subject|false|false||high schoolnull|High Schools|Entity|false|false||high schoolnull|Message Waiting Priority - High|Finding|false|false||high
null|high - ActExposureLevelCode|Finding|false|false||high
null|IPSS Risk Category High|Finding|false|false||high
null|IPSS-R Risk Category High|Finding|false|false||high
null|High (finding)|Finding|false|false||highnull|Observation Value - High|Modifier|false|false||high
null|High|Modifier|false|false||high
null|Abnormally high|Modifier|false|false||highnull|School|Device|false|false||schoolnull|School|Entity|false|false||schoolnull|School type - Graduate|Finding|false|false||graduatenull|Graduate (person)|Subject|false|false||graduatenull|Current (present time)|Time|false|false||Currentlynull|Academic Research Enhancement Awards|Event|false|false||areanull|Geographic Locations|Entity|false|false||areanull|Area|Modifier|false|false||areanull|Mental concentration|Finding|false|false||concentrationnull|Concentration measurement|LabModifier|false|false||concentrationnull|Difficult (qualifier value)|Finding|false|false||difficultnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Table Frame - above|Finding|false|false||abovenull|Upper|Modifier|false|false||abovenull|Living Alone|Finding|false|false||alonenull|alone - group size|Subject|false|false||alonenull|Singular|LabModifier|false|false||alonenull|student|Subject|false|false||studentnull|Housing Device|Device|false|false||housing
null|Housing|Device|false|false||housingnull|Electrical Current|Phenomenon|true|false||currentnull|Current (present time)|Time|true|false||currentnull|Romantic relationships|Finding|true|false||romantic relationshipsnull|romantic|Finding|true|false||romanticnull|Relationships|Modifier|true|false||relationshipsnull|Female child|Subject|false|false||girl
null|Woman|Subject|false|false||girlnull|Concept Relationship|Finding|true|false||relationship
null|Object Relationship|Finding|true|false||relationshipnull|Relationships|Modifier|true|false||relationshipnull|Female child|Subject|true|false||girl
null|Woman|Subject|true|false||girlnull|Organization Name Type - Legal|Finding|true|false||legal
null|Entity Name Use - Legal|Finding|true|false||legal
null|Legal|Finding|true|false||legalnull|Problems - What subject filter|Finding|true|false||problemsnull|Role Class - access|Finding|true|false||accessnull|Access|Modifier|true|false||accessnull|Guns|Device|true|false||gunsnull|Family Medical History|Finding|false|false||Family Historynull|Entity Name Part Type - family|Finding|false|false||Family
null|Last Name|Finding|false|false||Family
null|Living Arrangement - Family|Finding|false|false||Family
null|Family (taxonomic)|Finding|false|false||Family
null|Family Collection|Finding|false|false||Familynull|Family|Subject|false|false||Familynull|History of present illness (finding)|Finding|false|true||History
null|History of previous events|Finding|false|true||History
null|Historical aspects qualifier|Finding|false|true||History
null|Medical History|Finding|false|true||History
null|Concept History|Finding|false|true||Historynull|History|Subject|false|false||Historynull|Family Medical History|Finding|false|true||Family historynull|Entity Name Part Type - family|Finding|false|false||Family
null|Last Name|Finding|false|false||Family
null|Living Arrangement - Family|Finding|false|false||Family
null|Family (taxonomic)|Finding|false|false||Family
null|Family Collection|Finding|false|false||Familynull|Family|Subject|false|false||Familynull|History of present illness (finding)|Finding|false|true||history
null|History of previous events|Finding|false|true||history
null|Historical aspects qualifier|Finding|false|true||history
null|Medical History|Finding|false|true||history
null|Concept History|Finding|false|true||historynull|History|Subject|false|false||historynull|Indirect exposure mechanism - Father|Finding|false|true||father
null|Relationship - Father|Finding|false|true||father
null|Father - courtesy title|Finding|false|true||fathernull|Father (person)|Subject|false|false||fathernull|Alcohol Problem|Disorder|false|true||alcohol problemsnull|Alcohols|Drug|false|false||alcohol
null|Alcohols|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcoholnull|Alcohol - Recreational Drug Use Code|Finding|false|false||alcoholnull|Problems - What subject filter|Finding|false|true||problemsnull|Cancer Remission|Disorder|false|false||remissionnull|Disease remission|Finding|false|false||remissionnull|Relationship - Mother|Finding|false|false||mothernull|Mother (person)|Subject|false|false||mothernull|Hypothyroidism|Disorder|false|false||hypothyroidismnull|Entity Name Part Type - family|Finding|true|false||family
null|Last Name|Finding|true|false||family
null|Living Arrangement - Family|Finding|true|false||family
null|Family (taxonomic)|Finding|true|false||family
null|Family Collection|Finding|true|false||familynull|Family|Subject|true|false||familynull|Medical referral type|Finding|true|false||medical
null|Medical|Finding|true|false||medical
null|Medical school type|Finding|true|false||medicalnull|Medical service|Procedure|true|false||medicalnull|Psychiatric problem|Disorder|true|false||psychiatric problemsnull|Referral type - Psychiatric|Finding|true|false||psychiatric
null|Psychiatric|Finding|true|false||psychiatricnull|Psychiatric service|Procedure|true|false||psychiatricnull|Psychiatry Specialty|Title|true|false||psychiatricnull|Problems - What subject filter|Finding|true|false||problemsnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|physical examination (physical finding)|Finding|false|false||Physical Examnull|Physical Examination|Procedure|false|false||Physical Examnull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|MYELINATING SCHWANN CELL ELEMENT|Finding|false|false||MSE
null|ENO3 gene|Finding|false|false||MSEnull|White (population group)|Subject|false|false||white
null|Caucasian|Subject|false|false||white
null|Caucasians|Subject|false|false||whitenull|White color|Modifier|false|false||whitenull|Male Gender|Finding|false|false||malenull|Male, Self-Reported|Subject|false|false||male
null|Males|Subject|false|false||malenull|Male Phenotype|Modifier|false|false||malenull|Hospitals|Device|false|false||in hospitalnull|Hospitals|Entity|false|false||in hospitalnull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Anxiety|Disorder|false|false||anxiousnull|Panic Attacks|Disorder|false|false||panic attacknull|Panic|Finding|false|false||panicnull|Attack (finding)|Finding|false|false||attack
null|Attack behavior|Finding|false|false||attacknull|Attack device|Device|false|false||attacknull|Published Interview|Finding|false|false||interviewnull|Interview|Event|false|false||interviewnull|null|Finding|false|false||Speech normalnull|Speech|Finding|false|false||Speechnull|Speech assessment|Procedure|false|false||Speechnull|Amount type - Rate|Finding|false|false||ratenull|Rating (action)|Event|false|false||ratenull|Rate|LabModifier|false|false||ratenull|Volume (publication)|Finding|false|false||volumenull|Volume|LabModifier|false|false||volumenull|Programming Languages|Finding|false|false||languagenull|null|Attribute|false|false||languagenull|Languages|Entity|false|false||languagenull|Mood (psychological function)|Finding|false|false||Mood
null|mood (physical finding)|Finding|false|false||Mood
null|Mood (attribute)|Finding|false|false||Moodnull|null|Attribute|false|false||Moodnull|Depressed mood|Disorder|false|false||depressednull|Constricting sensation quality|Finding|false|false||constrictednull|Concept model range (foundation metadata concept)|Finding|false|false||rangenull|Sample Range|LabModifier|false|false||range
null|Range|LabModifier|false|false||rangenull|Anxiety|Disorder|false|false||anxiousnull|Realm|Finding|false|false||realmnull|null|Finding|false|false||Thoughts
null|Thought|Finding|false|false||Thoughtsnull|Organized|Finding|false|false||organizednull|Guilt|Finding|false|false||guiltnull|Suicidal thoughts|Finding|false|false||suicidal ideationnull|null|Attribute|false|false||suicidal ideationnull|Suicidal|Disorder|false|false||suicidalnull|ideation|Finding|false|false||ideationnull|Infantile Neuroaxonal Dystrophy|Disorder|false|false||plannull|Treatment Plan|Finding|false|false||plan
null|Planned|Finding|false|false||plan
null|null|Finding|false|false||plannull|Commit Lozenge|Drug|false|false||commit
null|Commit Lozenge|Drug|false|false||commitnull|Commit Operation|Procedure|false|false||commitnull|Cancer patients and suicide and depression|Disorder|false|false||suicidenull|Suicide|Finding|false|false||suicidenull|knife|Device|false|false||knifenull|Act Mood - intent|Finding|false|false||intent
null|null|Finding|false|false||intentnull|intent|Modifier|false|false||intentnull|null|Finding|true|false||thoughts
null|Thought|Finding|true|false||thoughtsnull|Insight|Finding|false|false||Insightnull|Patient need for (contextual qualifier)|Finding|false|false||neednull|Needs|Modifier|false|false||neednull|Help document|Finding|false|false||helpnull|Assisted (qualifier value)|Modifier|false|false||helpnull|Language Ability Proficiency - Good|Finding|false|false||good
null|Language Proficiency - Good|Finding|false|false||goodnull|Specimen Quality - Good|Modifier|false|false||good
null|Good|Modifier|false|false||goodnull|Judgment|Finding|false|false||judgmentnull|Fair - language proficiency|Modifier|false|false||fair
null|Fair (qualifier value)|Modifier|false|false||fair
null|Fair Specimen Quality|Modifier|false|false||fairnull|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSEnull|Glucose measurement|Procedure|false|false||GLUCOSEnull|Glucose^1.5H post dose glucagon|Lab|false|false||GLUCOSEnull|urea|Drug|false|false||UREA
null|urea|Drug|false|false||UREA
null|urea|Drug|false|false||UREAnull|Urea measurement|Procedure|false|false||UREAnull|Sodium supplements|Drug|false|false||SODIUM
null|sodium|Drug|false|false||SODIUM
null|sodium|Drug|false|false||SODIUM
null|Sodium Drug Class|Drug|false|false||SODIUMnull|Sodium metabolic function|Finding|false|false||SODIUMnull|Sodium measurement|Procedure|false|false||SODIUMnull|Potassium Drug Class|Drug|false|false||POTASSIUM
null|Dietary Potassium|Drug|false|false||POTASSIUM
null|potassium|Drug|false|false||POTASSIUM
null|potassium|Drug|false|false||POTASSIUM
null|potassium|Drug|false|false||POTASSIUM
null|Potassium supplement|Drug|false|false||POTASSIUM
null|Potassium supplement|Drug|false|false||POTASSIUMnull|Potassium metabolic function|Finding|false|false||POTASSIUMnull|Potassium measurement|Procedure|false|false||POTASSIUMnull|chloride ion|Drug|false|false||CHLORIDE
null|Chlorides|Drug|false|false||CHLORIDEnull|Chloride metabolic function|Finding|false|false||CHLORIDEnull|Chloride measurement|Procedure|false|false||CHLORIDEnull|Total|Modifier|false|false||TOTALnull|carbon dioxide|Drug|false|false||CO2
null|carbon dioxide|Drug|false|false||CO2null|MT-CO2 gene|Finding|false|false||CO2
null|null|Finding|false|false||CO2
null|C2 wt Allele|Finding|false|false||CO2null|blood anion gap (lab test)|Procedure|false|false||ANION GAP
null|Anion gap measurement|Procedure|false|false||ANION GAPnull|Anion Gap|Attribute|false|false||ANION GAPnull|Anion gap result|Lab|false|false||ANION GAPnull|Anions|Drug|false|false||ANIONnull|Ras GTPase-Activating Protein 1, Human|Drug|false|false||GAP
null|Ras GTPase-Activating Protein 1, Human|Drug|false|false||GAP
null|GTPase-Activating Proteins|Drug|false|false||GAP
null|GTPase-Activating Proteins|Drug|false|false||GAPnull|RASA1 wt Allele|Finding|false|false||GAP
null|RASA1 gene|Finding|false|false||GAPnull|Gap (space)|Modifier|false|false||GAPnull|thyrotropin|Drug|false|false||TSH
null|thyrotropin|Drug|false|false||TSH
null|thyrotropin|Drug|false|false||TSHnull|Thyroid stimulating hormone measurement|Procedure|false|false||TSHnull|null|Attribute|false|false||TSHnull|Arylsulfatase A, human|Drug|false|false||ASA
null|Arylsulfatase A, human|Drug|false|false||ASA
null|aspirin|Drug|false|false||ASA
null|aspirin|Drug|false|false||ASAnull|ARSA gene|Finding|false|false||ASAnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|CNS depressants ethanol|Drug|false|false||ETHANOL
null|CNS depressants ethanol|Drug|false|false||ETHANOL
null|antiseptics ethanol|Drug|false|false||ETHANOL
null|antiseptics ethanol|Drug|false|false||ETHANOL
null|ethanol|Drug|false|false||ETHANOL
null|ethanol|Drug|false|false||ETHANOLnull|Toxic effect of ethyl alcohol|Disorder|false|false||ETHANOLnull|Ethanol measurement|Procedure|false|false||ETHANOLnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Hour|Time|false|false||HOURSnull|Random|Modifier|false|false||RANDOMnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Hour|Time|false|false||HOURSnull|Random|Modifier|false|false||RANDOMnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Hold - dosing instruction fragment|Finding|false|false||HOLD
null|hold - Data Operation|Finding|false|false||HOLDnull|Hold (action)|Event|false|false||HOLDnull|Hold - dosing instruction fragment|Finding|false|false||HOLD
null|hold - Data Operation|Finding|false|false||HOLDnull|Hold (action)|Event|false|false||HOLDnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Opiates|Drug|false|false||opiates
null|Opiates|Drug|false|false||opiates
null|Opiates|Drug|false|false||opiates
null|Opiate Alkaloids|Drug|false|false||opiates
null|Opiate Alkaloids|Drug|false|false||opiates
null|Opiate Alkaloids|Drug|false|false||opiatesnull|Opiate Measurement|Procedure|false|false||opiatesnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|cocaine|Drug|false|false||cocaine
null|cocaine|Drug|false|false||cocaine
null|cocaine|Drug|false|false||cocaine
null|cocaine|Drug|false|false||cocainenull|Poisoning by cocaine|Disorder|false|false||cocainenull|Cocaine measurement|Procedure|false|false||cocainenull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||HGB
null|Hemoglobin|Drug|false|false||HGBnull|CYGB gene|Finding|false|false||HGBnull|Hemoglobin concentration|Lab|false|false||HGBnull|Hemopoietic stem cell transplant|Procedure|false|false||HCT
null|Hematocrit Measurement|Procedure|false|false||HCTnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Monos|Drug|false|false||MONOS
null|Mono-S|Drug|false|false||MONOS
null|Monos|Drug|false|false||MONOSnull|SARCOIDOSIS, EARLY-ONSET|Disorder|false|false||EOS
null|Familial eosinophilia|Disorder|false|false||EOSnull|PRSS33 gene|Finding|false|false||EOS
null|IKZF4 gene|Finding|false|false||EOSnull|Eos <Loriini>|Entity|false|false||EOSnull|Primed lymphocyte test|Procedure|false|false||PLTnull|Count Dosing Unit|LabModifier|false|false||COUNT
null|Count|LabModifier|false|false||COUNTnull|Color of urine|Finding|false|false||URINE  COLORnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|color additive|Drug|false|false||COLOR
null|Coloring Excipient|Drug|false|false||COLORnull|color - solid dosage form|Modifier|false|false||COLOR
null|Color|Modifier|false|false||COLORnull|Color quantity|LabModifier|false|false||COLORnull|Yellow color|Modifier|false|false||Yellownull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Hematuria|Disorder|false|false||URINE  BLOODnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|nitrite ion|Drug|false|false||NITRITE
null|Nitrites|Drug|false|false||NITRITE
null|Nitrites|Drug|false|false||NITRITE
null|Nitrites|Drug|false|false||NITRITE
null|nitrite ion|Drug|false|false||NITRITE
null|nitrite ion|Drug|false|false||NITRITEnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Proteins|Drug|false|false||PROTEIN
null|Proteins|Drug|false|false||PROTEINnull|Protein Info|Finding|false|false||PROTEINnull|Protein measurement|Procedure|false|false||PROTEINnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSEnull|Glucose measurement|Procedure|false|false||GLUCOSEnull|Glucose^1.5H post dose glucagon|Lab|false|false||GLUCOSEnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Ketones|Drug|false|false||KETONEnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|bilirubin preparation|Drug|false|false||BILIRUBIN
null|bilirubin preparation|Drug|false|false||BILIRUBIN
null|Bilirubin|Drug|false|false||BILIRUBIN
null|Bilirubin|Drug|false|false||BILIRUBINnull|Bilirubin, total measurement|Procedure|false|false||BILIRUBIN
null|blood bilirubin level test|Procedure|false|false||BILIRUBINnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|BRIEF Health Literacy Screening Tool|Finding|false|false||Brief
null|Behavior Rating Inventory of Executive Function|Finding|false|false||Briefnull|Brief|Time|false|false||Briefnull|Shortened|Modifier|false|false||Briefnull|Hospital course|Finding|false|false||Hospital Coursenull|null|Attribute|false|false||Hospital Coursenull|Organization unit type - Hospital|Finding|false|false||Hospitalnull|Hospitals|Device|false|false||Hospitalnull|Hospitals|Entity|false|false||Hospitalnull|Hospital environment|Modifier|false|false||Hospitalnull|Course|Time|false|false||Coursenull|Referral type - Psychiatric|Finding|false|false||Psychiatric
null|Psychiatric|Finding|false|false||Psychiatricnull|Psychiatric service|Procedure|false|false||Psychiatricnull|Psychiatry Specialty|Title|false|false||Psychiatricnull|Floor (anatomic)|Anatomy|true|false||floornull|floor (object)|Device|true|false||floornull|Floor - story of building|Entity|true|false||floornull|Passive|Modifier|true|false||passivenull|Absence of Biallelic TCRgamma Deletion|Disorder|true|false||abdnull|ABD (body structure)|Anatomy|true|false||abd
null|Abdomen|Anatomy|true|false||abdnull|Act Mood - intent|Finding|true|false||intent
null|null|Finding|true|false||intentnull|intent|Modifier|true|false||intentnull|Infantile Neuroaxonal Dystrophy|Disorder|false|false||plannull|Treatment Plan|Finding|false|false||plan
null|Planned|Finding|false|false||plan
null|null|Finding|false|false||plannull|Still|Disorder|false|false||stillnull|Feeling depressed|Finding|false|false||feeling depressednull|null|Attribute|false|false||feeling depressednull|Depressed mood|Disorder|false|false||depressednull|Anxiety|Disorder|false|false||anxiousnull|Enthusiastic|Finding|false|false||eagernull|Biomaterial Treatment|Finding|false|false||treatment
null|Treating|Finding|false|false||treatment
null|therapeutic aspects|Finding|false|false||treatmentnull|treatment - ActInformationManagementReason|Procedure|false|false||treatment
null|Administration (procedure)|Procedure|false|false||treatment
null|Therapeutic procedure|Procedure|false|false||treatmentnull|MICROCEPHALY, EPILEPSY, AND DIABETES SYNDROME 1|Disorder|false|false||medsnull|Medications|Finding|false|false||medsnull|Celexa|Drug|false|false||celexa
null|Celexa|Drug|false|false||celexanull|Klonopin|Drug|false|false||klonopin
null|Klonopin|Drug|false|false||klonopinnull|Once a day, at bedtime|Time|false|false||QHSnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Anxiety Disorders|Disorder|false|false||anxiety
null|Anxiety|Disorder|false|false||anxietynull|Anxiety symptoms|Finding|false|false||anxietynull|Side|Modifier|true|false||sidenull|Effect|Modifier|true|false||effectsnull|Significant|Finding|true|false||significantnull|Event Seriousness - Significant|Modifier|true|false||significantnull|Alleviating anxiety|Procedure|false|false||anxiety reductionnull|Anxiety Disorders|Disorder|false|false||anxiety
null|Anxiety|Disorder|false|false||anxietynull|Anxiety symptoms|Finding|false|false||anxietynull|Reduced|Finding|false|false||reductionnull|Reduction procedure|Procedure|false|false||reduction
null|Surgical reduction|Procedure|false|false||reductionnull|Reduction (chemical)|Phenomenon|false|false||reductionnull|physiologic resolution|Finding|false|false||resolution
null|Resolution|Finding|false|false||resolutionnull|Resolution Property|LabModifier|false|false||resolutionnull|Depressive Symptoms|Disorder|false|false||depressive symptomsnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Night time|Time|false|false||nightnull|Sibling|Subject|false|false||SIBnull|day|Time|false|false||daysnull|arrival - ActRelationshipType|Finding|false|false||arrivalnull|null|Event|false|false||arrivalnull|Patient's teacher when immunized|Finding|false|false||teachernull|Teacher|Subject|false|false||teachernull|School|Device|false|false||schoolnull|School|Entity|false|false||schoolnull|counselor|Finding|false|false||counselornull|Counselors|Subject|false|false||counselornull|Academic title|Finding|false|false||Academicnull|Academia (organization)|Entity|false|false||Academicnull|Impulsive Behavior|Disorder|false|false||impulsivitynull|apparently|Finding|false|false||apparentlynull|Fighting|Finding|false|false||fightnull|student|Subject|false|false||studentnull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|Housemate|Subject|false|false||roommatenull|Throat Homeopathic Medication|Drug|false|false||throatnull|Specimen Type - Throat|Finding|false|false||throat
null|null|Finding|false|false||throatnull|Throat|Anatomy|false|false||throat
null|Anterior portion of neck|Anatomy|false|false||throat
null|Pharyngeal structure|Anatomy|false|false||throatnull|Very Much|Finding|false|false||a lotnull|Stock (in-store merchandise)|Finding|false|false||lotnull|nucleus of the lateral olfactory tract|Anatomy|false|false||lot
null|Olfactory tract|Anatomy|false|false||lotnull|Lot (entire collection)|Modifier|false|false||lotnull|More|LabModifier|false|false||morenull|Type of bridge device|Device|false|false||bridgesnull|Patient's teacher when immunized|Finding|false|false||teachernull|Teacher|Subject|false|false||teachernull|Teacher|Subject|false|false||teachersnull|Still|Disorder|false|false||stillnull|Unwilling|Finding|false|false||unwillingnull|student|Subject|false|false||studentnull|reputation|Modifier|false|false||reputationnull|Impulsive character (finding)|Disorder|false|false||impulsive
null|Impulsive Behavior|Disorder|false|false||impulsivenull|Necrotizing enterocolitis in fetus OR newborn|Disorder|false|false||NEC
null|Carcinoma, Neuroendocrine|Disorder|false|false||NECnull|null|Finding|false|false||NECnull|null|Modifier|false|false||NECnull|null|LabModifier|false|false||NECnull|REST protein, human|Drug|false|false||rest
null|REST protein, human|Drug|false|false||restnull|REST gene|Finding|false|false||rest
null|site-specific telomere resolvase activity|Finding|false|false||rest
null|Rest|Finding|false|false||restnull|Semester|Time|false|false||semesternull|Medical Leave|Time|false|false||medical leavenull|Medical referral type|Finding|false|false||medical
null|Medical|Finding|false|false||medical
null|Medical school type|Finding|false|false||medicalnull|Medical service|Procedure|false|false||medicalnull|Leave from Employment|Finding|false|false||leavenull|null|Event|false|false||leavenull|Meetings|Event|false|false||meetingnull|Team|Subject|false|false||teamnull|Academic title|Finding|false|false||academicnull|Academia (organization)|Entity|false|false||academicnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|REST protein, human|Drug|false|false||rest
null|REST protein, human|Drug|false|false||restnull|REST gene|Finding|false|false||rest
null|site-specific telomere resolvase activity|Finding|false|false||rest
null|Rest|Finding|false|false||restnull|Semester|Time|false|false||semesternull|Medical leave of absence|Finding|false|false||medical leave of absencenull|Medical Leave|Time|false|false||medical leavenull|Medical referral type|Finding|false|false||medical
null|Medical|Finding|false|false||medical
null|Medical school type|Finding|false|false||medicalnull|Medical service|Procedure|false|false||medicalnull|Leave of Absence - Inactive Reason Code|Finding|false|false||leave of absencenull|Leave of Absence Supply|Procedure|false|false||leave of absencenull|Leave from Employment|Finding|false|false||leavenull|null|Event|false|false||leavenull|Absence (morphologic abnormality)|Disorder|false|false||absencenull|Absent|Finding|false|false||absencenull|next - HtmlLinkType|Finding|false|false||nextnull|Following|Time|false|false||next
null|Then|Time|false|false||nextnull|Adjacent|Modifier|false|false||nextnull|Transaction counts and value totals - year|Finding|false|false||year
null|Precision - year|Finding|false|false||yearnull|year|Time|false|false||yearnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Entity Name Part Type - family|Finding|false|false||family
null|Last Name|Finding|false|false||family
null|Living Arrangement - Family|Finding|false|false||family
null|Family (taxonomic)|Finding|false|false||family
null|Family Collection|Finding|false|false||familynull|Family|Subject|false|false||familynull|Stat (do immediately)|Time|false|false||immediatelynull|Close|Finding|false|false||close
null|Closed|Finding|false|false||closenull|Entity Name Part Type - family|Finding|false|false||family
null|Last Name|Finding|false|false||family
null|Living Arrangement - Family|Finding|false|false||family
null|Family (taxonomic)|Finding|false|false||family
null|Family Collection|Finding|false|false||familynull|Family|Subject|false|false||familynull|Support brand of multivitamin|Drug|false|false||support
null|Support brand of multivitamin|Drug|false|false||support
null|Support brand of multivitamin|Drug|false|false||supportnull|Supportive assistance|Finding|false|false||supportnull|Supportive care|Procedure|false|false||supportnull|Support - dental|Attribute|false|false||supportnull|null|Device|false|false||supportnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Medical referral type|Finding|false|false||medical
null|Medical|Finding|false|false||medical
null|Medical school type|Finding|false|false||medicalnull|Medical service|Procedure|false|false||medicalnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|follow-up|Procedure|false|false||followupnull|Psychiatric therapeutic procedure|Procedure|false|false||psychiatric carenull|Referral type - Psychiatric|Finding|false|false||psychiatric
null|Psychiatric|Finding|false|false||psychiatricnull|Psychiatric service|Procedure|false|false||psychiatricnull|Psychiatry Specialty|Title|false|false||psychiatricnull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|School|Device|false|false||The schoolnull|School|Entity|false|false||The schoolnull|School|Device|false|false||schoolnull|School|Entity|false|false||schoolnull|Satisfied|Finding|false|false||satisfied
null|Satisfaction|Finding|false|false||satisfiednull|Mental state|Finding|false|false||mental statusnull|null|Attribute|false|false||mental status
null|null|Attribute|false|false||mental statusnull|Psyche structure|Finding|false|false||mentalnull|What subject filter - Status|Finding|false|false||statusnull|null|Attribute|false|false||statusnull|Social status|Modifier|false|false||status
null|Status|Modifier|false|false||statusnull|Joint problem|Finding|false|false||jointnull|null|Anatomy|false|false||joint
null|Joints|Anatomy|false|false||joint
null|Articular system|Anatomy|false|false||jointnull|Joint Device|Device|false|false||jointnull|Meetings|Event|false|false||meetingnull|SAFE-Biopharma Standard|Finding|true|false||safenull|Deny (action)|Event|false|false||denynull|Cancer patients and suicide and depression|Disorder|true|false||depression
null|Mental Depression|Disorder|true|false||depression
null|Depressive disorder|Disorder|true|false||depression
null|Depressed mood|Disorder|true|false||depressionnull|Depression - motion|Finding|true|false||depression
null|null|Finding|true|false||depressionnull|Depression - recess|Modifier|true|false||depressionnull|Sibling|Subject|true|false||SIBnull|Future|Time|false|false||futurenull|objective (goal)|Finding|false|false||goal
null|Act Mood - Goal|Finding|false|false||goalnull|SAFE-Biopharma Standard|Finding|false|false||safenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Medical referral type|Finding|false|false||Medical
null|Medical|Finding|false|false||Medical
null|Medical school type|Finding|false|false||Medicalnull|Medical service|Procedure|false|false||Medicalnull|Hospital Stay|Time|true|false||hospital staynull|Organization unit type - Hospital|Finding|true|false||hospitalnull|Hospitals|Device|true|false||hospitalnull|Hospitals|Entity|true|false||hospitalnull|Hospital environment|Modifier|true|false||hospitalnull|Table Rules - groups|Finding|false|false||Groups
null|Groups|Finding|false|false||Groupsnull|Social group|Subject|false|false||Groupsnull|Behavior|Finding|false|false||Behavioralnull|Table Rules - groups|Finding|false|false||groups
null|Groups|Finding|false|false||groupsnull|Social group|Subject|false|false||groupsnull|Visible|Modifier|false|false||visiblenull|Calmodulin 1|Drug|false|false||calm
null|Calmodulin 1|Drug|false|false||calmnull|Feeling calm|Finding|false|false||calm
null|PICALM wt Allele|Finding|false|false||calm
null|SNAP91 gene|Finding|false|false||calm
null|PICALM gene|Finding|false|false||calm
null|SNAP91 wt Allele|Finding|false|false||calmnull|Cancer and Living Meaningfully Therapy|Procedure|false|false||calmnull|Storage Unit|Device|false|false||unit
null|Unit device|Device|false|false||unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||unit
null|Unit of Measure|LabModifier|false|false||unit
null|Unit|LabModifier|false|false||unit
null|Enzyme Unit|LabModifier|false|false||unitnull|Threatening behavior|Finding|true|false||threatening behaviornull|Behavior|Finding|true|false||behaviornull|null|Attribute|true|false||behaviornull|Quiet|Modifier|true|false||quietnull|Room - Patient location type|Modifier|true|false||room
null|Room|Modifier|true|false||roomnull|physical examination (physical finding)|Finding|true|false||physical
null|Physical|Finding|true|false||physicalnull|Physical Examination|Procedure|true|false||physicalnull|Chemical restraint (procedure)|Procedure|true|false||chemical restraintsnull|Chemicals|Drug|true|false||chemicalnull|null|Attribute|true|false||restraintsnull|null|Device|true|false||restraintsnull|null|Time|false|false||at any timenull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|true|false||time
null|Time (foundation metadata concept)|Finding|true|false||time
null|Value type - Time|Finding|true|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|true|false||time
null|Data types - Time|Finding|true|false||time
null|null|Finding|true|false||timenull|Time|Time|true|false||timenull|Organization Name Type - Legal|Finding|false|false||Legal
null|Entity Name Use - Legal|Finding|false|false||Legal
null|Legal|Finding|false|false||Legalnull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|Medication.discharge|Finding|true|false||Discharge Medicationsnull|Body Substance Discharge|Finding|true|false||Discharge
null|Discharge Body Fluid|Finding|true|false||Discharge
null|Body Fluid Discharge|Finding|true|false||Discharge
null|null|Finding|true|false||Dischargenull|Patient Discharge|Procedure|true|false||Dischargenull|Pharmaceutical Preparations|Drug|true|false||Medicationsnull|Medications|Finding|true|false||Medicationsnull|null|Attribute|true|false||Medications
null|null|Attribute|true|false||Medicationsnull|citalopram|Drug|false|false||Citalopram
null|citalopram|Drug|false|false||Citalopramnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|clonazepam|Drug|false|false||Clonazepam
null|clonazepam|Drug|false|false||Clonazepamnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Every morning|Time|false|false||QAMnull|Once a day, at bedtime|Time|false|false||QHSnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|axis i|Finding|false|false||Axis Inull|Fracture of second cervical vertebra|Disorder|false|false||Axisnull|Axis vertebra|Anatomy|false|false||Axisnull|Genus Axis|Entity|false|false||Axisnull|Axis|Modifier|false|false||Axisnull|Major Depressive Disorder|Disorder|true|false||Major depressive disorder
null|Unipolar Depression|Disorder|true|false||Major depressive disordernull|United States Military Commissioned Officer O4 (qualifier value)|Finding|true|false||Majornull|Major <Sympycninae>|Entity|true|false||Majornull|Major|Modifier|true|false||Majornull|Depressive disorder|Disorder|true|false||depressive disordernull|Disease|Disorder|true|false||disordernull|Severe - Severity of Illness Code|Finding|true|false||severe
null|Intensity and Distress 5|Finding|true|false||severe
null|Severe - Triage Code|Finding|true|false||severe
null|Severe (severity modifier)|Finding|true|false||severe
null|Allergy Severity - Severe|Finding|true|false||severenull|Psychotic features|Finding|true|false||psychotic featuresnull|Psychotic Disorders|Disorder|true|false||psychoticnull|Psychotic symptom present|Finding|true|false||psychoticnull|Anxiety Disorders|Disorder|true|false||Anxiety disordernull|Anxiety Disorders|Disorder|true|false||Anxiety
null|Anxiety|Disorder|true|false||Anxietynull|Anxiety symptoms|Finding|true|false||Anxietynull|Disease|Disorder|true|false||disordernull|Specific (qualifier value)|Modifier|true|false||specifiednull|Query Priority - Deferred|Finding|true|false||deferred
null|deferred - ResponseMode|Finding|true|false||deferred
null|Protocol Deferred|Finding|true|false||deferrednull|Deferred|Time|true|false||deferrednull|Status post|Time|false|false||status post
null|Post|Time|false|false||status postnull|What subject filter - Status|Finding|false|false||statusnull|null|Attribute|false|false||statusnull|Social status|Modifier|false|false||status
null|Status|Modifier|false|false||statusnull|Repair of meniscus|Procedure|false|false||meniscus repairnull|Meniscus structure of joint|Anatomy|false|false||meniscusnull|Genus Meniscus|Entity|false|false||meniscusnull|Repair|Finding|false|false||repair
null|Wound Healing|Finding|false|false||repairnull|Repair - Remedial Action|Procedure|false|false||repair
null|Surgical repair|Procedure|false|false||repairnull|Examination of knee joint|Procedure|false|false||kneenull|Knee region structure|Anatomy|false|false||knee
null|Knee|Anatomy|false|false||knee
null|Lower extremity>Knee|Anatomy|false|false||knee
null|Knee joint|Anatomy|false|false||kneenull|Moderate Response|Finding|false|false||moderately
null|Moderate|Finding|false|false||moderately
null|Moderate Effect|Finding|false|false||moderatelynull|Moderate (severity modifier)|Modifier|false|false||moderately
null|Moderation|Modifier|false|false||moderatelynull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|psychosocial stressor|Disorder|false|false||psychosocial stressorsnull|Psychosocial problem|Disorder|false|false||psychosocialnull|Psychosocial|Finding|false|false||psychosocialnull|Stressor|Finding|false|false||stressorsnull|FGF9 protein, human|Drug|false|false||GAF
null|FGF9 protein, human|Drug|false|false||GAFnull|FGF9 wt Allele|Finding|false|false||GAF
null|FGF9 gene|Finding|false|false||GAFnull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Disease|Disorder|false|false||Conditionnull|Logical Condition|Finding|false|false||Conditionnull|null|Attribute|false|false||Conditionnull|Condition|Modifier|false|false||Conditionnull|MYELINATING SCHWANN CELL ELEMENT|Finding|false|false||MSE
null|ENO3 gene|Finding|false|false||MSEnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||generalnull|General medical service|Procedure|false|false||generalnull|Generalized|Modifier|false|false||generalnull|Thin (qualifier value)|Modifier|false|false||thinnull|Caucasian|Subject|false|false||caucasian
null|Caucasians|Subject|false|false||caucasiannull|Caucasian Languages|Entity|false|false||caucasiannull|Male population group|Subject|false|false||man
null|Homo sapiens|Subject|false|false||man
null|Males|Subject|false|false||mannull|Mandinka Language|Entity|false|false||mannull|nicotinamide adenine dinucleotide (NAD)|Drug|true|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|true|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|true|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|true|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|true|false||NAD
null|Dysplastic Nevus|Disorder|true|false||NAD
null|Neuroaxonal Dystrophies|Disorder|true|false||NADnull|patient appears in no acute distress (physical finding)|Finding|true|false||NADnull|Behavior|Finding|true|false||behaviornull|null|Attribute|true|false||behaviornull|Calmodulin 1|Drug|true|false||calm
null|Calmodulin 1|Drug|true|false||calmnull|Feeling calm|Finding|true|false||calm
null|PICALM wt Allele|Finding|true|false||calm
null|SNAP91 gene|Finding|true|false||calm
null|PICALM gene|Finding|true|false||calm
null|SNAP91 wt Allele|Finding|true|false||calmnull|Cancer and Living Meaningfully Therapy|Procedure|true|false||calmnull|Tremor|Finding|true|false||tremorsnull|Tetradecanoylphorbol Acetate|Drug|true|false||PMA
null|4-methoxyamphetamine|Drug|true|false||PMA
null|4-methoxyamphetamine|Drug|true|false||PMA
null|4-methoxyamphetamine|Drug|true|false||PMA
null|Tetradecanoylphorbol Acetate|Drug|true|false||PMA
null|Tetradecanoylphorbol Acetate|Drug|true|false||PMAnull|Progressive Muscular Atrophy|Disorder|true|false||PMAnull|Premarket Device Application|Finding|true|false||PMAnull|null|Finding|true|false||speech- normalnull|Speech|Finding|true|false||speechnull|Speech assessment|Procedure|true|false||speechnull|Affect (mental function)|Finding|true|false||affectnull|assessment of affect|Procedure|true|false||affectnull|More|LabModifier|false|false||morenull|Reactive Therapy|Procedure|false|false||reactivenull|Reactive|Modifier|false|false||reactivenull|null|Time|false|false||priornull|Smiles (finding)|Finding|false|false||smiles
null|Simplified Molecular Input Line Entry Specification|Finding|false|false||smilesnull|Delusions|Disorder|true|false||delusionsnull|Linear|Modifier|false|false||linearnull|objective (goal)|Finding|false|false||goal
null|Act Mood - Goal|Finding|false|false||goalnull|Safety|Phenomenon|true|false||safetynull|Sibling|Subject|true|false||SIBnull|Act Mood - intent|Finding|true|false||intent
null|null|Finding|true|false||intentnull|intent|Modifier|true|false||intentnull|Infantile Neuroaxonal Dystrophy|Disorder|true|false||plannull|Treatment Plan|Finding|true|false||plan
null|Planned|Finding|true|false||plan
null|null|Finding|true|false||plannull|Clusters of Orthologous Groups of Genes|Finding|false|false||cognull|Children's Oncology Group|Entity|false|false||cognull|Fair - language proficiency|Modifier|false|false||fair
null|Fair (qualifier value)|Modifier|false|false||fair
null|Fair Specimen Quality|Modifier|false|false||fairnull|Fair - language proficiency|Modifier|false|false||fair
null|Fair (qualifier value)|Modifier|false|false||fair
null|Fair Specimen Quality|Modifier|false|false||fairnull|Discharge instructions|Finding|false|false||Discharge Instructionsnull|hospital discharge instructions (treatment)|Procedure|false|false||Discharge Instructionsnull|null|Attribute|false|false||Discharge Instructionsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructionsnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|Appointments|Event|false|false||appointmentsnull|feeling unsafe|Finding|false|false||feeling unsafenull|Disease|Disorder|false|false||conditionnull|Logical Condition|Finding|false|false||conditionnull|null|Attribute|false|false||conditionnull|Condition|Modifier|false|false||conditionnull|Patient Outcome - Worsening|Finding|false|false||worseningnull|Worsening (qualifier value)|Modifier|false|false||worseningnull|Call - dosing instruction fragment|Finding|false|false||call
null|Call (Instruction)|Finding|false|false||call
null|Decision|Finding|false|false||call
null|CHL1 gene|Finding|false|false||callnull|Proximal|Modifier|false|false||nearestnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions