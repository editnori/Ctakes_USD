CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Pharmaceutical Preparations|Drug|false|false||MEDICINEnull|Medicine|Title|false|false||MEDICINEnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|codeine|Drug|false|false||Codeine
null|codeine|Drug|false|false||Codeinenull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Chief complaint (finding)|Finding|false|false||Chief Complaintnull|Complaint (finding)|Finding|false|false||Complaintnull|null|Attribute|false|false||Complaintnull|Chest pressure|Finding|false|false|C1527391;C0817096|chest pressurenull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0438716;C0741025|chest
null|Anterior thoracic region|Anatomy|false|false|C0438716;C0741025|chestnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Cardiac attachment|Finding|false|false|C0018787|Cardiacnull|Heart|Anatomy|false|false|C1314974|Cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||Cardiacnull|History of present illness (finding)|Finding|false|false||History of Present Illnessnull|null|Attribute|false|false||History of Present Illnessnull|Medical History|Finding|false|false||History ofnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Present illness|Finding|false|false||Present Illnessnull|Present|Finding|false|false||Present
null|Presentation|Finding|false|false||Presentnull|Illness (finding)|Finding|false|false||Illnessnull|Females|Subject|false|false||female
null|Woman|Subject|false|false||femalenull|Female, Self-Report|Modifier|false|false||female
null|Female Phenotype|Modifier|false|false||femalenull|PMH - past medical history|Finding|false|false||past medical history
null|Medical History|Finding|false|false||past medical historynull|Medical History|Finding|false|false||medical history ofnull|Medical History|Finding|false|false||medical historynull|Medical referral type|Finding|false|false||medical
null|Medical|Finding|false|false||medical
null|Medical school type|Finding|false|false||medicalnull|Medical service|Procedure|false|false||medicalnull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Vessel Positions|Anatomy|false|false||vessel
null|Blood Vessel|Anatomy|false|false||vesselnull|Vessel (unit of presentation)|LabModifier|false|false||vesselnull|Coronary Artery Bypass Surgery|Procedure|false|false||CABGnull|Scalable Vector Graphics|Entity|false|false||SVGnull|Leukocyte adhesion deficiency type 1|Disorder|false|false|C0226032|LAD
null|Leukocyte adhesion deficiency|Disorder|false|false|C0226032|LADnull|ITGB2 wt Allele|Finding|false|false|C0226032|LAD
null|DLD gene|Finding|false|false|C0226032|LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false|C5550999;C0398738;C1414063;C1706333|LADnull|Ladino Language|Entity|false|false||LADnull|Chest pressure|Finding|false|false|C1527391;C0817096|chest pressurenull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0741025;C0438716|chest
null|Anterior thoracic region|Anatomy|false|false|C0741025;C0438716|chestnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0741025|chest
null|Anterior thoracic region|Anatomy|false|false|C0741025|chestnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Initially|Time|false|false||initiallynull|GLAUCOMA, NORMAL TENSION, SUSCEPTIBILITY TO|Finding|false|false||NTG
null|OPA1 wt Allele|Finding|false|false||NTG
null|OPA1 gene|Finding|false|false||NTGnull|Relief brand of phenylephrine|Drug|false|false||relief
null|Relief brand of phenylephrine|Drug|false|false||reliefnull|Feeling relief|Finding|false|false||reliefnull|Short menstrual periods|Finding|false|false||short periodnull|Shortened|Modifier|false|false||shortnull|Short Value|LabModifier|false|false||short
null|Short|LabModifier|false|false||shortnull|Menstruation|Finding|false|false||periodnull|Clinical Trial Period|Procedure|false|false||periodnull|per period (qualifier value)|Time|false|false||period
null|Time periods|Time|false|false||periodnull|Transaction counts and value totals - Period|LabModifier|false|false||periodnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Radiating to|Finding|false|false||radiatednull|RIGHT SIDE (USED TO IDENTIFY PROCEDURES PERFORMED ON THE RIGHT SIDE OF THE BODY)|Modifier|false|false||right side
null|Right|Modifier|false|false||right sidenull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Side|Modifier|false|false||sidenull|Both upper arms|Anatomy|false|false|C5575339;C2681631;C5782111;C0206655|both armsnull|Alveolar rhabdomyosarcoma|Disorder|false|false|C0446516;C0230348|armsnull|Adherence to Refills and Medications Scale|Finding|false|false|C0230348;C0446516|arms
null|KIDINS220 gene|Finding|false|false|C0230348;C0446516|armsnull|Upper arm|Anatomy|false|false|C5782111;C0206655;C5575339;C2681631|armsnull|null|Attribute|false|false|C0446516;C0230348|armsnull|Increased sweating|Finding|false|false||diaphoresisnull|Associated with|Modifier|false|false||associatednull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|Vomiting|Finding|true|false||vomitingnull|Lightheadedness|Finding|false|false||lightheadednessnull|Dizziness|Finding|false|false||dizziness
null|Vertigo|Finding|false|false||dizzinessnull|MILDLY|Modifier|false|false||mildly
null|Mild (qualifier value)|Modifier|false|false||mildlynull|Dyspnea|Finding|false|false||SOBnull|Recent|Time|false|false||recentnull|Pneumonia|Disorder|false|false||pneumonianull|Firstly|Modifier|false|false||firstnull|First (number)|LabModifier|false|false||firstnull|week|Time|false|false||weeksnull|FBXW7 wt Allele|Finding|false|false||ago
null|FBXW7 gene|Finding|false|false||agonull|null|Finding|false|false||dyspnea
null|Dyspnea|Finding|false|false||dyspneanull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|Very|Modifier|false|false||verynull|Minimal|Modifier|false|false||minimal
null|Mild (qualifier value)|Modifier|false|false||minimal
null|Minimum|Modifier|false|false||minimalnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|Address type - Office|Finding|false|false||officenull|Office|Device|false|false||officenull|Organization unit type - Office|Entity|false|false||officenull|New LBBB|Finding|false|false||new LBBBnull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|Left Bundle-Branch Block|Disorder|false|false||LBBBnull|null|Lab|false|false||LBBBnull|Adenohypophyseal Diseases|Disorder|false|false||anteriornull|Anterior|Modifier|false|false||anteriornull|Elevation|Modifier|false|false||elevationsnull|Plavix|Drug|false|false||Plavix
null|Plavix|Drug|false|false||Plavixnull|aspirin|Drug|false|false||Aspirin
null|aspirin|Drug|false|false||Aspirinnull|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparinnull|ST segment elevation myocardial infarction|Disorder|false|false||STEMInull|ST Elevation Myocardial Infarction by ECG Finding|Finding|false|false||STEMInull|Catheterization|Procedure|false|false||cathnull|AML Lab Table|Finding|false|false||lab
null|LAT2 gene|Finding|false|false||lab
null|EWS Lab Table|Finding|false|false||labnull|Laboratory|Device|false|false||labnull|Labrador retriever|Entity|false|false||lab
null|Laboratory|Entity|false|false||labnull|Catheterization|Procedure|false|false||Cathnull|Occluded|Finding|false|false||occluded
null|Obstruction|Finding|false|false||occludednull|Scalable Vector Graphics|Entity|false|false||SVGnull|Native (qualifier value)|Finding|false|false||Nativenull|Occluded|Finding|false|false|C0226032|occluded
null|Obstruction|Finding|false|false|C0226032|occludednull|Proximal Resection Margin|Attribute|false|false||proximalnull|Proximal|Modifier|false|false||proximalnull|Leukocyte adhesion deficiency type 1|Disorder|false|false|C0226032|LAD
null|Leukocyte adhesion deficiency|Disorder|false|false|C0226032|LADnull|ITGB2 wt Allele|Finding|false|false|C0226032|LAD
null|DLD gene|Finding|false|false|C0226032|LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false|C0028778;C1947917;C5550999;C0398738;C1414063;C1706333|LADnull|Ladino Language|Entity|false|false||LADnull|Leukocyte adhesion deficiency type 1|Disorder|false|false|C0226032|LAD
null|Leukocyte adhesion deficiency|Disorder|false|false|C0226032|LADnull|ITGB2 wt Allele|Finding|false|false|C0226032|LAD
null|DLD gene|Finding|false|false|C0226032|LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false|C5550999;C0398738;C1414063;C1706333|LADnull|Ladino Language|Entity|false|false||LADnull|Difficult (qualifier value)|Finding|false|false||difficultnull|Concern|Finding|false|false||concernnull|Possible|Finding|false|false||possiblenull|Possible diagnosis|Modifier|false|false||possible
null|Possibly Related to Intervention|Modifier|false|false||possiblenull|Dissecting hemorrhage|Finding|false|false||dissectionnull|Tissue Dissection|Procedure|false|false||dissectionnull|Burning Mouth Syndrome|Disorder|false|false|C0226032|BMSnull|Proximal Resection Margin|Attribute|false|false||proximalnull|Proximal|Modifier|false|false||proximalnull|Leukocyte adhesion deficiency type 1|Disorder|false|false|C0226032|LAD
null|Leukocyte adhesion deficiency|Disorder|false|false|C0226032|LADnull|ITGB2 wt Allele|Finding|false|false|C0226032|LAD
null|DLD gene|Finding|false|false|C0226032|LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false|C1414063;C1706333;C5550999;C0398738;C0006430|LADnull|Ladino Language|Entity|false|false||LADnull|Distal Resection Margin|Attribute|false|false|C0226032|Distalnull|Distal (qualifier value)|Modifier|false|false||Distalnull|Leukocyte adhesion deficiency type 1|Disorder|false|false|C0226032|LAD
null|Leukocyte adhesion deficiency|Disorder|false|false|C0226032|LADnull|ITGB2 wt Allele|Finding|false|false|C0226032|LAD
null|DLD gene|Finding|false|false|C0226032|LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false|C1704338;C5550999;C0398738;C0011900;C4522154;C3842384;C1414063;C1706333|LADnull|Ladino Language|Entity|false|false||LADnull|Diminutive|Finding|false|false|C0226032|diminutivenull|Septal|Modifier|false|false||septalnull|diagnosis aspects|Finding|false|false|C0226032|diagnull|Diagnosis|Procedure|false|false|C0226032|diagnull|Hemodynamically stable|Finding|false|false||hemodynamically stablenull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Androgen Binding Protein|Drug|false|false||SBP
null|Androgen Binding Protein|Drug|false|false||SBPnull|CCHCR1 wt Allele|Finding|false|false||SBP
null|SHBG wt Allele|Finding|false|false||SBPnull|Systolic blood pressure measurement|Procedure|false|false||SBPnull|Systolic Pressure|Attribute|false|false||SBPnull|Floor (anatomic)|Anatomy|false|false|C0008031;C0741025;C1549543;C0030193|floornull|floor (object)|Device|false|false||floornull|Floor - story of building|Entity|false|false||floornull|Current (present time)|Time|false|false||currentlynull|Chest Pain|Finding|false|false|C1527391;C0817096;C3714591|chest painnull|null|Attribute|false|false|C1527391;C0817096|chest painnull|Chest problem|Finding|false|false|C1527391;C0817096;C3714591|chestnull|Chest|Anatomy|false|false|C0741025;C2926613;C0008031|chest
null|Anterior thoracic region|Anatomy|false|false|C0741025;C2926613;C0008031|chestnull|Pain-Free|Drug|false|false||pain freenull|Administration Method - Pain|Finding|false|false|C3714591|pain
null|Pain|Finding|false|false|C3714591|painnull|null|Attribute|false|false||painnull|Free of (attribute)|Finding|false|false||freenull|Empty (qualifier)|Modifier|false|false||freenull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Review of systems (procedure)|Procedure|false|false||review of systemsnull|null|Attribute|false|false||review of systems
null|null|Attribute|false|false||review of systemsnull|Review of|Finding|false|false||review ofnull|Review (Publication Type)|Finding|false|false||review
null|Act Class - review|Finding|false|false||reviewnull|System|Finding|false|false||systemsnull|null|Time|false|false||priornull|Medical History|Finding|true|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Deep Resection Margin|Attribute|true|false||deepnull|Deep (qualifier value)|Modifier|false|false||deepnull|Venous thrombosis after immobility|Finding|false|false|C0042449|venous thrombosis
null|Venous Thrombosis|Finding|false|false|C0042449|venous thrombosisnull|Veins|Anatomy|false|false|C0517555;C0042487|venousnull|Venous|Modifier|false|false||venousnull|Thrombosis|Finding|false|false||thrombosisnull|Pulmonary Embolism|Finding|false|false|C0024109|pulmonary embolismnull|Pulmonary (intended site)|Finding|false|false|C0024109|pulmonarynull|Lung|Anatomy|false|false|C0034065;C1704212;C0013922;C4522268;C2707265|pulmonarynull|null|Attribute|false|false|C0024109|pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Embolism|Finding|false|false|C0024109|embolism
null|Embolus|Finding|false|false|C0024109|embolismnull|Hemorrhage|Finding|false|false||bleedingnull|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Myalgia|Finding|false|false||myalgiasnull|Arthralgia|Finding|false|false|C0392905;C1269611;C0022417|joint painsnull|Joint problem|Finding|false|false|C0392905;C1269611;C0022417|jointnull|null|Anatomy|false|false|C0003862;C0575044;C0030193|joint
null|Joints|Anatomy|false|false|C0003862;C0575044;C0030193|joint
null|Articular system|Anatomy|false|false|C0003862;C0575044;C0030193|jointnull|Joint Device|Device|false|false||jointnull|Pain|Finding|false|false|C0392905;C1269611;C0022417|painsnull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|Hemoptysis|Finding|false|false||hemoptysisnull|null|Finding|false|false||black stools
null|Melena|Finding|false|false||black stoolsnull|Black - ethnic group (ethnic group)|Subject|false|false||black
null|Black race|Subject|false|false||black
null|African|Subject|false|false||blacknull|Black - Structured Product Labeling Color|Modifier|false|false||black
null|Black color|Modifier|false|false||blacknull|Feces|Finding|false|false||stoolsnull|null|Attribute|false|false||stoolsnull|Stool seat|Device|false|false||stoolsnull|Red stools|Finding|false|false||red stoolsnull|DYRK3 gene|Finding|false|false||red
null|Redness|Finding|false|false||red
null|IK gene|Finding|false|false||rednull|Radiological Exposure Device|Device|false|false||rednull|Red color|Modifier|false|false||rednull|Feces|Finding|false|false||stoolsnull|null|Attribute|false|false||stoolsnull|Stool seat|Device|false|false||stoolsnull|Recent|Time|false|false||recentnull|Fever|Finding|true|false||feversnull|Chills|Finding|true|false||chillsnull|Rigor - Temperature-associated observation|Finding|true|false||rigorsnull|Review of systems (procedure)|Procedure|false|false||review of systemsnull|null|Attribute|false|false||review of systems
null|null|Attribute|false|false||review of systemsnull|Review of|Finding|false|false||review ofnull|Review (Publication Type)|Finding|false|false||review
null|Act Class - review|Finding|false|false||reviewnull|System|Finding|false|false||systemsnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Cardiac attachment|Finding|false|false|C0018787|Cardiacnull|Heart|Anatomy|false|false|C1314974;C1552617;C0282443;C0699752;C0489633;C0449913|Cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||Cardiacnull|Review of systems (procedure)|Procedure|false|false|C0018787|review of systemsnull|null|Attribute|false|false||review of systems
null|null|Attribute|false|false||review of systemsnull|Review of|Finding|false|false|C0018787|review ofnull|Review (Publication Type)|Finding|false|false|C0018787|review
null|Act Class - review|Finding|false|false|C0018787|reviewnull|System|Finding|false|false|C0018787|systemsnull|Absent|Finding|false|false||absence ofnull|Absence (morphologic abnormality)|Disorder|false|false||absencenull|Absent|Finding|false|false||absencenull|Chest Pain|Finding|false|false|C1527391;C0817096|chest painnull|null|Attribute|false|false|C1527391;C0817096|chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0741025;C2926613;C0008031|chest
null|Anterior thoracic region|Anatomy|false|false|C0741025;C2926613;C0008031|chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Dyspnea on exertion|Finding|false|false||dyspnea on exertionnull|null|Finding|false|false||dyspnea
null|Dyspnea|Finding|false|false||dyspneanull|Exertion|Finding|false|false||exertionnull|Paroxysmal nocturnal dyspnea|Disorder|false|false||paroxysmal nocturnal dyspneanull|Paroxysmal|Time|false|false||paroxysmalnull|null|Finding|false|false||dyspnea
null|Dyspnea|Finding|false|false||dyspneanull|sleeping upright or using specific number of extra pillows (orthopnea)|Finding|false|false||orthopnea
null|Orthopnea|Finding|false|false||orthopneanull|Ankle edema (finding)|Finding|false|false|C0003086;C0003087;C4284979|ankle edemanull|Lower extremity>Ankle|Anatomy|false|false|C0013604;C0235439|ankle
null|Ankle|Anatomy|false|false|C0013604;C0235439|ankle
null|Ankle joint structure|Anatomy|false|false|C0013604;C0235439|anklenull|Edema|Finding|false|false|C0003086;C0003087;C4284979|edemanull|null|Attribute|false|false||edemanull|Palpitations|Finding|false|false||palpitationsnull|Presyncope or syncope|Finding|false|false||syncope or presyncopenull|Syncope|Finding|false|false||syncopenull|Syncope <Gastrophryninae>|Entity|false|false||syncopenull|Presyncope|Finding|false|false||presyncopenull|PMH - past medical history|Finding|false|false||Past Medical History
null|Medical History|Finding|false|false||Past Medical Historynull|Medical History|Finding|false|false||Medical Historynull|Medical referral type|Finding|false|false||Medical
null|Medical|Finding|false|false||Medical
null|Medical school type|Finding|false|false||Medicalnull|Medical service|Procedure|false|false||Medicalnull|Medical History|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|History of present illness (finding)|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|cardiac risk factors|Finding|false|false|C0018787|CARDIAC RISK FACTORSnull|CARD.RISK|Finding|false|false|C0018787|CARDIAC RISKnull|Cardiac attachment|Finding|false|false|C0018787|CARDIACnull|Heart|Anatomy|false|false|C1830376;C1314974;C2024776;C1553898;C0455624;C0035648;C0035647;C3176821|CARDIACnull|Cardiac - anatomy qualifier|Modifier|false|false||CARDIACnull|risk factors - observation list|Finding|false|false|C0018787|RISK FACTORS
null|risk factors|Finding|false|false|C0018787|RISK FACTORS
null|History of - risk factor|Finding|false|false|C0018787|RISK FACTORSnull|null|Attribute|false|false|C0018787|RISK FACTORSnull|Risk|Finding|false|false|C0018787|RISKnull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||Diabetes
null|Diabetes|Disorder|false|false||Diabetes
null|Diabetes Mellitus|Disorder|false|false||Diabetesnull|Dyslipidemias|Disorder|false|false||Dyslipidemianull|Hypertensive disease|Disorder|false|false||Hypertensionnull|Cardiac attachment|Finding|true|false|C0018787|CARDIACnull|Heart|Anatomy|false|false|C0262926;C1705255;C0019665;C0262512;C2004062;C1314974|CARDIACnull|Cardiac - anatomy qualifier|Modifier|false|false||CARDIACnull|History of present illness (finding)|Finding|false|false|C0018787|HISTORY
null|History of previous events|Finding|false|false|C0018787|HISTORY
null|Historical aspects qualifier|Finding|false|false|C0018787|HISTORY
null|Medical History|Finding|false|false|C0018787|HISTORY
null|Concept History|Finding|false|false|C0018787|HISTORYnull|History|Subject|false|false||HISTORYnull|Coronary Artery Bypass Surgery|Procedure|false|false||CABGnull|Following|Time|false|false||subsequentnull|Vessel Positions|Anatomy|false|false||vessel
null|Blood Vessel|Anatomy|false|false||vesselnull|Vessel (unit of presentation)|LabModifier|false|false||vesselnull|Coronary Artery Bypass Surgery|Procedure|false|false||CABGnull|Scalable Vector Graphics|Entity|false|false||SVGnull|Leukocyte adhesion deficiency type 1|Disorder|false|false|C0226032|LAD
null|Leukocyte adhesion deficiency|Disorder|false|false|C0226032|LADnull|ITGB2 wt Allele|Finding|false|false|C0226032|LAD
null|DLD gene|Finding|false|false|C0226032|LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false|C5550999;C0398738;C1414063;C1706333|LADnull|Ladino Language|Entity|false|false||LADnull|Percutaneous Coronary Intervention|Procedure|false|false|C0018787|PERCUTANEOUS CORONARY INTERVENTIONSnull|Percutaneous Route of Drug Administration|Finding|false|false|C0018787|PERCUTANEOUSnull|Percutaneous|Modifier|false|false||PERCUTANEOUSnull|Heart|Anatomy|false|false|C1522243;C0886296;C1273869;C1532338|CORONARYnull|Coronary|Modifier|false|false||CORONARYnull|Nursing interventions|Procedure|false|false|C0018787|INTERVENTIONS
null|Intervention regimes|Procedure|false|false|C0018787|INTERVENTIONSnull|null|Attribute|false|false||INTERVENTIONSnull|Pacing up and down|Finding|false|false||PACINGnull|Disruptive, Impulse Control, and Conduct Disorders|Disorder|false|false||ICD
null|Type II Mucolipidosis|Disorder|false|false||ICDnull|International Classification of Diseases|Finding|false|false||ICD
null|GNPTAB wt Allele|Finding|false|false||ICDnull|Icd Regimen|Procedure|false|false||ICDnull|between lunch and dinner|Time|false|false||ICDnull|PMH - past medical history|Finding|false|false||PAST MEDICAL HISTORY
null|Medical History|Finding|false|false||PAST MEDICAL HISTORYnull|Medical History|Finding|false|false||MEDICAL HISTORYnull|Medical referral type|Finding|false|false||MEDICAL
null|Medical|Finding|false|false||MEDICAL
null|Medical school type|Finding|false|false||MEDICALnull|Medical service|Procedure|false|false||MEDICALnull|Medical History|Finding|false|false||HISTORY
null|History of previous events|Finding|false|false||HISTORY
null|Historical aspects qualifier|Finding|false|false||HISTORY
null|History of present illness (finding)|Finding|false|false||HISTORY
null|Concept History|Finding|false|false||HISTORYnull|History|Subject|false|false||HISTORYnull|Cyclophosphamide/Doxorubicin/Vincristine|Drug|false|false||CVAnull|Acute ill-defined cerebrovascular disease|Disorder|false|false||CVA
null|Cerebrovascular accident|Disorder|false|false||CVAnull|Small|LabModifier|false|false||smallnull|Left posterior|Modifier|false|false||left posteriornull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Posterior pituitary disease|Disorder|false|false||posteriornull|Dorsal|Modifier|false|false||posteriornull|Coronal (qualifier value)|Modifier|false|false||frontalnull|Infarction|Finding|false|false||infarctnull|Tablet Dosage Form|Drug|false|false||tabnull|Tablet Dosing Unit|LabModifier|false|false||tabnull|Plavix|Drug|false|false||plavix
null|Plavix|Drug|false|false||plavixnull|Daily|Time|false|false||dailynull|Hypercholesterolemia|Disorder|false|false||hypercholesterolemianull|Hypercholesterolemia result|Finding|false|false||hypercholesterolemianull|Small|LabModifier|false|false||smallnull|macular|Modifier|false|false||Macularnull|Social and personal history|Finding|false|false||Social History
null|Social History|Finding|false|false||Social Historynull|Social|Finding|false|false||Socialnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Family Medical History|Finding|false|false||Family Historynull|Entity Name Part Type - family|Finding|false|false||Family
null|Last Name|Finding|false|false||Family
null|Living Arrangement - Family|Finding|false|false||Family
null|Family (taxonomic)|Finding|false|false||Family
null|Family Collection|Finding|false|false||Familynull|Family|Subject|false|false||Familynull|History of present illness (finding)|Finding|false|true||History
null|History of previous events|Finding|false|true||History
null|Historical aspects qualifier|Finding|false|true||History
null|Medical History|Finding|false|true||History
null|Concept History|Finding|false|true||Historynull|History|Subject|false|false||Historynull|Indirect exposure mechanism - Father|Finding|false|false||father
null|Relationship - Father|Finding|false|false||father
null|Father - courtesy title|Finding|false|false||fathernull|Father (person)|Subject|false|false||fathernull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Glycation End Products, Advanced|Drug|false|false||age
null|Glycation End Products, Advanced|Drug|false|false||agenull|null|Attribute|false|false||agenull|Age|Subject|false|false||agenull|Relationship - Mother|Finding|false|false||mothernull|Mother (person)|Subject|false|false||mothernull|Malignant neoplasm of stomach|Disorder|false|false|C3714551;C0038351;C4266636|stomach cancer
null|Stomach Carcinoma|Disorder|false|false|C3714551;C0038351;C4266636|stomach cancernull|Neoplasm of uncertain or unknown behavior of stomach|Disorder|false|false|C3714551;C0038351;C4266636|stomach
null|Stomach Diseases|Disorder|false|false|C3714551;C0038351;C4266636|stomach
null|Benign neoplasm of stomach|Disorder|false|false|C3714551;C0038351;C4266636|stomach
null|Carcinoma in situ of stomach|Disorder|false|false|C3714551;C0038351;C4266636|stomachnull|Stomach problem|Finding|false|false|C3714551;C0038351;C4266636|stomachnull|Procedure on stomach|Procedure|false|false|C3714551;C0038351;C4266636|stomachnull|Stomach structure|Anatomy|false|false|C0038354;C0496905;C0153943;C0154060;C0024623;C0699791;C0577027;C0872393;C0585442;C0279530;C0006826;C0006826;C1546560;C1550616|stomach
null|Abdomen>Stomach|Anatomy|false|false|C0038354;C0496905;C0153943;C0154060;C0024623;C0699791;C0577027;C0872393;C0585442;C0279530;C0006826;C0006826;C1546560;C1550616|stomach
null|Stomach|Anatomy|false|false|C0038354;C0496905;C0153943;C0154060;C0024623;C0699791;C0577027;C0872393;C0585442;C0279530;C0006826;C0006826;C1546560;C1550616|stomachnull|Malignant Neoplasms|Disorder|false|false|C3714551;C0038351;C4266636|cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Malignant Bone Neoplasm|Disorder|false|false|C1442209;C0262950;C3714551;C0038351;C4266636|bone cancer
null|Osteosarcoma of bone|Disorder|false|false|C1442209;C0262950;C3714551;C0038351;C4266636|bone cancernull|Specimen Type - Bone|Finding|false|false|C1442209;C0262950;C3714551;C0038351;C4266636|bone
null|null|Finding|false|false|C1442209;C0262950;C3714551;C0038351;C4266636|bonenull|Skeletal bone|Anatomy|false|false|C1546560;C1550616;C0585442;C0279530|bone
null|XXX bone|Anatomy|false|false|C1546560;C1550616;C0585442;C0279530|bonenull|Malignant Neoplasms|Disorder|false|false|C3714551;C0038351;C4266636|cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|physical examination (physical finding)|Finding|false|false||Physical Examnull|Physical Examination|Procedure|false|false||Physical Examnull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||GENERALnull|General medical service|Procedure|false|false||GENERALnull|Generalized|Modifier|false|false||GENERALnull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|Oriented to place|Finding|false|false||Orientednull|Orientation, Spatial|Modifier|false|false||Orientednull|Mood (psychological function)|Finding|false|false||Mood
null|mood (physical finding)|Finding|false|false||Mood
null|Mood (attribute)|Finding|false|false||Moodnull|null|Attribute|false|false||Moodnull|Appropriate|Modifier|false|false||appropriatenull|HEENT|Anatomy|false|false||HEENTnull|Scleral Diseases|Disorder|false|false|C0036410|Scleranull|examination of sclera|Procedure|false|false|C0036410|Scleranull|Sclera|Anatomy|false|false|C0036412;C0205180;C2228481|Scleranull|Anicteric|Finding|false|false|C0036410|anictericnull|Pupil equal round and reacting to light|Finding|false|false||PERRLnull|Malignant neoplasm of conjunctiva|Disorder|false|false|C0229274;C0009758|Conjunctiva
null|Benign neoplasm of conjunctiva|Disorder|false|false|C0229274;C0009758|Conjunctiva
null|Conjunctival Diseases|Disorder|false|false|C0229274;C0009758|Conjunctivanull|Specimen Type - Conjunctiva|Finding|false|false|C0229274;C0009758|Conjunctiva
null|null|Finding|false|false|C0229274;C0009758|Conjunctivanull|examination of conjunctiva|Procedure|false|false|C0229274;C0009758|Conjunctiva
null|Procedure on conjunctiva|Procedure|false|false|C0229274;C0009758|Conjunctivanull|Structure of palpebral conjunctiva|Anatomy|false|false|C0872390;C2228431;C1550624;C1546576;C0153628;C0154025;C0009759|Conjunctiva
null|conjunctiva|Anatomy|false|false|C0872390;C2228431;C1550624;C1546576;C0153628;C0154025;C0009759|Conjunctivanull|Pink color|Modifier|false|false||pinknull|Pallor of skin|Finding|true|false|C0026724;C0026639|pallornull|Cyanosis|Finding|true|false|C0026639;C0026724|cyanosisnull|Oral mucous membrane structure|Anatomy|false|false|C1561514;C1527415;C4521986;C1272919;C0010520;C0241137|oral mucosanull|Oral Dosage Form|Drug|false|false|C0026724;C0026639;C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0026639;C0226896;C0026724|oral
null|Oral (intended site)|Finding|false|false|C0026639;C0226896;C0026724|oralnull|Oral cavity|Anatomy|false|false|C1561514;C1272919;C1527415;C4521986|oralnull|Oral|Modifier|false|false||oralnull|null|Finding|false|false|C0226896;C0026639;C0026724|mucosanull|Mucous Membrane|Anatomy|false|false|C1272919;C0241137;C0010520;C1561514;C1527415;C4521986|mucosanull|Passive joint movement of neck (finding)|Finding|false|false|C0027530;C3159206|NECK
null|Neck problem|Finding|false|false|C0027530;C3159206|NECKnull|dendritic spine neck|Anatomy|false|false|C0812434;C0684335|NECK
null|Neck|Anatomy|false|false|C0812434;C0684335|NECKnull|Supple|Finding|false|false||Supplenull|Jugular venous pressure|Finding|false|false||JVPnull|Cardiac attachment|Finding|false|false|C0018787|CARDIACnull|Heart|Anatomy|false|false|C1314974|CARDIACnull|Cardiac - anatomy qualifier|Modifier|false|false||CARDIACnull|Point of Maximum Impulse|Finding|false|false|C4085247;C0230136|PMI
null|TMEM11 gene|Finding|false|false|C4085247;C0230136|PMI
null|PMM2 wt Allele|Finding|false|false|C4085247;C0230136|PMI
null|PMM2 gene|Finding|false|false|C4085247;C0230136|PMI
null|MPI gene|Finding|false|false|C4085247;C0230136|PMInull|Prostate Mechanical Imager|Device|false|false||PMInull|Space of intercostal compartment|Anatomy|false|false|C0282173;C1823304;C5780972;C5238618;C1418674;C1417244|intercostal space
null|Structure of intercostal space|Anatomy|false|false|C0282173;C1823304;C5780972;C5238618;C1418674;C1417244|intercostal spacenull|Intercostal|Modifier|false|false||intercostalnull|Space (Astronomy)|Phenomenon|false|false|C4085247;C0230136|spacenull|Space - property|Modifier|false|false||spacenull|Midclavicular|Modifier|false|false||midclavicularnull|Line Specimen|Drug|false|false||line
null|Long Interspersed Elements|Drug|false|false||line
null|Long Interspersed Elements|Drug|false|false||linenull|line source specimen code|Finding|false|false||linenull|Intravascular line|Device|false|false||linenull|Linear|Modifier|false|false||linenull|Line Unit of Length|LabModifier|false|false||linenull|Cardiac thrill (finding)|Finding|true|false||thrillsnull|hoist [device]|Device|true|false||liftsnull|Lung|Anatomy|false|false||LUNGSnull|Deformity of chest wall|Disorder|true|false|C0205076;C4266615;C1527391;C0817096|chest wall deformitiesnull|Chest wall structure|Anatomy|false|false|C3164427|chest wall
null|Chest>Chest wall|Anatomy|false|false|C3164427|chest wallnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0741025;C3164427|chest
null|Anterior thoracic region|Anatomy|false|false|C0741025;C3164427|chestnull|Walls of a building|Device|false|false||wallnull|Congenital Abnormality|Disorder|true|false||deformitiesnull|deformities qualifier|Modifier|false|false||deformitiesnull|Congenital scoliosis|Disorder|true|false||scoliosis
null|null|Disorder|true|false||scoliosis
null|Acquired scoliosis|Disorder|true|false||scoliosisnull|Kyphosis deformity of spine|Disorder|true|false||kyphosis
null|Acquired kyphosis|Disorder|true|false||kyphosis
null|Congenital kyphosis|Disorder|true|false||kyphosisnull|kyphosis|Finding|true|false||kyphosisnull|Respiratory, thoracic and mediastinal disorders|Disorder|false|false||Respnull|Respiratory rate|Attribute|false|false||Respnull|Unlabored|Finding|false|false||unlaborednull|Use of accessory muscles|Finding|true|false|C4083049;C0026845|accessory muscle usenull|Accessory skeletal muscle|Disorder|true|false|C4083049;C0026845|accessory musclenull|Accessory|Device|true|false||accessorynull|Muscle (organ)|Anatomy|false|false|C1821466;C0158784;C1947944;C0042153;C0457083|muscle
null|Muscle Tissue|Anatomy|false|false|C1821466;C0158784;C1947944;C0042153;C0457083|musclenull|Use - dosing instruction imperative|Finding|true|false|C4083049;C0026845|use
null|utilization qualifier|Finding|true|false|C4083049;C0026845|use
null|Usage|Finding|true|false|C4083049;C0026845|usenull|Cancer/Testis Antigen|Drug|false|false||CTAnull|PCYT1A wt Allele|Finding|false|false||CTA
null|CERNA3 gene|Finding|false|false||CTAnull|Cardiac Computerized Tomographic Angiography|Procedure|false|false||CTAnull|Basilar Rales|Finding|false|false||crackles
null|Rales|Finding|false|false||cracklesnull|Wheezing|Finding|false|false||wheezesnull|Rhonchi|Finding|false|false||rhonchinull|Malignant neoplasm of abdomen|Disorder|false|false|C0230168;C0000726|ABDOMENnull|Abdomen problem|Finding|false|false|C0230168;C0000726|ABDOMENnull|Abdomen|Anatomy|false|false|C0941288;C0153662|ABDOMEN
null|Abdominal Cavity|Anatomy|false|false|C0941288;C0153662|ABDOMENnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||Softnull|Soft|Modifier|false|false||Softnull|LRRC4B gene|Finding|true|false||HSMnull|Emotional tenderness|Finding|true|false||tenderness
null|Sore to touch|Finding|true|false||tendernessnull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false|C0449202;C0000726;C4037978;C0003483|Abdnull|ABD (body structure)|Anatomy|false|false|C3811055;C0869784|Abd
null|Abdomen|Anatomy|false|false|C3811055;C0869784|Abdnull|Procedure on aorta|Procedure|false|false|C4037978;C0003483;C0449202;C0000726|aortanull|Chest+Abdomen>Aorta|Anatomy|false|false|C3811055;C0869784|aorta
null|Aorta|Anatomy|false|false|C3811055;C0869784|aortanull|Palpation|Procedure|false|false||palpationnull|Bruit|Finding|true|false||bruitsnull|All extremities|Anatomy|false|false||EXTREMITIES
null|Limb structure|Anatomy|false|false||EXTREMITIESnull|Femur|Anatomy|false|false||Femoralnull|Foreskin of penis|Anatomy|false|false|C1533810;C1882509;C1552823;C1704765|sheathnull|Condoms, Male|Device|false|false||sheathnull|Place - dosing instruction imperative|Finding|false|false|C0816951;C4266533;C0018246;C0227952|placenull|null|Procedure|false|false|C0816951;C4266533;C0018246;C0227952|placenull|put - instruction imperative|Event|false|false|C0816951;C4266533;C0018246;C0227952|placenull|Place|Modifier|false|false||placenull|Table Cell Horizontal Align - right|Finding|false|false|C0816951;C4266533;C0018246;C0227952|rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Pelvis>Groin|Anatomy|false|false|C1882509;C1533810;C1552823;C1704765|groin
null|Inguinal region|Anatomy|false|false|C1882509;C1533810;C1552823;C1704765|groin
null|Inguinal part of abdomen|Anatomy|false|false|C1882509;C1533810;C1552823;C1704765|groinnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false|C1123023;C4520765|SKIN
null|Skin and subcutaneous tissue disorders|Disorder|false|false|C1123023;C4520765|SKINnull|Skin Specimen Source Code|Finding|false|false|C1123023;C4520765|SKIN
null|Skin Specimen|Finding|false|false|C1123023;C4520765|SKINnull|Skin, Human|Anatomy|false|false|C1546781;C0444099;C0178298;C0496955|SKIN
null|Skin|Anatomy|false|false|C1546781;C0444099;C0178298;C0496955|SKINnull|Stasis dermatitis|Disorder|true|false||stasis dermatitisnull|Stasis|Finding|false|false||stasisnull|Dermatitis|Disorder|true|false||dermatitisnull|Ulcer|Finding|true|false||ulcersnull|Scar Tissue|Finding|true|false||scars
null|Cicatrix|Finding|true|false||scarsnull|Xanthoma|Disorder|true|false||xanthomasnull|null|Drug|false|false||PULSESnull|Physiologic pulse|Finding|false|false||PULSESnull|Pulse taking|Procedure|false|false||PULSESnull|Table Cell Horizontal Align - right|Finding|false|false||Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|Carotid Arteries|Anatomy|false|false||Carotidnull|Table Cell Horizontal Align - left|Finding|false|false||Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|Carotid Arteries|Anatomy|false|false||Carotidnull|Electrocardiogram image|Finding|false|false||EKG
null|Electrocardiogram|Finding|false|false||EKGnull|Electrocardiography|Procedure|false|false||EKGnull|New LBBB|Finding|false|false||new LBBBnull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|Left Bundle-Branch Block|Disorder|false|false||LBBBnull|null|Lab|false|false||LBBBnull|SULT1E1 wt Allele|Finding|false|false||STE
null|SULT1E1 gene|Finding|false|false||STEnull|Lead Device|Device|false|false||leadsnull|Telemetry|Procedure|false|false||TELEMETRYnull|null|Finding|false|false||NSR
null|Neutral Sidebent Rotated|Finding|false|false||NSRnull|Echocardiography|Procedure|false|false||ECHOCARDIOGRAMnull|Pending - Allergy Clinical Status|Finding|false|false||pending
null|Pending - referral status|Finding|false|false||pendingnull|Pending - status|Time|false|false||pendingnull|pending - ManagedParticipationStatus|Modifier|false|false||pending
null|pending - RoleStatus|Modifier|false|false||pending
null|Pending - Day type|Modifier|false|false||pendingnull|Trophoblastic tumor, epithelioid|Disorder|false|false||ETTnull|Cardiac Catheterization Procedures|Procedure|false|false|C0018787|CARDIAC CATHnull|Cardiac attachment|Finding|false|false|C0018787|CARDIACnull|Heart|Anatomy|false|false|C1314974;C0018795;C0007430|CARDIACnull|Cardiac - anatomy qualifier|Modifier|false|false||CARDIACnull|Catheterization|Procedure|false|false|C0018787|CATHnull|levomefolate calcium|Drug|false|false||LMCA
null|levomefolate calcium|Drug|false|false||LMCA
null|levomefolate calcium|Drug|false|false||LMCAnull|Distal Resection Margin|Attribute|false|false||distalnull|Distal (qualifier value)|Modifier|false|false||distalnull|Leukocyte adhesion deficiency type 1|Disorder|false|false|C0226032|LAD
null|Leukocyte adhesion deficiency|Disorder|false|false|C0226032|LADnull|ITGB2 wt Allele|Finding|false|false|C0226032|LAD
null|DLD gene|Finding|false|false|C0226032|LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false|C1414063;C1706333;C5550999;C0398738|LADnull|Ladino Language|Entity|false|false||LADnull|Occluded|Finding|false|false||Occluded
null|Obstruction|Finding|false|false||Occludednull|Difficult (qualifier value)|Finding|false|false||difficultnull|Proximal Resection Margin|Attribute|false|false||proximalnull|Proximal|Modifier|false|false||proximalnull|Leukocyte adhesion deficiency type 1|Disorder|false|false|C0226032|LAD
null|Leukocyte adhesion deficiency|Disorder|false|false|C0226032|LADnull|ITGB2 wt Allele|Finding|false|false|C0226032|LAD
null|DLD gene|Finding|false|false|C0226032|LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false|C1414063;C1706333;C5550999;C0398738|LADnull|Ladino Language|Entity|false|false||LADnull|Distal Resection Margin|Attribute|false|false||Distalnull|Distal (qualifier value)|Modifier|false|false||Distalnull|Leukocyte adhesion deficiency type 1|Disorder|false|false|C0226032|LAD
null|Leukocyte adhesion deficiency|Disorder|false|false|C0226032|LADnull|ITGB2 wt Allele|Finding|false|false|C0226032|LAD
null|DLD gene|Finding|false|false|C0226032|LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false|C5550999;C0398738;C1414063;C1706333|LADnull|Ladino Language|Entity|false|false||LADnull|Diffuse|Modifier|false|false||diffusenull|Diseased|Modifier|false|false||diseasednull|Methylcytosine Dioxygenase TET1|Drug|false|false||LCX
null|Methylcytosine Dioxygenase TET1|Drug|false|false||LCXnull|TET1 wt Allele|Finding|false|false||LCX
null|TET1 gene|Finding|false|false||LCXnull|Occluded|Finding|false|false||occluded
null|Obstruction|Finding|false|false||occludednull|Methylcytosine Dioxygenase TET1|Drug|false|false||LCX
null|Methylcytosine Dioxygenase TET1|Drug|false|false||LCXnull|TET1 wt Allele|Finding|false|false||LCX
null|TET1 gene|Finding|false|false||LCXnull|Occluded|Finding|false|false||Occluded
null|Obstruction|Finding|false|false||Occludednull|BRIEF Health Literacy Screening Tool|Finding|false|false||Brief
null|Behavior Rating Inventory of Executive Function|Finding|false|false||Briefnull|Brief|Time|false|false||Briefnull|Shortened|Modifier|false|false||Briefnull|Hospital course|Finding|false|false||Hospital Coursenull|null|Attribute|false|false||Hospital Coursenull|Organization unit type - Hospital|Finding|false|false||Hospitalnull|Hospitals|Device|false|false||Hospitalnull|Hospitals|Entity|false|false||Hospitalnull|Hospital environment|Modifier|false|false||Hospitalnull|Course|Time|false|false||Coursenull|Females|Subject|false|false||female
null|Woman|Subject|false|false||femalenull|Female, Self-Report|Modifier|false|false||female
null|Female Phenotype|Modifier|false|false||femalenull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|ST segment elevation myocardial infarction|Disorder|false|false||STEMInull|ST Elevation Myocardial Infarction by ECG Finding|Finding|false|false||STEMInull|Catheterization|Procedure|false|false||catheterizationnull|Multiple Pulmonary Nodules|Finding|false|false|C0024109|multiple pulmonary nodulesnull|Numerous|LabModifier|false|false||multiplenull|Multiple Pulmonary Nodules|Finding|false|false|C0024109|pulmonary nodulesnull|Pulmonary (intended site)|Finding|false|false|C0024109|pulmonarynull|Lung|Anatomy|false|false|C2707265;C0748164;C4522268;C0332290;C0332290;C0748164|pulmonarynull|null|Attribute|false|false|C0024109|pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Consistent with|Finding|false|false|C0024109|consistent withnull|Compatible|Modifier|false|false||consistent withnull|Consistent with|Finding|false|false|C0024109|consistentnull|Adenocarcinoma|Disorder|false|false||adenocarcinoma
null|Malignant adenomatous neoplasm|Disorder|false|false||adenocarcinomanull|ST segment elevation myocardial infarction|Disorder|false|false||STEMInull|ST Elevation Myocardial Infarction by ECG Finding|Finding|false|false||STEMInull|Adenohypophyseal Diseases|Disorder|false|false||anteriornull|Anterior|Modifier|false|false||anteriornull|ST segment elevation myocardial infarction|Disorder|false|false||STEMInull|ST Elevation Myocardial Infarction by ECG Finding|Finding|false|false||STEMInull|Risk|Finding|false|false||risknull|Score|Finding|false|false||scorenull|Risk|Finding|false|false||risknull|14 days|Time|false|false||14 daysnull|day|Time|false|false||daysnull|Aspects of mortality statistics|LabModifier|false|false||mortality
null|Mortality Vital Statistics|LabModifier|false|false||mortalitynull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|Recurrent|Time|false|false||recurrent
null|Episodic|Time|false|false||recurrentnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Recurrent|Time|false|false||recurrent
null|Episodic|Time|false|false||recurrentnull|Ischemia|Finding|false|false||ischemianull|Ischemia Procedure|Procedure|false|false||ischemianull|Certification patient type - Urgent|Finding|false|false||urgent
null|Admission Type - Urgent|Finding|false|false||urgent
null|Triage Code - Urgent|Finding|false|false||urgent
null|Visit Priority Code - Urgent|Finding|false|false||urgentnull|Act Priority - urgent|Time|false|false||urgentnull|Urgent|Modifier|false|false||urgentnull|urgent - premium|LabModifier|false|false||urgentnull|null|Procedure|false|false||revascularizationnull|Scalable Vector Graphics|Entity|false|false||SVGnull|Completely - dosing instruction fragment|Finding|false|false||completelynull|Complete|Modifier|false|false||completelynull|Occluded|Finding|false|false||occluded
null|Obstruction|Finding|false|false||occludednull|Burning Mouth Syndrome|Disorder|false|false|C0226032|BMSnull|Proximal Resection Margin|Attribute|false|false||proximalnull|Proximal|Modifier|false|false||proximalnull|Leukocyte adhesion deficiency type 1|Disorder|false|false|C0226032|LAD
null|Leukocyte adhesion deficiency|Disorder|false|false|C0226032|LADnull|ITGB2 wt Allele|Finding|false|false|C0226032|LAD
null|DLD gene|Finding|false|false|C0226032|LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false|C5550999;C0398738;C1414063;C1706333;C0006430|LADnull|Ladino Language|Entity|false|false||LADnull|Timing, LOINC Axis 3|Finding|false|false||timingnull|Timing|Time|false|false||timingnull|Scalable Vector Graphics|Entity|false|false||SVGnull|null|Procedure|false|false||placement
null|Implantation procedure|Procedure|false|false||placement
null|Clinical act of insertion|Procedure|false|false||placementnull|Placement|Modifier|false|false||placementnull|year|Time|false|false||yearsnull|FBXW7 wt Allele|Finding|false|false||ago
null|FBXW7 gene|Finding|false|false||agonull|Leukocyte adhesion deficiency type 1|Disorder|false|false|C0226032|LAD
null|Leukocyte adhesion deficiency|Disorder|false|false|C0226032|LADnull|ITGB2 wt Allele|Finding|false|false|C0226032|LAD
null|DLD gene|Finding|false|false|C0226032|LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false|C5550999;C0398738;C1414063;C1706333|LADnull|Ladino Language|Entity|false|false||LADnull|subscriber - self|Finding|false|false||self
null|Self|Finding|false|false||selfnull|Extended Priority Codes - Routine|Finding|false|false||routine
null|Report priority - Routine|Finding|false|false||routine
null|Admission Type - Routine|Finding|false|false||routine
null|Level of Care - Routine|Finding|false|false||routine
null|Processing priority - Routine|Finding|false|false||routine
null|Referral priority - Routine|Finding|false|false||routinenull|Routine coag|Procedure|false|false||routinenull|Priority - Routine|Time|false|false||routinenull|Routine|Modifier|false|false||routinenull|ACSS2 protein, human|Drug|false|false|C0262187|ACS
null|ACSS2 protein, human|Drug|false|false|C0262187|ACSnull|Acrocallosal Syndrome|Disorder|false|false|C0262187|ACS
null|Acute Chest Syndrome|Disorder|false|false|C0262187|ACSnull|ACS - Activity Card Sort|Finding|false|false|C0262187|ACS
null|American Community Survey|Finding|false|false|C0262187|ACS
null|ACCS gene|Finding|false|false|C0262187|ACS
null|CO-methylating acetyl-CoA synthase activity|Finding|false|false|C0262187|ACS
null|PLA2G15 gene|Finding|false|false|C0262187|ACS
null|ACSS2 wt Allele|Finding|false|false|C0262187|ACS
null|ACSS2 gene|Finding|false|false|C0262187|ACS
null|acetate-CoA ligase activity|Finding|false|false|C0262187|ACSnull|anterior calcarine sulcus (human only)|Anatomy|false|false|C4042561;C0742343;C0796147;C1825842;C5400867;C4318612;C1842089;C1424787;C1150760;C2266615;C5551036|ACSnull|Alternate Care Site|Device|false|false||ACSnull|American College of Surgeons|Entity|false|false||ACS
null|American Cancer Society|Entity|false|false||ACS
null|Alternate Care Site|Entity|false|false||ACSnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|eptifibatide|Drug|false|false||eptifibatide
null|eptifibatide|Drug|false|false||eptifibatidenull|HGS protein, human|Drug|false|false||hrs
null|HGS protein, human|Drug|false|false||hrsnull|Dentatorubral-Pallidoluysian Atrophy|Disorder|false|false||hrsnull|HARS1 wt Allele|Finding|false|false||hrs
null|HARS1 gene|Finding|false|false||hrs
null|HGS wt Allele|Finding|false|false||hrs
null|HGS gene|Finding|false|false||hrs
null|ATN1 wt Allele|Finding|false|false||hrs
null|SRSF5 gene|Finding|false|false||hrsnull|Hour|Time|false|false||hrsnull|Plavix|Drug|false|false||plavix
null|Plavix|Drug|false|false||plavixnull|aspirin|Drug|false|false||aspirin
null|aspirin|Drug|false|false||aspirinnull|metoprolol|Drug|false|false||metoprolol
null|metoprolol|Drug|false|false||metoprololnull|captopril|Drug|false|false||captopril
null|captopril|Drug|false|false||captoprilnull|atorvastatin|Drug|false|false||atorvastatin
null|atorvastatin|Drug|false|false||atorvastatinnull|Cardiac enzymes|Drug|false|false|C0018787|Cardiac enzymes
null|Cardiac enzymes|Drug|false|false|C0018787|Cardiac enzymesnull|Cardiac enzymes/isoenzymes measurement|Procedure|false|false|C0018787|Cardiac enzymesnull|null|Attribute|false|false|C0018787|Cardiac enzymesnull|Cardiac attachment|Finding|false|false|C0018787|Cardiacnull|Heart|Anatomy|false|false|C0014445;C0443763;C0201934;C2926589;C1314974;C3540772;C0014442;C3540048;C3542456;C3540017;C3540790;C3541394|Cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||Cardiacnull|Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM|Drug|false|false|C0018787|enzymes
null|Enzymes, peripheral vasodilators|Drug|false|false|C0018787|enzymes
null|Enzymes, peripheral vasodilators|Drug|false|false|C0018787|enzymes
null|Enzymes, peripheral vasodilators|Drug|false|false|C0018787|enzymes
null|Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM|Drug|false|false|C0018787|enzymes
null|Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM|Drug|false|false|C0018787|enzymes
null|Enzymes, antithrombotic|Drug|false|false|C0018787|enzymes
null|Enzymes, antithrombotic|Drug|false|false|C0018787|enzymes
null|Enzymes, antithrombotic|Drug|false|false|C0018787|enzymes
null|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS|Drug|false|false|C0018787|enzymes
null|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS|Drug|false|false|C0018787|enzymes
null|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS|Drug|false|false|C0018787|enzymes
null|Enzymes, hematological|Drug|false|false|C0018787|enzymes
null|Enzymes, hematological|Drug|false|false|C0018787|enzymes
null|Enzymes, hematological|Drug|false|false|C0018787|enzymes
null|Enzymes|Drug|false|false|C0018787|enzymes
null|Enzymes|Drug|false|false|C0018787|enzymes
null|Enzymes for ALIMENTARY TRACT AND METABOLISM|Drug|false|false|C0018787|enzymes
null|Enzymes for ALIMENTARY TRACT AND METABOLISM|Drug|false|false|C0018787|enzymes
null|Enzymes for ALIMENTARY TRACT AND METABOLISM|Drug|false|false|C0018787|enzymesnull|enzymology|Finding|false|false|C0018787|enzymesnull|Peak level|Modifier|false|false||peaknull|Creatine Kinase MB Isoenzyme|Drug|false|false||CKMB
null|Creatine Kinase MB Isoenzyme|Drug|false|false||CKMBnull|Concern|Finding|false|false||concernnull|Acute heart failure|Disorder|false|false|C4037974;C0018787|acute heart failurenull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Congestive heart failure|Disorder|false|false|C4037974;C0018787|heart failure
null|Heart failure|Disorder|false|false|C4037974;C0018787|heart failurenull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787|heart
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787|heartnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|heartnull|Chest>Heart|Anatomy|false|false|C0795691;C0680095;C0231174;C5200924;C0153957;C0153500;C0018801;C0018802;C0264714;C0184633|heart
null|Heart|Anatomy|false|false|C0795691;C0680095;C0231174;C5200924;C0153957;C0153500;C0018801;C0018802;C0264714;C0184633|heartnull|Failure (biologic function)|Finding|false|false|C4037974;C0018787|failure
null|Failure|Finding|false|false|C4037974;C0018787|failure
null|Personal failure|Finding|false|false|C4037974;C0018787|failurenull|Ischemic|Finding|false|false||ischemicnull|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygennull|Oxygen Therapy Care|Procedure|false|false|C4037974;C0018787|oxygennull|Oxygen Equipment Location|Modifier|false|false||oxygennull|Requirement|Finding|false|false||requirementnull|Radiolucent Lines|Finding|false|false|C1261075|RLLnull|Structure of right lower lobe of lung|Anatomy|false|false|C0032285;C5703311|RLLnull|Pneumonia|Disorder|false|false|C1261075|pneumonianull|Significant|Finding|false|false|C0024109|significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|Pulmonary Edema|Finding|false|false|C0024109|pulmonary edemanull|Pulmonary (intended site)|Finding|false|false|C0024109|pulmonarynull|Lung|Anatomy|false|false|C4522268;C0750502;C0034063;C5575284;C0058928;C0013604;C2707265|pulmonarynull|null|Attribute|false|false|C0024109|pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Edema|Finding|false|false|C0024109|edemanull|null|Attribute|false|false||edemanull|ECHO protocol|Procedure|false|false|C0024109|ECHO
null|Extension for Community Healthcare Outcomes|Procedure|false|false|C0024109|ECHOnull|Echo <Calopterygidae>|Entity|false|false||ECHOnull|Moderate - Severity of Illness Code|Finding|false|false||moderate
null|Moderate|Finding|false|false||moderatenull|Moderate (severity modifier)|Modifier|false|false||moderate
null|Moderate - Allergy Severity|Modifier|false|false||moderate
null|Moderation|Modifier|false|false||moderatenull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|regional|Modifier|false|false||regional
null|Local|Modifier|false|false||regionalnull|Left ventricular systolic dysfunction|Disorder|false|false|C0018827|left ventricular systolic dysfunctionnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Heart Ventricle|Anatomy|false|false|C1277187;C3887505;C0749225|ventricularnull|Ventricular|Modifier|false|false||ventricularnull|Systolic dysfunction|Finding|false|false|C0018827|systolic dysfunctionnull|Systole|Finding|false|false||systolicnull|DYSFUNCTION - SKIN DISORDERS|Disorder|false|false|C0018827|dysfunctionnull|Dysfunction|Finding|false|false||dysfunction
null|physiopathological|Finding|false|false||dysfunction
null|Functional disorder|Finding|false|false||dysfunctionnull|Adenohypophyseal Diseases|Disorder|false|false||anteriornull|Anterior|Modifier|false|false||anteriornull|inferiority|Finding|false|false||inferiornull|Inferior|Modifier|false|false||inferiornull|Inferolateral|Modifier|false|false||inferolateralnull|Hypokinesia|Finding|false|false||hypokinesisnull|Initially|Time|false|false||Initiallynull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Coumadin|Drug|false|false||coumadin
null|Coumadin|Drug|false|false||coumadinnull|Cardiac ventricular thrombosis|Disorder|false|false|C0018827|ventricular thrombusnull|Heart Ventricle|Anatomy|false|false|C0302148;C0087086;C0876993;C0199176|ventricularnull|Ventricular|Modifier|false|false||ventricularnull|Thrombus|Finding|false|false|C0018827|thrombus
null|Blood Clot|Finding|false|false|C0018827|thrombusnull|Thrombus <Thrombidae>|Entity|false|false||thrombusnull|Prophylactic treatment|Procedure|false|false|C0018827|prophylaxisnull|prevention & control|Modifier|false|false||prophylaxisnull|Bleeding risk|Finding|false|false||risk of bleedingnull|Risk|Finding|false|false||risk ofnull|Risk|Finding|false|false||risknull|Hemorrhage|Finding|false|false||bleedingnull|Benefit|LabModifier|false|false||benefitnull|Hypoxia, CTCAE|Finding|false|false||Hypoxia
null|Hypoxia|Finding|false|false||Hypoxianull|Hospitalization|Procedure|false|false||hospitalizationnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Saturated|Phenomenon|false|false||saturationsnull|IPSS-R Risk Category Low|Finding|false|false||low
null|IPSS Risk Category Low|Finding|false|false||low
null|low confidentiality|Finding|false|false||lownull|Low - MessageWaitingPriority|Modifier|false|false||low
null|low|Modifier|false|false||low
null|low exposure|Modifier|false|false||lownull|null|LabModifier|false|false||lownull|BaseLine dental cement|Drug|false|false||baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|Plain chest X-ray|Procedure|false|false||CXRnull|Radiolucent Lines|Finding|false|false|C1261075|RLLnull|Structure of right lower lobe of lung|Anatomy|false|false|C5703311;C0032285|RLLnull|Pneumonia|Disorder|false|false|C1261075|pneumonianull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|ceftriaxone|Drug|false|false||ceftriaxone
null|ceftriaxone|Drug|false|false||ceftriaxonenull|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED|Drug|false|false||azithromycin
null|azithromycin|Drug|false|false||azithromycin
null|azithromycin|Drug|false|false||azithromycinnull|metronidazole|Drug|false|false||metronidazole
null|metronidazole|Drug|false|false||metronidazolenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Recurrent|Time|false|false||recurrent
null|Episodic|Time|false|false||recurrentnull|Radiolucent Lines|Finding|false|false|C1261075|RLLnull|Structure of right lower lobe of lung|Anatomy|false|false|C5703311;C0032285|RLLnull|Pneumonia|Disorder|false|false|C1261075|pneumonianull|X-Ray Computed Tomography|Procedure|false|false||CT scannull|Radionuclide Imaging|Procedure|false|false||scan
null|Scanning|Procedure|false|false||scannull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Structure of right lower lobe of lung|Anatomy|false|false|C1552823;C3539671;C1428707;C0521530|right lower lobenull|Table Cell Horizontal Align - right|Finding|false|false|C0225758;C1261075|rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Structure of lower lobe of lung|Anatomy|false|false|C1552823;C3539671;C1428707;C0521530|lower lobenull|Body Site Modifier - Lower|Anatomy|false|false|C2003888;C3539671;C1428707|lowernull|Lower (action)|Event|false|false|C1548802|lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|AKT1S1 wt Allele|Finding|false|false|C0225758;C0796494;C1261075;C1548802|lobe
null|AKT1S1 gene|Finding|false|false|C0225758;C0796494;C1261075;C1548802|lobenull|lobe|Anatomy|false|false|C0521530;C3539671;C1428707|lobenull|Lung consolidation|Disorder|false|false|C0796494;C1261075;C0225758|consolidationnull|Consolidation|Modifier|false|false||consolidationnull|Extensive|Modifier|false|false||extensivenull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|Diffuse|Modifier|false|false||diffusenull|null|Finding|false|false|C4037972;C0024109|lung nodulesnull|Lung diseases|Disorder|false|false|C4037972;C0024109|lungnull|Lung Problem|Finding|false|false|C4037972;C0024109|lungnull|Chest>Lung|Anatomy|false|false|C0034079;C0024115;C0740941|lung
null|Lung|Anatomy|false|false|C0034079;C0024115;C0740941|lungnull|Abnormality detected in sputum by cytology|Lab|false|false||sputum cytology positivenull|Sputum cytology (finding)|Finding|false|false||sputum cytologynull|Sputum Cytology Screening|Procedure|false|false||sputum cytologynull|Specimen Type - Sputum|Finding|false|false||sputum
null|null|Finding|false|false||sputum
null|Sputum|Finding|false|false||sputumnull|Cytology--Technique|Procedure|false|false||cytology
null|Cytological Techniques|Procedure|false|false||cytologynull|Cytology|Title|false|false||cytologynull|cellular aspects|Modifier|false|false||cytologynull|Positive|Finding|false|false||positive fornull|BRAF Gene Rearrangement|Disorder|false|false||positivenull|Rh Positive Blood Group|Finding|false|false||positive
null|Positive Finding|Finding|false|false||positive
null|Positive|Finding|false|false||positivenull|Positive Charge|Modifier|false|false||positivenull|Positive Number|LabModifier|false|false||positivenull|Adenocarcinoma|Disorder|false|false||adenocarcinoma
null|Malignant adenomatous neoplasm|Disorder|false|false||adenocarcinomanull|Hypoxia, CTCAE|Finding|false|false||Hypoxia
null|Hypoxia|Finding|false|false||Hypoxianull|Initially|Time|false|false||initiallynull|combination - answer to question|Finding|false|false||combinationnull|combination of objects|Entity|false|false||combinationnull|Combined|Modifier|false|false||combinationnull|Postobstructive pneumonia|Disorder|false|false||postobstructive pneumonianull|Pneumonia|Disorder|false|false||pneumonianull|Tumor Burden|Procedure|false|false||tumor burdennull|Neoplasms|Disorder|false|false||tumornull|Tumor Mass|Finding|false|false||tumor
null|null|Finding|false|false||tumornull|Burden|Finding|false|false||burdennull|Adenocarcinoma|Disorder|false|false||adenocarcinoma
null|Malignant adenomatous neoplasm|Disorder|false|false||adenocarcinomanull|Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE|Drug|false|false||Antibiotics
null|Antibiotics|Drug|false|false||Antibiotics
null|Antibiotics, ophthalmologic|Drug|false|false||Antibiotics
null|Antibiotics, Gynecological|Drug|false|false||Antibiotics
null|antibiotics, intestinal|Drug|false|false||Antibiotics
null|Antibiotic throat preparations|Drug|false|false||Antibiotics
null|Antibiotics, Antitubercular|Drug|false|false||Antibiotics
null|Antibiotics for systemic use|Drug|false|false||Antibiotics
null|Antifungal Antibiotics, Topical|Drug|false|false||Antibioticsnull|vancomycin|Drug|false|false||vancomycin
null|vancomycin|Drug|false|false||vancomycinnull|Vancomycin measurement|Procedure|false|false||vancomycinnull|levofloxacin|Drug|false|false||levofloxacin
null|levofloxacin|Drug|false|false||levofloxacinnull|Flagyl|Drug|false|false||flagyl
null|Flagyl|Drug|false|false||flagylnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Course|Time|false|false||coursenull|X-Ray Computed Tomography|Procedure|false|false||CT scannull|Radionuclide Imaging|Procedure|false|false||scan
null|Scanning|Procedure|false|false||scannull|Little's Disease|Disorder|false|false||littlenull|Only a Little|Finding|false|false||littlenull|Smallest|LabModifier|false|false||little
null|Small|LabModifier|false|false||littlenull|Parameterized Data Type - Interval|Finding|false|false|C1548802|intervalnull|Interval|Time|false|false||intervalnull|Improvement|Finding|false|false||improvementnull|Table Cell Horizontal Align - right|Finding|false|false|C1548802|rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Body Site Modifier - Lower|Anatomy|false|false|C2003888;C1552823;C1552654|lowernull|Lower (action)|Event|false|false|C1548802|lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|AKT1S1 wt Allele|Finding|false|false|C0796494|lobe
null|AKT1S1 gene|Finding|false|false|C0796494|lobenull|lobe|Anatomy|false|false|C0332448;C1549537;C1546677;C3539671;C1428707|lobenull|Administration Method - Infiltrate|Finding|false|false|C0796494|infiltrate
null|null|Finding|false|false|C0796494|infiltrate
null|Infiltration|Finding|false|false|C0796494|infiltratenull|Respiratory Status|Finding|false|false||Respiratory statusnull|null|Attribute|false|false||Respiratory statusnull|Respiratory attachment|Finding|false|false||Respiratory
null|respiratory|Finding|false|false||Respiratory
null|null|Finding|false|false||Respiratory
null|Respiratory specimen|Finding|false|false||Respiratorynull|Respiratory rate|Attribute|false|false||Respiratorynull|What subject filter - Status|Finding|false|false||statusnull|null|Attribute|false|false||statusnull|Social status|Modifier|false|false||status
null|Status|Modifier|false|false||statusnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Message Waiting Priority - High|Finding|false|false||high
null|high - ActExposureLevelCode|Finding|false|false||high
null|IPSS Risk Category High|Finding|false|false||high
null|IPSS-R Risk Category High|Finding|false|false||high
null|High (finding)|Finding|false|false||highnull|Observation Value - High|Modifier|false|false||high
null|High|Modifier|false|false||high
null|Abnormally high|Modifier|false|false||highnull|Flow|Phenomenon|false|false||flownull|Message Waiting Priority - High|Finding|false|false||high
null|high - ActExposureLevelCode|Finding|false|false||high
null|IPSS Risk Category High|Finding|false|false||high
null|IPSS-R Risk Category High|Finding|false|false||high
null|High (finding)|Finding|false|false||highnull|Observation Value - High|Modifier|false|false||high
null|High|Modifier|false|false||high
null|Abnormally high|Modifier|false|false||highnull|Activity (animal life circumstance)|Finding|false|false||activity
null|Physical activity|Finding|false|false||activitynull|Activities|Event|false|false||activitynull|null|Modifier|false|false||activitynull|null|Time|false|false||Prior tonull|null|Time|false|false||Priornull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Requirement|Finding|false|false||requirementnull|Oxygen nasal cannula|Device|false|false||nasal cannula
null|Nasal Cannula|Device|false|false||nasal cannulanull|Nasal brand of oxymetazoline|Drug|false|false|C1550232;C0028429|nasal
null|Nasal brand of oxymetazoline|Drug|false|false|C1550232;C0028429|nasal
null|Nasal dosage form|Drug|false|false|C1550232;C0028429|nasalnull|Nasal Route of Administration|Finding|false|false|C0028429;C1550232|nasal
null|Nasal (intended site)|Finding|false|false|C0028429;C1550232|nasalnull|null|Anatomy|false|false|C4520890;C1522019;C1550622;C1546577;C1272939;C0721966|nasalnull|Specimen Type - Cannula|Finding|false|false|C0028429;C1550232|cannula
null|null|Finding|false|false|C0028429;C1550232|cannulanull|Body Parts - Cannula|Anatomy|false|false|C1272939;C0721966;C4520890;C1522019;C1550622;C1546577|cannulanull|Cannula device|Device|false|false||cannulanull|Calamus <grasshoppers>|Entity|false|false||cannulanull|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygennull|Oxygen Therapy Care|Procedure|false|false||oxygennull|Oxygen Equipment Location|Modifier|false|false||oxygennull|Saturated|Phenomenon|false|false||saturationnull|IPSS-R Risk Category Low|Finding|false|false||low
null|IPSS Risk Category Low|Finding|false|false||low
null|low confidentiality|Finding|false|false||lownull|Low - MessageWaitingPriority|Modifier|false|false||low
null|low|Modifier|false|false||low
null|low exposure|Modifier|false|false||lownull|null|LabModifier|false|false||lownull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|masked - No information|Finding|false|false||mask
null|ANKHD1 gene|Finding|false|false||mask
null|STK26 gene|Finding|false|false||masknull|Protective Face Mask|Device|false|false||mask
null|Masks|Device|false|false||masknull|Helping Behavior|Finding|false|false||assistnull|Assisting (procedure)|Procedure|false|false||assistnull|American Stop Smoking Intervention for Cancer Prevention|Entity|false|false||assistnull|Assisted (qualifier value)|Modifier|false|false||assistnull|Alveolar ventilation function|Finding|false|false||oxygenation
null|Cell Respiration|Finding|false|false||oxygenationnull|null|Finding|false|false|C4037972;C0024109|Lung nodulesnull|Lung diseases|Disorder|false|false|C4037972;C0024109|Lungnull|Lung Problem|Finding|false|false|C4037972;C0024109|Lungnull|Chest>Lung|Anatomy|false|false|C0007097;C0740941;C0024115;C0034079|Lung
null|Lung|Anatomy|false|false|C0007097;C0740941;C0024115;C0034079|Lungnull|Carcinoma|Disorder|false|false|C4037972;C0024109|carcinomanull|X-Ray Computed Tomography|Procedure|false|false||CT scannull|Radionuclide Imaging|Procedure|false|false||scan
null|Scanning|Procedure|false|false||scannull|Diffuse|Modifier|false|false||diffusenull|Multiple Pulmonary Nodules|Finding|false|false|C0024109|pulmonary nodulesnull|Pulmonary (intended site)|Finding|false|false|C0024109|pulmonarynull|Lung|Anatomy|false|false|C4522268;C1521752;C0748164;C2707265;C0038056;C1576419;C1546789;C1305671;C0010818;C0551076|pulmonarynull|null|Attribute|false|false|C0024109|pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Abnormality detected in sputum by cytology|Lab|false|false||sputum cytology positivenull|Sputum cytology (finding)|Finding|false|false|C0024109|sputum cytologynull|Sputum Cytology Screening|Procedure|false|false|C0024109|sputum cytologynull|Specimen Type - Sputum|Finding|false|false|C0024109|sputum
null|null|Finding|false|false|C0024109|sputum
null|Sputum|Finding|false|false|C0024109|sputumnull|Cytology--Technique|Procedure|false|false|C0024109|cytology
null|Cytological Techniques|Procedure|false|false|C0024109|cytologynull|Cytology|Title|false|false||cytologynull|cellular aspects|Modifier|false|false||cytologynull|Positive|Finding|false|false||positive fornull|BRAF Gene Rearrangement|Disorder|false|false||positivenull|Rh Positive Blood Group|Finding|false|false||positive
null|Positive Finding|Finding|false|false||positive
null|Positive|Finding|false|false||positivenull|Positive Charge|Modifier|false|false||positivenull|Positive Number|LabModifier|false|false||positivenull|Adenocarcinoma|Disorder|false|false||adenocarcinoma
null|Malignant adenomatous neoplasm|Disorder|false|false||adenocarcinomanull|Science of Etiology|Finding|false|false||Etiology
null|Etiology aspects|Finding|false|false||Etiology
null|Etiology|Finding|false|false||Etiologynull|True primary (qualifier value)|Time|false|false||primarynull|Primary|Modifier|false|false||primarynull|metastatic qualifier|Finding|false|false||metastatic
null|Metastatic to|Finding|false|false||metastaticnull|THYROID DIAGNOSTIC RADIOPHARMACEUTICALS|Drug|false|false|C0040132|thyroid
null|THYROID|Drug|false|false|C0040132|thyroid
null|THYROID|Drug|false|false|C0040132|thyroid
null|thyroid (USP)|Drug|false|false|C0040132|thyroid
null|thyroid (USP)|Drug|false|false|C0040132|thyroid
null|thyroid (USP)|Drug|false|false|C0040132|thyroidnull|Thyroid Diseases|Disorder|false|false|C0040132|thyroidnull|examination of thyroid|Procedure|false|false|C0040132|thyroidnull|Thyroid Gland|Anatomy|false|false|C3540038;C0040134;C5781115;C0040128;C2228489|thyroidnull|null|Time|false|false||priornull|Possible|Finding|false|false||possiblenull|Possible diagnosis|Modifier|false|false||possible
null|Possibly Related to Intervention|Modifier|false|false||possiblenull|Carcinoma|Disorder|false|false||carcinomanull|Extended Priority Codes - Routine|Finding|false|false||routine
null|Report priority - Routine|Finding|false|false||routine
null|Admission Type - Routine|Finding|false|false||routine
null|Level of Care - Routine|Finding|false|false||routine
null|Processing priority - Routine|Finding|false|false||routine
null|Referral priority - Routine|Finding|false|false||routinenull|Routine coag|Procedure|false|false||routinenull|Priority - Routine|Time|false|false||routinenull|Routine|Modifier|false|false||routinenull|Screening for cancer|Procedure|false|false||cancer screeningnull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Screening - procedure intent|Finding|false|false||screening
null|Special screening finding|Finding|false|false||screening
null|Aspects of disease screening|Finding|false|false||screeningnull|Screening for cancer|Procedure|false|false||screening
null|Disease Screening|Procedure|false|false||screening
null|research subject screening|Procedure|false|false||screening
null|Screening|Procedure|false|false||screening
null|Screening procedure|Procedure|false|false||screeningnull|Tissue diagnosis|Finding|false|false|C0040300|tissue diagnosisnull|Tissue Specimen Code|Finding|false|false|C0040300|tissuenull|Body tissue|Anatomy|false|false|C1546899;C1704338;C1547928;C1546905;C0011900|tissuenull|Diagnosis Classification - Diagnosis|Finding|false|false|C0040300|diagnosis
null|diagnosis aspects|Finding|false|false|C0040300|diagnosisnull|Diagnosis|Procedure|false|false|C0040300|diagnosisnull|null|Attribute|false|false||diagnosisnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Message Waiting Priority - High|Finding|false|false||high
null|high - ActExposureLevelCode|Finding|false|false||high
null|IPSS Risk Category High|Finding|false|false||high
null|IPSS-R Risk Category High|Finding|false|false||high
null|High (finding)|Finding|false|false||highnull|Observation Value - High|Modifier|false|false||high
null|High|Modifier|false|false||high
null|Abnormally high|Modifier|false|false||highnull|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygennull|Oxygen Therapy Care|Procedure|false|false||oxygennull|Oxygen Equipment Location|Modifier|false|false||oxygennull|Requirement|Finding|false|false||requirementnull|ANTICOAGULATION (finding)|Finding|false|false||anticoagulation
null|Anticoagulation function|Finding|false|false||anticoagulation
null|Decreased Coagulation Activity [PE]|Finding|false|false||anticoagulationnull|Anticoagulation Therapy|Procedure|false|false||anticoagulationnull|Plavix|Drug|false|false||plavix
null|Plavix|Drug|false|false||plavixnull|Arylsulfatase A, human|Drug|false|false||asa
null|Arylsulfatase A, human|Drug|false|false||asa
null|aspirin|Drug|false|false||asa
null|aspirin|Drug|false|false||asanull|ARSA gene|Finding|false|false||asanull|contextual factors|Finding|false|false||settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|Recent|Time|false|false||recentnull|Clinical act of insertion|Procedure|false|false||placement
null|Implantation procedure|Procedure|false|false||placement
null|null|Procedure|false|false||placementnull|Placement|Modifier|false|false||placementnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Imaging problem|Finding|false|false|C0018670;C0152336|imagingnull|Diagnostic Imaging|Procedure|false|false|C0018670;C0152336|imaging
null|Imaging Techniques|Procedure|false|false|C0018670;C0152336|imagingnull|Imaging Technology|Title|false|false||imagingnull|Problems with head|Disorder|false|false|C0018670;C0152336|headnull|Procedure on head|Procedure|false|false|C0018670;C0152336|headnull|Structure of head of caudate nucleus|Anatomy|false|false|C0876917;C0740845;C0079595;C0011923;C0362076;C0332305|head
null|Head|Anatomy|false|false|C0876917;C0740845;C0079595;C0011923;C0362076;C0332305|headnull|Head Device|Device|false|false||headnull|With staging|Finding|false|false|C0018670;C0152336|stagingnull|Venezuelan equine encephalitis virus subtype IIIA|Disorder|false|false||IIIanull|Multiple Pulmonary Nodules|Finding|false|false|C0024109|pulmonary nodulesnull|Pulmonary (intended site)|Finding|false|false|C0024109|pulmonarynull|Lung|Anatomy|false|false|C2707265;C4522268;C0748164|pulmonarynull|null|Attribute|false|false|C0024109|pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Lung diseases|Disorder|false|false|C4037972;C0024109|lungnull|Lung Problem|Finding|false|false|C4037972;C0024109|lungnull|Chest>Lung|Anatomy|false|false|C0024115;C0740941|lung
null|Lung|Anatomy|false|false|C0024115;C0740941|lungnull|Obvious|Modifier|false|false||obviousnull|Distal Resection Margin|Attribute|false|false||distalnull|Distal (qualifier value)|Modifier|false|false||distalnull|Leukocyte adhesion deficiency type 1|Disorder|true|false|C0226032|LAD
null|Leukocyte adhesion deficiency|Disorder|true|false|C0226032|LADnull|ITGB2 wt Allele|Finding|true|false|C0226032|LAD
null|DLD gene|Finding|true|false|C0226032|LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false|C0027627;C2939419;C1414063;C1706333;C1513183;C4255448;C5550999;C0398738|LADnull|Ladino Language|Entity|true|false||LADnull|Neoplasm Metastasis|Disorder|false|false|C0226032|metastasis
null|Metastatic malignant neoplasm|Disorder|false|false|C0226032|metastasisnull|Metastasis|Finding|false|false|C0226032|metastasis
null|Metastatic Lesion|Finding|false|false|C0226032|metastasisnull|Empiric|Modifier|false|false||Empiricnull|Therapy Object (animal model)|Finding|false|false||therapy
null|therapeutic aspects|Finding|false|false||therapynull|Therapeutic procedure|Procedure|false|false||therapynull|Marital Status - Single|Finding|false|false||single
null|Unmarried|Finding|false|false||singlenull|Singular|LabModifier|false|false||singlenull|Agent|Drug|false|false||agent
null|Pharmacologic Substance|Drug|false|false||agentnull|GDC Therapeutic Agent Terminology|Finding|false|false||agent
null|agent - RoleClass|Finding|false|false||agent
null|Protocol Agent|Finding|false|false||agentnull|pharmacotherapeutic|Finding|false|false||chemotherapynull|Chemotherapy Regimen|Procedure|false|false||chemotherapy
null|Pharmacotherapy|Procedure|false|false||chemotherapy
null|Chemotherapy|Procedure|false|false||chemotherapynull|pemetrexed|Drug|false|false||Pemetrexed
null|pemetrexed|Drug|false|false||Pemetrexednull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|dexamethasone|Drug|false|false||dexamethasone
null|dexamethasone|Drug|false|false||dexamethasonenull|Eruption of skin (disorder)|Disorder|false|false||rashnull|Skin rash|Finding|false|false||rash
null|Eruptions|Finding|false|false||rash
null|Exanthema|Finding|false|false||rashnull|Chronic Kidney Insufficiency|Disorder|false|false|C0022646|Chronic renal insufficiencynull|Chronic - Admission Level of Care Code|Finding|false|false||Chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||Chronicnull|chronic|Time|false|false||Chronicnull|Renal Insufficiency|Disorder|false|false|C0022646|renal insufficiency
null|Kidney Failure|Disorder|false|false|C0022646|renal insufficiencynull|Urologic Diseases|Disorder|false|false|C0022646|renalnull|Kidney|Anatomy|false|false|C0042075;C0403447;C0035078;C1565489;C0231179|renalnull|Insufficiency|Finding|false|false|C0022646|insufficiencynull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|With glomerular filtration rate|Modifier|false|false||with GFRnull|RAPGEF5 gene|Finding|false|false||GFRnull|Glomerular Filtration Rate|LabModifier|false|false||GFRnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|Renal function|Finding|false|false|C0022646|renal functionnull|Kidney Function Tests|Procedure|false|false|C0022646|renal functionnull|Urologic Diseases|Disorder|false|false|C0022646|renalnull|Kidney|Anatomy|false|false|C0042075;C0232804;C0022662|renalnull|Function (attribute)|Finding|false|false||function
null|physiological aspects|Finding|false|false||function
null|Mathematical Operator|Finding|false|false||function
null|Functional Status|Finding|false|false||functionnull|Function Axis|Subject|false|false||functionnull|Mucomyst|Drug|false|false||mucomyst
null|Mucomyst|Drug|false|false||mucomystnull|null|Time|false|false||priornull|IV contrast|Drug|false|false||IV contrastnull|Contrast Media|Drug|false|false||contrastnull|Contrast|Modifier|false|false||contrastnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|creatinine|Drug|false|false||Creatinine
null|creatinine|Drug|false|false||Creatininenull|Creatinine metabolic function|Finding|false|false||Creatininenull|Creatinine measurement|Procedure|false|false||Creatininenull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Hyperkalemia|Finding|false|false||Hyperkalemia
null|Serum potassium level above reference range|Finding|false|false||Hyperkalemianull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|MILDLY|Modifier|false|false||mildly
null|Mild (qualifier value)|Modifier|false|false||mildlynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|null|Time|false|false||prior tonull|null|Time|false|false||priornull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Electrocardiogram image|Finding|false|false||EKG
null|Electrocardiogram|Finding|false|false||EKGnull|Electrocardiography|Procedure|false|false||EKGnull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|Kayexalate|Drug|false|false||kayexalate
null|Kayexalate|Drug|false|false||kayexalatenull|Electrolytes|Drug|false|false||Electrolytes
null|Electrolytes|Drug|false|false||Electrolytes
null|Electrolyte [EPC]|Drug|false|false||Electrolytesnull|Daily|Time|false|false||dailynull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Hypertensive disease|Disorder|false|false||HTNnull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|clopidogrel|Drug|false|false||Clopidogrel
null|clopidogrel|Drug|false|false||Clopidogrelnull|Plavix|Drug|false|false||Plavix
null|Plavix|Drug|false|false||Plavixnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Daily|Time|false|false||Dailynull|ezetimibe / simvastatin|Drug|false|false||Ezetimibe-Simvastatinnull|ezetimibe|Drug|false|false||Ezetimibe
null|ezetimibe|Drug|false|false||Ezetimibenull|simvastatin|Drug|false|false||Simvastatin
null|simvastatin|Drug|false|false||Simvastatinnull|Vytorin|Drug|false|false||Vytorin
null|Vytorin|Drug|false|false||Vytorinnull|Daily|Time|false|false||dailynull|nifedipine|Drug|false|false||Nifedipine
null|nifedipine|Drug|false|false||Nifedipinenull|nitroglycerin|Drug|false|false||Nitroglycerin
null|nitroglycerin|Drug|false|false||Nitroglycerinnull|/hour|Time|false|false||/hournull|Hour|Time|false|false||hournull|Patch - Extended Release Film|Drug|false|false||Patch
null|Human patch material|Drug|false|false||Patch
null|Body tissue patch material|Drug|false|false||Patchnull|Plaque (lesion)|Finding|false|false||Patchnull|Patch Dosage Form|Device|false|false||Patch
null|Surgical patch|Device|false|false||Patchnull|Patch (unit of presentation)|LabModifier|false|false||Patch
null|Patch Dosing Unit|LabModifier|false|false||Patchnull|Patch - Extended Release Film|Drug|false|false||patch
null|Human patch material|Drug|false|false||patch
null|Body tissue patch material|Drug|false|false||patchnull|Plaque (lesion)|Finding|false|false||patchnull|Patch Dosage Form|Device|false|false||patch
null|Surgical patch|Device|false|false||patchnull|Patch (unit of presentation)|LabModifier|false|false||patch
null|Patch Dosing Unit|LabModifier|false|false||patchnull|Once A Day|Drug|false|false||once a daynull|Once daily|Time|false|false||once a daynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Sublingual Route of Administration|Finding|false|false||sublingual
null|Sublingual (intended site)|Finding|false|false||sublingualnull|Sublingual location|Modifier|false|false||sublingualnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Recent|Time|false|false||recentlynull|null|Time|false|false||priornull|propranolol|Drug|false|false||Propranolol
null|propranolol|Drug|false|false||Propranololnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Once A Day|Drug|false|false||once a daynull|Once daily|Time|false|false||once a daynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Multivitamin preparation|Drug|false|false||Multivitamin
null|Multivitamin preparation|Drug|false|false||Multivitamin
null|Multivitamin preparation|Drug|false|false||Multivitaminnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|long-term care|Procedure|false|false||Extended Carenull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|In care (finding)|Finding|false|false||Care
null|Continuity Assessment Record and Evaluation|Finding|false|false||Carenull|care activity|Event|false|false||Carenull|ADMIN.FACILITY|Finding|false|false||Facilitynull|Facility (object)|Device|false|false||Facilitynull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|True primary (qualifier value)|Time|false|false||Primarynull|Primary|Modifier|false|false||Primarynull|ST segment elevation myocardial infarction|Disorder|false|false|C0027061|ST elevation myocardial infarctionnull|ST segment elevation (finding)|Finding|false|false|C0027061|ST elevationnull|Elevation procedure|Procedure|false|false|C0027061|elevationnull|Elevation|Modifier|false|false||elevationnull|Myocardial Infarction|Disorder|false|false|C0027061|myocardial infarctionnull|null|Attribute|false|false|C0027061|myocardial infarctionnull|Myocardium|Anatomy|false|false|C0021308;C2926063;C1536220;C0520886;C0439775;C0027051|myocardialnull|Myocardial|Modifier|false|false||myocardialnull|Infarction|Finding|false|false|C0027061|infarctionnull|Carcinoma|Disorder|false|false||carcinomanull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Disease|Disorder|false|false||Conditionnull|Logical Condition|Finding|false|false||Conditionnull|null|Attribute|false|false||Conditionnull|Condition|Modifier|false|false||Conditionnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygennull|Oxygen Therapy Care|Procedure|false|false||oxygennull|Oxygen Equipment Location|Modifier|false|false||oxygennull|Requirement|Finding|false|false||requirementnull|SAT1 protein, human|Drug|false|false||Sat
null|SAT1 protein, human|Drug|false|false||Satnull|College Entrance Examination Board Scholastic Aptitude Test|Finding|false|false||Sat
null|SAT1 wt Allele|Finding|false|false||Sat
null|SAT1 gene|Finding|false|false||Satnull|Santali language|Entity|false|false||Satnull|IPSS-R Risk Category Low|Finding|false|false||low
null|IPSS Risk Category Low|Finding|false|false||low
null|low confidentiality|Finding|false|false||lownull|Low - MessageWaitingPriority|Modifier|false|false||low
null|low|Modifier|false|false||low
null|low exposure|Modifier|false|false||lownull|null|LabModifier|false|false||lownull|Discharge instructions|Finding|false|false||Discharge Instructionsnull|hospital discharge instructions (treatment)|Procedure|false|false||Discharge Instructionsnull|null|Attribute|false|false||Discharge Instructionsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructionsnull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Chest pressure|Finding|false|false|C1527391;C0817096|chest pressurenull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0438716;C0741025|chest
null|Anterior thoracic region|Anatomy|false|false|C0438716;C0741025|chestnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|Present|Finding|false|false||foundnull|Myocardial Infarction|Disorder|false|false|C4037974;C0018787|heart attacknull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787|heart
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787|heartnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|heartnull|Chest>Heart|Anatomy|false|false|C0027051;C0153957;C0153500;C0795691;C1304680;C1261512|heart
null|Heart|Anatomy|false|false|C0027051;C0153957;C0153500;C0795691;C1304680;C1261512|heartnull|Attack (finding)|Finding|false|false|C4037974;C0018787|attack
null|Attack behavior|Finding|false|false|C4037974;C0018787|attacknull|Attack device|Device|false|false||attacknull|Cardiac catheterisation as the cause of abnormal reaction of the patient, or of later complication, without mention of misadventure at the time of the procedure|Disorder|false|false|C0018787|cardiac catheterizationnull|Diagnostic Service Section ID - Cardiac Catheterization|Finding|false|false|C0018787|cardiac catheterizationnull|Consent Type - Cardiac Catheterization|Procedure|false|false|C0018787|cardiac catheterization
null|Cardiac Catheterization Procedures|Procedure|false|false|C0018787|cardiac catheterizationnull|Cardiac attachment|Finding|false|false|C0018787|cardiacnull|Heart|Anatomy|false|false|C1547981;C1314974;C0018795;C1548828;C0261588|cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||cardiacnull|Catheterization|Procedure|false|false||catheterizationnull|Bare metal stent|Device|false|false||bare metal stentnull|null|Modifier|false|false||barenull|Metal stent|Device|false|false||metal stentnull|Metals|Drug|false|false||metalnull|null|Device|false|false||stentnull|outcomes otolaryngology breathing|Finding|false|false|C0024109|breathing
null|Inspiration (function)|Finding|false|false|C0024109|breathing
null|Respiration|Finding|false|false|C0024109|breathingnull|null|Attribute|false|false|C0024109|breathingnull|respiratory system process|Phenomenon|false|false|C0024109|breathingnull|Radionuclide Imaging|Procedure|false|false|C0024109|scan
null|Scanning|Procedure|false|false|C0024109|scannull|Lung|Anatomy|false|false|C1160636;C2015926;C0004048;C0035203;C5885990;C0034606;C0441633|lungsnull|Sputum specimen|Finding|false|false|C0334227|sputum samplenull|Specimen Type - Sputum|Finding|false|false||sputum
null|null|Finding|false|false||sputum
null|Sputum|Finding|false|false||sputumnull|Specimen|Drug|false|false||samplenull|Nucleotide Sequence Sample Name|Finding|false|false|C0334227|sample
null|Biospecimen|Finding|false|false|C0334227|samplenull|Tumor cells, malignant|Anatomy|false|false|C0444159;C5551027;C2347026|malignant cellsnull|Malignant (qualifier value)|Modifier|false|false||malignantnull|Cells|Anatomy|false|false||cellsnull|Malignant neoplasm of lung|Disorder|false|false|C4037972;C0024109|lung cancer
null|Carcinoma of lung|Disorder|false|false|C4037972;C0024109|lung cancernull|Lung diseases|Disorder|false|false|C4037972;C0024109|lungnull|Lung Problem|Finding|false|false|C4037972;C0024109|lungnull|Chest>Lung|Anatomy|false|false|C0024115;C0740941;C0242379;C0684249|lung
null|Lung|Anatomy|false|false|C0024115;C0740941;C0242379;C0684249|lungnull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|pharmacotherapeutic|Finding|false|false||chemotherapynull|Chemotherapy Regimen|Procedure|false|false||chemotherapy
null|Pharmacotherapy|Procedure|false|false||chemotherapy
null|Chemotherapy|Procedure|false|false||chemotherapynull|Further|Modifier|false|false||furthernull|Biomaterial Treatment|Finding|false|false||treatment
null|Treating|Finding|false|false||treatment
null|therapeutic aspects|Finding|false|false||treatmentnull|treatment - ActInformationManagementReason|Procedure|false|false||treatment
null|Administration (procedure)|Procedure|false|false||treatment
null|Therapeutic procedure|Procedure|false|false||treatmentnull|Every morning|Time|false|false||every morningnull|Morning|Time|false|false||morningnull|infant weight for previous delivery (history)|Finding|false|false||weight
null|Weight symptom (finding)|Finding|false|false||weightnull|Weighing patient|Procedure|false|false||weightnull|null|Attribute|false|false||weightnull|Body Weight|Subject|false|false||weightnull|Importance Weight|Modifier|false|false||weightnull|Weight|LabModifier|false|false||weightnull|More|LabModifier|false|false||morenull|liquid-based cytology (procedure)|Procedure|false|false||lbsnull|Pounds|LabModifier|false|false||lbsnull|Following|Time|false|false||following
null|Status post|Time|false|false||followingnull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Plavix|Drug|false|false||plavix
null|Plavix|Drug|false|false||plavixnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|1 Month|Time|false|false||1 monthnull|Transaction counts and value totals - month|Finding|false|false||month
null|Precision - month|Finding|false|false||monthnull|month|Time|false|false||month
null|Monthly (qualifier value)|Time|false|false||monthnull|Ensure (product)|Drug|false|false||ensurenull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787|heart
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787|heartnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|heartnull|Chest>Heart|Anatomy|false|false|C0795691;C0153957;C0153500|heart
null|Heart|Anatomy|false|false|C0795691;C0153957;C0153500|heartnull|null|Device|false|false||stentnull|Obstruction|Finding|false|false||blocked
null|Blocking|Finding|false|false||blockednull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions