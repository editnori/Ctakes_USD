 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
_|28,29
_|29,30
_|30,31
No|32,34
:|34,35
_|38,39
_|39,40
_|40,41
<EOL>|41,42
<EOL>|43,44
Admission|44,53
Date|54,58
:|58,59
_|61,62
_|62,63
_|63,64
Discharge|78,87
Date|88,92
:|92,93
_|96,97
_|97,98
_|98,99
<EOL>|99,100
<EOL>|101,102
Date|102,106
of|107,109
Birth|110,115
:|115,116
_|118,119
_|119,120
_|120,121
Sex|134,137
:|137,138
M|141,142
<EOL>|142,143
<EOL>|144,145
Service|145,152
:|152,153
MEDICINE|154,162
<EOL>|162,163
<EOL>|164,165
Allergies|165,174
:|174,175
<EOL>|176,177
No|177,179
Known|180,185
Allergies|186,195
/|196,197
Adverse|198,205
Drug|206,210
Reactions|211,220
<EOL>|220,221
<EOL>|222,223
Attending|223,232
:|232,233
_|234,235
_|235,236
_|236,237
.|237,238
<EOL>|238,239
<EOL>|240,241
Chief|241,246
Complaint|247,256
:|256,257
<EOL>|257,258
Lower|258,263
extremity|264,273
swelling|274,282
<EOL>|282,283
<EOL>|284,285
Major|285,290
Surgical|291,299
or|300,302
Invasive|303,311
Procedure|312,321
:|321,322
<EOL>|322,323
None|323,327
<EOL>|327,328
<EOL>|329,330
History|330,337
of|338,340
Present|341,348
Illness|349,356
:|356,357
<EOL>|357,358
_|358,359
_|359,360
_|360,361
with|362,366
AF|367,369
on|370,372
warfarin|373,381
,|381,382
DM|383,385
,|385,386
and|387,390
recent|391,397
steroid|398,405
pulse|406,411
p|412,413
/|413,414
w|414,415
<EOL>|416,417
bilaterally|417,428
swollen|429,436
and|437,440
painful|441,448
ankles|449,455
.|455,456
Pt|457,459
had|460,463
no|464,466
complaints|467,477
in|478,480
<EOL>|481,482
the|482,485
ED|486,488
,|488,489
but|490,493
his|494,497
wife|498,502
was|503,506
concerned|507,516
about|517,522
his|523,526
increasing|527,537
swelling|538,546
<EOL>|547,548
and|548,551
his|552,555
inability|556,565
to|566,568
walk|569,573
without|574,581
pain|582,586
.|586,587
He|588,590
had|591,594
a|595,596
fall|597,601
over|602,606
a|607,608
<EOL>|609,610
bathtub|610,617
one|618,621
week|622,626
ago|627,630
(|631,632
reports|632,639
no|640,642
head|643,647
strike|648,654
)|654,655
.|655,656
He|657,659
was|660,663
at|664,666
a|667,668
<EOL>|669,670
_|670,671
_|671,672
_|672,673
in|674,676
_|677,678
_|678,679
_|679,680
at|681,683
that|684,688
time|689,693
and|694,697
went|698,702
to|703,705
the|706,709
local|710,715
_|716,717
_|717,718
_|718,719
<EOL>|720,721
_|721,722
_|722,723
_|723,724
.|724,725
He|726,728
was|729,732
found|733,738
to|739,741
have|742,746
a|747,748
vertebral|749,758
fracture|759,767
and|768,771
was|772,775
<EOL>|776,777
given|777,782
a|783,784
back|785,789
brace|790,795
,|795,796
which|797,802
he|803,805
has|806,809
been|810,814
wearing|815,822
inconsistently|823,837
.|837,838
<EOL>|840,841
<EOL>|841,842
In|842,844
the|845,848
ED|849,851
,|851,852
exam|853,857
was|858,861
remarkable|862,872
for|873,876
bilateral|877,886
ankle|887,892
swelling|893,901
with|902,906
<EOL>|907,908
3|908,909
+|909,910
pitting|911,918
edema|919,924
,|924,925
cold|926,930
and|931,934
mottled|935,942
toes|943,947
,|947,948
+|949,950
dopplerable|951,962
dorsalis|963,971
<EOL>|972,973
pedis|973,978
pulses|979,985
with|986,990
no|991,993
sensory|994,1001
disturbances|1002,1014
.|1014,1015
BNP|1016,1019
was|1020,1023
elevated|1024,1032
at|1033,1035
<EOL>|1036,1037
6310|1037,1041
.|1041,1042
CXR|1043,1046
showed|1047,1053
pulmonary|1054,1063
edema|1064,1069
.|1069,1070
LENIs|1071,1076
were|1077,1081
negative|1082,1090
for|1091,1094
DVT|1095,1098
.|1098,1099
<EOL>|1100,1101
ED|1101,1103
bedside|1104,1111
US|1112,1114
showed|1115,1121
no|1122,1124
evidence|1125,1133
of|1134,1136
pericardial|1137,1148
effusion|1149,1157
or|1158,1160
IVC|1161,1164
<EOL>|1165,1166
volume|1166,1172
depletion|1173,1182
<EOL>|1184,1185
<EOL>|1185,1186
He|1186,1188
was|1189,1192
given|1193,1198
40mg|1199,1203
IV|1204,1206
Lasix|1207,1212
.|1212,1213
Nursing|1214,1221
in|1222,1224
the|1225,1228
ED|1229,1231
noted|1232,1237
that|1238,1242
pt|1243,1245
able|1246,1250
<EOL>|1251,1252
to|1252,1254
stand|1255,1260
and|1261,1264
weight|1265,1271
bear|1272,1276
but|1277,1280
unsteady|1281,1289
,|1289,1290
fall|1291,1295
risk|1296,1300
.|1300,1301
T|1302,1303
-|1303,1304
spine|1304,1309
film|1310,1314
<EOL>|1315,1316
was|1316,1319
also|1320,1324
done|1325,1329
in|1330,1332
the|1333,1336
ED|1337,1339
and|1340,1343
was|1344,1347
without|1348,1355
fractures|1356,1365
or|1366,1368
<EOL>|1369,1370
dislocations|1370,1382
.|1382,1383
<EOL>|1385,1386
<EOL>|1386,1387
He|1387,1389
triggered|1390,1399
for|1400,1403
hypotension|1404,1415
to|1416,1418
mid|1419,1422
_|1423,1424
_|1424,1425
_|1425,1426
and|1427,1430
bradycardia|1431,1442
to|1443,1445
mid|1446,1449
<EOL>|1450,1451
_|1451,1452
_|1452,1453
_|1453,1454
x|1455,1456
2|1457,1458
,|1458,1459
responded|1460,1469
well|1470,1474
to|1475,1477
250cc|1478,1483
fluid|1484,1489
boluses|1490,1497
.|1497,1498
Vitals|1499,1505
prior|1506,1511
to|1512,1514
<EOL>|1515,1516
transfer|1516,1524
:|1524,1525
T|1526,1527
98.8|1528,1532
,|1532,1533
HR|1534,1536
63|1537,1539
,|1539,1540
RR|1541,1543
15|1544,1546
,|1546,1547
BP|1548,1550
118|1551,1554
/|1554,1555
85|1555,1557
,|1557,1558
02|1559,1561
100|1562,1565
%|1565,1566
on|1567,1569
RA|1570,1572
<EOL>|1574,1575
<EOL>|1575,1576
<EOL>|1577,1578
Past|1578,1582
Medical|1583,1590
History|1591,1598
:|1598,1599
<EOL>|1599,1600
DM|1600,1602
II|1603,1605
,|1605,1606
HTN|1607,1610
,|1610,1611
HL|1612,1614
,|1614,1615
MI|1616,1618
(|1619,1620
in|1620,1622
past|1623,1627
)|1627,1628
,|1628,1629
AF|1630,1632
on|1633,1635
coumadin|1636,1644
,|1644,1645
prostate|1646,1654
CA|1655,1657
<EOL>|1658,1659
treated|1659,1666
non-operatively|1667,1682
<EOL>|1682,1683
<EOL>|1683,1684
<EOL>|1685,1686
Social|1686,1692
History|1693,1700
:|1700,1701
<EOL>|1701,1702
_|1702,1703
_|1703,1704
_|1704,1705
<EOL>|1705,1706
Family|1706,1712
History|1713,1720
:|1720,1721
<EOL>|1721,1722
Non-contributory|1722,1738
<EOL>|1739,1740
<EOL>|1741,1742
Physical|1742,1750
Exam|1751,1755
:|1755,1756
<EOL>|1756,1757
VS|1757,1759
:|1759,1760
T|1761,1762
96.6|1763,1767
,|1767,1768
BP|1769,1771
140|1772,1775
/|1775,1776
palp|1776,1780
,|1780,1781
HR|1782,1784
64|1785,1787
,|1787,1788
RR|1789,1791
24|1792,1794
,|1794,1795
98|1796,1798
%|1798,1799
on|1800,1802
RA|1803,1805
<EOL>|1807,1808
GENERAL|1808,1815
:|1815,1816
Well|1817,1821
-|1821,1822
appearing|1822,1831
man|1832,1835
in|1836,1838
NAD|1839,1842
,|1842,1843
comfortable|1844,1855
,|1855,1856
appropriate|1857,1868
.|1868,1869
<EOL>|1871,1872
HEENT|1872,1877
:|1877,1878
NC|1879,1881
/|1881,1882
AT|1882,1884
,|1884,1885
sclerae|1886,1893
anicteric|1894,1903
,|1903,1904
MMM|1905,1908
<EOL>|1910,1911
HEART|1911,1916
:|1916,1917
irregularly|1918,1929
irregular|1930,1939
,|1939,1940
III|1941,1944
/|1944,1945
VI|1945,1947
systolic|1948,1956
ejection|1957,1965
murmur|1966,1972
<EOL>|1973,1974
loudest|1974,1981
at|1982,1984
the|1985,1988
LUS|1989,1992
boarder|1993,2000
,|2000,2001
nl|2002,2004
S1|2005,2007
-|2007,2008
S2|2008,2010
.|2010,2011
<EOL>|2013,2014
LUNGS|2014,2019
:|2019,2020
CTA|2021,2024
bilat|2025,2030
,|2030,2031
no|2032,2034
r|2035,2036
/|2036,2037
rh|2037,2039
/|2039,2040
wh|2040,2042
,|2042,2043
good|2044,2048
air|2049,2052
movement|2053,2061
,|2061,2062
resp|2063,2067
unlabored|2068,2077
.|2077,2078
<EOL>|2079,2080
<EOL>|2081,2082
ABDOMEN|2082,2089
:|2089,2090
Normoactive|2091,2102
BS|2103,2105
,|2105,2106
soft|2107,2111
/|2111,2112
NT|2112,2114
/|2114,2115
ND|2115,2117
,|2117,2118
no|2119,2121
masses|2122,2128
or|2129,2131
HSM|2132,2135
,|2135,2136
no|2137,2139
<EOL>|2140,2141
rebound|2141,2148
/|2148,2149
guarding|2149,2157
.|2157,2158
<EOL>|2160,2161
EXTREMITIES|2161,2172
:|2172,2173
Bruising|2174,2182
of|2183,2185
the|2186,2189
toes|2190,2194
of|2195,2197
the|2198,2201
left|2202,2206
foot|2207,2211
.|2211,2212
B|2213,2214
/|2214,2215
L|2215,2216
edema|2217,2222
,|2222,2223
<EOL>|2224,2225
most|2225,2229
pronounced|2230,2240
at|2241,2243
the|2244,2247
feet|2248,2252
/|2252,2253
ankles|2253,2259
,|2259,2260
3|2261,2262
+|2262,2263
to|2264,2266
the|2267,2270
thighs|2271,2277
.|2277,2278
<EOL>|2280,2281
NEURO|2281,2286
:|2286,2287
Awake|2288,2293
,|2293,2294
alert|2295,2300
,|2300,2301
conversant|2302,2312
,|2312,2313
grossly|2314,2321
intact|2322,2328
<EOL>|2330,2331
<EOL>|2331,2332
<EOL>|2333,2334
Pertinent|2334,2343
Results|2344,2351
:|2351,2352
<EOL>|2352,2353
ADMISSION|2353,2362
LABS|2363,2367
<EOL>|2367,2368
_|2368,2369
_|2369,2370
_|2370,2371
06|2372,2374
:|2374,2375
30PM|2375,2379
BLOOD|2380,2385
WBC|2386,2389
-|2389,2390
6|2390,2391
.|2391,2392
2|2392,2393
#|2393,2394
RBC|2395,2398
-|2398,2399
4|2399,2400
.|2400,2401
17|2401,2403
*|2403,2404
Hgb|2405,2408
-|2408,2409
13|2409,2411
.|2411,2412
3|2412,2413
*|2413,2414
Hct|2415,2418
-|2418,2419
40.3|2419,2423
<EOL>|2424,2425
MCV|2425,2428
-|2428,2429
97|2429,2431
MCH|2432,2435
-|2435,2436
32.0|2436,2440
MCHC|2441,2445
-|2445,2446
33.1|2446,2450
RDW|2451,2454
-|2454,2455
14.8|2455,2459
Plt|2460,2463
_|2464,2465
_|2465,2466
_|2466,2467
<EOL>|2467,2468
_|2468,2469
_|2469,2470
_|2470,2471
06|2472,2474
:|2474,2475
30PM|2475,2479
BLOOD|2480,2485
_|2486,2487
_|2487,2488
_|2488,2489
PTT|2490,2493
-|2493,2494
35|2494,2496
.|2496,2497
9|2497,2498
*|2498,2499
_|2500,2501
_|2501,2502
_|2502,2503
<EOL>|2503,2504
_|2504,2505
_|2505,2506
_|2506,2507
06|2508,2510
:|2510,2511
30PM|2511,2515
BLOOD|2516,2521
Glucose|2522,2529
-|2529,2530
210|2530,2533
*|2533,2534
UreaN|2535,2540
-|2540,2541
56|2541,2543
*|2543,2544
Creat|2545,2550
-|2550,2551
1|2551,2552
.|2552,2553
6|2553,2554
*|2554,2555
Na|2556,2558
-|2558,2559
141|2559,2562
<EOL>|2563,2564
K|2564,2565
-|2565,2566
3.6|2566,2569
Cl|2570,2572
-|2572,2573
99|2573,2575
HCO3|2576,2580
-|2580,2581
33|2581,2583
*|2583,2584
AnGap|2585,2590
-|2590,2591
13|2591,2593
<EOL>|2593,2594
_|2594,2595
_|2595,2596
_|2596,2597
06|2598,2600
:|2600,2601
30PM|2601,2605
BLOOD|2606,2611
ALT|2612,2615
-|2615,2616
49|2616,2618
*|2618,2619
AST|2620,2623
-|2623,2624
46|2624,2626
*|2626,2627
LD|2628,2630
(|2630,2631
LDH|2631,2634
)|2634,2635
-|2635,2636
440|2636,2639
*|2639,2640
CK|2641,2643
(|2643,2644
CPK|2644,2647
)|2647,2648
-|2648,2649
173|2649,2652
<EOL>|2653,2654
AlkPhos|2654,2661
-|2661,2662
66|2662,2664
TotBili|2665,2672
-|2672,2673
0.8|2673,2676
<EOL>|2676,2677
_|2677,2678
_|2678,2679
_|2679,2680
06|2681,2683
:|2683,2684
30PM|2684,2688
BLOOD|2689,2694
CK|2695,2697
-|2697,2698
MB|2698,2700
-|2700,2701
10|2701,2703
MB|2704,2706
Indx|2707,2711
-|2711,2712
5.8|2712,2715
proBNP|2716,2722
-|2722,2723
6310|2723,2727
*|2727,2728
<EOL>|2728,2729
<EOL>|2730,2731
DISCHARGE|2731,2740
LABS|2741,2745
<EOL>|2745,2746
_|2746,2747
_|2747,2748
_|2748,2749
06|2750,2752
:|2752,2753
07AM|2753,2757
BLOOD|2758,2763
WBC|2764,2767
-|2767,2768
4.9|2768,2771
RBC|2772,2775
-|2775,2776
4|2776,2777
.|2777,2778
10|2778,2780
*|2780,2781
Hgb|2782,2785
-|2785,2786
12|2786,2788
.|2788,2789
9|2789,2790
*|2790,2791
Hct|2792,2795
-|2795,2796
39|2796,2798
.|2798,2799
3|2799,2800
*|2800,2801
<EOL>|2802,2803
MCV|2803,2806
-|2806,2807
96|2807,2809
MCH|2810,2813
-|2813,2814
31.5|2814,2818
MCHC|2819,2823
-|2823,2824
32.9|2824,2828
RDW|2829,2832
-|2832,2833
14.6|2833,2837
Plt|2838,2841
Ct|2842,2844
-|2844,2845
95|2845,2847
*|2847,2848
<EOL>|2848,2849
_|2849,2850
_|2850,2851
_|2851,2852
08|2853,2855
:|2855,2856
05AM|2856,2860
BLOOD|2861,2866
_|2867,2868
_|2868,2869
_|2869,2870
<EOL>|2870,2871
_|2871,2872
_|2872,2873
_|2873,2874
08|2875,2877
:|2877,2878
05AM|2878,2882
BLOOD|2883,2888
UreaN|2889,2894
-|2894,2895
40|2895,2897
*|2897,2898
Creat|2899,2904
-|2904,2905
1|2905,2906
.|2906,2907
4|2907,2908
*|2908,2909
Na|2910,2912
-|2912,2913
140|2913,2916
K|2917,2918
-|2918,2919
3.5|2919,2922
Cl|2923,2925
-|2925,2926
103|2926,2929
<EOL>|2930,2931
HCO3|2931,2935
-|2935,2936
28|2936,2938
AnGap|2939,2944
-|2944,2945
13|2945,2947
<EOL>|2947,2948
_|2948,2949
_|2949,2950
_|2950,2951
06|2952,2954
:|2954,2955
07AM|2955,2959
BLOOD|2960,2965
CK|2966,2968
-|2968,2969
MB|2969,2971
-|2971,2972
7|2972,2973
cTropnT|2974,2981
-|2981,2982
0|2982,2983
.|2983,2984
01|2984,2986
<EOL>|2986,2987
<EOL>|2987,2988
CXR|2988,2991
_|2992,2993
_|2993,2994
_|2994,2995
:|2995,2996
1.|2997,2999
Mild|3000,3004
congestive|3005,3015
heart|3016,3021
failure|3022,3029
.|3029,3030
<EOL>|3032,3033
2.|3033,3035
Widened|3036,3043
superior|3044,3052
mediastinum|3053,3064
with|3065,3069
leftward|3070,3078
deviation|3079,3088
of|3089,3091
the|3092,3095
<EOL>|3096,3097
trachea|3097,3104
,|3104,3105
similar|3106,3113
when|3114,3118
compared|3119,3127
to|3128,3130
the|3131,3134
prior|3135,3140
study|3141,3146
.|3146,3147
Findings|3148,3156
may|3157,3160
<EOL>|3161,3162
reflect|3162,3169
the|3170,3173
presence|3174,3182
of|3183,3185
a|3186,3187
thyroid|3188,3195
goiter|3196,3202
,|3202,3203
and|3204,3207
clinical|3208,3216
<EOL>|3217,3218
correlation|3218,3229
is|3230,3232
recommended|3233,3244
,|3244,3245
and|3246,3249
if|3250,3252
indicated|3253,3262
,|3262,3263
this|3264,3268
could|3269,3274
be|3275,3277
<EOL>|3278,3279
confirmed|3279,3288
with|3289,3293
a|3294,3295
CT|3296,3298
of|3299,3301
the|3302,3305
chest|3306,3311
.|3311,3312
<EOL>|3314,3315
<EOL>|3317,3318
L|3318,3319
-|3319,3320
spine|3320,3325
film|3326,3330
_|3331,3332
_|3332,3333
_|3333,3334
:|3334,3335
Five|3336,3340
non-rib|3341,3348
-|3348,3349
bearing|3349,3356
lumbar|3357,3363
-|3363,3364
type|3364,3368
vertebral|3369,3378
<EOL>|3379,3380
<EOL>|3381,3382
bodies|3382,3388
are|3389,3392
present|3393,3400
.|3400,3401
There|3402,3407
are|3408,3411
multilevel|3412,3422
degenerative|3423,3435
changes|3436,3443
,|3443,3444
<EOL>|3445,3446
with|3446,3450
loss|3451,3455
of|3456,3458
intervertebral|3459,3473
disc|3474,3478
height|3479,3485
at|3486,3488
multiple|3489,3497
levels|3498,3504
,|3504,3505
<EOL>|3506,3507
endplate|3507,3515
sclerotic|3516,3525
changes|3526,3533
,|3533,3534
and|3535,3538
anterior|3539,3547
osteophyte|3548,3558
formation|3559,3568
.|3568,3569
<EOL>|3570,3571
There|3571,3576
is|3577,3579
no|3580,3582
fracture|3583,3591
or|3592,3594
vertebral|3595,3604
compression|3605,3616
deformity|3617,3626
<EOL>|3627,3628
identified|3628,3638
.|3638,3639
There|3640,3645
is|3646,3648
likely|3649,3655
mild|3656,3660
grade|3661,3666
1|3667,3668
L5|3669,3671
on|3672,3674
S1|3675,3677
<EOL>|3678,3679
anterolisthesis|3679,3694
,|3694,3695
which|3696,3701
is|3702,3704
likely|3705,3711
degenerative|3712,3724
in|3725,3727
etiology|3728,3736
.|3736,3737
Facet|3738,3743
<EOL>|3744,3745
hypertrophic|3745,3757
changes|3758,3765
are|3766,3769
noted|3770,3775
within|3776,3782
the|3783,3786
lower|3787,3792
lumbar|3793,3799
spine|3800,3805
<EOL>|3806,3807
primarily|3807,3816
affecting|3817,3826
L3|3827,3829
through|3830,3837
L5|3838,3840
levels|3841,3847
.|3847,3848
Vascular|3849,3857
<EOL>|3858,3859
calcifications|3859,3873
are|3874,3877
visualized|3878,3888
.|3888,3889
The|3890,3893
sacroiliac|3894,3904
joints|3905,3911
are|3912,3915
not|3916,3919
<EOL>|3920,3921
diastatic|3921,3930
.|3930,3931
<EOL>|3933,3934
IMPRESSION|3934,3944
:|3944,3945
No|3946,3948
fracture|3949,3957
identified|3958,3968
.|3968,3969
<EOL>|3971,3972
<EOL>|3972,3973
CT|3973,3975
head|3976,3980
_|3981,3982
_|3982,3983
_|3983,3984
:|3984,3985
<EOL>|3985,3986
There|3986,3991
is|3992,3994
no|3995,3997
acute|3998,4003
intracranial|4004,4016
hemorrhage|4017,4027
,|4027,4028
edema|4029,4034
or|4035,4037
acute|4038,4043
<EOL>|4044,4045
vascular|4045,4053
<EOL>|4054,4055
territorial|4055,4066
infarction|4067,4077
.|4077,4078
Note|4079,4083
is|4084,4086
made|4087,4091
of|4092,4094
areas|4095,4100
of|4101,4103
<EOL>|4104,4105
encephalomalacia|4105,4121
involving|4122,4131
the|4132,4135
parietal|4136,4144
lobe|4145,4149
on|4150,4152
the|4153,4156
left|4157,4161
,|4161,4162
which|4163,4168
<EOL>|4169,4170
appear|4170,4176
unchanged|4177,4186
as|4187,4189
does|4190,4194
an|4195,4197
area|4198,4202
of|4203,4205
hypodensity|4206,4217
on|4218,4220
the|4221,4224
right|4225,4230
<EOL>|4231,4232
adjacent|4232,4240
to|4241,4243
the|4244,4247
caudat|4248,4254
.|4254,4255
.|4255,4256
Similarly|4257,4266
unchanged|4267,4276
are|4277,4280
two|4281,4284
left|4285,4289
<EOL>|4290,4291
frontal|4291,4298
meningiomas|4299,4310
,|4310,4311
the|4312,4315
larger|4316,4322
of|4323,4325
which|4326,4331
is|4332,4334
partially|4335,4344
calcified|4345,4354
,|4354,4355
<EOL>|4356,4357
and|4357,4360
better|4361,4367
depicted|4368,4376
on|4377,4379
the|4380,4383
prior|4384,4389
MRI|4390,4393
(|4394,4395
2|4395,4396
:|4396,4397
24|4397,4399
,|4399,4400
601|4401,4404
:|4404,4405
19|4405,4407
)|4407,4408
.|4408,4409
Ventricles|4410,4420
<EOL>|4421,4422
and|4422,4425
sulci|4426,4431
are|4432,4435
enlarged|4436,4444
,|4444,4445
reflecting|4446,4456
parenchymal|4457,4468
volume|4469,4475
loss|4476,4480
.|4480,4481
Note|4482,4486
<EOL>|4487,4488
is|4488,4490
made|4491,4495
of|4496,4498
atherosclerotic|4499,4514
calcification|4515,4528
at|4529,4531
the|4532,4535
carotid|4536,4543
siphons|4544,4551
<EOL>|4552,4553
bilaterally|4553,4564
as|4565,4567
well|4568,4572
as|4573,4575
of|4576,4578
both|4579,4583
V4|4584,4586
segments|4587,4595
.|4595,4596
There|4597,4602
is|4603,4605
no|4606,4608
<EOL>|4609,4610
fracture|4610,4618
.|4618,4619
The|4620,4623
mastoid|4624,4631
air|4632,4635
cells|4636,4641
are|4642,4645
clear|4646,4651
.|4651,4652
<EOL>|4653,4654
IMPRESSION|4654,4664
:|4664,4665
No|4666,4668
acute|4669,4674
intracranial|4675,4687
abnormality|4688,4699
,|4699,4700
and|4701,4704
unchanged|4705,4714
<EOL>|4715,4716
findings|4716,4724
of|4725,4727
<EOL>|4728,4729
previous|4729,4737
infarcts|4738,4746
and|4747,4750
meningiomas|4751,4762
.|4762,4763
<EOL>|4764,4765
<EOL>|4765,4766
LENIs|4766,4771
_|4772,4773
_|4773,4774
_|4774,4775
:|4775,4776
<EOL>|4776,4777
Waveforms|4777,4786
in|4787,4789
the|4790,4793
common|4794,4800
femoral|4801,4808
veins|4809,4814
are|4815,4818
symmetric|4819,4828
bilaterally|4829,4840
<EOL>|4841,4842
with|4842,4846
appropriate|4847,4858
responses|4859,4868
to|4869,4871
Valsalva|4872,4880
maneuvers|4881,4890
.|4890,4891
In|4892,4894
both|4895,4899
lower|4900,4905
<EOL>|4906,4907
extremities|4907,4918
,|4918,4919
the|4920,4923
common|4924,4930
femoral|4931,4938
,|4938,4939
proximal|4940,4948
greater|4949,4956
saphenous|4957,4966
,|4966,4967
<EOL>|4968,4969
superficial|4969,4980
femoral|4981,4988
and|4989,4992
popliteal|4993,5002
veins|5003,5008
are|5009,5012
normal|5013,5019
with|5020,5024
<EOL>|5025,5026
appropriate|5026,5037
compressibility|5038,5053
,|5053,5054
wall|5055,5059
-|5059,5060
to|5060,5062
-|5062,5063
wall|5063,5067
flow|5068,5072
on|5073,5075
color|5076,5081
Doppler|5082,5089
<EOL>|5090,5091
analysis|5091,5099
and|5100,5103
response|5104,5112
to|5113,5115
waveform|5116,5124
augmentation|5125,5137
.|5137,5138
Wall|5139,5143
-|5143,5144
to|5144,5146
-|5146,5147
wall|5147,5151
<EOL>|5152,5153
flow|5153,5157
is|5158,5160
also|5161,5165
visualized|5166,5176
in|5177,5179
the|5180,5183
posterior|5184,5193
tibial|5194,5200
and|5201,5204
peroneal|5205,5213
<EOL>|5214,5215
veins|5215,5220
of|5221,5223
both|5224,5228
calves|5229,5235
.|5235,5236
<EOL>|5236,5237
IMPRESSION|5237,5247
:|5247,5248
No|5249,5251
deep|5252,5256
venous|5257,5263
thrombosis|5264,5274
in|5275,5277
either|5278,5284
lower|5285,5290
extremity|5291,5300
.|5300,5301
<EOL>|5302,5303
<EOL>|5303,5304
<EOL>|5306,5307
<EOL>|5307,5308
MICROBIOLOGY|5308,5320
:|5320,5321
<EOL>|5322,5323
_|5323,5324
_|5324,5325
_|5325,5326
:|5326,5327
Blood|5328,5333
culture|5334,5341
-|5342,5343
no|5344,5346
growth|5347,5353
to|5354,5356
date|5357,5361
<EOL>|5361,5362
<EOL>|5362,5363
<EOL>|5364,5365
Brief|5365,5370
Hospital|5371,5379
Course|5380,5386
:|5386,5387
<EOL>|5387,5388
_|5388,5389
_|5389,5390
_|5390,5391
yo|5392,5394
M|5395,5396
with|5397,5401
DM|5402,5404
,|5404,5405
afib|5406,5410
,|5410,5411
and|5412,5415
CHF|5416,5419
presenting|5420,5430
with|5431,5435
pulm|5436,5440
edema|5441,5446
and|5447,5450
<EOL>|5451,5452
worsening|5452,5461
_|5462,5463
_|5463,5464
_|5464,5465
edema|5466,5471
.|5471,5472
<EOL>|5472,5473
<EOL>|5474,5475
#|5475,5476
CHF|5477,5480
:|5480,5481
Likely|5482,5488
an|5489,5491
acute|5492,5497
on|5498,5500
chronic|5501,5508
worsening|5509,5518
of|5519,5521
diastolic|5522,5531
<EOL>|5532,5533
congestive|5533,5543
heart|5544,5549
failure|5550,5557
(|5558,5559
most|5559,5563
recent|5564,5570
LVEF|5571,5575
>|5576,5577
55|5577,5579
%|5579,5580
)|5580,5581
and|5582,5585
recent|5586,5592
<EOL>|5593,5594
decrease|5594,5602
in|5603,5605
mobility|5606,5614
from|5615,5619
fall|5620,5624
.|5624,5625
Ruled|5626,5631
out|5632,5635
for|5636,5639
MI|5640,5642
.|5642,5643
Likely|5644,5650
his|5651,5654
<EOL>|5655,5656
worsening|5656,5665
edema|5666,5671
is|5672,5674
due|5675,5678
to|5679,5681
medication|5682,5692
non-compliance|5693,5707
versus|5708,5714
<EOL>|5715,5716
worsening|5716,5725
of|5726,5728
his|5729,5732
aortic|5733,5739
stenosis|5740,5748
.|5748,5749
His|5750,5753
most|5754,5758
recent|5759,5765
echo|5766,5770
is|5771,5773
from|5774,5778
<EOL>|5779,5780
_|5780,5781
_|5781,5782
_|5782,5783
,|5783,5784
and|5785,5788
it|5789,5791
was|5792,5795
recommended|5796,5807
this|5808,5812
be|5813,5815
repeated|5816,5824
as|5825,5827
an|5828,5830
outpatient|5831,5841
.|5841,5842
<EOL>|5843,5844
He|5844,5846
was|5847,5850
never|5851,5856
hypoxic|5857,5864
,|5864,5865
though|5866,5872
lung|5873,5877
exam|5878,5882
suggested|5883,5892
increased|5893,5902
pulm|5903,5907
<EOL>|5908,5909
edema|5909,5914
.|5914,5915
His|5916,5919
legs|5920,5924
were|5925,5929
elevated|5930,5938
and|5939,5942
compression|5943,5954
stockings|5955,5964
were|5965,5969
<EOL>|5970,5971
used|5971,5975
.|5975,5976
His|5977,5980
torsemide|5981,5990
was|5991,5994
dosed|5995,6000
at|6001,6003
10mg|6004,6008
daily|6009,6014
,|6014,6015
though|6016,6022
it|6023,6025
's|6025,6027
unclear|6028,6035
<EOL>|6036,6037
if|6037,6039
this|6040,6044
was|6045,6048
an|6049,6051
increase|6052,6060
from|6061,6065
5mg|6066,6069
or|6070,6072
the|6073,6076
same|6077,6081
dose|6082,6086
,|6086,6087
and|6088,6091
the|6092,6095
<EOL>|6096,6097
patient|6097,6104
and|6105,6108
wife|6109,6113
were|6114,6118
unable|6119,6125
to|6126,6128
clarify|6129,6136
.|6136,6137
There|6138,6143
was|6144,6147
slight|6148,6154
<EOL>|6155,6156
improvement|6156,6167
in|6168,6170
swelling|6171,6179
on|6180,6182
discharge|6183,6192
.|6192,6193
<EOL>|6193,6194
<EOL>|6195,6196
#|6196,6197
RECENT|6198,6204
FALLS|6205,6210
:|6210,6211
Patient|6212,6219
reports|6220,6227
falling|6228,6235
twice|6236,6241
recently|6242,6250
at|6251,6253
home|6254,6258
<EOL>|6259,6260
and|6260,6263
on|6264,6266
a|6267,6268
trip|6269,6273
.|6273,6274
He|6275,6277
was|6278,6281
evaluated|6282,6291
by|6292,6294
physical|6295,6303
therapy|6304,6311
,|6311,6312
who|6313,6316
felt|6317,6321
he|6322,6324
<EOL>|6325,6326
is|6326,6328
unsteady|6329,6337
on|6338,6340
his|6341,6344
feet|6345,6349
but|6350,6353
safe|6354,6358
for|6359,6362
discharge|6363,6372
home|6373,6377
with|6378,6382
_|6383,6384
_|6384,6385
_|6385,6386
and|6387,6390
<EOL>|6391,6392
a|6392,6393
walker|6394,6400
/|6400,6401
commode|6401,6408
.|6408,6409
The|6410,6413
wife|6414,6418
was|6419,6422
instructed|6423,6433
to|6434,6436
maintain|6437,6445
24|6446,6448
hour|6449,6453
<EOL>|6454,6455
care|6455,6459
for|6460,6463
him|6464,6467
in|6468,6470
the|6471,6474
home|6475,6479
to|6480,6482
help|6483,6487
prevent|6488,6495
further|6496,6503
falls|6504,6509
.|6509,6510
<EOL>|6511,6512
<EOL>|6512,6513
#|6513,6514
_|6515,6516
_|6516,6517
_|6517,6518
:|6518,6519
Cr|6520,6522
up|6523,6525
to|6526,6528
1.6|6529,6532
on|6533,6535
admission|6536,6545
.|6545,6546
Improved|6547,6555
to|6556,6558
1.3|6559,6562
the|6563,6566
next|6567,6571
day|6572,6575
,|6575,6576
<EOL>|6577,6578
likely|6578,6584
closer|6585,6591
to|6592,6594
baseline|6595,6603
.|6603,6604
<EOL>|6605,6606
<EOL>|6609,6610
#|6610,6611
DM|6612,6614
:|6614,6615
Glipizide|6616,6625
and|6626,6629
actos|6630,6635
held|6636,6640
while|6641,6646
in|6647,6649
hospital|6650,6658
.|6658,6659
Covered|6660,6667
with|6668,6672
<EOL>|6673,6674
an|6674,6676
insulin|6677,6684
sliding|6685,6692
scale|6693,6698
and|6699,6702
oral|6703,6707
medications|6708,6719
restarted|6720,6729
on|6730,6732
<EOL>|6733,6734
discharge|6734,6743
.|6743,6744
<EOL>|6744,6745
<EOL>|6747,6748
#|6748,6749
HTN|6750,6753
:|6753,6754
Continued|6755,6764
isosorbide|6765,6775
and|6776,6779
lisinopril|6780,6790
(|6791,6792
held|6792,6796
for|6797,6800
one|6801,6804
day|6805,6808
<EOL>|6809,6810
given|6810,6815
_|6816,6817
_|6817,6818
_|6818,6819
.|6819,6820
Metoprolol|6821,6831
dose|6832,6836
was|6837,6840
lowered|6841,6848
to|6849,6851
25mg|6852,6856
TID|6857,6860
given|6861,6866
his|6867,6870
<EOL>|6871,6872
bradycardia|6872,6883
.|6883,6884
<EOL>|6884,6885
<EOL>|6885,6886
#|6886,6887
Afib|6888,6892
:|6892,6893
INR|6894,6897
was|6898,6901
2.9|6902,6905
on|6906,6908
admission|6909,6918
,|6918,6919
and|6920,6923
unclear|6924,6931
if|6932,6934
he|6935,6937
had|6938,6941
taken|6942,6947
<EOL>|6948,6949
his|6949,6952
daily|6953,6958
coumadin|6959,6967
dose|6968,6972
.|6972,6973
He|6974,6976
was|6977,6980
restarted|6981,6990
at|6991,6993
2.5|6994,6997
mg|6997,6999
daily|7000,7005
.|7005,7006
His|7007,7010
<EOL>|7011,7012
wife|7012,7016
noted|7017,7022
that|7023,7027
he|7028,7030
had|7031,7034
been|7035,7039
switched|7040,7048
to|7049,7051
alternate|7052,7061
1.25|7062,7066
mg|7066,7068
with|7069,7073
<EOL>|7074,7075
2.5|7075,7078
mg|7078,7080
.|7080,7081
He|7082,7084
was|7085,7088
discharged|7089,7099
with|7100,7104
home|7105,7109
services|7110,7118
to|7119,7121
follow|7122,7128
INRs|7129,7133
.|7133,7134
<EOL>|7134,7135
<EOL>|7135,7136
TRANSITIONAL|7136,7148
ISSUES|7149,7155
:|7155,7156
<EOL>|7156,7157
Blood|7157,7162
culture|7163,7170
_|7171,7172
_|7172,7173
_|7173,7174
_|7175,7176
_|7176,7177
_|7177,7178
needs|7179,7184
to|7185,7187
be|7188,7190
follow|7191,7197
up|7198,7200
-|7201,7202
no|7203,7205
growth|7206,7212
to|7213,7215
<EOL>|7216,7217
date|7217,7221
.|7221,7222
<EOL>|7222,7223
<EOL>|7224,7225
Medications|7225,7236
on|7237,7239
Admission|7240,7249
:|7249,7250
<EOL>|7250,7251
-|7251,7252
Allopurinol|7252,7263
_|7264,7265
_|7265,7266
_|7266,7267
MG|7268,7270
(|7271,7272
100|7272,7275
MG|7276,7278
TABLET|7279,7285
Take|7286,7290
1|7291,7292
)|7292,7293
PO|7294,7296
QD|7297,7299
_|7300,7301
_|7301,7302
_|7302,7303
<EOL>|7305,7306
-|7306,7307
Cyanocobalamin|7307,7321
1000|7322,7326
MCG|7327,7330
(|7331,7332
1000MCG|7332,7339
/|7339,7340
ML|7340,7342
VIAL|7343,7347
Take|7348,7352
1|7353,7354
ML|7355,7357
)|7357,7358
IM|7359,7361
QMONTH|7362,7368
<EOL>|7369,7370
_|7370,7371
_|7371,7372
_|7372,7373
<EOL>|7375,7376
-|7376,7377
Dexamethasone|7377,7390
0.5|7391,7394
MG|7395,7397
(|7398,7399
0.5|7399,7402
MG|7403,7405
TABLET|7406,7412
Take|7413,7417
1|7418,7419
)|7419,7420
PO|7421,7423
QD|7424,7426
_|7427,7428
_|7428,7429
_|7429,7430
<EOL>|7432,7433
-|7433,7434
Glipizide|7434,7443
10|7444,7446
MG|7447,7449
(|7450,7451
10|7451,7453
MG|7454,7456
TABLET|7457,7463
Take|7464,7468
1|7469,7470
)|7470,7471
PO|7472,7474
BID|7475,7478
_|7479,7480
_|7480,7481
_|7481,7482
<EOL>|7484,7485
-|7485,7486
Goserelin|7486,7495
acetate|7496,7503
10.8|7504,7508
MG|7509,7511
(|7512,7513
10.8|7513,7517
MG|7517,7519
IMPLANT|7520,7527
Take|7528,7532
1|7533,7534
)|7534,7535
SC|7536,7538
QMONTH|7539,7545
<EOL>|7546,7547
_|7547,7548
_|7548,7549
_|7549,7550
<EOL>|7552,7553
-|7553,7554
Isosorbide|7554,7564
dinitrate|7565,7574
10|7575,7577
MG|7578,7580
(|7581,7582
10|7582,7584
MG|7585,7587
TABLET|7588,7594
Take|7595,7599
1|7600,7601
)|7601,7602
PO|7603,7605
BID|7606,7609
<EOL>|7610,7611
_|7611,7612
_|7612,7613
_|7613,7614
<EOL>|7616,7617
-|7617,7618
Lisinopril|7618,7628
20|7629,7631
MG|7632,7634
(|7635,7636
20|7636,7638
MG|7639,7641
TABLET|7642,7648
Take|7649,7653
1|7654,7655
)|7655,7656
PO|7657,7659
QD|7660,7662
_|7663,7664
_|7664,7665
_|7665,7666
<EOL>|7668,7669
-|7669,7670
Memantine|7670,7679
PO|7680,7682
_|7683,7684
_|7684,7685
_|7685,7686
<EOL>|7688,7689
-|7689,7690
Metoprolol|7690,7700
tartrate|7701,7709
50|7710,7712
MG|7713,7715
(|7716,7717
50|7717,7719
MG|7720,7722
TABLET|7723,7729
Take|7730,7734
1|7735,7736
)|7736,7737
PO|7738,7740
TID|7741,7744
_|7745,7746
_|7746,7747
_|7747,7748
<EOL>|7749,7750
<EOL>|7751,7752
-|7752,7753
Nilutamide|7753,7763
150|7764,7767
MG|7768,7770
(|7771,7772
150|7772,7775
MG|7776,7778
TABLET|7779,7785
Take|7786,7790
1|7791,7792
)|7792,7793
PO|7794,7796
QD|7797,7799
_|7800,7801
_|7801,7802
_|7802,7803
<EOL>|7805,7806
-|7806,7807
Nitroglycerin|7807,7820
PO|7821,7823
_|7824,7825
_|7825,7826
_|7826,7827
<EOL>|7829,7830
-|7830,7831
Oxycodone|7831,7840
5|7841,7842
MG|7843,7845
(|7846,7847
5MG|7847,7850
TABLET|7851,7857
Take|7858,7862
1|7863,7864
)|7864,7865
PO|7866,7868
Q6H|7869,7872
PRN|7873,7876
pain|7877,7881
_|7882,7883
_|7883,7884
_|7884,7885
<EOL>|7887,7888
-|7888,7889
Prednisone|7889,7899
Taper|7900,7905
(|7906,7907
10|7907,7909
MG|7910,7912
TABLET|7913,7919
Take|7920,7924
1|7925,7926
)|7926,7927
PO|7928,7930
x|7931,7932
19|7933,7935
days|7936,7940
_|7941,7942
_|7942,7943
_|7943,7944
<EOL>|7946,7947
-|7947,7948
Simvastatin|7948,7959
20|7960,7962
MG|7963,7965
(|7966,7967
20|7967,7969
MG|7970,7972
TABLET|7973,7979
Take|7980,7984
1|7985,7986
)|7986,7987
PO|7988,7990
QPM|7991,7994
_|7995,7996
_|7996,7997
_|7997,7998
<EOL>|8000,8001
-|8001,8002
Torsemide|8002,8011
5|8012,8013
MG|8014,8016
(|8017,8018
5|8018,8019
MG|8020,8022
TABLET|8023,8029
Take|8030,8034
1|8035,8036
)|8036,8037
PO|8038,8040
QD|8041,8043
_|8044,8045
_|8045,8046
_|8046,8047
<EOL>|8049,8050
-|8050,8051
Warfarin|8051,8059
sodium|8060,8066
2.5|8067,8070
MG|8071,8073
(|8074,8075
2.5|8075,8078
MG|8079,8081
TABLET|8082,8088
Take|8089,8093
1|8094,8095
)|8095,8096
PO|8097,8099
as|8100,8102
directed|8103,8111
<EOL>|8113,8114
<EOL>|8114,8115
<EOL>|8116,8117
Discharge|8117,8126
Medications|8127,8138
:|8138,8139
<EOL>|8139,8140
1.|8140,8142
dexamethasone|8143,8156
0.5|8157,8160
mg|8161,8163
Tablet|8164,8170
Sig|8171,8174
:|8174,8175
One|8176,8179
(|8180,8181
1|8181,8182
)|8182,8183
Tablet|8184,8190
PO|8191,8193
once|8194,8198
a|8199,8200
<EOL>|8201,8202
day|8202,8205
.|8205,8206
<EOL>|8208,8209
2.|8209,8211
glipizide|8212,8221
10|8222,8224
mg|8225,8227
Tablet|8228,8234
Sig|8235,8238
:|8238,8239
One|8240,8243
(|8244,8245
1|8245,8246
)|8246,8247
Tablet|8248,8254
PO|8255,8257
once|8258,8262
a|8263,8264
day|8265,8268
.|8268,8269
<EOL>|8271,8272
3.|8272,8274
goserelin|8275,8284
10.8|8285,8289
mg|8290,8292
Implant|8293,8300
Sig|8301,8304
:|8304,8305
One|8306,8309
(|8310,8311
1|8311,8312
)|8312,8313
implant|8314,8321
Subcutaneous|8322,8334
<EOL>|8335,8336
as|8336,8338
directed|8339,8347
.|8347,8348
<EOL>|8350,8351
4.|8351,8353
isosorbide|8354,8364
dinitrate|8365,8374
10|8375,8377
mg|8378,8380
Tablet|8381,8387
Sig|8388,8391
:|8391,8392
One|8393,8396
(|8397,8398
1|8398,8399
)|8399,8400
Tablet|8401,8407
PO|8408,8410
<EOL>|8411,8412
twice|8412,8417
a|8418,8419
day|8420,8423
.|8423,8424
<EOL>|8426,8427
5.|8427,8429
lisinopril|8430,8440
20|8441,8443
mg|8444,8446
Tablet|8447,8453
Sig|8454,8457
:|8457,8458
One|8459,8462
(|8463,8464
1|8464,8465
)|8465,8466
Tablet|8467,8473
PO|8474,8476
once|8477,8481
a|8482,8483
day|8484,8487
.|8487,8488
<EOL>|8490,8491
6.|8491,8493
metoprolol|8494,8504
tartrate|8505,8513
25|8514,8516
mg|8517,8519
Tablet|8520,8526
Sig|8527,8530
:|8530,8531
One|8532,8535
(|8536,8537
1|8537,8538
)|8538,8539
Tablet|8540,8546
PO|8547,8549
three|8550,8555
<EOL>|8556,8557
times|8557,8562
a|8563,8564
day|8565,8568
.|8568,8569
<EOL>|8569,8570
Disp|8570,8574
:|8574,8575
*|8575,8576
90|8576,8578
Tablet|8579,8585
(|8585,8586
s|8586,8587
)|8587,8588
*|8588,8589
Refills|8590,8597
:|8597,8598
*|8598,8599
0|8599,8600
*|8600,8601
<EOL>|8601,8602
7.|8602,8604
nilutamide|8605,8615
150|8616,8619
mg|8620,8622
Tablet|8623,8629
Sig|8630,8633
:|8633,8634
One|8635,8638
(|8639,8640
1|8640,8641
)|8641,8642
Tablet|8643,8649
PO|8650,8652
once|8653,8657
a|8658,8659
day|8660,8663
.|8663,8664
<EOL>|8666,8667
8.|8667,8669
oxycodone|8670,8679
5|8680,8681
mg|8682,8684
Tablet|8685,8691
Sig|8692,8695
:|8695,8696
One|8697,8700
(|8701,8702
1|8702,8703
)|8703,8704
Tablet|8705,8711
PO|8712,8714
every|8715,8720
six|8721,8724
(|8725,8726
6|8726,8727
)|8727,8728
<EOL>|8729,8730
hours|8730,8735
as|8736,8738
needed|8739,8745
for|8746,8749
pain|8750,8754
.|8754,8755
<EOL>|8757,8758
9.|8758,8760
simvastatin|8761,8772
40|8773,8775
mg|8776,8778
Tablet|8779,8785
Sig|8786,8789
:|8789,8790
0.5|8791,8794
Tablet|8795,8801
PO|8802,8804
DAILY|8805,8810
(|8811,8812
Daily|8812,8817
)|8817,8818
.|8818,8819
<EOL>|8821,8822
10.|8822,8825
torsemide|8826,8835
10|8836,8838
mg|8839,8841
Tablet|8842,8848
Sig|8849,8852
:|8852,8853
One|8854,8857
(|8858,8859
1|8859,8860
)|8860,8861
Tablet|8862,8868
PO|8869,8871
once|8872,8876
a|8877,8878
day|8879,8882
.|8882,8883
<EOL>|8883,8884
Disp|8884,8888
:|8888,8889
*|8889,8890
30|8890,8892
Tablet|8893,8899
(|8899,8900
s|8900,8901
)|8901,8902
*|8902,8903
Refills|8904,8911
:|8911,8912
*|8912,8913
0|8913,8914
*|8914,8915
<EOL>|8915,8916
11.|8916,8919
cyanocobalamin|8920,8934
(|8935,8936
vitamin|8936,8943
B|8944,8945
-|8945,8946
12|8946,8948
)|8948,8949
1,000|8950,8955
mcg|8956,8959
/|8959,8960
15|8960,8962
mL|8963,8965
Liquid|8966,8972
Sig|8973,8976
:|8976,8977
<EOL>|8978,8979
One|8979,8982
(|8983,8984
1|8984,8985
)|8985,8986
dose|8987,8991
PO|8992,8994
once|8995,8999
a|9000,9001
week|9002,9006
.|9006,9007
<EOL>|9009,9010
12.|9010,9013
memantine|9014,9023
10|9024,9026
mg|9027,9029
Tablet|9030,9036
Sig|9037,9040
:|9040,9041
One|9042,9045
(|9046,9047
1|9047,9048
)|9048,9049
Tablet|9050,9056
PO|9057,9059
twice|9060,9065
a|9066,9067
day|9068,9071
.|9071,9072
<EOL>|9074,9075
13.|9075,9078
allopurinol|9079,9090
_|9091,9092
_|9092,9093
_|9093,9094
mg|9095,9097
Tablet|9098,9104
Sig|9105,9108
:|9108,9109
Two|9110,9113
(|9114,9115
2|9115,9116
)|9116,9117
Tablet|9118,9124
PO|9125,9127
once|9128,9132
a|9133,9134
day|9135,9138
.|9138,9139
<EOL>|9140,9141
<EOL>|9142,9143
14.|9143,9146
warfarin|9147,9155
2.5|9156,9159
mg|9160,9162
Tablet|9163,9169
Sig|9170,9173
:|9173,9174
One|9175,9178
(|9179,9180
1|9180,9181
)|9181,9182
Tablet|9183,9189
PO|9190,9192
_|9193,9194
_|9194,9195
_|9195,9196
,|9196,9197
Th|9198,9200
,|9200,9201
Sa|9202,9204
:|9204,9205
<EOL>|9206,9207
and|9207,9210
0.5|9211,9214
tablets|9215,9222
on|9223,9225
Mo|9226,9228
,|9228,9229
We|9230,9232
,|9232,9233
Fr|9234,9236
and|9237,9240
_|9241,9242
_|9242,9243
_|9243,9244
.|9244,9245
<EOL>|9247,9248
15|9248,9250
.|9250,9251
Vitamin|9252,9259
D|9260,9261
1,000|9262,9267
unit|9268,9272
Tablet|9273,9279
Sig|9280,9283
:|9283,9284
One|9285,9288
(|9289,9290
1|9290,9291
)|9291,9292
Tablet|9293,9299
PO|9300,9302
once|9303,9307
a|9308,9309
<EOL>|9310,9311
day|9311,9314
.|9314,9315
<EOL>|9317,9318
16.|9318,9321
insulin|9322,9329
glargine|9330,9338
100|9339,9342
unit|9343,9347
/|9347,9348
mL|9348,9350
Cartridge|9351,9360
Sig|9361,9364
:|9364,9365
Ten|9366,9369
(|9370,9371
10|9371,9373
)|9373,9374
units|9375,9380
<EOL>|9381,9382
Subcutaneous|9382,9394
at|9395,9397
bedtime|9398,9405
.|9405,9406
<EOL>|9408,9409
<EOL>|9409,9410
<EOL>|9411,9412
Discharge|9412,9421
Disposition|9422,9433
:|9433,9434
<EOL>|9434,9435
Home|9435,9439
With|9440,9444
Service|9445,9452
<EOL>|9452,9453
<EOL>|9454,9455
Facility|9455,9463
:|9463,9464
<EOL>|9464,9465
_|9465,9466
_|9466,9467
_|9467,9468
<EOL>|9468,9469
<EOL>|9470,9471
Discharge|9471,9480
Diagnosis|9481,9490
:|9490,9491
<EOL>|9491,9492
PRIMARY|9492,9499
<EOL>|9499,9500
Acute|9500,9505
on|9506,9508
chronic|9509,9516
diastolic|9517,9526
congestive|9527,9537
heart|9538,9543
failure|9544,9551
<EOL>|9551,9552
<EOL>|9552,9553
SECONDARY|9553,9562
<EOL>|9562,9563
Atrial|9563,9569
fibrillation|9570,9582
<EOL>|9582,9583
Diabetes|9583,9591
<EOL>|9591,9592
Hypertension|9592,9604
<EOL>|9604,9605
<EOL>|9606,9607
Discharge|9607,9616
Condition|9617,9626
:|9626,9627
<EOL>|9627,9628
Mental|9628,9634
Status|9635,9641
:|9641,9642
Clear|9643,9648
and|9649,9652
coherent|9653,9661
.|9661,9662
<EOL>|9662,9663
Level|9663,9668
of|9669,9671
Consciousness|9672,9685
:|9685,9686
Alert|9687,9692
and|9693,9696
interactive|9697,9708
.|9708,9709
<EOL>|9709,9710
Activity|9710,9718
Status|9719,9725
:|9725,9726
Ambulatory|9727,9737
-|9738,9739
requires|9740,9748
assistance|9749,9759
or|9760,9762
aid|9763,9766
(|9767,9768
walker|9768,9774
<EOL>|9775,9776
or|9776,9778
cane|9779,9783
)|9783,9784
.|9784,9785
<EOL>|9785,9786
<EOL>|9787,9788
Discharge|9788,9797
Instructions|9798,9810
:|9810,9811
<EOL>|9811,9812
Mr.|9812,9815
_|9816,9817
_|9817,9818
_|9818,9819
,|9819,9820
<EOL>|9820,9821
<EOL>|9822,9823
You|9823,9826
were|9827,9831
admitted|9832,9840
to|9841,9843
the|9844,9847
hospital|9848,9856
for|9857,9860
swelling|9861,9869
in|9870,9872
your|9873,9877
legs|9878,9882
,|9882,9883
<EOL>|9884,9885
likely|9885,9891
due|9892,9895
to|9896,9898
your|9899,9903
heart|9904,9909
failure|9910,9917
.|9917,9918
We|9919,9921
increased|9922,9931
your|9932,9936
diuretic|9937,9945
<EOL>|9946,9947
dosing|9947,9953
and|9954,9957
had|9958,9961
you|9962,9965
work|9966,9970
with|9971,9975
physical|9976,9984
therapy|9985,9992
.|9992,9993
<EOL>|9993,9994
<EOL>|9994,9995
Please|9995,10001
weigh|10002,10007
yourself|10008,10016
daily|10017,10022
and|10023,10026
notify|10027,10033
your|10034,10038
doctor|10039,10045
if|10046,10048
your|10049,10053
<EOL>|10054,10055
weight|10055,10061
increases|10062,10071
by|10072,10074
more|10075,10079
than|10080,10084
3|10085,10086
pounds|10087,10093
<EOL>|10093,10094
<EOL>|10094,10095
Medication|10095,10105
changes|10106,10113
:|10113,10114
<EOL>|10114,10115
#|10115,10116
CONTINUE|10117,10125
torsemide|10126,10135
10mg|10136,10140
daily|10141,10146
to|10147,10149
help|10150,10154
remove|10155,10161
fluid|10162,10167
<EOL>|10167,10168
#|10168,10169
REDUCE|10170,10176
metoprolol|10177,10187
to|10188,10190
25mg|10191,10195
daily|10196,10201
as|10202,10204
your|10205,10209
blood|10210,10215
pressure|10216,10224
has|10225,10228
<EOL>|10229,10230
been|10230,10234
low|10235,10238
while|10239,10244
you|10245,10248
were|10249,10253
hospitalized|10254,10266
.|10266,10267
Your|10269,10273
doctor|10274,10280
may|10281,10284
decide|10285,10291
to|10292,10294
<EOL>|10295,10296
increase|10296,10304
it|10305,10307
again|10308,10313
at|10314,10316
your|10317,10321
office|10322,10328
visit|10329,10334
.|10334,10335
<EOL>|10335,10336
<EOL>|10337,10338
Followup|10338,10346
Instructions|10347,10359
:|10359,10360
<EOL>|10360,10361
_|10361,10362
_|10362,10363
_|10363,10364
<EOL>|10364,10365

