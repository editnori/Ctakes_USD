 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
_|27,28
_|28,29
_|29,30
No|31,33
:|33,34
_|37,38
_|38,39
_|39,40
<EOL>|40,41
<EOL>|42,43
Admission|43,52
Date|53,57
:|57,58
_|60,61
_|61,62
_|62,63
Discharge|77,86
Date|87,91
:|91,92
_|95,96
_|96,97
_|97,98
<EOL>|98,99
<EOL>|100,101
Date|101,105
of|106,108
Birth|109,114
:|114,115
_|117,118
_|118,119
_|119,120
Sex|133,136
:|136,137
F|140,141
<EOL>|141,142
<EOL>|143,144
Service|144,151
:|151,152
MEDICINE|153,161
<EOL>|161,162
<EOL>|163,164
meropenem|176,185
/|186,187
Penicillins|188,199
<EOL>|199,200
<EOL>|201,202
Attending|202,211
:|211,212
_|213,214
_|214,215
_|215,216
.|216,217
<EOL>|217,218
<EOL>|219,220
BRBPR|237,242
<EOL>|242,243
<EOL>|244,245
Major|245,250
Surgical|251,259
or|260,262
Invasive|263,271
Procedure|272,281
:|281,282
<EOL>|282,283
aborted|283,290
flexible|291,299
sigmoidoscopy|300,313
attempt|314,321
(|322,323
due|323,326
to|327,329
stool|330,335
in|336,338
vault|339,344
)|344,345
<EOL>|346,347
_|347,348
_|348,349
_|349,350
<EOL>|350,351
Flexible|351,359
sigmoidoscopy|360,373
_|374,375
_|375,376
_|376,377
<EOL>|377,378
<EOL>|378,379
<EOL>|380,381
This|409,413
is|414,416
an|417,419
_|420,421
_|421,422
_|422,423
year|424,428
old|429,432
female|433,439
with|440,444
past|445,449
medical|450,457
history|458,465
of|466,468
<EOL>|468,469
sjogrens|469,477
,|477,478
hypothyroidism|479,493
,|493,494
recent|495,501
diagnosis|502,511
of|512,514
L1|515,517
compression|518,529
<EOL>|529,530
fracture|530,538
,|538,539
prior|540,545
cdiff|546,551
infection|552,561
,|561,562
presenting|563,573
with|574,578
bright|579,585
red|586,589
<EOL>|590,591
blood|591,596
<EOL>|596,597
per|597,600
rectum|601,607
.|607,608
Patient|610,617
reports|618,625
that|626,630
on|631,633
morning|634,641
of|642,644
presentation|645,657
,|657,658
<EOL>|659,660
she|660,663
<EOL>|663,664
awoke|664,669
in|670,672
her|673,676
normal|677,683
state|684,689
of|690,692
health|693,699
.|699,700
Her|702,705
home|706,710
health|711,717
aid|718,721
helped|722,728
<EOL>|728,729
her|729,732
to|733,735
the|736,739
commode|740,747
and|748,751
she|752,755
suddenly|756,764
had|765,768
a|769,770
large|771,776
volume|777,783
over|784,788
<EOL>|789,790
blood|790,795
<EOL>|795,796
per|796,799
rectum|800,806
.|806,807
Over|809,813
the|814,817
next|818,822
_|823,824
_|824,825
_|825,826
minutes|827,834
she|835,838
then|839,843
had|844,847
2|848,849
subsequent|850,860
<EOL>|860,861
episodes|861,869
.|869,870
Home|872,876
health|877,883
aid|884,887
consulted|888,897
with|898,902
family|903,909
and|910,913
then|914,918
called|919,925
<EOL>|925,926
_|926,927
_|927,928
_|928,929
.|929,930
<EOL>|932,933
<EOL>|933,934
In|934,936
the|937,940
ED|941,943
VS|944,946
were|947,951
97.2|952,956
98|957,959
158|960,963
/|963,964
89|964,966
14|967,969
98|970,972
%|972,973
RA|973,975
_|976,977
_|977,978
_|978,979
99.|980,983
Labs|985,989
were|990,994
<EOL>|994,995
notable|995,1002
for|1003,1006
WBC|1007,1010
10.1|1011,1015
,|1015,1016
Hgb|1017,1020
9.8|1021,1024
,|1024,1025
Plt|1026,1029
245|1030,1033
;|1033,1034
K|1035,1036
4.4|1037,1040
,|1040,1041
Cr|1042,1044
0.6|1045,1048
;|1048,1049
lactate|1050,1057
<EOL>|1057,1058
1.0|1058,1061
;|1061,1062
UA|1063,1065
neg|1066,1069
leuk|1070,1074
,|1074,1075
nitr|1076,1080
.|1080,1081
Exam|1083,1087
reported|1088,1096
as|1097,1099
tachycardia|1100,1111
,|1111,1112
grossly|1113,1120
<EOL>|1120,1121
blood|1121,1126
rectum|1127,1133
without|1134,1141
large|1142,1147
hemorrhoids|1148,1159
.|1159,1160
PEG|1161,1164
lavage|1165,1171
reported|1172,1180
as|1181,1183
<EOL>|1183,1184
negative|1184,1192
for|1193,1196
blood|1197,1202
.|1202,1203
<EOL>|1203,1204
<EOL>|1204,1205
GI|1205,1207
note|1208,1212
on|1213,1215
the|1216,1219
ED|1220,1222
dashboard|1223,1232
stated|1233,1239
_|1240,1241
_|1241,1242
_|1242,1243
with|1244,1248
C|1249,1250
.|1250,1251
diff|1251,1255
on|1256,1258
flagyl|1259,1265
,|1265,1266
<EOL>|1266,1267
presenting|1267,1277
with|1278,1282
maroon|1283,1289
colored|1290,1297
GIB|1298,1301
.|1301,1302
HDS|1303,1306
.|1306,1307
HCT|1308,1311
30.7|1312,1316
with|1317,1321
normal|1322,1328
<EOL>|1328,1329
Coag|1329,1333
.|1333,1334
Please|1335,1341
continue|1342,1350
with|1351,1355
supportive|1356,1366
care|1367,1371
with|1372,1376
fluids|1377,1383
and|1384,1387
<EOL>|1387,1388
transfusion|1388,1399
as|1400,1402
needed|1403,1409
.|1409,1410
If|1411,1413
on|1414,1416
-|1416,1417
going|1417,1422
bleeding|1423,1431
or|1432,1434
hemodynamic|1435,1446
<EOL>|1446,1447
changes|1447,1454
,|1454,1455
please|1456,1462
get|1463,1466
CTA|1467,1470
.|1470,1471
If|1472,1474
concern|1475,1482
of|1483,1485
upper|1486,1491
GI|1492,1494
bleeding|1495,1503
,|1503,1504
can|1505,1508
<EOL>|1508,1509
lavage|1509,1515
via|1516,1519
PEG|1520,1523
.|1523,1524
Please|1525,1531
give|1532,1536
PPI|1537,1540
if|1541,1543
positive|1544,1552
.|1552,1553
"|1553,1554
<EOL>|1554,1555
<EOL>|1555,1556
Patient|1556,1563
was|1564,1567
given|1568,1573
1L|1574,1576
normal|1577,1583
saline|1584,1590
and|1591,1594
was|1595,1598
admitted|1599,1607
to|1608,1610
medicine|1611,1619
.|1619,1620
<EOL>|1620,1621
On|1621,1623
arrival|1624,1631
to|1632,1634
the|1635,1638
floor|1639,1644
patient|1645,1652
reported|1653,1661
above|1662,1667
.|1667,1668
Reported|1670,1678
recent|1679,1685
<EOL>|1685,1686
diagnosis|1686,1695
of|1696,1698
L1|1699,1701
compression|1702,1713
fracture|1714,1722
and|1723,1726
intermittent|1727,1739
difficulty|1740,1750
<EOL>|1750,1751
with|1751,1755
flushing|1756,1764
her|1765,1768
PEG|1769,1772
tube|1773,1777
at|1778,1780
home|1781,1785
.|1785,1786
Full|1788,1792
10|1793,1795
point|1796,1801
review|1802,1808
of|1809,1811
<EOL>|1811,1812
systems|1812,1819
positive|1820,1828
where|1829,1834
noted|1835,1840
,|1840,1841
otherwise|1842,1851
negative|1852,1860
.|1860,1861
<EOL>|1862,1863
<EOL>|1863,1864
<EOL>|1865,1866
Sjogrens|1888,1896
<EOL>|1896,1897
Hypothyroidism|1897,1911
<EOL>|1911,1912
h|1912,1913
/|1913,1914
o|1914,1915
severe|1916,1922
Cdiff|1923,1928
<EOL>|1928,1929
Protein|1929,1936
calorie|1937,1944
malnutrition|1945,1957
s|1958,1959
/|1959,1960
p|1960,1961
PEG|1962,1965
<EOL>|1965,1966
Osteoporosis|1966,1978
s|1979,1980
/|1980,1981
p|1981,1982
L1|1983,1985
compression|1986,1997
fracture|1998,2006
<EOL>|2006,2007
Depression|2007,2017
<EOL>|2017,2018
Hemorrhoids|2018,2029
<EOL>|2029,2030
Normocytic|2030,2040
anemia|2041,2047
<EOL>|2048,2049
Bronchiectasis|2049,2063
<EOL>|2064,2065
h|2065,2066
/|2066,2067
o|2067,2068
Shingles|2069,2077
<EOL>|2078,2079
Dementia|2079,2087
(|2088,2089
_|2089,2090
_|2090,2091
_|2091,2092
_|2093,2094
_|2094,2095
_|2095,2096
<EOL>|2097,2098
Mitral|2098,2104
regurgitation|2105,2118
<EOL>|2120,2121
<EOL>|2122,2123
:|2137,2138
<EOL>|2138,2139
_|2139,2140
_|2140,2141
_|2141,2142
<EOL>|2142,2143
:|2157,2158
<EOL>|2158,2159
Has|2159,2162
2|2163,2164
children|2165,2173
.|2173,2174
Father|2176,2182
had|2183,2186
hemorrhoids|2187,2198
.|2198,2199
No|2201,2203
history|2204,2211
of|2212,2214
cancer|2215,2221
,|2221,2222
<EOL>|2222,2223
GI|2223,2225
bleeding|2226,2234
.|2234,2235
<EOL>|2237,2238
<EOL>|2239,2240
ADMISSION|2255,2264
<EOL>|2264,2265
VS|2265,2267
:|2267,2268
187|2269,2272
-|2272,2273
106|2273,2276
(|2277,2278
128|2278,2281
/|2281,2282
78|2282,2284
on|2285,2287
recheck|2288,2295
)|2295,2296
112|2297,2300
16|2301,2303
96|2304,2306
%|2306,2307
RA|2307,2309
<EOL>|2309,2310
Gen|2310,2313
-|2314,2315
supine|2316,2322
in|2323,2325
bed|2326,2329
,|2329,2330
comfortable|2331,2342
,|2342,2343
pale|2344,2348
<EOL>|2348,2349
Eyes|2349,2353
-|2354,2355
EOMI|2356,2360
<EOL>|2360,2361
ENT|2361,2364
-|2365,2366
OP|2367,2369
clear|2370,2375
,|2375,2376
MMM|2377,2380
<EOL>|2380,2381
Heart|2381,2386
-|2387,2388
regularly|2389,2398
tachycardic|2399,2410
;|2410,2411
II|2412,2414
/|2414,2415
VI|2415,2417
systolic|2418,2426
murmur|2427,2433
loudest|2434,2441
at|2442,2444
<EOL>|2444,2445
axilla|2445,2451
;|2451,2452
<EOL>|2453,2454
Lungs|2454,2459
-|2460,2461
CTA|2462,2465
bilaterally|2466,2477
<EOL>|2477,2478
Abd|2478,2481
-|2482,2483
soft|2484,2488
nontender|2489,2498
,|2498,2499
normoactive|2500,2511
bowel|2512,2517
sounds|2518,2524
;|2524,2525
PEG|2526,2529
in|2530,2532
place|2533,2538
<EOL>|2538,2539
Rectum|2539,2545
-|2546,2547
dark|2548,2552
maroon|2553,2559
blood|2560,2565
in|2566,2568
vault|2569,2574
,|2574,2575
no|2576,2578
large|2579,2584
hemorrhoids|2585,2596
<EOL>|2596,2597
palpated|2597,2605
<EOL>|2605,2606
Ext|2606,2609
-|2610,2611
trace|2612,2617
edema|2618,2623
to|2624,2626
mid-shin|2627,2635
<EOL>|2635,2636
Skin|2636,2640
-|2641,2642
+|2643,2644
pale|2644,2648
;|2648,2649
no|2650,2652
rashes|2653,2659
<EOL>|2659,2660
Vasc|2660,2664
-|2665,2666
2|2667,2668
+|2668,2669
DP|2670,2672
/|2672,2673
radial|2673,2679
pulses|2680,2686
<EOL>|2686,2687
Neuro|2687,2692
-|2693,2694
AOx2|2695,2699
-|2699,2700
3|2700,2701
(|2702,2703
full|2703,2707
name|2708,2712
,|2712,2713
_|2714,2715
_|2715,2716
_|2716,2717
"|2717,2718
,|2718,2719
_|2720,2721
_|2721,2722
_|2722,2723
,|2723,2724
<EOL>|2724,2725
moving|2725,2731
all|2732,2735
extremities|2736,2747
<EOL>|2747,2748
Psych|2748,2753
-|2754,2755
appropriate|2756,2767
<EOL>|2767,2768
<EOL>|2768,2769
DISCHARGE|2769,2778
<EOL>|2778,2779
VS|2779,2781
:|2781,2782
98.1|2783,2787
135|2788,2791
/|2791,2792
64|2792,2794
103|2795,2798
20|2799,2801
95|2802,2804
%|2804,2805
RA|2805,2807
<EOL>|2807,2808
Gen|2808,2811
-|2812,2813
supine|2814,2820
in|2821,2823
bed|2824,2827
,|2827,2828
comfortable|2829,2840
appearing|2841,2850
<EOL>|2850,2851
Eyes|2851,2855
-|2856,2857
EOMI|2858,2862
<EOL>|2862,2863
ENT|2863,2866
-|2867,2868
OP|2869,2871
clear|2872,2877
,|2877,2878
MMM|2879,2882
<EOL>|2882,2883
Heart|2883,2888
-|2889,2890
RRR|2891,2894
,|2894,2895
II|2896,2898
/|2898,2899
VI|2899,2901
systolic|2902,2910
murmur|2911,2917
loudest|2918,2925
at|2926,2928
axilla|2929,2935
;|2935,2936
<EOL>|2937,2938
Lungs|2938,2943
-|2944,2945
CTA|2946,2949
bilaterally|2950,2961
,|2961,2962
unchanged|2963,2972
from|2973,2977
day|2978,2981
prior|2982,2987
<EOL>|2987,2988
Abd|2988,2991
-|2992,2993
soft|2994,2998
nontender|2999,3008
,|3008,3009
normoactive|3010,3021
bowel|3022,3027
sounds|3028,3034
;|3034,3035
PEG|3036,3039
in|3040,3042
place|3043,3048
;|3048,3049
<EOL>|3050,3051
unchanged|3051,3060
from|3061,3065
yesterday|3066,3075
<EOL>|3076,3077
Ext|3077,3080
-|3081,3082
no|3083,3085
edema|3086,3091
<EOL>|3092,3093
Skin|3093,3097
-|3098,3099
no|3100,3102
rashes|3103,3109
<EOL>|3109,3110
Vasc|3110,3114
-|3115,3116
2|3117,3118
+|3118,3119
DP|3120,3122
/|3122,3123
radial|3123,3129
pulses|3130,3136
<EOL>|3136,3137
Neuro|3137,3142
-|3143,3144
AOx3|3145,3149
(|3150,3151
full|3151,3155
name|3156,3160
,|3160,3161
_|3162,3163
_|3163,3164
_|3164,3165
,|3165,3166
_|3167,3168
_|3168,3169
_|3169,3170
,|3170,3171
<EOL>|3172,3173
moving|3173,3179
all|3180,3183
extremities|3184,3195
<EOL>|3195,3196
Psych|3196,3201
-|3202,3203
appropriate|3204,3215
<EOL>|3215,3216
<EOL>|3217,3218
Pertinent|3218,3227
Results|3228,3235
:|3235,3236
<EOL>|3236,3237
ADMISSION|3237,3246
<EOL>|3246,3247
_|3247,3248
_|3248,3249
_|3249,3250
10|3251,3253
:|3253,3254
37AM|3254,3258
BLOOD|3259,3264
WBC|3265,3268
-|3268,3269
10|3269,3271
.|3271,3272
1|3272,3273
*|3273,3274
RBC|3275,3278
-|3278,3279
3|3279,3280
.|3280,3281
15|3281,3283
*|3283,3284
Hgb|3285,3288
-|3288,3289
9|3289,3290
.|3290,3291
8|3291,3292
*|3292,3293
Hct|3294,3297
-|3297,3298
30|3298,3300
.|3300,3301
7|3301,3302
*|3302,3303
<EOL>|3304,3305
MCV|3305,3308
-|3308,3309
98|3309,3311
MCH|3312,3315
-|3315,3316
31.1|3316,3320
MCHC|3321,3325
-|3325,3326
31|3326,3328
.|3328,3329
9|3329,3330
*|3330,3331
RDW|3332,3335
-|3335,3336
13.6|3336,3340
RDWSD|3341,3346
-|3346,3347
48|3347,3349
.|3349,3350
4|3350,3351
*|3351,3352
Plt|3353,3356
_|3357,3358
_|3358,3359
_|3359,3360
<EOL>|3360,3361
_|3361,3362
_|3362,3363
_|3363,3364
10|3365,3367
:|3367,3368
37AM|3368,3372
BLOOD|3373,3378
Glucose|3379,3386
-|3386,3387
96|3387,3389
UreaN|3390,3395
-|3395,3396
27|3396,3398
*|3398,3399
Creat|3400,3405
-|3405,3406
0.6|3406,3409
Na|3410,3412
-|3412,3413
136|3413,3416
<EOL>|3417,3418
K|3418,3419
-|3419,3420
4.4|3420,3423
Cl|3424,3426
-|3426,3427
97|3427,3429
HCO3|3430,3434
-|3434,3435
30|3435,3437
AnGap|3438,3443
-|3443,3444
13|3444,3446
<EOL>|3446,3447
_|3447,3448
_|3448,3449
_|3449,3450
06|3451,3453
:|3453,3454
00AM|3454,3458
BLOOD|3459,3464
ALT|3465,3468
-|3468,3469
12|3469,3471
AST|3472,3475
-|3475,3476
19|3476,3478
AlkPhos|3479,3486
-|3486,3487
81|3487,3489
TotBili|3490,3497
-|3497,3498
0.3|3498,3501
<EOL>|3501,3502
<EOL>|3502,3503
DISCHARGE|3503,3512
<EOL>|3512,3513
_|3513,3514
_|3514,3515
_|3515,3516
06|3517,3519
:|3519,3520
20AM|3520,3524
BLOOD|3525,3530
WBC|3531,3534
-|3534,3535
8.9|3535,3538
RBC|3539,3542
-|3542,3543
3|3543,3544
.|3544,3545
35|3545,3547
*|3547,3548
Hgb|3549,3552
-|3552,3553
10|3553,3555
.|3555,3556
5|3556,3557
*|3557,3558
Hct|3559,3562
-|3562,3563
32|3563,3565
.|3565,3566
7|3566,3567
*|3567,3568
<EOL>|3569,3570
MCV|3570,3573
-|3573,3574
98|3574,3576
MCH|3577,3580
-|3580,3581
31.3|3581,3585
MCHC|3586,3590
-|3590,3591
32.1|3591,3595
RDW|3596,3599
-|3599,3600
13.4|3600,3604
RDWSD|3605,3610
-|3610,3611
47|3611,3613
.|3613,3614
7|3614,3615
*|3615,3616
Plt|3617,3620
_|3621,3622
_|3622,3623
_|3623,3624
<EOL>|3624,3625
_|3625,3626
_|3626,3627
_|3627,3628
06|3629,3631
:|3631,3632
20AM|3632,3636
BLOOD|3637,3642
Glucose|3643,3650
-|3650,3651
106|3651,3654
*|3654,3655
UreaN|3656,3661
-|3661,3662
18|3662,3664
Creat|3665,3670
-|3670,3671
0.7|3671,3674
Na|3675,3677
-|3677,3678
137|3678,3681
<EOL>|3682,3683
K|3683,3684
-|3684,3685
3.8|3685,3688
Cl|3689,3691
-|3691,3692
100|3692,3695
HCO3|3696,3700
-|3700,3701
28|3701,3703
AnGap|3704,3709
-|3709,3710
13|3710,3712
<EOL>|3712,3713
<EOL>|3713,3714
Flexible|3714,3722
Sigmoidoscopy|3723,3736
-|3737,3738
_|3739,3740
_|3740,3741
_|3741,3742
<EOL>|3742,3743
Mucosa|3743,3749
:|3749,3750
Normal|3751,3757
mucosa|3758,3764
was|3765,3768
noted|3769,3774
in|3775,3777
the|3778,3781
rectum|3782,3788
and|3789,3792
sigmoid|3793,3800
colon|3801,3806
.|3806,3807
<EOL>|3808,3809
<EOL>|3810,3811
Other|3811,3816
No|3817,3819
bleeding|3820,3828
sources|3829,3836
or|3837,3839
blood|3840,3845
identified|3846,3856
,|3856,3857
though|3858,3864
extent|3865,3871
of|3872,3874
<EOL>|3875,3876
sigmoid|3876,3883
colon|3884,3889
evaluated|3890,3899
was|3900,3903
limited|3904,3911
by|3912,3914
poor|3915,3919
prep|3920,3924
.|3924,3925
<EOL>|3927,3928
Impression|3928,3938
:|3938,3939
Normal|3940,3946
mucosa|3947,3953
in|3954,3956
the|3957,3960
rectum|3961,3967
and|3968,3971
sigmoid|3972,3979
colon|3980,3985
<EOL>|3985,3986
No|3986,3988
bleeding|3989,3997
sources|3998,4005
or|4006,4008
blood|4009,4014
identified|4015,4025
,|4025,4026
though|4027,4033
extent|4034,4040
of|4041,4043
<EOL>|4044,4045
sigmoid|4045,4052
colon|4053,4058
evaluated|4059,4068
was|4069,4072
limited|4073,4080
by|4081,4083
poor|4084,4088
prep|4089,4093
.|4093,4094
<EOL>|4094,4095
Otherwise|4095,4104
normal|4105,4111
sigmoidoscopy|4112,4125
to|4126,4128
sigmoid|4129,4136
colon|4137,4142
at|4143,4145
25|4146,4148
cm|4149,4151
<EOL>|4152,4153
Recommendations|4153,4168
:|4168,4169
If|4170,4172
bleeding|4173,4181
recurs|4182,4188
,|4188,4189
would|4190,4195
recommend|4196,4205
full|4206,4210
<EOL>|4211,4212
colonoscopy|4212,4223
with|4224,4228
prep|4229,4233
.|4233,4234
<EOL>|4235,4236
<EOL>|4236,4237
<EOL>|4238,4239
This|4262,4266
is|4267,4269
an|4270,4272
_|4273,4274
_|4274,4275
_|4275,4276
year|4277,4281
old|4282,4285
female|4286,4292
with|4293,4297
past|4298,4302
medical|4303,4310
history|4311,4318
of|4319,4321
<EOL>|4322,4323
sjogrens|4323,4331
,|4331,4332
hemorrhoids|4333,4344
,|4344,4345
prior|4346,4351
cdiff|4352,4357
infection|4358,4367
,|4367,4368
admitted|4369,4377
_|4378,4379
_|4379,4380
_|4380,4381
<EOL>|4382,4383
with|4383,4387
bright|4388,4394
red|4395,4398
blood|4399,4404
per|4405,4408
rectum|4409,4415
thought|4416,4423
to|4424,4426
be|4427,4429
acute|4430,4435
lower|4436,4441
GI|4442,4444
<EOL>|4445,4446
bleed|4446,4451
,|4451,4452
subsequently|4453,4465
stabilizing|4466,4477
without|4478,4485
intervention|4486,4498
,|4498,4499
status|4500,4506
<EOL>|4507,4508
post|4508,4512
flexible|4513,4521
sigmoidoscopy|4522,4535
without|4536,4543
identifiable|4544,4556
source|4557,4563
,|4563,4564
<EOL>|4565,4566
remaining|4566,4575
stable|4576,4582
x|4583,4584
greater|4585,4592
than|4593,4597
4|4598,4599
days|4600,4604
,|4604,4605
able|4606,4610
to|4611,4613
be|4614,4616
discharged|4617,4627
to|4628,4630
<EOL>|4631,4632
rehab|4632,4637
facility|4638,4646
.|4646,4647
<EOL>|4647,4648
<EOL>|4648,4649
#|4649,4650
Acute|4651,4656
GI|4657,4659
Bleed|4660,4665
NOS|4666,4669
-|4670,4671
Patient|4672,4679
presented|4680,4689
with|4690,4694
acute|4695,4700
episode|4701,4708
of|4709,4711
<EOL>|4712,4713
BRBPR|4713,4718
concerning|4719,4729
for|4730,4733
lower|4734,4739
GI|4740,4742
source|4743,4749
.|4749,4750
Patient|4752,4759
subsequently|4760,4772
<EOL>|4773,4774
monitored|4774,4783
without|4784,4791
new|4792,4795
or|4796,4798
worsening|4799,4808
anemia|4809,4815
.|4815,4816
After|4818,4823
discussion|4824,4834
<EOL>|4835,4836
with|4836,4840
family|4841,4847
and|4848,4851
patient|4852,4859
regarding|4860,4869
whether|4870,4877
or|4878,4880
not|4881,4884
to|4885,4887
further|4888,4895
<EOL>|4896,4897
workup|4897,4903
,|4903,4904
they|4905,4909
opted|4910,4915
for|4916,4919
flexible|4920,4928
sigmoidoscopy|4929,4942
(|4943,4944
felt|4944,4948
colonoscopy|4949,4960
<EOL>|4961,4962
might|4962,4967
be|4968,4970
too|4971,4974
invasive|4975,4983
)|4983,4984
.|4984,4985
Patient|4987,4994
underwent|4995,5004
aborted|5005,5012
flexible|5013,5021
<EOL>|5022,5023
sigmoidoscopy|5023,5036
on|5037,5039
_|5040,5041
_|5041,5042
_|5042,5043
due|5044,5047
to|5048,5050
pressence|5051,5060
of|5061,5063
copious|5064,5071
stool|5072,5077
in|5078,5080
<EOL>|5081,5082
rectal|5082,5088
vault|5089,5094
,|5094,5095
and|5096,5099
then|5100,5104
underwent|5105,5114
successful|5115,5125
flexible|5126,5134
<EOL>|5135,5136
sigmoidoscopy|5136,5149
on|5150,5152
_|5153,5154
_|5154,5155
_|5155,5156
without|5157,5164
identifiable|5165,5177
source|5178,5184
for|5185,5188
her|5189,5192
<EOL>|5193,5194
bleeding|5194,5202
.|5202,5203
From|5205,5209
admission|5210,5219
Hgb|5220,5223
9.8|5224,5227
,|5227,5228
discharge|5229,5238
hemoglobin|5239,5249
was|5250,5253
<EOL>|5254,5255
10.5|5255,5259
.|5259,5260
Per|5262,5265
GI|5266,5268
,|5268,5269
could|5270,5275
consider|5276,5284
outpatient|5285,5295
colonoscopy|5296,5307
if|5308,5310
<EOL>|5311,5312
consistent|5312,5322
with|5323,5327
patient|5328,5335
's|5335,5337
wishes|5338,5344
.|5344,5345
<EOL>|5347,5348
<EOL>|5348,5349
#|5349,5350
Osteoporosis|5351,5363
/|5364,5365
chronic|5366,5373
L1|5374,5376
compression|5377,5388
fracture|5389,5397
/|5398,5399
<EOL>|5400,5401
deconditioning|5401,5415
-|5416,5417
patient|5418,5425
with|5426,5430
recent|5431,5437
L1|5438,5440
compression|5441,5452
fracture|5453,5461
as|5462,5464
<EOL>|5465,5466
outpatient|5466,5476
prior|5477,5482
to|5483,5485
admission|5486,5495
;|5495,5496
patient|5497,5504
noted|5505,5510
to|5511,5513
be|5514,5516
significantly|5517,5530
<EOL>|5531,5532
deconditioned|5532,5545
this|5546,5550
admission|5551,5560
,|5560,5561
requiring|5562,5571
assistance|5572,5582
with|5583,5587
ADLs|5588,5592
;|5592,5593
<EOL>|5594,5595
patient|5595,5602
seen|5603,5607
by|5608,5610
_|5611,5612
_|5612,5613
_|5613,5614
and|5615,5618
recommended|5619,5630
for|5631,5634
rehab|5635,5640
.|5640,5641
Continued|5643,5652
home|5653,5657
<EOL>|5658,5659
Calcium|5659,5666
500|5667,5670
+|5671,5672
vitamin|5673,5680
D|5681,5682
,|5682,5683
calcitonin|5684,5694
.|5694,5695
Placed|5697,5703
on|5704,5706
Tylenol|5707,5714
and|5715,5718
<EOL>|5719,5720
tramadol|5720,5728
for|5729,5732
pain|5733,5737
control|5738,5745
with|5746,5750
good|5751,5755
effect|5756,5762
<EOL>|5763,5764
<EOL>|5764,5765
#|5765,5766
Chronic|5767,5774
Severe|5775,5781
Protein|5782,5789
Calorie|5790,5797
Malnutrition|5798,5810
-|5811,5812
per|5813,5816
discussion|5817,5827
<EOL>|5828,5829
with|5829,5833
family|5834,5840
and|5841,5844
review|5845,5851
of|5852,5854
chart|5855,5860
,|5860,5861
patient|5862,5869
has|5870,5873
lost|5874,5878
weight|5879,5885
despite|5886,5893
<EOL>|5894,5895
PEG|5895,5898
placement|5899,5908
and|5909,5912
bolus|5913,5918
tube|5919,5923
feeds|5924,5929
(|5930,5931
has|5931,5934
had|5935,5938
difficulty|5939,5949
<EOL>|5950,5951
maintaining|5951,5962
PO|5963,5965
intake|5966,5972
due|5973,5976
to|5977,5979
her|5980,5983
Sjogrens|5984,5992
)|5992,5993
.|5993,5994
At|5996,5998
home|5999,6003
patient|6004,6011
has|6012,6015
<EOL>|6016,6017
not|6017,6020
be|6021,6023
using|6024,6029
full|6030,6034
recommended|6035,6046
2|6047,6048
cans|6049,6053
of|6054,6056
Nutren|6057,6063
2.0|6064,6067
,|6067,6068
500|6069,6072
<EOL>|6073,6074
Cal|6074,6077
/|6077,6078
250ml|6078,6083
BID|6084,6087
.|6087,6088
Here|6090,6094
patient|6095,6102
seen|6103,6107
by|6108,6110
nutrition|6111,6120
,|6120,6121
continued|6122,6131
on|6132,6134
<EOL>|6135,6136
above|6136,6141
2|6142,6143
cans|6144,6148
,|6148,6149
and|6150,6153
was|6154,6157
given|6158,6163
oral|6164,6168
supplementation|6169,6184
with|6185,6189
her|6190,6193
PO|6194,6196
<EOL>|6197,6198
meals|6198,6203
as|6204,6206
well|6207,6211
.|6211,6212
<EOL>|6215,6216
<EOL>|6216,6217
#|6217,6218
Depression|6219,6229
-|6230,6231
continued|6232,6241
home|6242,6246
BuPROPion|6247,6256
and|6257,6260
mirtazapine|6261,6272
<EOL>|6273,6274
<EOL>|6274,6275
#|6275,6276
Hypothryoidism|6277,6291
-|6292,6293
continued|6294,6303
levothyroxine|6304,6317
<EOL>|6318,6319
<EOL>|6319,6320
Transitional|6320,6332
Issues|6333,6339
<EOL>|6339,6340
-|6340,6341
Code|6342,6346
status|6347,6353
-|6354,6355
DNR|6356,6359
/|6359,6360
DNI|6360,6363
<EOL>|6363,6364
-|6364,6365
Discharged|6366,6376
to|6377,6379
rehab|6380,6385
<EOL>|6385,6386
-|6386,6387
No|6388,6390
source|6391,6397
for|6398,6401
bleeding|6402,6410
identified|6411,6421
this|6422,6426
admission|6427,6436
;|6436,6437
can|6438,6441
consider|6442,6450
<EOL>|6451,6452
future|6452,6458
colonoscopy|6459,6470
to|6471,6473
look|6474,6478
for|6479,6482
source|6483,6489
of|6490,6492
bleeding|6493,6501
,|6501,6502
but|6503,6506
would|6507,6512
<EOL>|6513,6514
first|6514,6519
discuss|6520,6527
if|6528,6530
consistent|6531,6541
with|6542,6546
patient|6547,6554
's|6554,6556
goals|6557,6562
of|6563,6565
care|6566,6570
<EOL>|6570,6571
-|6571,6572
Would|6573,6578
consider|6579,6587
encouragement|6588,6601
of|6602,6604
PO|6605,6607
intake|6608,6614
and|6615,6618
PEG|6619,6622
-|6622,6623
tube|6623,6627
<EOL>|6628,6629
supplementation|6629,6644
given|6645,6650
her|6651,6654
malnutrition|6655,6667
<EOL>|6668,6669
<EOL>|6670,6671
Medications|6671,6682
on|6683,6685
Admission|6686,6695
:|6695,6696
<EOL>|6696,6697
The|6697,6700
Preadmission|6701,6713
Medication|6714,6724
list|6725,6729
is|6730,6732
accurate|6733,6741
and|6742,6745
complete|6746,6754
.|6754,6755
<EOL>|6755,6756
1.|6756,6758
BuPROPion|6759,6768
XL|6769,6771
(|6772,6773
Once|6773,6777
Daily|6778,6783
)|6783,6784
150|6785,6788
mg|6789,6791
PO|6792,6794
DAILY|6795,6800
<EOL>|6801,6802
2|6802,6803
.|6803,6804
Calcium|6805,6812
500|6813,6816
+|6817,6818
D|6819,6820
(|6821,6822
calcium|6822,6829
carbonate|6830,6839
-|6839,6840
vitamin|6840,6847
D3|6848,6850
)|6850,6851
500|6852,6855
<EOL>|6856,6857
mg|6857,6859
(|6859,6860
1,250|6860,6865
mg|6865,6867
)|6867,6868
-|6869,6870
400|6870,6873
unit|6874,6878
oral|6879,6883
DAILY|6884,6889
<EOL>|6890,6891
3.|6891,6893
Levothyroxine|6894,6907
Sodium|6908,6914
75|6915,6917
mcg|6918,6921
PO|6922,6924
DAILY|6925,6930
<EOL>|6931,6932
4.|6932,6934
Mirtazapine|6935,6946
30|6947,6949
mg|6950,6952
PO|6953,6955
QHS|6956,6959
<EOL>|6960,6961
5.|6961,6963
TraMADol|6964,6972
50|6973,6975
mg|6976,6978
PO|6979,6981
BID|6982,6985
:|6985,6986
PRN|6986,6989
back|6990,6994
pain|6995,6999
<EOL>|7000,7001
6.|7001,7003
Acetaminophen|7004,7017
500|7018,7021
mg|7022,7024
PO|7025,7027
Q6H|7028,7031
:|7031,7032
PRN|7032,7035
back|7036,7040
pain|7041,7045
<EOL>|7046,7047
7.|7047,7049
Alendronate|7050,7061
Sodium|7062,7068
70|7069,7071
mg|7072,7074
PO|7075,7077
QSUN|7078,7082
<EOL>|7083,7084
8.|7084,7086
Calcitonin|7087,7097
Salmon|7098,7104
200|7105,7108
UNIT|7109,7113
NAS|7114,7117
DAILY|7118,7123
<EOL>|7124,7125
9.|7125,7127
Multivitamins|7128,7141
1|7142,7143
TAB|7144,7147
PO|7148,7150
DAILY|7151,7156
<EOL>|7157,7158
10.|7158,7161
TraMADol|7162,7170
100|7171,7174
mg|7175,7177
PO|7178,7180
QHS|7181,7184
:|7184,7185
PRN|7185,7188
back|7189,7193
pain|7194,7198
<EOL>|7199,7200
11|7200,7202
.|7202,7203
Artificial|7204,7214
Tears|7215,7220
_|7221,7222
_|7222,7223
_|7223,7224
DROP|7225,7229
BOTH|7230,7234
EYES|7235,7239
QID|7240,7243
<EOL>|7244,7245
<EOL>|7245,7246
<EOL>|7247,7248
Discharge|7248,7257
Medications|7258,7269
:|7269,7270
<EOL>|7270,7271
1.|7271,7273
Acetaminophen|7274,7287
1000|7288,7292
mg|7293,7295
PO|7296,7298
Q8H|7299,7302
:|7302,7303
PRN|7303,7306
pain|7307,7311
<EOL>|7312,7313
2.|7313,7315
BuPROPion|7316,7325
XL|7326,7328
(|7329,7330
Once|7330,7334
Daily|7335,7340
)|7340,7341
150|7342,7345
mg|7346,7348
PO|7349,7351
DAILY|7352,7357
<EOL>|7358,7359
3.|7359,7361
Calcitonin|7362,7372
Salmon|7373,7379
200|7380,7383
UNIT|7384,7388
NAS|7389,7392
DAILY|7393,7398
<EOL>|7399,7400
4.|7400,7402
Levothyroxine|7403,7416
Sodium|7417,7423
75|7424,7426
mcg|7427,7430
PO|7431,7433
DAILY|7434,7439
<EOL>|7440,7441
5.|7441,7443
Mirtazapine|7444,7455
30|7456,7458
mg|7459,7461
PO|7462,7464
QHS|7465,7468
<EOL>|7469,7470
6.|7470,7472
Multivitamins|7473,7486
1|7487,7488
TAB|7489,7492
PO|7493,7495
DAILY|7496,7501
<EOL>|7502,7503
7.|7503,7505
TraMADol|7506,7514
50|7515,7517
mg|7518,7520
PO|7521,7523
BID|7524,7527
:|7527,7528
PRN|7528,7531
back|7532,7536
pain|7537,7541
<EOL>|7542,7543
8.|7543,7545
Alendronate|7546,7557
Sodium|7558,7564
70|7565,7567
mg|7568,7570
PO|7571,7573
QSUN|7574,7578
<EOL>|7579,7580
9.|7580,7582
Calcium|7583,7590
500|7591,7594
+|7595,7596
D|7597,7598
(|7599,7600
calcium|7600,7607
carbonate|7608,7617
-|7617,7618
vitamin|7618,7625
D3|7626,7628
)|7628,7629
500|7630,7633
<EOL>|7634,7635
mg|7635,7637
(|7637,7638
1,250|7638,7643
mg|7643,7645
)|7645,7646
-|7647,7648
400|7648,7651
unit|7652,7656
oral|7657,7661
DAILY|7662,7667
<EOL>|7668,7669
10.|7669,7672
TraMADol|7673,7681
100|7682,7685
mg|7686,7688
PO|7689,7691
QHS|7692,7695
:|7695,7696
PRN|7696,7699
back|7700,7704
pain|7705,7709
<EOL>|7710,7711
11|7711,7713
.|7713,7714
Artificial|7715,7725
Tears|7726,7731
_|7732,7733
_|7733,7734
_|7734,7735
DROP|7736,7740
BOTH|7741,7745
EYES|7746,7750
QID|7751,7754
<EOL>|7755,7756
<EOL>|7756,7757
<EOL>|7758,7759
Discharge|7759,7768
Disposition|7769,7780
:|7780,7781
<EOL>|7781,7782
Extended|7782,7790
Care|7791,7795
<EOL>|7795,7796
<EOL>|7797,7798
Facility|7798,7806
:|7806,7807
<EOL>|7807,7808
_|7808,7809
_|7809,7810
_|7810,7811
<EOL>|7811,7812
<EOL>|7813,7814
Discharge|7814,7823
Diagnosis|7824,7833
:|7833,7834
<EOL>|7834,7835
#|7835,7836
Acute|7837,7842
GI|7843,7845
Bleed|7846,7851
NOS|7852,7855
<EOL>|7856,7857
#|7857,7858
Depression|7859,7869
<EOL>|7869,7870
#|7870,7871
Osteoporosis|7872,7884
/|7885,7886
chronic|7887,7894
L1|7895,7897
compression|7898,7909
fracture|7910,7918
<EOL>|7918,7919
#|7919,7920
Hypothryoidism|7921,7935
<EOL>|7935,7936
#|7936,7937
Chronic|7938,7945
Severe|7946,7952
Protein|7953,7960
Calorie|7961,7968
Malnutrition|7969,7981
<EOL>|7981,7982
#|7982,7983
Dementia|7984,7992
<EOL>|7992,7993
<EOL>|7993,7994
<EOL>|7995,7996
Mental|8017,8023
Status|8024,8030
:|8030,8031
Confused|8032,8040
-|8041,8042
sometimes|8043,8052
.|8052,8053
<EOL>|8053,8054
Level|8054,8059
of|8060,8062
Consciousness|8063,8076
:|8076,8077
Alert|8078,8083
and|8084,8087
interactive|8088,8099
.|8099,8100
<EOL>|8100,8101
Activity|8101,8109
Status|8110,8116
:|8116,8117
Ambulatory|8118,8128
-|8129,8130
requires|8131,8139
assistance|8140,8150
or|8151,8153
aid|8154,8157
(|8158,8159
walker|8159,8165
<EOL>|8166,8167
or|8167,8169
cane|8170,8174
)|8174,8175
.|8175,8176
<EOL>|8176,8177
<EOL>|8177,8178
<EOL>|8179,8180
Ms.|8204,8207
_|8208,8209
_|8209,8210
_|8210,8211
:|8211,8212
<EOL>|8213,8214
<EOL>|8214,8215
It|8215,8217
was|8218,8221
a|8222,8223
pleasure|8224,8232
caring|8233,8239
for|8240,8243
you|8244,8247
at|8248,8250
_|8251,8252
_|8252,8253
_|8253,8254
.|8254,8255
You|8257,8260
were|8261,8265
admitted|8266,8274
<EOL>|8275,8276
with|8276,8280
gastrointestinal|8281,8297
bleeding|8298,8306
.|8306,8307
You|8309,8312
were|8313,8317
seen|8318,8322
by|8323,8325
GI|8326,8328
specialists|8329,8340
<EOL>|8341,8342
and|8342,8345
underwent|8346,8355
a|8356,8357
flexible|8358,8366
sigmoidiscopy|8367,8380
without|8381,8388
signs|8389,8394
of|8395,8397
a|8398,8399
source|8400,8406
<EOL>|8407,8408
of|8408,8410
your|8411,8415
bleeding|8416,8424
.|8424,8425
You|8427,8430
were|8431,8435
monitored|8436,8445
and|8446,8449
your|8450,8454
blood|8455,8460
levels|8461,8467
were|8468,8472
<EOL>|8473,8474
stable|8474,8480
.|8480,8481
You|8483,8486
are|8487,8490
now|8491,8494
ready|8495,8500
for|8501,8504
discharge|8505,8514
home|8515,8519
.|8519,8520
<EOL>|8520,8521
<EOL>|8521,8522
In|8522,8524
the|8525,8528
future|8529,8535
you|8536,8539
may|8540,8543
wish|8544,8548
to|8549,8551
consider|8552,8560
a|8561,8562
colonoscopy|8563,8574
to|8575,8577
look|8578,8582
for|8583,8586
<EOL>|8587,8588
the|8588,8591
source|8592,8598
of|8599,8601
your|8602,8606
bleeding|8607,8615
,|8615,8616
especially|8617,8627
if|8628,8630
it|8631,8633
occurs|8634,8640
again|8641,8646
.|8646,8647
You|8649,8652
<EOL>|8653,8654
should|8654,8660
discuss|8661,8668
with|8669,8673
your|8674,8678
family|8679,8685
and|8686,8689
primary|8690,8697
care|8698,8702
doctor|8703,8709
<EOL>|8710,8711
regarding|8711,8720
if|8721,8723
this|8724,8728
is|8729,8731
within|8732,8738
your|8739,8743
goals|8744,8749
of|8750,8752
care|8753,8757
.|8757,8758
<EOL>|8758,8759
<EOL>|8760,8761
Followup|8761,8769
Instructions|8770,8782
:|8782,8783
<EOL>|8783,8784
_|8784,8785
_|8785,8786
_|8786,8787
<EOL>|8787,8788

