 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Procedure|Health Care Activity|SIMPLE_SEGMENT|43,52|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|43,57|false|false|false|C2598112||Admission Date
Finding|Body Substance|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|77,86|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|77,91|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|133,136|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|144,151|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|144,151|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Antibiotic|Allergies|180,189|false|false|false|C0066005;C1314417|INJECTION, MEROPENEM, 100 MG ADMINISTERED;meropenem|meropenem
Drug|Clinical Drug|Allergies|180,189|false|false|false|C0066005;C1314417|INJECTION, MEROPENEM, 100 MG ADMINISTERED;meropenem|meropenem
Drug|Organic Chemical|Allergies|180,189|false|false|false|C0066005;C1314417|INJECTION, MEROPENEM, 100 MG ADMINISTERED;meropenem|meropenem
Finding|Functional Concept|Allergies|192,201|false|false|false|C1999232|Attending (action)|Attending
Finding|Functional Concept|Chief Complaint|227,231|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|Chief Complaint|227,235|false|false|false|C0524471|Left hip region structure|left hip
Finding|Sign or Symptom|Chief Complaint|227,240|false|false|false|C2141922|Pain of left hip joint|left hip pain
Anatomy|Body Part, Organ, or Organ Component|Chief Complaint|232,235|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|hip
Drug|Amino Acid, Peptide, or Protein|Chief Complaint|232,235|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Biologically Active Substance|Chief Complaint|232,235|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Pharmacologic Substance|Chief Complaint|232,235|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Finding|Gene or Genome|Chief Complaint|232,235|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|hip
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|232,235|false|false|false|C1292890|Procedure on hip|hip
Attribute|Clinical Attribute|Chief Complaint|232,240|false|false|false|C1716793||hip pain
Finding|Sign or Symptom|Chief Complaint|232,240|false|false|false|C0019559;C4551516|Hip joint pain;Hip pain|hip pain
Attribute|Clinical Attribute|Chief Complaint|236,240|false|false|false|C2598155||pain
Finding|Functional Concept|Chief Complaint|236,240|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Chief Complaint|236,240|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Classification|Chief Complaint|243,248|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|249,257|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|249,257|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|261,279|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|270,279|false|false|false|C0945766||Procedure
Event|Occupational Activity|Chief Complaint|270,279|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|270,279|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|270,279|false|false|false|C0184661|Interventional procedure|Procedure
Finding|Finding|Chief Complaint|288,297|false|false|false|C0392756|Reduced|reduction
Phenomenon|Natural Phenomenon or Process|Chief Complaint|288,297|false|false|false|C0301630|Reduction (chemical)|reduction
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|288,297|false|false|false|C1293152;C4551656|Reduction procedure;Surgical reduction|reduction
Finding|Functional Concept|Chief Complaint|302,314|false|false|false|C1522243|Percutaneous Route of Drug Administration|percutaneous
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|315,322|false|false|false|C0021885|Intramedullary Nailing|pinning
Finding|Functional Concept|Chief Complaint|324,328|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Chief Complaint|329,336|false|false|false|C0015811|Femur|femoral
Anatomy|Body Part, Organ, or Organ Component|Chief Complaint|329,341|false|false|false|C0015815|Structure of neck of femur|femoral neck
Disorder|Injury or Poisoning|Chief Complaint|329,350|false|false|false|C0015806|Femoral Neck Fractures|femoral neck fracture
Anatomy|Body Location or Region|Chief Complaint|337,341|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|Chief Complaint|337,341|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|Chief Complaint|337,341|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Disorder|Injury or Poisoning|Chief Complaint|337,350|false|false|false|C0262414|Fracture of cervical spine|neck fracture
Disorder|Injury or Poisoning|Chief Complaint|342,350|false|false|false|C0016658|Fracture|fracture
Finding|Idea or Concept|History of Present Illness|427,430|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|History of Present Illness|427,430|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Idea or Concept|History of Present Illness|434,446|false|false|false|C0449450|Presentation|presentation
Finding|Functional Concept|History of Present Illness|469,479|false|false|false|C0443254|mechanical method|mechanical
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|469,479|false|false|false|C0699886|Mechanical Treatments|mechanical
Finding|Finding|History of Present Illness|480,484|false|false|false|C0085639|Falls|fall
Finding|Functional Concept|History of Present Illness|494,498|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|History of Present Illness|499,504|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|History of Present Illness|499,504|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|506,515|false|false|false|C0015385|Limb structure|extremity
Finding|Idea or Concept|History of Present Illness|521,530|false|false|false|C1548167;C1697779|Query Priority - Immediate;immediate - ResponseCode|immediate
Finding|Intellectual Product|History of Present Illness|521,530|false|false|false|C1548167;C1697779|Query Priority - Immediate;immediate - ResponseCode|immediate
Attribute|Clinical Attribute|History of Present Illness|531,535|false|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|531,535|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|531,535|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|History of Present Illness|537,558|false|false|false|C5436357|Inability to ambulate|inability to ambulate
Finding|Finding|History of Present Illness|550,558|false|false|false|C4036205|Ambulate|ambulate
Finding|Body Substance|History of Present Illness|566,573|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|566,573|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|566,573|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|History of Present Illness|598,606|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|History of Present Illness|598,606|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Anatomy|Body Space or Junction|History of Present Illness|611,614|false|false|false|C0262327|rostral sulcus|ROS
Drug|Biologically Active Substance|History of Present Illness|611,614|false|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Drug|Element, Ion, or Isotope|History of Present Illness|611,614|false|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Drug|Organic Chemical|History of Present Illness|611,614|false|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Drug|Pharmacologic Substance|History of Present Illness|611,614|false|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Finding|Gene or Genome|History of Present Illness|611,614|false|false|false|C0812281;C1709820|ROS1 gene;ROS1 wt Allele|ROS
Procedure|Health Care Activity|History of Present Illness|611,614|false|false|false|C0489633|Review of systems (procedure)|ROS
Drug|Biomedical or Dental Material|History of Present Illness|632,640|false|false|false|C0168634|BaseLine dental cement|baseline
Finding|Idea or Concept|History of Present Illness|632,640|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Disorder|Disease or Syndrome|Past Medical History|668,674|false|false|false|C0002871|Anemia|Anemia
Lab|Laboratory or Test Result|Past Medical History|677,699|false|false|false|C0694540|borderline cholesterol|Borderline cholesterol
Drug|Biologically Active Substance|Past Medical History|688,699|false|false|false|C0008377|cholesterol|cholesterol
Drug|Organic Chemical|Past Medical History|688,699|false|false|false|C0008377|cholesterol|cholesterol
Procedure|Laboratory Procedure|Past Medical History|688,699|false|false|false|C0201950|Cholesterol measurement|cholesterol
Finding|Sign or Symptom|Past Medical History|722,732|false|false|false|C0016204|Flatulence|Flatulence
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|735,740|false|false|false|C0018787;C4037974|Chest>Heart;Heart|Heart
Disorder|Neoplastic Process|Past Medical History|735,740|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|Heart
Finding|Sign or Symptom|Past Medical History|735,740|false|false|false|C0795691|HEART PROBLEM|Heart
Finding|Finding|Past Medical History|735,747|false|false|false|C0018808|Heart murmur|Heart Murmur
Finding|Finding|Past Medical History|741,747|false|false|false|C0018808|Heart murmur|Murmur
Disorder|Disease or Syndrome|Past Medical History|750,762|false|false|false|C0020538|Hypertensive disease|Hypertension
Disorder|Disease or Syndrome|Past Medical History|765,779|false|false|false|C0020676|Hypothyroidism|Hypothyroidism
Disorder|Disease or Syndrome|Past Medical History|782,802|false|false|false|C0026266|Mitral Valve Insufficiency|Mitral Regurgitation
Finding|Finding|Past Medical History|789,802|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|Regurgitation
Finding|Sign or Symptom|Past Medical History|789,802|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|Regurgitation
Phenomenon|Biologic Function|Past Medical History|789,802|false|false|false|C0460152|Regurgitation - mechanism|Regurgitation
Disorder|Disease or Syndrome|Past Medical History|805,817|false|false|false|C0029456|Osteoporosis|Osteoporosis
Finding|Finding|Past Medical History|805,817|false|false|false|C2911643|Encounter due to family history of osteoporosis|Osteoporosis
Disorder|Disease or Syndrome|Past Medical History|820,829|false|false|false|C0032285|Pneumonia|Pneumonia
Disorder|Disease or Syndrome|Past Medical History|832,841|false|false|false|C0037199|Sinusitis|Sinusitis
Finding|Conceptual Entity|Family Medical History|896,903|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|896,903|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Family Medical History|896,903|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|896,906|false|false|false|C0262926|Medical History|history of
Finding|Finding|Family Medical History|896,919|false|false|false|C0455527||history of hypertension
Disorder|Disease or Syndrome|Family Medical History|907,919|false|false|false|C0020538|Hypertensive disease|hypertension
Drug|Amino Acid, Peptide, or Protein|Family Medical History|923,933|false|false|false|C3812393|ErbB Receptors|her family
Drug|Enzyme|Family Medical History|923,933|false|false|false|C3812393|ErbB Receptors|her family
Finding|Receptor|Family Medical History|923,933|false|false|false|C3812393|ErbB Receptors|her family
Finding|Classification|Family Medical History|927,933|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|Family Medical History|927,933|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|Family Medical History|927,933|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|Family Medical History|927,933|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|Family Medical History|936,942|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Idea or Concept|Family Medical History|936,942|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Classification|Family Medical History|945,951|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|Family Medical History|945,951|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|Family Medical History|945,951|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|Family Medical History|945,951|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|Family Medical History|959,966|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|959,966|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Family Medical History|959,966|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|959,969|false|false|false|C0262926|Medical History|history of
Disorder|Neoplastic Process|Family Medical History|979,986|false|false|false|C0006826|Malignant Neoplasms|cancers
Finding|Conceptual Entity|Family Medical History|1019,1026|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|1019,1026|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Family Medical History|1019,1026|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|1019,1029|false|false|false|C0262926|Medical History|history of
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1030,1037|false|false|false|C0038351;C3714551;C4266636|Abdomen>Stomach;Stomach;Stomach structure|stomach
Disorder|Disease or Syndrome|Family Medical History|1030,1037|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Disorder|Neoplastic Process|Family Medical History|1030,1037|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Finding|Finding|Family Medical History|1030,1037|false|false|false|C0577027|Stomach problem|stomach
Procedure|Therapeutic or Preventive Procedure|Family Medical History|1030,1037|false|false|false|C0872393|Procedure on stomach|stomach
Disorder|Neoplastic Process|Family Medical History|1030,1044|false|false|false|C0024623;C0699791|Malignant neoplasm of stomach;Stomach Carcinoma|stomach cancer
Disorder|Neoplastic Process|Family Medical History|1038,1044|false|false|false|C0006826|Malignant Neoplasms|cancer
Finding|Conceptual Entity|Family Medical History|1065,1072|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|1065,1072|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Family Medical History|1065,1072|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|1065,1075|false|false|false|C0262926|Medical History|history of
Anatomy|Body Location or Region|Family Medical History|1076,1082|false|false|false|C0031354;C0230069;C3665375|Anterior portion of neck;Pharyngeal structure;Throat|throat
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1076,1082|false|false|false|C0031354;C0230069;C3665375|Anterior portion of neck;Pharyngeal structure;Throat|throat
Drug|Pharmacologic Substance|Family Medical History|1076,1082|false|false|false|C1950455|Throat Homeopathic Medication|throat
Finding|Body Substance|Family Medical History|1076,1082|false|false|false|C1547926;C1550663|Specimen Type - Throat|throat
Finding|Intellectual Product|Family Medical History|1076,1082|false|false|false|C1547926;C1550663|Specimen Type - Throat|throat
Disorder|Neoplastic Process|Family Medical History|1084,1090|false|false|false|C0006826|Malignant Neoplasms|cancer
Finding|Conceptual Entity|Family Medical History|1096,1103|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|1096,1103|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Family Medical History|1096,1103|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|1096,1106|true|false|false|C0262926|Medical History|history of
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1107,1112|false|false|false|C0009368;C4071907|Abdomen+Pelvis>Colon;Colon structure (body structure)|colon
Disorder|Disease or Syndrome|Family Medical History|1107,1112|true|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Disorder|Neoplastic Process|Family Medical History|1107,1112|true|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Finding|Finding|Family Medical History|1107,1112|true|false|false|C0750873|COLON PROBLEM|colon
Disorder|Neoplastic Process|Family Medical History|1107,1120|true|false|false|C0007102|Malignant tumor of colon|colon cancers
Disorder|Neoplastic Process|Family Medical History|1113,1120|true|false|false|C0006826|Malignant Neoplasms|cancers
Finding|Conceptual Entity|Family Medical History|1122,1128|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Idea or Concept|Family Medical History|1122,1128|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Disorder|Disease or Syndrome|Family Medical History|1133,1139|false|false|false|C0038454|Cerebrovascular accident|stroke
Finding|Finding|Family Medical History|1133,1139|false|false|false|C5977286|Stroke (heart beat)|stroke
Finding|Classification|Family Medical History|1145,1151|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|Family Medical History|1145,1151|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|Family Medical History|1145,1151|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|Family Medical History|1145,1151|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|Family Medical History|1160,1166|false|false|false|C1546508|Relationship - Mother|Mother
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1173,1178|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Family Medical History|1173,1178|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Family Medical History|1173,1178|false|false|false|C0795691|HEART PROBLEM|heart
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1173,1184|false|false|false|C0018826;C1305961|Heart Valves|heart valve
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1179,1184|false|false|false|C1186983|Anatomical valve|valve
Procedure|Health Care Activity|General Exam|1216,1225|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Anatomy|Body Part, Organ, or Organ Component|General Exam|1228,1234|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|Pelvis
Anatomy|Body Space or Junction|General Exam|1228,1234|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|Pelvis
Disorder|Neoplastic Process|General Exam|1228,1234|false|false|false|C0153663|Malignant neoplasm of pelvis|Pelvis
Finding|Finding|General Exam|1228,1234|false|false|false|C0812455|Pelvis problem|Pelvis
Finding|Intellectual Product|General Exam|1235,1241|false|false|false|C1547311|Patient Condition Code - Stable|stable
Finding|Functional Concept|General Exam|1260,1271|false|false|false|C0332459;C4551657|Compressed structure|compression
Phenomenon|Natural Phenomenon or Process|General Exam|1260,1271|false|false|false|C0728907|Compression|compression
Procedure|Machine Activity|General Exam|1260,1271|false|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Procedure|Therapeutic or Preventive Procedure|General Exam|1260,1271|false|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Anatomy|Body System|General Exam|1279,1283|false|false|false|C1123023;C4520765|Skin;Skin, Human|skin
Disorder|Disease or Syndrome|General Exam|1279,1283|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Disorder|Neoplastic Process|General Exam|1279,1283|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Finding|Body Substance|General Exam|1279,1283|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Finding|Intellectual Product|General Exam|1279,1283|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Finding|Finding|General Exam|1279,1289|false|false|false|C0574729|Skin clean|skin clean
Event|Activity|General Exam|1284,1289|false|false|false|C1947930|Cleaning (activity)|clean
Finding|Finding|General Exam|1294,1300|false|false|false|C1554187|Gender Status - Intact|intact
Finding|Sign or Symptom|General Exam|1340,1347|false|false|false|C0030193|Pain|painful
Anatomy|Body Location or Region|General Exam|1366,1374|false|false|false|C1548801|Body Site Modifier - External|external
Finding|Functional Concept|General Exam|1366,1374|false|false|false|C0521134|External route|external
Finding|Functional Concept|General Exam|1366,1383|false|false|false|C0231462|External rotation|external rotation
Disorder|Anatomical Abnormality|General Exam|1375,1383|false|false|false|C3669037|Rotation (malposition) (morphologic abnormality)|rotation
Finding|Finding|General Exam|1375,1383|false|false|false|C0035868;C0677597;C2117331|Musculoskeletal rotation;Rotation|rotation
Finding|Functional Concept|General Exam|1375,1383|false|false|false|C0035868;C0677597;C2117331|Musculoskeletal rotation;Rotation|rotation
Anatomy|Body Part, Organ, or Organ Component|General Exam|1391,1394|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|hip
Drug|Amino Acid, Peptide, or Protein|General Exam|1391,1394|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Biologically Active Substance|General Exam|1391,1394|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Pharmacologic Substance|General Exam|1391,1394|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Finding|Gene or Genome|General Exam|1391,1394|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|hip
Procedure|Therapeutic or Preventive Procedure|General Exam|1391,1394|false|false|false|C1292890|Procedure on hip|hip
Anatomy|Body Location or Region|General Exam|1398,1404|false|false|false|C0039866|Thigh structure|Thighs
Anatomy|Body Part, Organ, or Organ Component|General Exam|1409,1412|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Finding|Intellectual Product|General Exam|1413,1425|false|false|false|C1185625|Anatomical compartments|compartments
Phenomenon|Natural Phenomenon or Process|General Exam|1413,1425|false|false|false|C1382196|Compartments [PK]|compartments
Disorder|Disease or Syndrome|General Exam|1426,1430|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Drug|Pharmacologic Substance|General Exam|1443,1448|false|false|false|C0626053|sural|Sural
Attribute|Clinical Attribute|General Exam|1450,1454|false|false|false|C4318566|Deep Resection Margin|Deep
Event|Event|Family Medical History|1517,1521|false|false|false|C0016141|fire disaster|Fire
Finding|Gene or Genome|Family Medical History|1517,1521|false|false|false|C1426107|ADGRE4P gene|Fire
Phenomenon|Human-caused Phenomenon or Process|Family Medical History|1517,1521|false|false|false|C0000912;C0700614;C0702194|Accident caused by unspecified fire;Fire (physical force);Fire as a heat source|Fire
Phenomenon|Natural Phenomenon or Process|Family Medical History|1517,1521|false|false|false|C0000912;C0700614;C0702194|Accident caused by unspecified fire;Fire (physical force);Fire as a heat source|Fire
Phenomenon|Phenomenon or Process|Family Medical History|1517,1521|false|false|false|C0000912;C0700614;C0702194|Accident caused by unspecified fire;Fire (physical force);Fire as a heat source|Fire
Drug|Food|Family Medical History|1537,1543|false|false|false|C5890763||pulses
Finding|Physiologic Function|Family Medical History|1537,1543|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|Family Medical History|1537,1543|false|false|false|C0034107|Pulse taking|pulses
Anatomy|Body Location or Region|Family Medical History|1545,1549|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|Knee
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1545,1549|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|Knee
Anatomy|Body Space or Junction|Family Medical History|1545,1549|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|Knee
Procedure|Diagnostic Procedure|Family Medical History|1545,1549|false|false|false|C0562271|Examination of knee joint|Knee
Finding|Intellectual Product|Family Medical History|1550,1556|false|false|false|C1547311|Patient Condition Code - Stable|stable
Disorder|Anatomical Abnormality|Family Medical History|1570,1576|false|false|false|C0042282|Valgus deformity|valgus
Attribute|Clinical Attribute|Family Medical History|1577,1583|false|false|false|C1718621|W stress|stress
Drug|Organic Chemical|Family Medical History|1577,1583|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|Family Medical History|1577,1583|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Finding|Finding|Family Medical History|1577,1583|false|false|false|C0038435|Stress|stress
Finding|Classification|Family Medical History|1588,1596|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|Negative
Finding|Finding|Family Medical History|1588,1596|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|Negative
Lab|Laboratory or Test Result|Family Medical History|1588,1596|false|false|false|C5237010|Expression Negative|Negative
Disorder|Disease or Syndrome|Family Medical History|1597,1605|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Disorder|Disease or Syndrome|Family Medical History|1607,1616|false|false|false|C0751438|Posterior pituitary disease|posterior
Finding|Finding|Family Medical History|1624,1629|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|Family Medical History|1624,1629|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Body Substance|Family Medical History|1637,1646|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Family Medical History|1637,1646|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Family Medical History|1637,1646|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Family Medical History|1637,1646|false|false|false|C0030685|Patient Discharge|discharge
Disorder|Disease or Syndrome|Family Medical History|1649,1652|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|Family Medical History|1649,1652|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|Family Medical History|1649,1652|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Family Medical History|1649,1652|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|Family Medical History|1649,1652|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Finding|Finding|Family Medical History|1649,1652|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Location or Region|Family Medical History|1660,1668|false|false|false|C2338258|Cranial incision point|INcision
Disorder|Injury or Poisoning|Family Medical History|1660,1668|false|false|false|C0332803|Surgical wound|INcision
Procedure|Therapeutic or Preventive Procedure|Family Medical History|1660,1668|false|false|false|C0184898|Surgical incisions|INcision
Drug|Biomedical or Dental Material|Family Medical History|1670,1678|false|false|false|C1705365|Dressing Dosage Form|dressing
Finding|Daily or Recreational Activity|Family Medical History|1670,1678|false|false|false|C0518459;C1305428|Ability to dress|dressing
Finding|Finding|Family Medical History|1670,1678|false|false|false|C0518459;C1305428|Ability to dress|dressing
Procedure|Health Care Activity|Family Medical History|1670,1678|false|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|dressing
Procedure|Therapeutic or Preventive Procedure|Family Medical History|1670,1678|false|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|dressing
Finding|Finding|Family Medical History|1715,1721|false|false|false|C1554187|Gender Status - Intact|intact
Finding|Finding|Family Medical History|1732,1738|false|false|false|C1554187|Gender Status - Intact|intact
Attribute|Clinical Attribute|Family Medical History|1783,1788|false|false|false|C0232117|Pulse Rate|pulse
Finding|Physiologic Function|Family Medical History|1783,1788|false|false|false|C0391850|Physiologic pulse|pulse
Phenomenon|Phenomenon or Process|Family Medical History|1783,1788|false|false|false|C1947910|Pulse phenomenon|pulse
Procedure|Health Care Activity|Family Medical History|1783,1788|false|false|false|C0034107|Pulse taking|pulse
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1811,1814|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|Hip
Drug|Amino Acid, Peptide, or Protein|Family Medical History|1811,1814|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|Hip
Drug|Biologically Active Substance|Family Medical History|1811,1814|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|Hip
Drug|Pharmacologic Substance|Family Medical History|1811,1814|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|Hip
Finding|Gene or Genome|Family Medical History|1811,1814|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|Hip
Procedure|Therapeutic or Preventive Procedure|Family Medical History|1811,1814|false|false|false|C1292890|Procedure on hip|Hip
Finding|Intellectual Product|Family Medical History|1823,1833|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|Family Medical History|1823,1833|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Disorder|Disease or Syndrome|Family Medical History|1836,1844|false|false|false|C0040456|Impacted tooth|Impacted
Finding|Functional Concept|Family Medical History|1836,1844|false|false|false|C0333125|Impacted|Impacted
Finding|Functional Concept|Family Medical History|1845,1849|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1861,1868|false|false|false|C0015811|Femur|femoral
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1861,1873|false|false|false|C0015815|Structure of neck of femur|femoral neck
Anatomy|Body Location or Region|Family Medical History|1869,1873|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|Family Medical History|1869,1873|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|Family Medical History|1869,1873|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Disorder|Injury or Poisoning|Family Medical History|1875,1883|false|false|false|C0016658|Fracture|fracture
Finding|Idea or Concept|Hospital Course|1944,1949|false|false|false|C0812371|Ortho-|ortho
Disorder|Injury or Poisoning|Hospital Course|1950,1956|false|false|false|C1368081;C3263723;C3714660|Physical trauma;Trauma;Traumatic injury|trauma
Procedure|Health Care Activity|Hospital Course|1950,1956|false|false|false|C0548346|Trauma assessment and care|trauma
Event|Occupational Activity|Hospital Course|1957,1964|false|false|false|C0557854|Services|service
Finding|Idea or Concept|Hospital Course|1957,1964|false|false|false|C3245478|ActInformationPrivacyReason - service|service
Disorder|Anatomical Abnormality|Hospital Course|1986,1992|false|false|false|C0042282|Valgus deformity|valgus
Finding|Functional Concept|Hospital Course|2002,2006|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|2002,2019|false|false|false|C0833290|Neck of left femur|left femoral neck
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|2007,2014|false|false|false|C0015811|Femur|femoral
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|2007,2019|false|false|false|C0015815|Structure of neck of femur|femoral neck
Anatomy|Body Location or Region|Hospital Course|2015,2019|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|Hospital Course|2015,2019|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|Hospital Course|2015,2019|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|2020,2023|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|hip
Drug|Amino Acid, Peptide, or Protein|Hospital Course|2020,2023|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Biologically Active Substance|Hospital Course|2020,2023|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Pharmacologic Substance|Hospital Course|2020,2023|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Finding|Gene or Genome|Hospital Course|2020,2023|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|hip
Procedure|Therapeutic or Preventive Procedure|Hospital Course|2020,2023|false|false|false|C1292890|Procedure on hip|hip
Disorder|Injury or Poisoning|Hospital Course|2020,2032|false|false|false|C0019557;C0149531|Fracture of pelvis;Hip Fractures|hip fracture
Disorder|Injury or Poisoning|Hospital Course|2024,2032|false|false|false|C0016658|Fracture|fracture
Finding|Finding|Hospital Course|2066,2075|false|false|false|C0392756|Reduced|reduction
Phenomenon|Natural Phenomenon or Process|Hospital Course|2066,2075|false|false|false|C0301630|Reduction (chemical)|reduction
Procedure|Therapeutic or Preventive Procedure|Hospital Course|2066,2075|false|false|false|C1293152;C4551656|Reduction procedure;Surgical reduction|reduction
Finding|Functional Concept|Hospital Course|2080,2092|false|false|false|C1522243|Percutaneous Route of Drug Administration|percutaneous
Procedure|Therapeutic or Preventive Procedure|Hospital Course|2094,2101|false|false|false|C0021885|Intramedullary Nailing|pinning
Finding|Functional Concept|Hospital Course|2103,2107|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|2108,2115|false|false|false|C0015811|Femur|femoral
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|2108,2120|false|false|false|C0015815|Structure of neck of femur|femoral neck
Disorder|Injury or Poisoning|Hospital Course|2108,2129|false|false|false|C0015806|Femoral Neck Fractures|femoral neck fracture
Anatomy|Body Location or Region|Hospital Course|2116,2120|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|Hospital Course|2116,2120|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|Hospital Course|2116,2120|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Disorder|Injury or Poisoning|Hospital Course|2116,2129|false|false|false|C0262414|Fracture of cervical spine|neck fracture
Disorder|Injury or Poisoning|Hospital Course|2121,2129|false|false|false|C0016658|Fracture|fracture
Finding|Body Substance|Hospital Course|2153,2160|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|2153,2160|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|2153,2160|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Finding|Hospital Course|2188,2192|false|false|false|C5575035|Well (answer to question)|well
Finding|Finding|Hospital Course|2199,2206|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|Hospital Course|2199,2206|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|Hospital Course|2199,2206|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|Hospital Course|2199,2206|false|false|false|C0543467|Operative Surgical Procedures|surgery
Finding|Pathologic Function|Hospital Course|2219,2230|false|false|false|C0857353|Hypotensive|hypotensive
Finding|Finding|Hospital Course|2236,2244|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Finding|Functional Concept|Hospital Course|2236,2244|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Procedure|Health Care Activity|Hospital Course|2236,2244|false|false|false|C0031809|Physical Examination|physical
Finding|Intellectual Product|Hospital Course|2236,2252|false|false|false|C1547999|Diagnostic Service Section ID - Physical Therapy|physical therapy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|2236,2252|false|false|false|C0949766|Physical therapy|physical therapy
Finding|Finding|Hospital Course|2245,2252|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|Hospital Course|2245,2252|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|2245,2252|false|false|false|C0087111|Therapeutic procedure|therapy
Finding|Daily or Recreational Activity|Hospital Course|2287,2295|false|false|false|C0015259|Exercise|exercise
Procedure|Therapeutic or Preventive Procedure|Hospital Course|2287,2295|false|false|false|C1522704|Exercise Pain Management|exercise
Finding|Body Substance|Hospital Course|2310,2317|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|2310,2317|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|2310,2317|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Finding|Hospital Course|2334,2338|false|false|false|C5575035|Well (answer to question)|well
Finding|Finding|Hospital Course|2357,2365|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Finding|Functional Concept|Hospital Course|2357,2365|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Procedure|Health Care Activity|Hospital Course|2357,2365|false|false|false|C0031809|Physical Examination|physical
Finding|Intellectual Product|Hospital Course|2357,2373|false|false|false|C1547999|Diagnostic Service Section ID - Physical Therapy|physical therapy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|2357,2373|false|false|false|C0949766|Physical therapy|physical therapy
Finding|Finding|Hospital Course|2366,2373|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|Hospital Course|2366,2373|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|2366,2373|false|false|false|C0087111|Therapeutic procedure|therapy
Finding|Body Substance|Hospital Course|2390,2399|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|2390,2399|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|2390,2399|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|2390,2399|false|false|false|C0030685|Patient Discharge|discharge
Procedure|Therapeutic or Preventive Procedure|Hospital Course|2405,2410|false|false|false|C0034991|Rehabilitation therapy|rehab
Finding|Intellectual Product|Hospital Course|2411,2419|false|false|false|C4695111|ADMIN.FACILITY|facility
Finding|Functional Concept|Hospital Course|2422,2428|false|false|false|C0728831|Social|SOcial
Event|Occupational Activity|Hospital Course|2429,2433|false|false|false|C0043227|Work|work
Finding|Finding|Hospital Course|2449,2459|false|false|false|C1299586|Has difficulty doing (qualifier value)|difficulty
Finding|Finding|Hospital Course|2449,2466|false|false|false|C0582154|Difficulty coping|difficulty coping
Finding|Finding|Hospital Course|2460,2466|false|true|false|C0009967;C0517270|Child coping with hospitalization;Coping Behavior|coping
Finding|Individual Behavior|Hospital Course|2460,2466|false|true|false|C0009967;C0517270|Child coping with hospitalization;Coping Behavior|coping
Procedure|Therapeutic or Preventive Procedure|Hospital Course|2460,2466|false|true|false|C2700390;C3502819|COPING - Dental Restorative Procedure;COPING - Fixed Prosthodontics|coping
Finding|Finding|Hospital Course|2472,2481|false|false|false|C0392756;C0442797|Decreasing;Reduced|decreased
Attribute|Clinical Attribute|Hospital Course|2483,2491|false|false|false|C0080078|Range of Motion, Articular|mobility
Finding|Finding|Hospital Course|2483,2491|false|false|false|C0425245|Mobility finding|mobility
Lab|Laboratory or Test Result|Hospital Course|2497,2501|false|false|false|C0587081|Laboratory test finding|labs
Drug|Biologically Active Substance|Hospital Course|2509,2515|false|true|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Element, Ion, or Isotope|Hospital Course|2509,2515|false|true|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Pharmacologic Substance|Hospital Course|2509,2515|false|true|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Finding|Physiologic Function|Hospital Course|2509,2515|false|true|false|C4553025|Sodium metabolic function|sodium
Procedure|Laboratory Procedure|Hospital Course|2509,2515|false|true|false|C0337443|Sodium measurement|sodium
Lab|Laboratory or Test Result|Hospital Course|2509,2521|false|false|false|C0428291|Finding of sodium level|sodium level
Procedure|Laboratory Procedure|Hospital Course|2509,2521|false|false|false|C0337443|Sodium measurement|sodium level
Finding|Finding|Hospital Course|2530,2539|false|false|false|C0442739||unchanged
Procedure|Health Care Activity|Hospital Course|2572,2581|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Attribute|Clinical Attribute|Hospital Course|2597,2609|false|false|false|C3263700||instructions
Finding|Intellectual Product|Hospital Course|2597,2609|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|instructions
Drug|Organic Chemical|Hospital Course|2669,2676|false|false|false|C0728963|Lovenox|lovenox
Drug|Pharmacologic Substance|Hospital Course|2669,2676|false|false|false|C0728963|Lovenox|lovenox
Attribute|Clinical Attribute|Hospital Course|2714,2725|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|2714,2725|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|Hospital Course|2714,2725|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|2714,2738|false|false|false|C1627937|Medications on admission|Medications on Admission
Procedure|Health Care Activity|Hospital Course|2729,2738|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|Hospital Course|2757,2767|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|Hospital Course|2757,2767|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|Hospital Course|2757,2772|false|false|false|C0746470|MEDICATION LIST|Medication list
Finding|Intellectual Product|Hospital Course|2768,2772|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Drug|Organic Chemical|Hospital Course|2789,2797|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|Hospital Course|2789,2797|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|Hospital Course|2789,2797|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Finding|Functional Concept|Hospital Course|2789,2797|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|Hospital Course|2789,2797|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Amino Acid, Peptide, or Protein|Hospital Course|2802,2815|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Hormone|Hospital Course|2802,2815|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Organic Chemical|Hospital Course|2802,2815|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Pharmacologic Substance|Hospital Course|2802,2815|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Amino Acid, Peptide, or Protein|Hospital Course|2802,2822|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Hormone|Hospital Course|2802,2822|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Pharmacologic Substance|Hospital Course|2802,2822|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Biologically Active Substance|Hospital Course|2816,2822|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|2816,2822|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|2816,2822|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Finding|Physiologic Function|Hospital Course|2816,2822|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|2816,2822|false|false|false|C0337443|Sodium measurement|Sodium
Drug|Amino Acid, Peptide, or Protein|Hospital Course|2843,2853|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Pharmacologic Substance|Hospital Course|2843,2853|false|false|false|C0065374|lisinopril|Lisinopril
Disorder|Injury or Poisoning|Hospital Course|2872,2887|false|false|false|C2878629|Poisoning by, adverse effect of and underdosing of methylphenidate|MethylPHENIDATE
Drug|Organic Chemical|Hospital Course|2872,2887|false|false|false|C0025810|methylphenidate|MethylPHENIDATE
Drug|Pharmacologic Substance|Hospital Course|2872,2887|false|false|false|C0025810|methylphenidate|MethylPHENIDATE
Procedure|Laboratory Procedure|Hospital Course|2872,2887|false|false|false|C0524188|Methylphenidate measurement|MethylPHENIDATE
Drug|Organic Chemical|Hospital Course|2889,2896|false|false|false|C0728759|Ritalin|Ritalin
Drug|Pharmacologic Substance|Hospital Course|2889,2896|false|false|false|C0728759|Ritalin|Ritalin
Disorder|Mental or Behavioral Dysfunction|Hospital Course|2908,2911|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|2908,2911|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|2908,2911|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|2908,2911|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|2916,2927|false|false|false|C0049506|mirtazapine|mirtazapine
Drug|Pharmacologic Substance|Hospital Course|2916,2927|false|false|false|C0049506|mirtazapine|mirtazapine
Anatomy|Body Space or Junction|Hospital Course|2934,2938|false|false|false|C0226896|Oral cavity|Oral
Drug|Biomedical or Dental Material|Hospital Course|2934,2938|false|false|false|C1272919|Oral Dosage Form|Oral
Finding|Finding|Hospital Course|2934,2938|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Finding|Functional Concept|Hospital Course|2934,2938|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Finding|Body Substance|Hospital Course|2947,2956|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|2947,2956|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|2947,2956|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|2947,2956|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|2947,2968|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|2957,2968|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|2957,2968|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|Hospital Course|2957,2968|false|false|false|C4284232|Medications|Medications
Drug|Amino Acid, Peptide, or Protein|Hospital Course|2973,2986|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Hormone|Hospital Course|2973,2986|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Organic Chemical|Hospital Course|2973,2986|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Pharmacologic Substance|Hospital Course|2973,2986|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Amino Acid, Peptide, or Protein|Hospital Course|2973,2993|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Hormone|Hospital Course|2973,2993|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Pharmacologic Substance|Hospital Course|2973,2993|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Biologically Active Substance|Hospital Course|2987,2993|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|2987,2993|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|2987,2993|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Finding|Physiologic Function|Hospital Course|2987,2993|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|2987,2993|false|false|false|C0337443|Sodium measurement|Sodium
Drug|Amino Acid, Peptide, or Protein|Hospital Course|3014,3024|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Pharmacologic Substance|Hospital Course|3014,3024|false|false|false|C0065374|lisinopril|Lisinopril
Disorder|Injury or Poisoning|Hospital Course|3043,3058|false|false|false|C2878629|Poisoning by, adverse effect of and underdosing of methylphenidate|MethylPHENIDATE
Drug|Organic Chemical|Hospital Course|3043,3058|false|false|false|C0025810|methylphenidate|MethylPHENIDATE
Drug|Pharmacologic Substance|Hospital Course|3043,3058|false|false|false|C0025810|methylphenidate|MethylPHENIDATE
Procedure|Laboratory Procedure|Hospital Course|3043,3058|false|false|false|C0524188|Methylphenidate measurement|MethylPHENIDATE
Drug|Organic Chemical|Hospital Course|3060,3067|false|false|false|C0728759|Ritalin|Ritalin
Drug|Pharmacologic Substance|Hospital Course|3060,3067|false|false|false|C0728759|Ritalin|Ritalin
Disorder|Mental or Behavioral Dysfunction|Hospital Course|3079,3082|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|3079,3082|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|3079,3082|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|3079,3082|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|3087,3098|false|false|false|C0049506|mirtazapine|mirtazapine
Drug|Pharmacologic Substance|Hospital Course|3087,3098|false|false|false|C0049506|mirtazapine|mirtazapine
Anatomy|Body Space or Junction|Hospital Course|3105,3109|false|false|false|C0226896|Oral cavity|Oral
Drug|Biomedical or Dental Material|Hospital Course|3105,3109|false|false|false|C1272919|Oral Dosage Form|Oral
Finding|Finding|Hospital Course|3105,3109|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Finding|Functional Concept|Hospital Course|3105,3109|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Drug|Organic Chemical|Hospital Course|3118,3131|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Hospital Course|3118,3131|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Procedure|Laboratory Procedure|Hospital Course|3118,3131|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Drug|Element, Ion, or Isotope|Hospital Course|3151,3159|false|false|false|C0002367|aluminum|Aluminum
Drug|Pharmacologic Substance|Hospital Course|3151,3159|false|false|false|C0002367|aluminum|Aluminum
Procedure|Laboratory Procedure|Hospital Course|3151,3159|false|false|false|C0202311|Aluminum measurement|Aluminum
Drug|Biologically Active Substance|Hospital Course|3160,3169|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|Magnesium
Drug|Element, Ion, or Isotope|Hospital Course|3160,3169|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|Magnesium
Drug|Inorganic Chemical|Hospital Course|3160,3169|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|Magnesium
Drug|Pharmacologic Substance|Hospital Course|3160,3169|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|Magnesium
Procedure|Laboratory Procedure|Hospital Course|3160,3169|false|false|false|C0373675|Magnesium measurement|Magnesium
Drug|Organic Chemical|Hospital Course|3178,3189|false|false|false|C0037138|simethicone|Simethicone
Drug|Pharmacologic Substance|Hospital Course|3178,3189|false|false|false|C0037138|simethicone|Simethicone
Finding|Gene or Genome|Hospital Course|3204,3207|false|false|false|C1422467|CIAO3 gene|PRN
Finding|Sign or Symptom|Hospital Course|3209,3218|false|false|false|C0013395|Dyspepsia|Dyspepsia
Drug|Pharmacologic Substance|Hospital Course|3223,3239|false|false|false|C0003921;C2608262;C3853661|Artificial Tears;Lubricant Eye Drops;artificial tears (medication)|Artificial Tears
Finding|Body Substance|Hospital Course|3234,3239|false|false|false|C0039409;C1547924;C1611838|Tears (substance);Tears specimen|Tears
Finding|Intellectual Product|Hospital Course|3234,3239|false|false|false|C0039409;C1547924;C1611838|Tears (substance);Tears specimen|Tears
Drug|Biomedical or Dental Material|Hospital Course|3244,3248|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|Hospital Course|3244,3248|false|false|false|C1705648|Dropping|DROP
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|3249,3258|false|false|false|C0229118|Structure of both eyes|BOTH EYES
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|3254,3258|false|false|false|C0015392|Eye|EYES
Attribute|Clinical Attribute|Hospital Course|3254,3258|false|false|false|C5848506||EYES
Finding|Gene or Genome|Hospital Course|3259,3262|false|false|false|C1422467|CIAO3 gene|PRN
Disorder|Disease or Syndrome|Hospital Course|3263,3271|false|false|false|C0013238;C0022575|Dry Eye Syndromes;Keratoconjunctivitis Sicca|dry eyes
Drug|Pharmacologic Substance|Hospital Course|3263,3271|false|false|false|C0720056|Dry Eyes brand of ocular lubricant|dry eyes
Finding|Sign or Symptom|Hospital Course|3263,3271|false|false|false|C0314719|Dryness of eye|dry eyes
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|3267,3271|false|false|false|C0015392|Eye|eyes
Attribute|Clinical Attribute|Hospital Course|3267,3271|false|false|false|C5848506||eyes
Drug|Amino Acid, Peptide, or Protein|Hospital Course|3276,3283|false|false|false|C0673636|Biotene|Biotene
Drug|Enzyme|Hospital Course|3276,3283|false|false|false|C0673636|Biotene|Biotene
Drug|Pharmacologic Substance|Hospital Course|3276,3283|false|false|false|C0673636|Biotene|Biotene
Drug|Pharmacologic Substance|Hospital Course|3276,3293|false|false|false|C5762022|Biotene Dry Mouth|Biotene Dry Mouth
Disorder|Disease or Syndrome|Hospital Course|3284,3293|false|false|false|C0043352|Xerostomia|Dry Mouth
Anatomy|Body Location or Region|Hospital Course|3288,3293|false|false|false|C0226896;C0230028|Oral cavity;Oral region|Mouth
Anatomy|Body Space or Junction|Hospital Course|3288,3293|false|false|false|C0226896;C0230028|Oral cavity;Oral region|Mouth
Drug|Biomedical or Dental Material|Hospital Course|3288,3299|false|false|false|C0026647|Mouthwash|Mouth Rinse
Finding|Body Substance|Hospital Course|3288,3299|false|false|false|C5849077|Mouth Rinse Specimen|Mouth Rinse
Event|Activity|Hospital Course|3294,3299|false|false|false|C1882955|Rinsing|Rinse
Finding|Functional Concept|Hospital Course|3294,3299|false|false|false|C1701810|Rinse Dosage Form|Rinse
Finding|Body Substance|Hospital Course|3301,3307|false|false|false|C0036087;C0438730;C1546769|Saliva specimen;saliva|saliva
Finding|Intellectual Product|Hospital Course|3301,3307|false|false|false|C0036087;C0438730;C1546769|Saliva specimen;saliva|saliva
Event|Activity|Hospital Course|3308,3320|false|false|false|C1706204|Substitution - change|substitution
Finding|Idea or Concept|Hospital Course|3308,3320|false|false|false|C1555721|Substitution - ActClass|substitution
Finding|Functional Concept|Hospital Course|3336,3347|false|false|false|C0870325;C1547755;C1947919;C2347934;C4048755|Application Document;Apply;Computer Application;HL7 Version 2.5 - Application;Regulatory Application|application
Finding|Idea or Concept|Hospital Course|3336,3347|false|false|false|C0870325;C1547755;C1947919;C2347934;C4048755|Application Document;Apply;Computer Application;HL7 Version 2.5 - Application;Regulatory Application|application
Finding|Intellectual Product|Hospital Course|3336,3347|false|false|false|C0870325;C1547755;C1947919;C2347934;C4048755|Application Document;Apply;Computer Application;HL7 Version 2.5 - Application;Regulatory Application|application
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3336,3347|false|false|false|C0185125|Application procedure|application
Finding|Body Substance|Hospital Course|3348,3354|false|false|false|C0026727;C2753459|Mucus (substance);mucus layer|Mucous
Anatomy|Tissue|Hospital Course|3348,3363|false|false|false|C0026724|Mucous Membrane|Mucous Membrane
Disorder|Disease or Syndrome|Hospital Course|3348,3363|false|false|false|C0151785|Disease of mucous membrane|Mucous Membrane
Finding|Functional Concept|Hospital Course|3348,3363|false|false|false|C1549524|Route of Administration - Mucous Membrane|Mucous Membrane
Anatomy|Cell Component|Hospital Course|3355,3363|false|false|false|C0025255;C0596901|Membrane;Membrane Tissue|Membrane
Anatomy|Tissue|Hospital Course|3355,3363|false|false|false|C0025255;C0596901|Membrane;Membrane Tissue|Membrane
Drug|Organic Chemical|Hospital Course|3373,3382|false|false|false|C0005632|bisacodyl|Bisacodyl
Drug|Pharmacologic Substance|Hospital Course|3373,3382|false|false|false|C0005632|bisacodyl|Bisacodyl
Finding|Gene or Genome|Hospital Course|3401,3404|false|false|false|C1422467|CIAO3 gene|PRN
Finding|Sign or Symptom|Hospital Course|3405,3417|false|false|false|C0009806|Constipation|Constipation
Drug|Biologically Active Substance|Hospital Course|3423,3430|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|Hospital Course|3423,3430|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|Hospital Course|3423,3430|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|Hospital Course|3423,3430|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|Hospital Course|3423,3430|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Finding|Physiologic Function|Hospital Course|3423,3430|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|Hospital Course|3423,3430|false|false|false|C0201925|Calcium measurement|Calcium
Drug|Inorganic Chemical|Hospital Course|3423,3440|false|false|false|C0006681|calcium carbonate|Calcium Carbonate
Drug|Pharmacologic Substance|Hospital Course|3423,3440|false|false|false|C0006681|calcium carbonate|Calcium Carbonate
Drug|Element, Ion, or Isotope|Hospital Course|3431,3440|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|Carbonate
Drug|Organic Chemical|Hospital Course|3431,3440|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|Carbonate
Drug|Pharmacologic Substance|Hospital Course|3431,3440|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|Carbonate
Drug|Organic Chemical|Hospital Course|3461,3469|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|Hospital Course|3461,3469|false|false|false|C1692318|docusate|Docusate
Drug|Organic Chemical|Hospital Course|3461,3476|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|Hospital Course|3461,3476|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|Hospital Course|3470,3476|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|3470,3476|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|3470,3476|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Finding|Physiologic Function|Hospital Course|3470,3476|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|3470,3476|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|Hospital Course|3487,3490|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|3487,3490|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|3487,3490|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|3487,3490|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|3496,3506|false|false|false|C0206460|enoxaparin|Enoxaparin
Drug|Pharmacologic Substance|Hospital Course|3496,3506|false|false|false|C0206460|enoxaparin|Enoxaparin
Drug|Organic Chemical|Hospital Course|3496,3513|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Pharmacologic Substance|Hospital Course|3496,3513|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Biologically Active Substance|Hospital Course|3507,3513|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|3507,3513|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|3507,3513|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Finding|Physiologic Function|Hospital Course|3507,3513|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|3507,3513|false|false|false|C0337443|Sodium measurement|Sodium
Anatomy|Body Location or Region|Hospital Course|3529,3532|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|Hospital Course|3529,3532|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|Hospital Course|3529,3532|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3529,3544|false|false|false|C0853245|DVT prophylaxis|DVT prophylaxis
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3533,3544|false|false|false|C0199176|Prophylactic treatment|prophylaxis
Drug|Pharmacologic Substance|Hospital Course|3545,3553|false|false|false|C0720099|Duration brand of oxymetazoline|Duration
Finding|Idea or Concept|Hospital Course|3588,3592|false|false|false|C1552851|next - HtmlLinkType|Next
Finding|Idea or Concept|Hospital Course|3593,3600|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|Routine
Finding|Intellectual Product|Hospital Course|3593,3600|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|Routine
Procedure|Laboratory Procedure|Hospital Course|3593,3600|false|false|false|C1979801|Routine coag|Routine
Event|Occupational Activity|Hospital Course|3601,3615|false|false|false|C0001554|Administration occupational activities|Administration
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3601,3615|false|false|false|C1533734|Administration (procedure)|Administration
Finding|Finding|Hospital Course|3617,3621|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Finding|Idea or Concept|Hospital Course|3617,3621|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Finding|Intellectual Product|Hospital Course|3617,3621|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Drug|Organic Chemical|Hospital Course|3627,3637|false|false|false|C0206460|enoxaparin|enoxaparin
Drug|Pharmacologic Substance|Hospital Course|3627,3637|false|false|false|C0206460|enoxaparin|enoxaparin
Finding|Idea or Concept|Hospital Course|3687,3694|false|false|false|C0807726|refill|Refills
Drug|Food|Hospital Course|3702,3706|false|false|false|C0349374;C0444318;C1446647;C2702362;C2825079;C5551141;C5552693|Cow's milk;Milk Beverage;Milk Specimen;Milk antigen;Plant-Based Milk;cow milk allergenic extract|Milk
Drug|Immunologic Factor|Hospital Course|3702,3706|false|false|false|C0349374;C0444318;C1446647;C2702362;C2825079;C5551141;C5552693|Cow's milk;Milk Beverage;Milk Specimen;Milk antigen;Plant-Based Milk;cow milk allergenic extract|Milk
Drug|Pharmacologic Substance|Hospital Course|3702,3706|false|false|false|C0349374;C0444318;C1446647;C2702362;C2825079;C5551141;C5552693|Cow's milk;Milk Beverage;Milk Specimen;Milk antigen;Plant-Based Milk;cow milk allergenic extract|Milk
Drug|Substance|Hospital Course|3702,3706|false|false|false|C0349374;C0444318;C1446647;C2702362;C2825079;C5551141;C5552693|Cow's milk;Milk Beverage;Milk Specimen;Milk antigen;Plant-Based Milk;cow milk allergenic extract|Milk
Finding|Body Substance|Hospital Course|3702,3706|false|false|false|C0026131;C1546713|Milk (body substance);Milk Specimen Code|Milk
Finding|Intellectual Product|Hospital Course|3702,3706|false|false|false|C0026131;C1546713|Milk (body substance);Milk Specimen Code|Milk
Drug|Clinical Drug|Hospital Course|3702,3718|false|false|false|C0591789;C0782828|Milk of Magnesia (Brand Name);magnesium hydroxide Oral Suspension|Milk of Magnesia
Drug|Inorganic Chemical|Hospital Course|3702,3718|false|false|false|C0591789;C0782828|Milk of Magnesia (Brand Name);magnesium hydroxide Oral Suspension|Milk of Magnesia
Drug|Pharmacologic Substance|Hospital Course|3702,3718|false|false|false|C0591789;C0782828|Milk of Magnesia (Brand Name);magnesium hydroxide Oral Suspension|Milk of Magnesia
Drug|Inorganic Chemical|Hospital Course|3710,3718|false|false|false|C0024477|magnesium oxide|Magnesia
Drug|Pharmacologic Substance|Hospital Course|3710,3718|false|false|false|C0024477|magnesium oxide|Magnesia
Disorder|Mental or Behavioral Dysfunction|Hospital Course|3728,3731|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|3728,3731|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|3728,3731|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|3728,3731|false|false|false|C1332410|BID gene|BID
Finding|Gene or Genome|Hospital Course|3732,3735|false|false|false|C1422467|CIAO3 gene|PRN
Finding|Sign or Symptom|Hospital Course|3736,3745|false|false|false|C0013395|Dyspepsia|Dyspepsia
Drug|Organic Chemical|Hospital Course|3751,3764|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|Hospital Course|3751,3764|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|Hospital Course|3751,3764|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Disorder|Congenital Abnormality|Hospital Course|3767,3770|false|false|false|C1855179|CATARACT, ANTERIOR POLAR|CAP
Drug|Biomedical or Dental Material|Hospital Course|3767,3770|false|false|false|C0006935|capsule (pharmacologic)|CAP
Finding|Gene or Genome|Hospital Course|3767,3770|false|false|false|C1416891;C1418551;C1419093;C1422073;C1422760;C2985259;C4522312|BRD4 gene;BRD4 wt Allele;CAP1 gene;HACD1 gene;LNPEP gene;SERPINB6 gene;SORBS1 gene|CAP
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3767,3770|false|false|false|C0278651;C0280547;C1879916|CAP Regimen;cisplatin/cyclophosphamide/doxorubicin protocol;cyclophosphamide/doxorubicin/prednisone protocol|CAP
Drug|Organic Chemical|Hospital Course|3785,3794|false|false|false|C0030049|oxycodone|OxycoDONE
Drug|Pharmacologic Substance|Hospital Course|3785,3794|false|false|false|C0030049|oxycodone|OxycoDONE
Procedure|Laboratory Procedure|Hospital Course|3785,3794|false|false|false|C0524222|Oxycodone measurement|OxycoDONE
Finding|Idea or Concept|Hospital Course|3796,3805|false|false|false|C1548167;C1697779|Query Priority - Immediate;immediate - ResponseCode|Immediate
Finding|Intellectual Product|Hospital Course|3796,3805|false|false|false|C1548167;C1697779|Query Priority - Immediate;immediate - ResponseCode|Immediate
Drug|Biomedical or Dental Material|Hospital Course|3796,3813|false|false|false|C1708470|Immediate Release Dosage Form|Immediate Release
Finding|Functional Concept|Hospital Course|3806,3813|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|3806,3813|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3806,3813|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Finding|Gene or Genome|Hospital Course|3830,3833|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|3834,3838|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|3834,3838|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|3834,3838|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|Hospital Course|3844,3853|false|false|false|C0030049|oxycodone|oxycodone
Drug|Pharmacologic Substance|Hospital Course|3844,3853|false|false|false|C0030049|oxycodone|oxycodone
Procedure|Laboratory Procedure|Hospital Course|3844,3853|false|false|false|C0524222|Oxycodone measurement|oxycodone
Drug|Biomedical or Dental Material|Hospital Course|3863,3869|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|Hospital Course|3873,3881|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|3876,3881|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|3876,3881|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Event|Activity|Hospital Course|3899,3903|false|false|false|C1880359|Dispense (activity)|Disp
Finding|Gene or Genome|Hospital Course|3899,3903|false|false|false|C2828567|PRSS30P gene|Disp
Drug|Biomedical or Dental Material|Hospital Course|3910,3916|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|Hospital Course|3917,3924|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|3932,3944|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Pharmacologic Substance|Hospital Course|3932,3944|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Organic Chemical|Hospital Course|3964,3969|false|false|false|C3489575|sennosides, USP|Senna
Drug|Pharmacologic Substance|Hospital Course|3964,3969|false|false|false|C3489575|sennosides, USP|Senna
Drug|Biomedical or Dental Material|Hospital Course|3972,3975|false|false|false|C0039225|Tablet Dosage Form|TAB
Drug|Organic Chemical|Hospital Course|3987,3994|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|Hospital Course|3987,3994|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|Hospital Course|3987,3994|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|Hospital Course|3987,3996|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|Hospital Course|3987,3996|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|Hospital Course|3987,3996|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|Hospital Course|3987,3996|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|Hospital Course|3987,3996|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Finding|Body Substance|Hospital Course|4019,4028|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|4019,4028|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|4019,4028|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|4019,4028|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|4019,4040|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|4019,4040|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|4029,4040|false|false|false|C2926604||Disposition
Procedure|Health Care Activity|Hospital Course|4029,4040|false|false|false|C0184758|Patient disposition|Disposition
Finding|Finding|Hospital Course|4042,4050|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|4042,4050|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Procedure|Health Care Activity|Hospital Course|4042,4055|false|false|false|C0023977|long-term care|Extended Care
Event|Activity|Hospital Course|4051,4055|false|false|false|C1947933|care activity|Care
Finding|Finding|Hospital Course|4051,4055|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|Hospital Course|4051,4055|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|Hospital Course|4058,4066|false|false|false|C4695111|ADMIN.FACILITY|Facility
Finding|Body Substance|Hospital Course|4074,4083|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|4074,4083|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|4074,4083|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|4074,4083|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|4074,4093|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|4084,4093|false|false|false|C0945731||Diagnosis
Finding|Classification|Hospital Course|4084,4093|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|4084,4093|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|4084,4093|false|false|false|C0011900|Diagnosis|Diagnosis
Finding|Functional Concept|Hospital Course|4095,4099|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4095,4112|false|false|false|C0833290|Neck of left femur|left femoral neck
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4100,4107|false|false|false|C0015811|Femur|femoral
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4100,4112|false|false|false|C0015815|Structure of neck of femur|femoral neck
Disorder|Injury or Poisoning|Hospital Course|4100,4121|false|false|false|C0015806|Femoral Neck Fractures|femoral neck fracture
Anatomy|Body Location or Region|Hospital Course|4108,4112|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|Hospital Course|4108,4112|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|Hospital Course|4108,4112|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Disorder|Injury or Poisoning|Hospital Course|4108,4121|false|false|false|C0262414|Fracture of cervical spine|neck fracture
Disorder|Injury or Poisoning|Hospital Course|4113,4121|false|false|false|C0016658|Fracture|fracture
Finding|Mental Process|Discharge Condition|4146,4152|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|4146,4159|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|4146,4159|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|4153,4159|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|4153,4159|false|false|false|C1546481|What subject filter - Status|Status
Finding|Idea or Concept|Discharge Condition|4161,4166|false|false|false|C1550016|Remote control command - Clear|Clear
Finding|Finding|Discharge Condition|4171,4179|false|false|false|C4068804|Coherent|coherent
Attribute|Clinical Attribute|Discharge Condition|4181,4203|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|4181,4203|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Finding|Finding|Discharge Condition|4190,4203|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|4190,4203|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|4205,4210|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|4205,4210|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|4205,4210|false|false|false|C0718338|Alert brand of caffeine|Alert
Finding|Finding|Discharge Condition|4205,4210|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|4205,4210|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|4205,4210|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|4215,4226|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|4228,4236|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|4228,4236|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|4228,4236|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|4237,4243|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|4237,4243|false|false|false|C1546481|What subject filter - Status|Status
Disorder|Disease or Syndrome|Discharge Condition|4252,4255|false|false|false|C3159311|BORNHOLM EYE DISEASE|Bed
Finding|Intellectual Product|Discharge Condition|4252,4255|false|false|false|C2346952|Bachelor of Education|Bed
Finding|Social Behavior|Discharge Condition|4261,4271|false|false|false|C0018896|Helping Behavior|assistance
Finding|Finding|Discharge Condition|4285,4295|false|false|false|C2135586;C4321408|Wheelchair Usually Used;has wheelchair at home (history)|wheelchair
Attribute|Clinical Attribute|Medications|4356,4367|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Medications|4356,4367|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|Medications|4356,4367|false|false|false|C4284232|Medications|medications
Finding|Body Substance|Medications|4405,4414|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Medications|4405,4414|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Medications|4405,4414|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Medications|4405,4414|false|false|false|C0030685|Patient Discharge|discharge
Finding|Idea or Concept|Medications|4432,4436|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Medications|4432,4436|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Medications|4432,4436|false|false|false|C1553498|home health encounter|home
Attribute|Clinical Attribute|Medications|4437,4448|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Medications|4437,4448|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|Medications|4437,4448|false|false|false|C4284232|Medications|medications
Attribute|Clinical Attribute|Medications|4497,4504|false|false|false|C5444295||surgeon
Drug|Organic Chemical|Medications|4522,4529|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Drug|Pharmacologic Substance|Medications|4522,4529|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Finding|Intellectual Product|Medications|4522,4529|false|false|false|C1547288|Alcohol - Recreational Drug Use Code|alcohol
Finding|Functional Concept|Medications|4539,4544|false|false|false|C1513492|motor movement|motor
Drug|Biomedical or Dental Material|Medications|4545,4552|false|false|false|C0042444|Drug vehicle|vehicle
Finding|Functional Concept|Medications|4557,4564|false|false|false|C3242339|operate|operate
Disorder|Injury or Poisoning|Medications|4566,4575|false|false|false|C0337246|Contact with machinery|machinery
Drug|Hazardous or Poisonous Substance|Medications|4589,4597|false|false|false|C0027415|Narcotics|narcotic
Drug|Pharmacologic Substance|Medications|4589,4597|false|false|false|C0027415|Narcotics|narcotic
Attribute|Clinical Attribute|Medications|4598,4602|false|false|false|C2598155||pain
Finding|Functional Concept|Medications|4598,4602|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Medications|4598,4602|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Hazardous or Poisonous Substance|Medications|4598,4612|false|false|false|C0002771;C0722425|Analgesics;Pain Relieve brand of acetaminophen|pain relievers
Drug|Organic Chemical|Medications|4598,4612|false|false|false|C0002771;C0722425|Analgesics;Pain Relieve brand of acetaminophen|pain relievers
Drug|Pharmacologic Substance|Medications|4598,4612|false|false|false|C0002771;C0722425|Analgesics;Pain Relieve brand of acetaminophen|pain relievers
Drug|Hazardous or Poisonous Substance|Medications|4617,4625|false|false|false|C0027415|Narcotics|Narcotic
Drug|Pharmacologic Substance|Medications|4617,4625|false|false|false|C0027415|Narcotics|Narcotic
Attribute|Clinical Attribute|Medications|4626,4630|false|false|false|C2598155||pain
Finding|Functional Concept|Medications|4626,4630|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Medications|4626,4630|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Hazardous or Poisonous Substance|Medications|4626,4640|false|false|false|C0002771;C0722425|Analgesics;Pain Relieve brand of acetaminophen|pain relievers
Drug|Organic Chemical|Medications|4626,4640|false|false|false|C0002771;C0722425|Analgesics;Pain Relieve brand of acetaminophen|pain relievers
Drug|Pharmacologic Substance|Medications|4626,4640|false|false|false|C0002771;C0722425|Analgesics;Pain Relieve brand of acetaminophen|pain relievers
Finding|Sign or Symptom|Medications|4651,4663|false|false|false|C0009806|Constipation|constipation
Drug|Food|Medications|4680,4685|false|false|false|C0452428|Drink (dietary substance)|drink
Drug|Inorganic Chemical|Medications|4707,4712|false|false|false|C0043047;C1550678|Water Specimen;water|water
Drug|Pharmacologic Substance|Medications|4707,4712|false|false|false|C0043047;C1550678|Water Specimen;water|water
Finding|Intellectual Product|Medications|4707,4712|false|false|false|C1547961|Water - Specimen Source Codes|water
Procedure|Therapeutic or Preventive Procedure|Medications|4707,4712|false|false|false|C0020311|Hydrotherapy|water
Finding|Body Substance|Medications|4730,4735|false|false|false|C0015733|Feces|stool
Drug|Organic Chemical|Medications|4730,4744|false|false|false|C0301470;C1154263|Stool Softener;Stool Softener brand of docusate sodium|stool softener
Drug|Pharmacologic Substance|Medications|4730,4744|false|false|false|C0301470;C1154263|Stool Softener;Stool Softener brand of docusate sodium|stool softener
Drug|Organic Chemical|Medications|4747,4753|false|false|false|C0282139|Colace|colace
Drug|Pharmacologic Substance|Medications|4747,4753|false|false|false|C0282139|Colace|colace
Finding|Pathologic Function|Medications|4771,4782|false|false|false|C0879626|Adverse effects|side effect
Finding|Finding|Medications|4788,4803|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|ANTICOAGULATION
Finding|Physiologic Function|Medications|4788,4803|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|ANTICOAGULATION
Procedure|Therapeutic or Preventive Procedure|Medications|4788,4803|false|false|false|C0003281|Anticoagulation Therapy|ANTICOAGULATION
Drug|Organic Chemical|Medications|4820,4827|false|false|false|C0728963|Lovenox|lovenox
Drug|Pharmacologic Substance|Medications|4820,4827|false|false|false|C0728963|Lovenox|lovenox
Disorder|Injury or Poisoning|Medications|4855,4860|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|WOUND
Finding|Body Substance|Medications|4855,4860|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|WOUND
Finding|Functional Concept|Medications|4855,4860|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|WOUND
Finding|Intellectual Product|Medications|4855,4860|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|WOUND
Procedure|Therapeutic or Preventive Procedure|Medications|4855,4865|false|false|false|C0886052;C1272654|Wound care management;wound care|WOUND CARE
Event|Activity|Medications|4861,4865|false|false|false|C1947933|care activity|CARE
Finding|Finding|Medications|4861,4865|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|CARE
Finding|Intellectual Product|Medications|4861,4865|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|CARE
Disorder|Injury or Poisoning|Medications|4886,4891|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|wound
Finding|Body Substance|Medications|4886,4891|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Functional Concept|Medications|4886,4891|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Intellectual Product|Medications|4886,4891|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Daily or Recreational Activity|Medications|4896,4909|false|false|false|C2937301|take a shower|take a shower
Finding|Finding|Medications|4938,4945|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|Medications|4938,4945|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|Medications|4938,4945|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|Medications|4938,4945|false|false|false|C0543467|Operative Surgical Procedures|surgery
Drug|Biomedical or Dental Material|Medications|4973,4977|false|false|false|C1705308|Soap Dosage Form|soap
Drug|Inorganic Chemical|Medications|4982,4987|false|false|false|C0043047;C1550678|Water Specimen;water|water
Drug|Pharmacologic Substance|Medications|4982,4987|false|false|false|C0043047;C1550678|Water Specimen;water|water
Finding|Intellectual Product|Medications|4982,4987|false|false|false|C1547961|Water - Specimen Source Codes|water
Procedure|Therapeutic or Preventive Procedure|Medications|4982,4987|false|false|false|C0020311|Hydrotherapy|water
Disorder|Disease or Syndrome|Medications|4993,4996|false|false|false|C0030587|Paroxysmal atrial tachycardia|pat
Drug|Organic Chemical|Medications|4993,4996|false|false|false|C2825250|Fenamole|pat
Drug|Pharmacologic Substance|Medications|4993,4996|false|false|false|C2825250|Fenamole|pat
Finding|Molecular Function|Medications|4993,4996|false|false|false|C2247344;C2247346;C2248827|aspartate-prephenate aminotransferase activity;glutamate-prephenate aminotransferase activity;protein acetyltransferase activity|pat
Procedure|Diagnostic Procedure|Medications|4993,4996|false|false|false|C3897364|Thermoacoustic Computed Tomography|pat
Anatomy|Body Location or Region|Medications|5002,5010|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|Medications|5002,5010|false|false|false|C0332803|Surgical wound|incision
Procedure|Therapeutic or Preventive Procedure|Medications|5002,5010|false|false|false|C0184898|Surgical incisions|incision
Procedure|Health Care Activity|Medications|5040,5045|true|false|false|C0150141|Bathing|baths
Finding|Daily or Recreational Activity|Medications|5049,5057|true|false|false|C0039003;C2362608|Swimming;swimming (history)|swimming
Finding|Finding|Medications|5049,5057|true|false|false|C0039003;C2362608|Swimming;swimming (history)|swimming
Finding|Intellectual Product|Medications|5160,5164|false|false|false|C1561540|Transaction counts and value totals - week|week
Event|Activity|Medications|5175,5186|false|false|false|C0003629|Appointments|appointment
Drug|Biomedical or Dental Material|Medications|5194,5202|true|false|false|C1705365|Dressing Dosage Form|dressing
Finding|Daily or Recreational Activity|Medications|5194,5202|true|false|false|C0518459;C1305428|Ability to dress|dressing
Finding|Finding|Medications|5194,5202|true|false|false|C0518459;C1305428|Ability to dress|dressing
Procedure|Health Care Activity|Medications|5194,5202|true|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|dressing
Procedure|Therapeutic or Preventive Procedure|Medications|5194,5202|true|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|dressing
Disorder|Injury or Poisoning|Medications|5216,5221|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|wound
Finding|Body Substance|Medications|5216,5221|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Functional Concept|Medications|5216,5221|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Intellectual Product|Medications|5216,5221|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Event|Activity|Medications|5256,5264|false|false|false|C0441655|Activities|ACTIVITY
Finding|Daily or Recreational Activity|Medications|5256,5264|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|ACTIVITY
Finding|Finding|Medications|5256,5264|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|ACTIVITY
Attribute|Clinical Attribute|Medications|5269,5275|false|false|false|C0944911||WEIGHT
Finding|Finding|Medications|5269,5275|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|WEIGHT
Finding|Sign or Symptom|Medications|5269,5275|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|WEIGHT
Procedure|Health Care Activity|Medications|5269,5275|false|false|false|C1305866|Weighing patient|WEIGHT
Finding|Mental Process|Medications|5286,5291|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Finding|Organ or Tissue Function|Medications|5286,5291|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Procedure|Therapeutic or Preventive Procedure|Medications|5286,5291|false|false|false|C0152054|Therapeutic Touch|touch
Attribute|Clinical Attribute|Medications|5297,5303|false|false|false|C0944911||weight
Finding|Finding|Medications|5297,5303|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|Medications|5297,5303|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|Medications|5297,5303|false|false|false|C1305866|Weighing patient|weight
Finding|Finding|Medications|5316,5324|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|Medications|5316,5324|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|Medications|5316,5324|false|false|false|C0031809|Physical Examination|Physical
Finding|Intellectual Product|Medications|5316,5332|false|false|false|C1547999|Diagnostic Service Section ID - Physical Therapy|Physical Therapy
Procedure|Therapeutic or Preventive Procedure|Medications|5316,5332|false|false|false|C0949766|Physical therapy|Physical Therapy
Finding|Finding|Medications|5325,5332|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|Therapy
Finding|Functional Concept|Medications|5325,5332|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|Therapy
Procedure|Therapeutic or Preventive Procedure|Medications|5325,5332|false|false|false|C0087111|Therapeutic procedure|Therapy
Finding|Mental Process|Medications|5334,5339|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|Touch
Finding|Organ or Tissue Function|Medications|5334,5339|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|Touch
Procedure|Therapeutic or Preventive Procedure|Medications|5334,5339|false|false|false|C0152054|Therapeutic Touch|Touch
Attribute|Clinical Attribute|Medications|5345,5351|false|false|false|C0944911||weight
Finding|Finding|Medications|5345,5351|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|Medications|5345,5351|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|Medications|5345,5351|false|false|false|C1305866|Weighing patient|weight
Procedure|Therapeutic or Preventive Procedure|Medications|5364,5374|false|false|false|C0087111|Therapeutic procedure|Treatments
Finding|Intellectual Product|Medications|5375,5384|false|false|false|C3898838;C4321352|Frequency;How Often|Frequency
Disorder|Injury or Poisoning|Medications|5386,5391|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|WOUND
Finding|Body Substance|Medications|5386,5391|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|WOUND
Finding|Functional Concept|Medications|5386,5391|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|WOUND
Finding|Intellectual Product|Medications|5386,5391|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|WOUND
Procedure|Therapeutic or Preventive Procedure|Medications|5386,5396|false|false|false|C0886052;C1272654|Wound care management;wound care|WOUND CARE
Event|Activity|Medications|5392,5396|false|false|false|C1947933|care activity|CARE
Finding|Finding|Medications|5392,5396|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|CARE
Finding|Intellectual Product|Medications|5392,5396|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|CARE
Disorder|Injury or Poisoning|Medications|5417,5422|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|wound
Finding|Body Substance|Medications|5417,5422|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Functional Concept|Medications|5417,5422|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Intellectual Product|Medications|5417,5422|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Daily or Recreational Activity|Medications|5427,5440|false|false|false|C2937301|take a shower|take a shower
Finding|Finding|Medications|5469,5476|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|Medications|5469,5476|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|Medications|5469,5476|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|Medications|5469,5476|false|false|false|C0543467|Operative Surgical Procedures|surgery
Drug|Biomedical or Dental Material|Medications|5504,5508|false|false|false|C1705308|Soap Dosage Form|soap
Drug|Inorganic Chemical|Medications|5513,5518|false|false|false|C0043047;C1550678|Water Specimen;water|water
Drug|Pharmacologic Substance|Medications|5513,5518|false|false|false|C0043047;C1550678|Water Specimen;water|water
Finding|Intellectual Product|Medications|5513,5518|false|false|false|C1547961|Water - Specimen Source Codes|water
Procedure|Therapeutic or Preventive Procedure|Medications|5513,5518|false|false|false|C0020311|Hydrotherapy|water
Disorder|Disease or Syndrome|Medications|5524,5527|false|false|false|C0030587|Paroxysmal atrial tachycardia|pat
Drug|Organic Chemical|Medications|5524,5527|false|false|false|C2825250|Fenamole|pat
Drug|Pharmacologic Substance|Medications|5524,5527|false|false|false|C2825250|Fenamole|pat
Finding|Molecular Function|Medications|5524,5527|false|false|false|C2247344;C2247346;C2248827|aspartate-prephenate aminotransferase activity;glutamate-prephenate aminotransferase activity;protein acetyltransferase activity|pat
Procedure|Diagnostic Procedure|Medications|5524,5527|false|false|false|C3897364|Thermoacoustic Computed Tomography|pat
Anatomy|Body Location or Region|Medications|5533,5541|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|Medications|5533,5541|false|false|false|C0332803|Surgical wound|incision
Procedure|Therapeutic or Preventive Procedure|Medications|5533,5541|false|false|false|C0184898|Surgical incisions|incision
Procedure|Health Care Activity|Medications|5571,5576|true|false|false|C0150141|Bathing|baths
Finding|Daily or Recreational Activity|Medications|5580,5588|true|false|false|C0039003;C2362608|Swimming;swimming (history)|swimming
Finding|Finding|Medications|5580,5588|true|false|false|C0039003;C2362608|Swimming;swimming (history)|swimming
Finding|Intellectual Product|Medications|5691,5695|false|false|false|C1561540|Transaction counts and value totals - week|week
Event|Activity|Medications|5706,5717|false|false|false|C0003629|Appointments|appointment
Drug|Biomedical or Dental Material|Medications|5725,5733|true|false|false|C1705365|Dressing Dosage Form|dressing
Finding|Daily or Recreational Activity|Medications|5725,5733|true|false|false|C0518459;C1305428|Ability to dress|dressing
Finding|Finding|Medications|5725,5733|true|false|false|C0518459;C1305428|Ability to dress|dressing
Procedure|Health Care Activity|Medications|5725,5733|true|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|dressing
Procedure|Therapeutic or Preventive Procedure|Medications|5725,5733|true|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|dressing
Disorder|Injury or Poisoning|Medications|5747,5752|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|wound
Finding|Body Substance|Medications|5747,5752|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Functional Concept|Medications|5747,5752|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Intellectual Product|Medications|5747,5752|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Procedure|Health Care Activity|Medications|5786,5794|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Medications|5795,5807|false|false|false|C3263700||Instructions
Finding|Intellectual Product|Medications|5795,5807|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

