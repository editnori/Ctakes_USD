 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
_|27,28
_|28,29
_|29,30
No|31,33
:|33,34
_|37,38
_|38,39
_|39,40
<EOL>|40,41
<EOL>|42,43
Admission|43,52
Date|53,57
:|57,58
_|60,61
_|61,62
_|62,63
Discharge|77,86
Date|87,91
:|91,92
_|95,96
_|96,97
_|97,98
<EOL>|98,99
<EOL>|100,101
Date|101,105
of|106,108
Birth|109,114
:|114,115
_|117,118
_|118,119
_|119,120
Sex|133,136
:|136,137
F|140,141
<EOL>|141,142
<EOL>|143,144
Service|144,151
:|151,152
MEDICINE|153,161
<EOL>|161,162
<EOL>|163,164
No|176,178
Known|179,184
Allergies|185,194
/|195,196
Adverse|197,204
Drug|205,209
Reactions|210,219
<EOL>|219,220
<EOL>|221,222
Attending|222,231
:|231,232
_|233,234
_|234,235
_|235,236
.|236,237
<EOL>|237,238
<EOL>|239,240
Shortness|257,266
of|267,269
breath|270,276
,|276,277
altered|278,285
mental|286,292
status|293,299
<EOL>|299,300
<EOL>|301,302
Major|302,307
Surgical|308,316
or|317,319
Invasive|320,328
Procedure|329,338
:|338,339
<EOL>|339,340
None|340,344
<EOL>|344,345
<EOL>|345,346
<EOL>|347,348
Patient|376,383
is|384,386
an|387,389
_|390,391
_|391,392
_|392,393
year|394,398
-|398,399
old|399,402
patient|403,410
with|411,415
history|416,423
of|424,426
Sjogren|427,434
's|434,436
<EOL>|437,438
syndrome|438,446
,|446,447
moderate|448,456
MR|457,459
,|459,460
recent|461,467
hospitalization|468,483
for|484,487
sepsis|488,494
<EOL>|495,496
secondary|496,505
to|506,508
c.|509,511
diff|512,516
colitis|517,524
complicated|525,536
by|537,539
hypercarbic|540,551
<EOL>|552,553
respiratory|553,564
failure|565,572
requiring|573,582
intubation|583,593
,|593,594
who|595,598
is|599,601
presenting|602,612
from|613,617
<EOL>|618,619
_|619,620
_|620,621
_|621,622
with|623,627
worsening|628,637
dyspnea|638,645
for|646,649
one|650,653
day|654,657
.|657,658
Patient|660,667
was|668,671
<EOL>|672,673
discharged|673,683
from|684,688
_|689,690
_|690,691
_|691,692
yesterday|693,702
(|703,704
_|704,705
_|705,706
_|706,707
)|707,708
following|709,718
hospitalization|719,734
<EOL>|735,736
for|736,739
c.|740,742
diff|743,747
colitis|748,755
.|755,756
Patient|758,765
had|766,769
ABG|770,773
at|774,776
_|777,778
_|778,779
_|779,780
,|780,781
which|782,787
was|788,791
<EOL>|792,793
7.|793,795
_|795,796
_|796,797
_|797,798
.|798,799
Her|801,804
vitals|805,811
on|812,814
transfer|815,823
were|824,828
97.9|829,833
99|834,836
24|837,839
113|840,843
/|843,844
68|844,846
92|847,849
%|849,850
<EOL>|851,852
2L|852,854
.|854,855
She|856,859
reports|860,867
shortness|868,877
of|878,880
breath|881,887
associated|888,898
with|899,903
the|904,907
cough|908,913
.|913,914
<EOL>|915,916
She|916,919
denies|920,926
chest|927,932
pain|933,937
.|937,938
She|939,942
denies|943,949
nausea|950,956
or|957,959
vomiting|960,968
.|968,969
She|970,973
denies|974,980
<EOL>|981,982
abdominal|982,991
pain|992,996
.|996,997
<EOL>|997,998
<EOL>|998,999
In|999,1001
the|1002,1005
ED|1006,1008
,|1008,1009
initial|1010,1017
vitals|1018,1024
are|1025,1028
100.2|1029,1034
95|1035,1037
99|1038,1040
/|1040,1041
47|1041,1043
28|1044,1046
100|1047,1050
%|1050,1051
4L|1052,1054
nc|1055,1057
.|1057,1058
<EOL>|1060,1061
Exam|1061,1065
was|1066,1069
notable|1070,1077
for|1078,1081
tachypnea|1082,1091
with|1092,1096
respiratory|1097,1108
rates|1109,1114
in|1115,1117
the|1118,1121
<EOL>|1122,1123
_|1123,1124
_|1124,1125
_|1125,1126
.|1126,1127
While|1129,1134
in|1135,1137
ED|1138,1140
,|1140,1141
blood|1142,1147
pressure|1148,1156
dipped|1157,1163
to|1164,1166
_|1167,1168
_|1168,1169
_|1169,1170
,|1170,1171
but|1172,1175
improved|1176,1184
on|1185,1187
<EOL>|1188,1189
it|1189,1191
's|1191,1193
own|1194,1197
.|1197,1198
Given|1199,1204
the|1205,1208
tachypnea|1209,1218
,|1218,1219
cough|1220,1225
,|1225,1226
and|1227,1230
dyspnea|1231,1238
,|1238,1239
there|1240,1245
was|1246,1249
<EOL>|1250,1251
concern|1251,1258
for|1259,1262
pneumonia|1263,1272
.|1272,1273
Patient|1275,1282
received|1283,1291
vancomycin|1292,1302
and|1303,1306
<EOL>|1307,1308
levofloxacin|1308,1320
.|1320,1321
CXR|1323,1326
appeared|1327,1335
improved|1336,1344
from|1345,1349
most|1350,1354
recent|1355,1361
CXR|1362,1365
.|1365,1366
<EOL>|1368,1369
Patiwnt|1369,1376
was|1377,1380
started|1381,1388
on|1389,1391
BIPAP|1392,1397
.|1397,1398
Patient|1400,1407
underwent|1408,1417
CTA|1418,1421
to|1422,1424
evaluate|1425,1433
<EOL>|1434,1435
for|1435,1438
PE|1439,1441
prior|1442,1447
to|1448,1450
leaving|1451,1458
ED|1459,1461
.|1461,1462
On|1464,1466
transfer|1467,1475
vitals|1476,1482
are|1483,1486
,|1486,1487
HR|1488,1490
93|1491,1493
,|1493,1494
BP|1495,1497
<EOL>|1498,1499
109|1499,1502
/|1502,1503
45|1503,1505
,|1505,1506
O2|1507,1509
sat|1510,1513
100|1514,1517
%|1517,1518
on|1519,1521
BIPAP|1522,1527
.|1527,1528
<EOL>|1531,1532
<EOL>|1532,1533
On|1533,1535
arrival|1536,1543
to|1544,1546
the|1547,1550
MICU|1551,1555
,|1555,1556
patient|1557,1564
is|1565,1567
wearing|1568,1575
BiPAP|1576,1581
,|1581,1582
but|1583,1586
wants|1587,1592
it|1593,1595
<EOL>|1596,1597
removed|1597,1604
and|1605,1608
does|1609,1613
not|1614,1617
want|1618,1622
any|1623,1626
other|1627,1632
supplemental|1633,1645
oxygen|1646,1652
.|1652,1653
She|1655,1658
<EOL>|1659,1660
denies|1660,1666
pain|1667,1671
.|1671,1672
She|1673,1676
denies|1677,1683
cough|1684,1689
or|1690,1692
shortness|1693,1702
of|1703,1705
breath|1706,1712
.|1712,1713
<EOL>|1715,1716
<EOL>|1716,1717
Review|1717,1723
of|1724,1726
systems|1727,1734
:|1734,1735
<EOL>|1736,1737
Unable|1737,1743
to|1744,1746
obtain|1747,1753
,|1753,1754
patient|1755,1762
wearing|1763,1770
BiPAP|1771,1776
and|1777,1780
is|1781,1783
delerious|1784,1793
.|1793,1794
<EOL>|1796,1797
<EOL>|1797,1798
<EOL>|1799,1800
Anemia|1822,1828
<EOL>|1830,1831
Borderline|1831,1841
cholesterol|1842,1853
<EOL>|1855,1856
C.|1856,1858
Diff|1859,1863
<EOL>|1865,1866
Flatulence|1866,1876
<EOL>|1878,1879
Health|1879,1885
Maintenance|1886,1897
<EOL>|1899,1900
Heart|1900,1905
Murmur|1906,1912
<EOL>|1914,1915
Hypertension|1915,1927
<EOL>|1929,1930
Hypothyroidism|1930,1944
<EOL>|1946,1947
Mitral|1947,1953
Regurgitation|1954,1967
<EOL>|1969,1970
Osteoporosis|1970,1982
<EOL>|1984,1985
Pneumonia|1985,1994
<EOL>|1996,1997
Sinusitis|1997,2006
<EOL>|2008,2009
_|2009,2010
_|2010,2011
_|2011,2012
<EOL>|2014,2015
<EOL>|2015,2016
<EOL>|2017,2018
:|2032,2033
<EOL>|2033,2034
_|2034,2035
_|2035,2036
_|2036,2037
<EOL>|2037,2038
:|2052,2053
<EOL>|2053,2054
Long|2054,2058
history|2059,2066
of|2067,2069
hypertension|2070,2082
in|2083,2085
her|2086,2089
family|2090,2096
.|2096,2097
She|2099,2102
does|2103,2107
report|2108,2114
<EOL>|2115,2116
that|2116,2120
her|2121,2124
father|2125,2131
's|2131,2133
family|2134,2140
has|2141,2144
a|2145,2146
history|2147,2154
of|2155,2157
multiple|2158,2166
cancers|2167,2174
.|2174,2175
She|2177,2180
<EOL>|2181,2182
has|2182,2185
a|2186,2187
grandfather|2188,2199
with|2200,2204
a|2205,2206
history|2207,2214
of|2215,2217
stomach|2218,2225
cancer|2226,2232
and|2233,2236
an|2237,2239
uncle|2240,2245
<EOL>|2246,2247
with|2247,2251
a|2252,2253
history|2254,2261
of|2262,2264
throat|2265,2271
cancer|2272,2278
.|2278,2279
She|2281,2284
denies|2285,2291
any|2292,2295
history|2296,2303
of|2304,2306
<EOL>|2307,2308
colon|2308,2313
cancers|2314,2321
.|2321,2322
Father|2323,2329
had|2330,2333
stroke|2334,2340
.|2340,2341
No|2342,2344
family|2345,2351
h|2352,2353
/|2353,2354
o|2354,2355
MI|2356,2358
.|2358,2359
Mother|2360,2366
had|2367,2370
a|2371,2372
<EOL>|2373,2374
heart|2374,2379
valve|2380,2385
replaced|2386,2394
(|2395,2396
pt|2396,2398
not|2399,2402
sure|2403,2407
which|2408,2413
one|2414,2417
)|2417,2418
.|2418,2419
<EOL>|2419,2420
<EOL>|2420,2421
<EOL>|2422,2423
Exam|2438,2442
upon|2443,2447
admission|2448,2457
:|2457,2458
<EOL>|2458,2459
General|2459,2466
:|2466,2467
Awake|2468,2473
,|2473,2474
interactive|2475,2486
,|2486,2487
but|2488,2491
delerious|2492,2501
.|2501,2502
Not|2503,2506
oriented|2507,2515
to|2516,2518
<EOL>|2519,2520
place|2520,2525
or|2526,2528
time|2529,2533
,|2533,2534
calling|2535,2542
out|2543,2546
,|2546,2547
trying|2548,2554
to|2555,2557
get|2558,2561
out|2562,2565
of|2566,2568
bed|2569,2572
.|2572,2573
Cachetic|2574,2582
,|2582,2583
<EOL>|2584,2585
frail|2585,2590
,|2590,2591
elderly|2592,2599
female|2600,2606
.|2606,2607
<EOL>|2608,2609
HEENT|2609,2614
:|2614,2615
Sclera|2616,2622
anicteric|2623,2632
,|2632,2633
dry|2634,2637
mucus|2638,2643
membranes|2644,2653
.|2653,2654
<EOL>|2656,2657
Neck|2657,2661
:|2661,2662
supple|2663,2669
,|2669,2670
JVP|2671,2674
not|2675,2678
elevated|2679,2687
,|2687,2688
no|2689,2691
LAD|2692,2695
<EOL>|2697,2698
CV|2698,2700
:|2700,2701
Regular|2702,2709
rate|2710,2714
and|2715,2718
rhythm|2719,2725
,|2725,2726
normal|2727,2733
S1|2734,2736
+|2737,2738
S2|2739,2741
,|2741,2742
II|2743,2745
/|2745,2746
VI|2746,2748
systolic|2749,2757
<EOL>|2758,2759
murmur|2759,2765
at|2766,2768
apex|2769,2773
.|2773,2774
<EOL>|2774,2775
Lungs|2775,2780
:|2780,2781
Dull|2782,2786
at|2787,2789
bases|2790,2795
bilaterally|2796,2807
,|2807,2808
breathing|2809,2818
comfortably|2819,2830
,|2830,2831
no|2832,2834
<EOL>|2835,2836
accessory|2836,2845
muscle|2846,2852
use|2853,2856
.|2856,2857
<EOL>|2857,2858
Abdomen|2858,2865
:|2865,2866
soft|2867,2871
,|2871,2872
distended|2873,2882
,|2882,2883
non-tender|2884,2894
,|2894,2895
no|2896,2898
rebound|2899,2906
/|2906,2907
guarding|2907,2915
.|2915,2916
bowel|2917,2922
<EOL>|2923,2924
sounds|2924,2930
present|2931,2938
.|2938,2939
Flexiseal|2941,2950
draining|2951,2959
watery|2960,2966
stool|2967,2972
with|2973,2977
blood|2978,2983
in|2984,2986
<EOL>|2987,2988
it|2988,2990
.|2990,2991
<EOL>|2991,2992
GU|2992,2994
:|2994,2995
foley|2996,3001
in|3002,3004
place|3005,3010
foley|3011,3016
<EOL>|3017,3018
Ext|3018,3021
:|3021,3022
warm|3023,3027
,|3027,3028
1|3029,3030
+|3030,3031
DP|3032,3034
pulses|3035,3041
,|3041,3042
Diffuse|3043,3050
edema|3051,3056
<EOL>|3056,3057
Neuro|3057,3062
:|3062,3063
CNII|3064,3068
-|3068,3069
XII|3069,3072
intact|3073,3079
,|3079,3080
disoriented|3081,3092
,|3092,3093
inattentive|3094,3105
<EOL>|3105,3106
<EOL>|3106,3107
Discharge|3107,3116
exam|3117,3121
-|3122,3123
unchanged|3124,3133
from|3134,3138
above|3139,3144
,|3144,3145
except|3146,3152
as|3153,3155
below|3156,3161
:|3161,3162
<EOL>|3162,3163
General|3163,3170
:|3170,3171
Awake|3172,3177
,|3177,3178
sleepy|3179,3185
but|3186,3189
arousable|3190,3199
to|3200,3202
voice|3203,3208
,|3208,3209
NAD|3210,3213
<EOL>|3213,3214
GU|3214,3216
:|3216,3217
Foley|3218,3223
removed|3224,3231
<EOL>|3231,3232
Neuro|3232,3237
:|3237,3238
A|3239,3240
&|3240,3241
Ox2|3241,3244
(|3245,3246
name|3246,3250
and|3251,3254
date|3255,3259
)|3259,3260
,|3260,3261
MS|3262,3264
has|3265,3268
been|3269,3273
waxing|3274,3280
/|3280,3281
waning|3281,3287
,|3287,3288
no|3289,3291
<EOL>|3292,3293
focal|3293,3298
defecits|3299,3307
<EOL>|3307,3308
<EOL>|3309,3310
Pertinent|3310,3319
Results|3320,3327
:|3327,3328
<EOL>|3328,3329
Labs|3329,3333
upon|3334,3338
admission|3339,3348
:|3348,3349
<EOL>|3349,3350
_|3350,3351
_|3351,3352
_|3352,3353
07|3354,3356
:|3356,3357
30AM|3357,3361
BLOOD|3362,3367
WBC|3368,3371
-|3371,3372
7.1|3372,3375
RBC|3376,3379
-|3379,3380
3|3380,3381
.|3381,3382
11|3382,3384
*|3384,3385
Hgb|3386,3389
-|3389,3390
9|3390,3391
.|3391,3392
3|3392,3393
*|3393,3394
Hct|3395,3398
-|3398,3399
30|3399,3401
.|3401,3402
3|3402,3403
*|3403,3404
<EOL>|3405,3406
MCV|3406,3409
-|3409,3410
97|3410,3412
MCH|3413,3416
-|3416,3417
29.9|3417,3421
MCHC|3422,3426
-|3426,3427
30|3427,3429
.|3429,3430
7|3430,3431
*|3431,3432
RDW|3433,3436
-|3436,3437
14.0|3437,3441
Plt|3442,3445
_|3446,3447
_|3447,3448
_|3448,3449
<EOL>|3449,3450
_|3450,3451
_|3451,3452
_|3452,3453
07|3454,3456
:|3456,3457
10PM|3457,3461
BLOOD|3462,3467
Neuts|3468,3473
-|3473,3474
68.2|3474,3478
_|3479,3480
_|3480,3481
_|3481,3482
Monos|3483,3488
-|3488,3489
6.6|3489,3492
Eos|3493,3496
-|3496,3497
2.4|3497,3500
<EOL>|3501,3502
Baso|3502,3506
-|3506,3507
1.0|3507,3510
<EOL>|3510,3511
_|3511,3512
_|3512,3513
_|3513,3514
07|3515,3517
:|3517,3518
30AM|3518,3522
BLOOD|3523,3528
Glucose|3529,3536
-|3536,3537
122|3537,3540
*|3540,3541
UreaN|3542,3547
-|3547,3548
20|3548,3550
Creat|3551,3556
-|3556,3557
0|3557,3558
.|3558,3559
3|3559,3560
*|3560,3561
Na|3562,3564
-|3564,3565
133|3565,3568
<EOL>|3569,3570
K|3570,3571
-|3571,3572
4.0|3572,3575
Cl|3576,3578
-|3578,3579
92|3579,3581
*|3581,3582
HCO3|3583,3587
-|3587,3588
39|3588,3590
*|3590,3591
AnGap|3592,3597
-|3597,3598
6|3598,3599
*|3599,3600
<EOL>|3600,3601
_|3601,3602
_|3602,3603
_|3603,3604
07|3605,3607
:|3607,3608
10PM|3608,3612
BLOOD|3613,3618
ALT|3619,3622
-|3622,3623
32|3623,3625
AST|3626,3629
-|3629,3630
40|3630,3632
AlkPhos|3633,3640
-|3640,3641
129|3641,3644
*|3644,3645
TotBili|3646,3653
-|3653,3654
0.2|3654,3657
<EOL>|3657,3658
_|3658,3659
_|3659,3660
_|3660,3661
07|3662,3664
:|3664,3665
10PM|3665,3669
BLOOD|3670,3675
cTropnT|3676,3683
-|3683,3684
0|3684,3685
.|3685,3686
01|3686,3688
<EOL>|3688,3689
_|3689,3690
_|3690,3691
_|3691,3692
07|3693,3695
:|3695,3696
30AM|3696,3700
BLOOD|3701,3706
Calcium|3707,3714
-|3714,3715
7|3715,3716
.|3716,3717
8|3717,3718
*|3718,3719
Phos|3720,3724
-|3724,3725
2|3725,3726
.|3726,3727
4|3727,3728
*|3728,3729
Mg|3730,3732
-|3732,3733
1.9|3733,3736
<EOL>|3736,3737
_|3737,3738
_|3738,3739
_|3739,3740
11|3741,3743
:|3743,3744
05PM|3744,3748
BLOOD|3749,3754
Type|3755,3759
-|3759,3760
ART|3760,3763
Temp|3764,3768
-|3768,3769
36.7|3769,3773
Tidal|3774,3779
V|3780,3781
-|3781,3782
300|3782,3785
PEEP|3786,3790
-|3790,3791
5|3791,3792
<EOL>|3793,3794
FiO2|3794,3798
-|3798,3799
50|3799,3801
pO2|3802,3805
-|3805,3806
133|3806,3809
*|3809,3810
pCO2|3811,3815
-|3815,3816
78|3816,3818
*|3818,3819
pH|3820,3822
-|3822,3823
7.37|3823,3827
calTCO2|3828,3835
-|3835,3836
47|3836,3838
*|3838,3839
Base|3840,3844
XS|3845,3847
-|3847,3848
15|3848,3850
<EOL>|3851,3852
Intubat|3852,3859
-|3859,3860
NOT|3860,3863
INTUBA|3864,3870
<EOL>|3870,3871
_|3871,3872
_|3872,3873
_|3873,3874
07|3875,3877
:|3877,3878
16PM|3878,3882
BLOOD|3883,3888
Lactate|3889,3896
-|3896,3897
1.5|3897,3900
<EOL>|3900,3901
<EOL>|3901,3902
Discharge|3902,3911
labs|3912,3916
:|3916,3917
<EOL>|3917,3918
_|3918,3919
_|3919,3920
_|3920,3921
06|3922,3924
:|3924,3925
30AM|3925,3929
BLOOD|3930,3935
WBC|3936,3939
-|3939,3940
4.9|3940,3943
RBC|3944,3947
-|3947,3948
2|3948,3949
.|3949,3950
67|3950,3952
*|3952,3953
Hgb|3954,3957
-|3957,3958
8|3958,3959
.|3959,3960
2|3960,3961
*|3961,3962
Hct|3963,3966
-|3966,3967
26|3967,3969
.|3969,3970
4|3970,3971
*|3971,3972
<EOL>|3973,3974
MCV|3974,3977
-|3977,3978
99|3978,3980
*|3980,3981
MCH|3982,3985
-|3985,3986
30.8|3986,3990
MCHC|3991,3995
-|3995,3996
31.2|3996,4000
RDW|4001,4004
-|4004,4005
15.0|4005,4009
Plt|4010,4013
_|4014,4015
_|4015,4016
_|4016,4017
<EOL>|4017,4018
_|4018,4019
_|4019,4020
_|4020,4021
06|4022,4024
:|4024,4025
30AM|4025,4029
BLOOD|4030,4035
Glucose|4036,4043
-|4043,4044
113|4044,4047
*|4047,4048
UreaN|4049,4054
-|4054,4055
6|4055,4056
Creat|4057,4062
-|4062,4063
0|4063,4064
.|4064,4065
3|4065,4066
*|4066,4067
Na|4068,4070
-|4070,4071
136|4071,4074
<EOL>|4075,4076
K|4076,4077
-|4077,4078
3.5|4078,4081
Cl|4082,4084
-|4084,4085
95|4085,4087
*|4087,4088
HCO3|4089,4093
-|4093,4094
37|4094,4096
*|4096,4097
AnGap|4098,4103
-|4103,4104
8|4104,4105
<EOL>|4105,4106
<EOL>|4106,4107
Micro|4107,4112
:|4112,4113
<EOL>|4113,4114
-|4114,4115
BCx|4115,4118
x2|4119,4121
(|4122,4123
NGTD|4123,4127
)|4127,4128
<EOL>|4128,4129
-|4129,4130
UCx|4130,4133
_|4134,4135
_|4135,4136
_|4136,4137
-|4138,4139
Yeast|4140,4145
,|4145,4146
no|4147,4149
bacterial|4150,4159
growth|4160,4166
<EOL>|4166,4167
-|4167,4168
Midline|4168,4175
tip|4176,4179
-|4180,4181
NGTD|4182,4186
<EOL>|4186,4187
-|4187,4188
C.|4188,4190
diff|4191,4195
PCR|4196,4199
-|4200,4201
neg|4202,4205
<EOL>|4205,4206
<EOL>|4206,4207
Imaging|4207,4214
:|4214,4215
<EOL>|4215,4216
<EOL>|4216,4217
_|4217,4218
_|4218,4219
_|4219,4220
:|4220,4221
CXR|4222,4225
:|4225,4226
IMPRESSION|4227,4237
:|4237,4238
No|4240,4242
significant|4243,4254
interval|4255,4263
change|4264,4270
with|4271,4275
<EOL>|4276,4277
bilateral|4277,4286
pleural|4287,4294
effusions|4295,4304
with|4305,4309
right|4310,4315
pigtail|4316,4323
catheter|4324,4332
in|4333,4335
the|4336,4339
<EOL>|4340,4341
lower|4341,4346
chest|4347,4352
.|4352,4353
Possible|4355,4363
small|4364,4369
right|4370,4375
apical|4376,4382
pneumothorax|4383,4395
.|4395,4396
<EOL>|4397,4398
<EOL>|4398,4399
_|4399,4400
_|4400,4401
_|4401,4402
:|4402,4403
CT|4404,4406
-|4406,4407
A|4407,4408
IMPRESSION|4409,4419
:|4419,4420
<EOL>|4421,4422
1|4422,4423
.|4423,4424
No|4426,4428
evidence|4429,4437
of|4438,4440
pulmonary|4441,4450
embolism|4451,4459
.|4459,4460
<EOL>|4461,4462
2.|4462,4464
Bilateral|4466,4475
pleural|4476,4483
effusions|4484,4493
,|4493,4494
small|4495,4500
to|4501,4503
moderate|4504,4512
on|4513,4515
the|4516,4519
left|4520,4524
,|4524,4525
<EOL>|4526,4527
decreased|4527,4536
<EOL>|4537,4538
since|4538,4543
the|4544,4547
most|4548,4552
recent|4553,4559
prior|4560,4565
examination|4566,4577
and|4578,4581
trace|4582,4587
on|4588,4590
the|4591,4594
right|4595,4600
,|4600,4601
<EOL>|4602,4603
markedly|4603,4611
<EOL>|4612,4613
decreased|4613,4622
compared|4623,4631
to|4632,4634
_|4635,4636
_|4636,4637
_|4637,4638
with|4639,4643
pigtail|4644,4651
catheter|4652,4660
noted|4661,4666
<EOL>|4667,4668
in|4668,4670
place|4671,4676
on|4677,4679
the|4680,4683
right|4684,4689
.|4689,4690
<EOL>|4693,4694
3.|4694,4696
Ascites|4698,4705
.|4705,4706
<EOL>|4707,4708
<EOL>|4708,4709
<EOL>|4710,4711
_|4734,4735
_|4735,4736
_|4736,4737
year|4738,4742
old|4743,4746
woman|4747,4752
,|4752,4753
recently|4754,4762
hospitalized|4763,4775
for|4776,4779
C.|4780,4782
Difficile|4783,4792
sepsis|4793,4799
<EOL>|4800,4801
and|4801,4804
shock|4805,4810
,|4810,4811
re-admitted|4812,4823
to|4824,4826
_|4827,4828
_|4828,4829
_|4829,4830
from|4831,4835
_|4836,4837
_|4837,4838
_|4838,4839
with|4840,4844
altered|4845,4852
<EOL>|4853,4854
mental|4854,4860
status|4861,4867
,|4867,4868
tachypnea|4869,4878
and|4879,4882
a|4883,4884
mild|4885,4889
respiratory|4890,4901
acidosis|4902,4910
.|4910,4911
<EOL>|4911,4912
<EOL>|4912,4913
#|4913,4914
Hypoxia|4914,4921
/|4921,4922
hypercarbia|4922,4933
:|4933,4934
She|4935,4938
initially|4939,4948
required|4949,4957
BiPAP|4958,4963
and|4964,4967
was|4968,4971
<EOL>|4972,4973
admitted|4973,4981
to|4982,4984
the|4985,4988
MICU|4989,4993
for|4994,4997
monitoring|4998,5008
of|5009,5011
her|5012,5015
respiratory|5016,5027
status|5028,5034
.|5034,5035
<EOL>|5037,5038
She|5038,5041
was|5042,5045
able|5046,5050
to|5051,5053
be|5054,5056
weaned|5057,5063
from|5064,5068
BiPAP|5069,5074
on|5075,5077
ICU|5078,5081
day|5082,5085
2|5086,5087
and|5088,5091
remained|5092,5100
<EOL>|5101,5102
on|5102,5104
2L|5105,5107
NC|5108,5110
at|5111,5113
the|5114,5117
time|5118,5122
of|5123,5125
discharge|5126,5135
.|5135,5136
Cause|5138,5143
of|5144,5146
her|5147,5150
respiratory|5151,5162
<EOL>|5163,5164
symptoms|5164,5172
is|5173,5175
unclear|5176,5183
,|5183,5184
but|5185,5188
may|5189,5192
be|5193,5195
due|5196,5199
to|5200,5202
hypoventilation|5203,5218
from|5219,5223
<EOL>|5224,5225
somnolence|5225,5235
related|5236,5243
to|5244,5246
oversedation|5247,5259
with|5260,5264
Zyprexa|5265,5272
.|5272,5273
Zyprexa|5275,5282
was|5283,5286
<EOL>|5287,5288
held|5288,5292
at|5293,5295
the|5296,5299
time|5300,5304
of|5305,5307
discharge|5308,5317
.|5317,5318
CTA|5320,5323
Chest|5324,5329
was|5330,5333
negative|5334,5342
for|5343,5346
PE|5347,5349
<EOL>|5350,5351
and|5351,5354
showed|5355,5361
no|5362,5364
clear|5365,5370
evidence|5371,5379
of|5380,5382
pneumonia|5383,5392
.|5392,5393
She|5395,5398
was|5399,5402
initially|5403,5412
<EOL>|5413,5414
started|5414,5421
on|5422,5424
HCAP|5425,5429
antibiotics|5430,5441
with|5442,5446
vanc|5447,5451
/|5451,5452
cefepime|5452,5460
which|5461,5466
were|5467,5471
<EOL>|5472,5473
stopped|5473,5480
on|5481,5483
HD|5484,5486
4|5487,5488
prior|5489,5494
to|5495,5497
discharge|5498,5507
given|5508,5513
that|5514,5518
all|5519,5522
cultures|5523,5531
were|5532,5536
<EOL>|5537,5538
negative|5538,5546
and|5547,5550
there|5551,5556
was|5557,5560
no|5561,5563
consolidation|5564,5577
on|5578,5580
imaging|5581,5588
.|5588,5589
<EOL>|5590,5591
<EOL>|5591,5592
#|5592,5593
Delirium|5594,5602
:|5602,5603
Likely|5604,5610
multifactorial|5611,5625
,|5625,5626
but|5627,5630
thought|5631,5638
to|5639,5641
be|5642,5644
related|5645,5652
to|5653,5655
<EOL>|5656,5657
oversedation|5657,5669
from|5670,5674
Zyprexa|5675,5682
.|5682,5683
There|5685,5690
was|5691,5694
no|5695,5697
evidence|5698,5706
of|5707,5709
infection|5710,5719
<EOL>|5720,5721
and|5721,5724
antibiotics|5725,5736
were|5737,5741
quickly|5742,5749
stopped|5750,5757
as|5758,5760
described|5761,5770
above|5771,5776
.|5776,5777
UA|5779,5781
was|5782,5785
<EOL>|5786,5787
dirty|5787,5792
,|5792,5793
but|5794,5797
UCx|5798,5801
was|5802,5805
negative|5806,5814
x2|5815,5817
(|5818,5819
grew|5819,5823
only|5824,5828
yeast|5829,5834
)|5834,5835
and|5836,5839
she|5840,5843
had|5844,5847
no|5848,5850
<EOL>|5851,5852
urinary|5852,5859
symptoms|5860,5868
.|5868,5869
Most|5871,5875
of|5876,5878
her|5879,5882
mental|5883,5889
status|5890,5896
changes|5897,5904
were|5905,5909
<EOL>|5910,5911
probably|5911,5919
related|5920,5927
to|5928,5930
her|5931,5934
sedationg|5935,5944
medications|5945,5956
and|5957,5960
hypercarbia|5961,5972
at|5973,5975
<EOL>|5976,5977
admission|5977,5986
,|5986,5987
which|5988,5993
improved|5994,6002
with|6003,6007
BiPAP|6008,6013
and|6014,6017
holding|6018,6025
her|6026,6029
<EOL>|6030,6031
antipsychotics|6031,6045
.|6045,6046
<EOL>|6046,6047
<EOL>|6047,6048
#|6048,6049
C|6050,6051
Diff|6052,6056
Colitis|6057,6064
:|6064,6065
Recently|6066,6074
admitted|6075,6083
for|6084,6087
C.|6088,6090
diff|6091,6095
colitis|6096,6103
with|6104,6108
<EOL>|6109,6110
sepsis|6110,6116
.|6116,6117
Repeat|6118,6124
C|6125,6126
Diff|6127,6131
PCR|6132,6135
was|6136,6139
negative|6140,6148
during|6149,6155
this|6156,6160
<EOL>|6161,6162
hospitalization|6162,6177
.|6177,6178
She|6179,6182
continued|6183,6192
to|6193,6195
have|6196,6200
high|6201,6205
volume|6206,6212
stool|6213,6218
output|6219,6225
<EOL>|6226,6227
and|6227,6230
Flexiseal|6231,6240
is|6241,6243
in|6244,6246
place|6247,6252
for|6253,6256
skin|6257,6261
ulceration|6262,6272
.|6272,6273
ID|6275,6277
was|6278,6281
curbsided|6282,6291
<EOL>|6292,6293
regarding|6293,6302
vanco|6303,6308
course|6309,6315
given|6316,6321
that|6322,6326
she|6327,6330
received|6331,6339
a|6340,6341
few|6342,6345
days|6346,6350
of|6351,6353
<EOL>|6354,6355
HCAP|6355,6359
antibotics|6360,6370
and|6371,6374
her|6375,6378
PO|6379,6381
vanco|6382,6387
was|6388,6391
changed|6392,6399
to|6400,6402
125mg|6403,6408
q6h|6409,6412
for|6413,6416
7|6417,6418
<EOL>|6419,6420
days|6420,6424
after|6425,6430
stopping|6431,6439
IV|6440,6442
vanc|6443,6447
/|6447,6448
cefepime|6448,6456
(|6457,6458
D7|6458,6460
will|6461,6465
be|6466,6468
_|6469,6470
_|6470,6471
_|6471,6472
.|6472,6473
<EOL>|6475,6476
Flexiseal|6476,6485
in|6486,6488
place|6489,6494
at|6495,6497
discharge|6498,6507
.|6507,6508
<EOL>|6508,6509
<EOL>|6509,6510
#|6510,6511
Anemia|6512,6518
:|6518,6519
Patient|6520,6527
with|6528,6532
guaiac|6533,6539
positive|6540,6548
stools|6549,6555
this|6556,6560
admission|6561,6570
,|6570,6571
<EOL>|6572,6573
new|6573,6576
from|6577,6581
past|6582,6586
admission|6587,6596
.|6596,6597
Felt|6599,6603
to|6604,6606
be|6607,6609
secondary|6610,6619
to|6620,6622
sloughing|6623,6632
and|6633,6636
<EOL>|6637,6638
mucosal|6638,6645
oozing|6646,6652
secondary|6653,6662
to|6663,6665
C|6666,6667
diff|6668,6672
.|6672,6673
Normal|6674,6680
lactate|6681,6688
on|6689,6691
admission|6692,6701
<EOL>|6702,6703
and|6703,6706
benign|6707,6713
abdominal|6714,6723
exam|6724,6728
.|6728,6729
Hct|6731,6734
has|6735,6738
been|6739,6743
variable|6744,6752
recently|6753,6761
,|6761,6762
but|6763,6766
<EOL>|6767,6768
fairly|6768,6774
stable|6775,6781
,|6781,6782
although|6783,6791
still|6792,6797
markedly|6798,6806
below|6807,6812
her|6813,6816
baseline|6817,6825
of|6826,6828
low|6829,6832
<EOL>|6833,6834
to|6834,6836
mid|6837,6840
_|6841,6842
_|6842,6843
_|6843,6844
.|6844,6845
<EOL>|6845,6846
<EOL>|6846,6847
#|6847,6848
Bilateral|6849,6858
pleural|6859,6866
effusions|6867,6876
:|6876,6877
Noted|6878,6883
to|6884,6886
have|6887,6891
bilateral|6892,6901
pleural|6902,6909
<EOL>|6910,6911
effusions|6911,6920
last|6921,6925
hospitalization|6926,6941
in|6942,6944
setting|6945,6952
of|6953,6955
massive|6956,6963
fluid|6964,6969
<EOL>|6970,6971
resuscitation|6971,6984
,|6984,6985
right|6986,6991
pleural|6992,6999
pigtail|7000,7007
catheter|7008,7016
removed|7017,7024
this|7025,7029
<EOL>|7030,7031
admission|7031,7040
in|7041,7043
the|7044,7047
MICU|7048,7052
.|7052,7053
She|7054,7057
is|7058,7060
still|7061,7066
volume|7067,7073
overloaded|7074,7084
on|7085,7087
exam|7088,7092
,|7092,7093
<EOL>|7094,7095
but|7095,7098
her|7099,7102
bicarb|7103,7109
remained|7110,7118
elevated|7119,7127
,|7127,7128
and|7129,7132
she|7133,7136
was|7137,7140
not|7141,7144
given|7145,7150
any|7151,7154
<EOL>|7155,7156
further|7156,7163
diuresis|7164,7172
.|7172,7173
The|7175,7178
elevated|7179,7187
bicarb|7188,7194
is|7195,7197
also|7198,7202
be|7203,7205
partially|7206,7215
due|7216,7219
<EOL>|7220,7221
to|7221,7223
compensation|7224,7236
from|7237,7241
her|7242,7245
respiratory|7246,7257
acidosis|7258,7266
.|7266,7267
<EOL>|7267,7268
<EOL>|7268,7269
#|7269,7270
Volume|7271,7277
overload|7278,7286
:|7286,7287
She|7288,7291
has|7292,7295
some|7296,7300
diastolic|7301,7310
dysfunction|7311,7322
and|7323,7326
has|7327,7330
2|7331,7332
+|7332,7333
<EOL>|7334,7335
MR|7335,7337
on|7338,7340
_|7341,7342
_|7342,7343
_|7343,7344
.|7344,7345
She|7346,7349
continues|7350,7359
to|7360,7362
appear|7363,7369
total|7370,7375
body|7376,7380
overloaded|7381,7391
,|7391,7392
likely|7393,7399
<EOL>|7400,7401
in|7401,7403
setting|7404,7411
of|7412,7414
volume|7415,7421
resuscitation|7422,7435
on|7436,7438
prior|7439,7444
admission|7445,7454
for|7455,7458
<EOL>|7459,7460
sepsis|7460,7466
,|7466,7467
but|7468,7471
with|7472,7476
contraction|7477,7488
alkalosis|7489,7498
currently|7499,7508
,|7508,7509
so|7510,7512
further|7513,7520
<EOL>|7521,7522
diuresis|7522,7530
was|7531,7534
held|7535,7539
as|7540,7542
above|7543,7548
.|7548,7549
Consider|7551,7559
further|7560,7567
diuresis|7568,7576
once|7577,7581
<EOL>|7582,7583
hypercarbia|7583,7594
improves|7595,7603
and|7604,7607
bicarb|7608,7614
trends|7615,7621
down|7622,7626
.|7626,7627
<EOL>|7629,7630
<EOL>|7630,7631
#|7631,7632
Hypothyroidism|7633,7647
:|7647,7648
Continued|7649,7658
on|7659,7661
levothyroxine|7662,7675
50|7676,7678
mcg|7679,7682
daily|7683,7688
<EOL>|7689,7690
<EOL>|7691,7692
#|7692,7693
Hypertension|7694,7706
:|7706,7707
Patient|7708,7715
was|7716,7719
previously|7720,7730
on|7731,7733
lisinopril|7734,7744
which|7745,7750
was|7751,7754
<EOL>|7755,7756
held|7756,7760
since|7761,7766
last|7767,7771
admission|7772,7781
in|7782,7784
setting|7785,7792
of|7793,7795
sepsis|7796,7802
and|7803,7806
relative|7807,7815
<EOL>|7816,7817
hypotension|7817,7828
.|7828,7829
She|7831,7834
remained|7835,7843
normotensive|7844,7856
<EOL>|7856,7857
<EOL>|7857,7858
#|7858,7859
GERD|7860,7864
:|7864,7865
Patient|7866,7873
previously|7874,7884
on|7885,7887
omeprazole|7888,7898
last|7899,7903
hospitalization|7904,7919
,|7919,7920
<EOL>|7921,7922
which|7922,7927
was|7928,7931
stopped|7932,7939
after|7940,7945
C.|7946,7948
diff|7949,7953
came|7954,7958
back|7959,7963
positive|7964,7972
,|7972,7973
and|7974,7977
she|7978,7981
was|7982,7985
<EOL>|7986,7987
transitioned|7987,7999
to|8000,8002
H2|8003,8005
blocker|8006,8013
for|8014,8017
GI|8018,8020
prophylaxis|8021,8032
but|8033,8036
this|8037,8041
was|8042,8045
<EOL>|8046,8047
stopped|8047,8054
again|8055,8060
when|8061,8065
she|8066,8069
became|8070,8076
delirious|8077,8086
last|8087,8091
hospitalization|8092,8107
.|8107,8108
<EOL>|8110,8111
She|8111,8114
remains|8115,8122
off|8123,8126
H2|8127,8129
blocker|8130,8137
at|8138,8140
discharge|8141,8150
because|8151,8158
of|8159,8161
concern|8162,8169
that|8170,8174
<EOL>|8175,8176
it|8176,8178
may|8179,8182
be|8183,8185
contributing|8186,8198
to|8199,8201
her|8202,8205
AMS|8206,8209
.|8209,8210
<EOL>|8210,8211
<EOL>|8211,8212
#|8212,8213
Code|8214,8218
status|8219,8225
this|8226,8230
admission|8231,8240
:|8240,8241
FULL|8242,8246
<EOL>|8246,8247
<EOL>|8247,8248
#|8248,8249
Transitional|8250,8262
issues|8263,8269
:|8269,8270
<EOL>|8270,8271
-|8271,8272
Foley|8272,8277
was|8278,8281
removed|8282,8289
_|8290,8291
_|8291,8292
_|8292,8293
and|8294,8297
she|8298,8301
has|8302,8305
not|8306,8309
voided|8310,8316
as|8317,8319
of|8320,8322
discharge|8323,8332
,|8332,8333
<EOL>|8334,8335
may|8335,8338
need|8339,8343
Foley|8344,8349
replaced|8350,8358
if|8359,8361
she|8362,8365
is|8366,8368
unable|8369,8375
to|8376,8378
void|8379,8383
<EOL>|8383,8384
-|8384,8385
Would|8385,8390
restart|8391,8398
diuresis|8399,8407
when|8408,8412
bicarb|8413,8419
trends|8420,8426
down|8427,8431
<EOL>|8431,8432
-|8432,8433
Continue|8433,8441
PO|8442,8444
vanco|8445,8450
125mg|8451,8456
q6h|8457,8460
through|8461,8468
_|8469,8470
_|8470,8471
_|8471,8472
<EOL>|8472,8473
-|8473,8474
Please|8474,8480
follow|8481,8487
Hct|8488,8491
daily|8492,8497
given|8498,8503
melanotic|8504,8513
stools|8514,8520
,|8520,8521
should|8522,8528
resolve|8529,8536
<EOL>|8537,8538
as|8538,8540
her|8541,8544
C.|8545,8547
diff|8548,8552
resolves|8553,8561
<EOL>|8561,8562
-|8562,8563
Midline|8563,8570
removed|8571,8578
_|8579,8580
_|8580,8581
_|8581,8582
<EOL>|8582,8583
-|8583,8584
Pigtail|8584,8591
catheter|8592,8600
removed|8601,8608
this|8609,8613
admission|8614,8623
<EOL>|8623,8624
-|8624,8625
F|8625,8626
/|8626,8627
u|8627,8628
pending|8629,8636
BCx|8637,8640
,|8640,8641
catheter|8642,8650
tip|8651,8654
cx|8655,8657
<EOL>|8657,8658
<EOL>|8659,8660
Medications|8660,8671
on|8672,8674
Admission|8675,8684
:|8684,8685
<EOL>|8685,8686
Medications|8686,8697
at|8698,8700
_|8701,8702
_|8702,8703
_|8703,8704
:|8704,8705
<EOL>|8705,8706
fluticasone|8706,8717
50|8718,8720
mcg|8721,8724
nasal|8725,8730
spray|8731,8736
_|8737,8738
_|8738,8739
_|8739,8740
puffs|8741,8746
BID|8747,8750
PRN|8751,8754
<EOL>|8755,8756
levothyroxine|8756,8769
50|8770,8772
mcg|8773,8776
dialy|8777,8782
<EOL>|8782,8783
acetaminophen|8783,8796
650|8797,8800
mg|8801,8803
Q4H|8804,8807
PRN|8808,8811
pain|8812,8816
<EOL>|8816,8817
polyvinyl|8817,8826
alcohol|8827,8834
1.4|8835,8838
%|8838,8839
drops|8840,8845
every|8846,8851
4H|8852,8854
PRN|8855,8858
dry|8859,8862
eyes|8863,8867
<EOL>|8867,8868
heparin|8868,8875
line|8876,8880
flush|8881,8886
<EOL>|8886,8887
Humalog|8887,8894
insulin|8895,8902
sliding|8903,8910
scale|8911,8916
<EOL>|8916,8917
Miconazole|8917,8927
nitrate|8928,8935
2|8936,8937
%|8937,8938
powder|8939,8945
,|8945,8946
1|8947,8948
application|8949,8960
TID|8961,8964
PRN|8965,8968
rash|8969,8973
<EOL>|8973,8974
ondansetron|8974,8985
4|8986,8987
mg|8988,8990
IV|8991,8993
Q8H|8994,8997
PRN|8998,9001
nausea|9002,9008
<EOL>|9008,9009
Olanzapine|9009,9019
2.5|9020,9023
mg|9024,9026
PO|9027,9029
daily|9030,9035
and|9036,9039
qHS|9040,9043
PRN|9044,9047
anxiety|9048,9055
/|9055,9056
insomnia|9056,9064
<EOL>|9064,9065
Vancomycin|9065,9075
500|9076,9079
mg|9080,9082
Q6H|9083,9086
planned|9087,9094
through|9095,9102
_|9103,9104
_|9104,9105
_|9105,9106
<EOL>|9106,9107
<EOL>|9107,9108
<EOL>|9109,9110
Discharge|9110,9119
Medications|9120,9131
:|9131,9132
<EOL>|9132,9133
1.|9133,9135
fluticasone|9136,9147
50|9148,9150
mcg|9151,9154
/|9154,9155
actuation|9155,9164
Spray|9165,9170
,|9170,9171
Suspension|9172,9182
Sig|9183,9186
:|9186,9187
_|9188,9189
_|9189,9190
_|9190,9191
puffs|9192,9197
<EOL>|9198,9199
Nasal|9199,9204
twice|9205,9210
a|9211,9212
day|9213,9216
as|9217,9219
needed|9220,9226
for|9227,9230
allergies|9231,9240
.|9240,9241
<EOL>|9243,9244
2.|9244,9246
levothyroxine|9247,9260
50|9261,9263
mcg|9264,9267
Tablet|9268,9274
Sig|9275,9278
:|9278,9279
One|9280,9283
(|9284,9285
1|9285,9286
)|9286,9287
Tablet|9288,9294
PO|9295,9297
DAILY|9298,9303
<EOL>|9304,9305
(|9305,9306
Daily|9306,9311
)|9311,9312
.|9312,9313
<EOL>|9315,9316
3.|9316,9318
acetaminophen|9319,9332
325|9333,9336
mg|9337,9339
Tablet|9340,9346
Sig|9347,9350
:|9350,9351
_|9352,9353
_|9353,9354
_|9354,9355
Tablets|9356,9363
PO|9364,9366
every|9367,9372
four|9373,9377
<EOL>|9378,9379
(|9379,9380
4|9380,9381
)|9381,9382
hours|9383,9388
as|9389,9391
needed|9392,9398
for|9399,9402
fever|9403,9408
or|9409,9411
pain|9412,9416
.|9416,9417
<EOL>|9419,9420
4.|9420,9422
polyvinyl|9423,9432
alcohol|9433,9440
1.4|9441,9444
%|9445,9446
Drops|9447,9452
Sig|9453,9456
:|9456,9457
One|9458,9461
(|9462,9463
1|9463,9464
)|9464,9465
drop|9466,9470
Ophthalmic|9471,9481
<EOL>|9482,9483
every|9483,9488
four|9489,9493
(|9494,9495
4|9495,9496
)|9496,9497
hours|9498,9503
as|9504,9506
needed|9507,9513
for|9514,9517
dry|9518,9521
eyes|9522,9526
.|9526,9527
<EOL>|9529,9530
5.|9530,9532
insulin|9533,9540
lispro|9541,9547
100|9548,9551
unit|9552,9556
/|9556,9557
mL|9557,9559
Solution|9560,9568
Sig|9569,9572
:|9572,9573
Sliding|9574,9581
scale|9582,9587
units|9588,9593
<EOL>|9594,9595
Subcutaneous|9595,9607
three|9608,9613
times|9614,9619
a|9620,9621
day|9622,9625
:|9625,9626
150|9627,9630
-|9630,9631
200|9631,9634
-|9635,9636
2|9637,9638
units|9639,9644
;|9644,9645
201|9646,9649
-|9649,9650
250|9650,9653
-|9654,9655
4|9656,9657
<EOL>|9658,9659
units|9659,9664
;|9664,9665
251|9666,9669
-|9669,9670
300|9670,9673
-|9674,9675
6|9676,9677
units|9678,9683
;|9683,9684
301|9685,9688
-|9688,9689
350|9689,9692
-|9693,9694
8|9695,9696
units|9697,9702
;|9702,9703
351|9704,9707
-|9707,9708
400|9708,9711
-|9712,9713
10|9714,9716
units|9717,9722
;|9722,9723
<EOL>|9724,9725
over|9725,9729
400|9730,9733
-|9734,9735
10|9736,9738
units|9739,9744
and|9745,9748
call|9749,9753
MD|9754,9756
.|9756,9757
<EOL>|9759,9760
6.|9760,9762
miconazole|9763,9773
nitrate|9774,9781
2|9782,9783
%|9784,9785
Powder|9786,9792
Sig|9793,9796
:|9796,9797
One|9798,9801
(|9802,9803
1|9803,9804
)|9804,9805
application|9806,9817
<EOL>|9818,9819
Topical|9819,9826
three|9827,9832
times|9833,9838
a|9839,9840
day|9841,9844
as|9845,9847
needed|9848,9854
for|9855,9858
rash|9859,9863
.|9863,9864
<EOL>|9866,9867
7.|9867,9869
vancomycin|9870,9880
125|9881,9884
mg|9885,9887
Capsule|9888,9895
Sig|9896,9899
:|9899,9900
One|9901,9904
(|9905,9906
1|9906,9907
)|9907,9908
Capsule|9909,9916
PO|9917,9919
Q6H|9920,9923
(|9924,9925
every|9925,9930
<EOL>|9931,9932
6|9932,9933
hours|9934,9939
)|9939,9940
for|9941,9944
7|9945,9946
days|9947,9951
:|9951,9952
Last|9953,9957
dose|9958,9962
on|9963,9965
_|9966,9967
_|9967,9968
_|9968,9969
.|9969,9970
<EOL>|9972,9973
8.|9973,9975
heparin|9976,9983
(|9984,9985
porcine|9985,9992
)|9992,9993
5,000|9994,9999
unit|10000,10004
/|10004,10005
mL|10005,10007
Solution|10008,10016
Sig|10017,10020
:|10020,10021
5000|10022,10026
(|10027,10028
5000|10028,10032
)|10032,10033
<EOL>|10034,10035
units|10035,10040
Injection|10041,10050
three|10051,10056
times|10057,10062
a|10063,10064
day|10065,10068
.|10068,10069
<EOL>|10071,10072
9.|10072,10074
albuterol|10075,10084
sulfate|10085,10092
2.5|10093,10096
mg|10097,10099
/|10100,10101
3|10101,10102
mL|10103,10105
(|10106,10107
0.083|10107,10112
%|10113,10114
)|10114,10115
Solution|10116,10124
for|10125,10128
<EOL>|10129,10130
Nebulization|10130,10142
Sig|10143,10146
:|10146,10147
One|10148,10151
(|10152,10153
1|10153,10154
)|10154,10155
neb|10156,10159
Inhalation|10160,10170
every|10171,10176
four|10177,10181
(|10182,10183
4|10183,10184
)|10184,10185
hours|10186,10191
as|10192,10194
<EOL>|10195,10196
needed|10196,10202
for|10203,10206
shortness|10207,10216
of|10217,10219
breath|10220,10226
or|10227,10229
wheezing|10230,10238
.|10238,10239
<EOL>|10241,10242
10.|10242,10245
ipratropium|10246,10257
bromide|10258,10265
0.02|10266,10270
%|10271,10272
Solution|10273,10281
Sig|10282,10285
:|10285,10286
One|10287,10290
(|10291,10292
1|10292,10293
)|10293,10294
neb|10295,10298
<EOL>|10299,10300
Inhalation|10300,10310
every|10311,10316
six|10317,10320
(|10321,10322
6|10322,10323
)|10323,10324
hours|10325,10330
as|10331,10333
needed|10334,10340
for|10341,10344
shortness|10345,10354
of|10355,10357
breath|10358,10364
<EOL>|10365,10366
or|10366,10368
wheezing|10369,10377
.|10377,10378
<EOL>|10380,10381
<EOL>|10381,10382
<EOL>|10383,10384
Discharge|10384,10393
Disposition|10394,10405
:|10405,10406
<EOL>|10406,10407
Extended|10407,10415
Care|10416,10420
<EOL>|10420,10421
<EOL>|10422,10423
Facility|10423,10431
:|10431,10432
<EOL>|10432,10433
_|10433,10434
_|10434,10435
_|10435,10436
<EOL>|10436,10437
<EOL>|10438,10439
Discharge|10439,10448
Diagnosis|10449,10458
:|10458,10459
<EOL>|10459,10460
Altered|10479,10486
mental|10487,10493
status|10494,10500
<EOL>|10500,10501
Hypoxia|10501,10508
<EOL>|10508,10509
<EOL>|10509,10510
Secondary|10510,10519
diagnoses|10520,10529
:|10529,10530
<EOL>|10530,10531
Clostridium|10531,10542
difficule|10543,10552
<EOL>|10552,10553
<EOL>|10553,10554
<EOL>|10555,10556
Mental|10577,10583
Status|10584,10590
:|10590,10591
Confused|10592,10600
-|10601,10602
sometimes|10603,10612
.|10612,10613
<EOL>|10613,10614
Level|10614,10619
of|10620,10622
Consciousness|10623,10636
:|10636,10637
Lethargic|10638,10647
but|10648,10651
arousable|10652,10661
.|10661,10662
<EOL>|10662,10663
Activity|10663,10671
Status|10672,10678
:|10678,10679
Out|10680,10683
of|10684,10686
Bed|10687,10690
with|10691,10695
assistance|10696,10706
to|10707,10709
chair|10710,10715
or|10716,10718
<EOL>|10719,10720
wheelchair|10720,10730
.|10730,10731
<EOL>|10731,10732
<EOL>|10732,10733
<EOL>|10734,10735
Dear|10759,10763
Ms.|10764,10767
_|10768,10769
_|10769,10770
_|10770,10771
,|10771,10772
<EOL>|10772,10773
<EOL>|10773,10774
It|10774,10776
was|10777,10780
a|10781,10782
pleasure|10783,10791
taking|10792,10798
care|10799,10803
of|10804,10806
you|10807,10810
during|10811,10817
your|10818,10822
admission|10823,10832
to|10833,10835
<EOL>|10836,10837
_|10837,10838
_|10838,10839
_|10839,10840
for|10841,10844
hypoxia|10845,10852
/|10852,10853
hypercarbia|10853,10864
and|10865,10868
altered|10869,10876
mental|10877,10883
status|10884,10890
.|10890,10891
Your|10893,10897
<EOL>|10898,10899
mental|10899,10905
status|10906,10912
improved|10913,10921
once|10922,10926
we|10927,10929
stopped|10930,10937
your|10938,10942
Zyprexa|10943,10950
and|10951,10954
your|10955,10959
<EOL>|10960,10961
breathing|10961,10970
improved|10971,10979
.|10979,10980
We|10982,10984
looked|10985,10991
for|10992,10995
an|10996,10998
infection|10999,11008
but|11009,11012
were|11013,11017
not|11018,11021
<EOL>|11022,11023
able|11023,11027
to|11028,11030
find|11031,11035
a|11036,11037
clear|11038,11043
source|11044,11050
.|11050,11051
You|11053,11056
received|11057,11065
a|11066,11067
few|11068,11071
days|11072,11076
of|11077,11079
<EOL>|11080,11081
antibiotics|11081,11092
while|11093,11098
your|11099,11103
cultures|11104,11112
were|11113,11117
pending|11118,11125
.|11125,11126
You|11128,11131
will|11132,11136
continue|11137,11145
<EOL>|11146,11147
PO|11147,11149
vanco|11150,11155
for|11156,11159
an|11160,11162
additional|11163,11173
7|11174,11175
days|11176,11180
.|11180,11181
<EOL>|11181,11182
<EOL>|11182,11183
The|11183,11186
following|11187,11196
changes|11197,11204
were|11205,11209
made|11210,11214
to|11215,11217
your|11218,11222
medications|11223,11234
:|11234,11235
<EOL>|11235,11236
CHANGE|11236,11242
vancomycin|11243,11253
125mg|11254,11259
by|11260,11262
mouth|11263,11268
every|11269,11274
6|11275,11276
hours|11277,11282
for|11283,11286
7|11287,11288
days|11289,11293
(|11294,11295
last|11295,11299
<EOL>|11300,11301
dose|11301,11305
_|11306,11307
_|11307,11308
_|11308,11309
<EOL>|11309,11310
START|11310,11315
albuterol|11316,11325
neb|11326,11329
every|11330,11335
4|11336,11337
hours|11338,11343
as|11344,11346
needed|11347,11353
for|11354,11357
SOB|11358,11361
/|11361,11362
wheezing|11362,11370
<EOL>|11370,11371
START|11371,11376
ipratropium|11377,11388
neb|11389,11392
every|11393,11398
6|11399,11400
hours|11401,11406
as|11407,11409
needed|11410,11416
for|11417,11420
SOB|11421,11424
/|11424,11425
wheezing|11425,11433
<EOL>|11433,11434
STOP|11434,11438
Zyprexa|11439,11446
<EOL>|11446,11447
<EOL>|11448,11449
Followup|11449,11457
Instructions|11458,11470
:|11470,11471
<EOL>|11471,11472
_|11472,11473
_|11473,11474
_|11474,11475
<EOL>|11475,11476

