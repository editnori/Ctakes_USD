CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Pharmaceutical Preparations|Drug|false|false||MEDICINEnull|Medicine|Title|false|false||MEDICINEnull|Known|Modifier|false|false||Knownnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|Adverse reaction to drug|Finding|true|false||Adverse Drug Reactionsnull|Adverse reaction to drug|Finding|true|false||Drug Reactionsnull|Pharmaceutical Preparations|Drug|false|false||Drug
null|Pharmacologic Substance|Drug|false|false||Drugnull|Drug problem|Finding|false|false||Drugnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Swelling of lower limb|Finding|false|false|C0015385;C0023216;C1548802|Lower extremity swellingnull|Lower Extremity|Anatomy|false|false|C0013604;C0038999;C0581394;C0158369;C2003888|Lower extremitynull|Body Site Modifier - Lower|Anatomy|false|false|C2003888;C0013604;C0038999;C0158369;C0581394|Lowernull|Lower (action)|Event|false|false|C1548802;C0023216|Lowernull|Lower - spatial qualifier|Modifier|false|false||Lowernull|Swelling of limb|Finding|false|false|C0015385;C0023216;C1548802|extremity swellingnull|Limb structure|Anatomy|false|false|C0581394;C0158369;C0013604;C0038999|extremitynull|Swelling|Finding|false|false|C0023216;C1548802;C0015385|swelling
null|Edema|Finding|false|false|C0023216;C1548802;C0015385|swellingnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|on warfarin|Procedure|false|false||on warfarinnull|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarinnull|Recent|Time|false|false||recentnull|Steroid [EPC]|Drug|false|false||steroid
null|Steroids|Drug|false|false||steroid
null|Steroids|Drug|false|false||steroidnull|Physiologic pulse|Finding|false|false||pulsenull|Pulse taking|Procedure|false|false||pulsenull|Pulse Rate|Attribute|false|false||pulsenull|Pulse phenomenon|Phenomenon|false|false||pulsenull|Swelling|Finding|false|false||swollennull|Pain|Finding|false|false|C0003086|painfulnull|Ankle|Anatomy|false|false|C0030193|anklesnull|Complaint (finding)|Finding|true|false||complaintsnull|wife|Subject|false|false||wifenull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|Unable to walk (finding)|Finding|false|false||inability to walknull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|History of fall|Finding|false|false||a fallnull|Falls|Finding|false|false||fallnull|Autumn|Time|false|false||fallnull|Bathtub|Device|false|false||bathtubnull|1 Week|Time|false|false||one weeknull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|FBXW7 wt Allele|Finding|false|false||ago
null|FBXW7 gene|Finding|false|false||agonull|Problems with head|Disorder|true|false|C0018670;C0152336|headnull|Procedure on head|Procedure|true|false|C0018670;C0152336|headnull|Structure of head of caudate nucleus|Anatomy|false|false|C0362076;C0038452;C0876917|head
null|Head|Anatomy|false|false|C0362076;C0038452;C0876917|headnull|Head Device|Device|true|false||headnull|Strikes, Employee|Event|true|false|C0018670;C0152336|strikenull|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Local Remote Control State - Local|Finding|false|false||localnull|Local|Modifier|false|false||localnull|Spinal Fractures|Disorder|false|false|C0549207|vertebral fracturenull|Bone structure of spine|Anatomy|false|false|C0016658;C0080179|vertebralnull|Fracture|Disorder|false|false|C0549207|fracturenull|Back braces|Device|false|false||back bracenull|Application of brace (procedure)|Procedure|false|false||bracenull|Braces - Orthopedic appliances|Device|false|false||brace
null|Braces - garment|Device|false|false||bracenull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|swelling of both ankles|Finding|false|false|C0003086;C0003087;C4284979|bilateral ankle swellingnull|Bilateral|Modifier|false|false||bilateralnull|Ankle edema (finding)|Finding|false|false|C0003086;C0003087;C4284979|ankle swellingnull|Lower extremity>Ankle|Anatomy|false|false|C0235439;C2109101|ankle
null|Ankle|Anatomy|false|false|C0235439;C2109101|ankle
null|Ankle joint structure|Anatomy|false|false|C0235439;C2109101|anklenull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|3+ pitting edema|Finding|false|false||3+ pitting edemanull|Pitting edema|Finding|false|false||pitting edemanull|Pitting|Finding|false|false||pittingnull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Cold brand of chlorpheniramine-phenylpropanolamine|Drug|false|false||cold
null|Cold brand of chlorpheniramine-phenylpropanolamine|Drug|false|false||coldnull|Common Cold|Disorder|false|false||cold
null|Chronic Obstructive Airway Disease|Disorder|false|false||coldnull|Cold Sensation|Finding|false|false||coldnull|Cold Therapy|Procedure|false|false||coldnull|Cold Temperature|Phenomenon|false|false||coldnull|Mottling|Finding|false|false|C0040357;C4299090|mottlednull|Lower extremity>Toes|Anatomy|false|false|C0302133|toes
null|Toes|Anatomy|false|false|C0302133|toesnull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false||pulsesnull|Sensory Disorders|Disorder|true|false||sensory disturbancesnull|Sensory (qualifier value)|Modifier|false|false||sensorynull|NPPB protein, human|Drug|false|false||BNP
null|NPPB protein, human|Drug|false|false||BNP
null|nesiritide|Drug|false|false||BNP
null|nesiritide|Drug|false|false||BNP
null|nesiritide|Drug|false|false||BNPnull|NPPB wt Allele|Finding|false|false||BNP
null|NPPB gene|Finding|false|false||BNPnull|Brain natriuretic peptide measurement|Procedure|false|false||BNPnull|Plain chest X-ray|Procedure|false|false||CXRnull|Pulmonary Edema|Finding|false|false|C0024109|pulmonary edemanull|Pulmonary (intended site)|Finding|false|false|C0024109|pulmonarynull|Lung|Anatomy|false|false|C4522268;C2707265;C0013604;C0034063|pulmonarynull|null|Attribute|false|false|C0024109|pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Edema|Finding|false|false|C0024109|edemanull|null|Attribute|false|false||edemanull|Negative|Finding|false|false|C5239664|negative fornull|Rh Negative Blood Group|Finding|false|false|C5239664|negative
null|Negative|Finding|false|false|C5239664|negative
null|Negative Finding|Finding|false|false|C5239664|negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Deep thrombophlebitis|Disorder|false|false|C5239664|DVT
null|Deep Vein Thrombosis|Disorder|false|false|C5239664|DVTnull|area DVT|Anatomy|false|false|C2926618;C0205160;C0149871;C0151950;C2699077;C0205160;C1513916|DVTnull|null|Attribute|false|false|C5239664|DVTnull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Pericardial effusion|Disorder|true|false|C0031050;C0442031;C3498924|pericardial effusionnull|Pericardial effusion body substance|Finding|true|false|C0031050;C0442031|pericardial effusionnull|Pericardial (qualifier value)|Anatomy|false|false|C2317432;C1546613;C0013687;C1253937;C0031039|pericardial
null|Pericardial sac structure|Anatomy|false|false|C2317432;C1546613;C0013687;C1253937;C0031039|pericardialnull|Effusion (substance)|Finding|true|false|C0031050;C0442031;C3498924|effusion
null|null|Finding|true|false|C0031050;C0442031;C3498924|effusion
null|effusion|Finding|true|false|C0031050;C0442031;C3498924|effusionnull|Inspiratory Vital Capacity Test|Procedure|true|false|C3498924|IVCnull|lamina IVC|Anatomy|false|false|C2317432;C1546613;C0013687;C0031039;C4085887|IVCnull|Hypovolemia|Finding|false|false||volume depletionnull|Volume (publication)|Finding|false|false||volumenull|Volume|LabModifier|false|false||volumenull|Depletion|Finding|false|false||depletionnull|Lasix|Drug|false|false||Lasix
null|Lasix|Drug|false|false||Lasixnull|Breast Feeding|Finding|false|false||Nursingnull|RNAx nursing therapy actions|Procedure|false|false||Nursingnull|Discipline of Nursing|Title|false|false||Nursingnull|Able (qualifier value)|Finding|false|false||ablenull|Ability|Subject|false|false||ablenull|Does stand|Finding|false|false||stand
null|standards characteristics|Finding|false|false||standnull|Stand (physical object)|Device|false|false||stand
null|Stand Device|Device|false|false||standnull|Weight-Bearing state|Subject|false|false||weight bearnull|infant weight for previous delivery (history)|Finding|false|false||weight
null|Weight symptom (finding)|Finding|false|false||weightnull|Weighing patient|Procedure|false|false||weightnull|null|Attribute|false|false||weightnull|Body Weight|Subject|false|false||weightnull|Importance Weight|Modifier|false|false||weightnull|Weight|LabModifier|false|false||weightnull|Ursidae <Caniformia>|Entity|false|false||bearnull|Unsteady|Modifier|false|false||unsteadynull|At increased risk for falls|Finding|false|false||fall risknull|Falls|Finding|false|false||fallnull|Autumn|Time|false|false||fallnull|Risk|Finding|false|false||risknull|Spine Problem|Finding|false|false|C2752558;C0037949|spinenull|Neuron spine|Anatomy|false|false|C0150920;C4019020|spine
null|Vertebral column|Anatomy|false|false|C0150920;C4019020|spinenull|Film Dosage Form|Drug|false|false||film
null|film - layer|Drug|false|false||filmnull|null|Finding|false|false|C2752558;C0037949|filmnull|film (photographic)|Device|false|false||film
null|Film Device|Device|false|false||film
null|Film Container Cap|Device|false|false||filmnull|Film (unit of presentation)|LabModifier|false|false||film
null|Film Dosing Unit|LabModifier|false|false||filmnull|Fracture|Disorder|true|false||fracturesnull|Fractured|Finding|true|false||fracturesnull|Dislocations|Disorder|false|false||dislocationsnull|Hypotension|Finding|false|false||hypotensionnull|Middle|Modifier|false|false||midnull|Bradycardia by ECG Finding|Finding|false|false||bradycardia
null|Bradycardia|Finding|false|false||bradycardianull|Middle|Modifier|false|false||midnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|null|Time|false|false||prior tonull|null|Time|false|false||priornull|Transfer - product ownership|Finding|false|false||transfer
null|Transfer Technique|Finding|false|false||transfer
null|ActClass - transfer|Finding|false|false||transfer
null|null|Finding|false|false||transfernull|Transfer (immobility management)|Procedure|false|false||transfernull|elongation factor DmS-II|Drug|false|false||DM IInull|Hypertensive disease|Disorder|false|false||HTNnull|Coumadin|Drug|false|false||coumadin
null|Coumadin|Drug|false|false||coumadinnull|Malignant neoplasm of prostate|Disorder|false|false|C0033572;C4266527|prostate CAnull|Carcinoma in situ of prostate|Disorder|false|false|C0033572;C4266527|prostate
null|Prostatic Diseases|Disorder|false|false|C0033572;C4266527|prostate
null|Benign neoplasm of prostate|Disorder|false|false|C0033572;C4266527|prostate
null|Neoplasm of uncertain or unknown behavior of prostate|Disorder|false|false|C0033572;C4266527|prostatenull|Structure of prostate (body structure)|Anatomy|false|false|C0376358;C0496923;C0154088;C0033575;C0154009|prostate
null|Prostate|Anatomy|false|false|C0376358;C0496923;C0154088;C0033575;C0154009|prostatenull|Palp - CHV concept|Finding|false|false||palp
null|ALPP gene|Finding|false|false||palp
null|ALPP wt Allele|Finding|false|false||palpnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||GENERALnull|General medical service|Procedure|false|false||GENERALnull|Generalized|Modifier|false|false||GENERALnull|Well (answer to question)|Finding|false|false||Wellnull|Well (container)|Device|false|false||Wellnull|Microplate Well|Modifier|false|false||Well
null|Good|Modifier|false|false||Well
null|Healthy|Modifier|false|false||Wellnull|Male population group|Subject|false|false||man
null|Homo sapiens|Subject|false|false||man
null|Males|Subject|false|false||mannull|Mandinka Language|Entity|false|false||mannull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|Feeling comfortable|Finding|false|false||comfortablenull|Appropriate|Modifier|false|false||appropriatenull|HEENT|Anatomy|false|false||HEENTnull|Anicteric|Finding|false|false||anictericnull|Myelofibrosis|Disorder|false|false|C0694605|MMMnull|Medial part of medial mammillary nucleus|Anatomy|false|false|C0026987|MMMnull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787|HEART
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787|HEARTnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|HEARTnull|Chest>Heart|Anatomy|false|false|C0795691;C0153957;C0153500|HEART
null|Heart|Anatomy|false|false|C0795691;C0153957;C0153500|HEARTnull|Irregular|Modifier|false|false||irregularnull|SYSTOLIC EJECTION MURMUR|Finding|false|false||systolic ejection murmurnull|Systole|Finding|false|false||systolicnull|Ejection Murmurs|Finding|false|false||ejection murmurnull|Ejection as a Sports activity|Finding|false|false||ejectionnull|Ejection time|Attribute|false|false||ejectionnull|Ejection as a Circumstance of Injury|Phenomenon|false|false||ejectionnull|Heart murmur|Finding|false|false||murmurnull|lunate sulcus of the macaque|Anatomy|false|false||LUS
null|Lunate Sulcus|Anatomy|false|false||LUSnull|Lushai Language|Entity|false|false||LUSnull|Lung|Anatomy|false|false||LUNGSnull|Cancer/Testis Antigen|Drug|false|false||CTAnull|PCYT1A wt Allele|Finding|false|false||CTA
null|CERNA3 gene|Finding|false|false||CTAnull|Cardiac Computerized Tomographic Angiography|Procedure|false|false||CTAnull|Language Ability Proficiency - Good|Finding|false|false||good
null|Language Proficiency - Good|Finding|false|false||goodnull|Specimen Quality - Good|Modifier|false|false||good
null|Good|Modifier|false|false||goodnull|Air Movements|Phenomenon|false|false||air movementnull|Air (substance)|Drug|false|false||air
null|air|Drug|false|false||air
null|air|Drug|false|false||airnull|ACUTE INSULIN RESPONSE|Finding|false|false||air
null|AIRN gene|Finding|false|false||air
null|AI/RHEUM|Finding|false|false||airnull|Movement|Finding|false|false||movementnull|Respiratory, thoracic and mediastinal disorders|Disorder|false|false||respnull|Respiratory rate|Attribute|false|false||respnull|Unlabored|Finding|false|false||unlaborednull|Malignant neoplasm of abdomen|Disorder|false|false|C0230168;C0000726|ABDOMENnull|Abdomen problem|Finding|false|false|C0230168;C0000726|ABDOMENnull|Abdomen|Anatomy|false|false|C0941288;C0153662|ABDOMEN
null|Abdominal Cavity|Anatomy|false|false|C0941288;C0153662|ABDOMENnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||softnull|Soft|Modifier|false|false||softnull|LRRC4B gene|Finding|true|false||HSMnull|Protective muscle spasm|Finding|false|false||guardingnull|All extremities|Anatomy|false|false||EXTREMITIES
null|Limb structure|Anatomy|false|false||EXTREMITIESnull|Contusions|Disorder|false|false|C0040357;C4299090;C0230461;C4299097;C0016504|Bruisingnull|reported bruising (history)|Finding|false|false|C0230461;C4299097;C0016504;C0040357;C4299090|Bruisingnull|Lower extremity>Toes|Anatomy|false|false|C0555980;C1552822;C0009938;C2136686|toes
null|Toes|Anatomy|false|false|C0555980;C1552822;C0009938;C2136686|toesnull|Structure of left foot|Anatomy|false|false|C2136686;C0555980;C1552822;C0009938|left footnull|Table Cell Horizontal Align - left|Finding|false|false|C0040357;C4299090;C0230461;C4299097;C0016504|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Foot problem|Finding|false|false|C0040357;C4299090;C4299097;C0016504;C0230461|footnull|Lower extremity>Foot|Anatomy|false|false|C0555980;C2136686;C1552822;C0009938|foot
null|Foot|Anatomy|false|false|C0555980;C2136686;C1552822;C0009938|footnull|Foot Unit of Length|LabModifier|false|false||footnull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Foot|Anatomy|false|false||feetnull|Foot Unit of Length|LabModifier|false|false||feetnull|Ankle|Anatomy|false|false||anklesnull|Thigh structure|Anatomy|false|false||thighsnull|Neurology speciality|Title|false|false||NEUROnull|Neurologic (qualifier value)|Modifier|false|false||NEUROnull|Alert brand of caffeine|Drug|false|false||alert
null|Alert brand of caffeine|Drug|false|false||alertnull|Mentally alert|Finding|false|false||alert
null|Consciousness clear|Finding|false|false||alert
null|Alert note|Finding|false|false||alert
null|Alert|Finding|false|false||alertnull|null|Attribute|false|false||alertnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|Laboratory test finding|Lab|false|false||LABSnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0851353;C0005768;C0229664;C0005767|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C0014792;C1114281|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Mandibular right first molar mesial prosthesis|Device|false|false||30PMnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Mandibular right first molar mesial prosthesis|Device|false|false||30PMnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Alanine Transaminase|Drug|false|false||ALT
null|Alanine Transaminase|Drug|false|false||ALTnull|Liposarcoma, well differentiated|Disorder|false|false||ALT
null|Atypical Lipoma|Disorder|false|false||ALTnull|null|Finding|false|false||ALT
null|Alternative Billing Concepts|Finding|false|false||ALT
null|GPT gene|Finding|false|false||ALTnull|Antibiotic Lock Therapy|Procedure|false|false||ALTnull|Southern Altai Language|Entity|false|false||ALTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false|C1185650|AST
null|Aspartate Transaminase|Drug|false|false|C1185650|AST
null|Aspartate Transaminase|Drug|false|false|C1185650|AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false|C1185650|AST
null|SLC17A5 protein, human|Drug|false|false|C1185650|AST
null|SLC17A5 protein, human|Drug|false|false|C1185650|ASTnull|Atypical Spitz Nevus|Disorder|false|false|C1185650|ASTnull|SLC17A5 wt Allele|Finding|false|false|C1185650|AST
null|SLC17A5 gene|Finding|false|false|C1185650|AST
null|GOT1 gene|Finding|false|false|C1185650|ASTnull|Asterion|Anatomy|false|false|C0004002;C0242192;C1121182;C1415181;C1420113;C5960784;C4522245|ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|Lactate Dehydrogenase|Drug|false|false||LDH
null|Lactate Dehydrogenase|Drug|false|false||LDHnull|Lifetime Drinking History|Finding|false|false||LDHnull|Lactate dehydrogenase measurement|Procedure|false|false||LDHnull|Creatine Kinase|Drug|false|false||CPK
null|Creatine Kinase|Drug|false|false||CPKnull|PIK3C2A gene|Finding|false|false||CPKnull|Creatine kinase measurement|Procedure|false|false||CPKnull|Alkaline Phosphatase|Drug|false|false||AlkPhos
null|Alkaline Phosphatase|Drug|false|false||AlkPhosnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MB
null|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MBnull|creatine kinase activity|Finding|false|false||CK-MBnull|Serum creatine phosphokinase MB isoenzyme measurement|Procedure|false|false||CK-MB
null|Creatine kinase MB measurement|Procedure|false|false||CK-MBnull|Natriuretic Peptides B, human|Drug|false|false||proBNP
null|Natriuretic Peptides B, human|Drug|false|false||proBNPnull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|Laboratory test finding|Lab|false|false||LABSnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0005768;C0229664;C0005767;C0851353|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C0014792;C1114281|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MB
null|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MBnull|creatine kinase activity|Finding|false|false||CK-MBnull|Serum creatine phosphokinase MB isoenzyme measurement|Procedure|false|false||CK-MB
null|Creatine kinase MB measurement|Procedure|false|false||CK-MBnull|Plain chest X-ray|Procedure|false|false||CXRnull|Mild Severity of Illness Code|Finding|false|false||Mildnull|Mild (qualifier value)|Modifier|false|false||Mild
null|Mild Allergy Severity|Modifier|false|false||Mildnull|Congestive heart failure|Disorder|false|false|C4037974;C0018787|congestive heart failurenull|Congestive|Modifier|false|false||congestivenull|Congestive heart failure|Disorder|false|false|C4037974;C0018787|heart failure
null|Heart failure|Disorder|false|false|C4037974;C0018787|heart failurenull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787|heart
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787|heartnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|heartnull|Chest>Heart|Anatomy|false|false|C0795691;C0153957;C0153500;C0018802;C0018801;C0018802|heart
null|Heart|Anatomy|false|false|C0795691;C0153957;C0153500;C0018802;C0018801;C0018802|heartnull|Failure (biologic function)|Finding|false|false||failure
null|Failure|Finding|false|false||failure
null|Personal failure|Finding|false|false||failurenull|Widening|Modifier|false|false||Widenednull|Chest>Mediastinum.superior|Anatomy|false|false|C0153956;C0496915|superior mediastinum
null|Superior mediastinum|Anatomy|false|false|C0153956;C0496915|superior mediastinumnull|Upper|Modifier|false|false||superiornull|Neoplasm of uncertain or unknown behavior of mediastinum|Disorder|false|false|C4299144;C0230147;C0025066;C4037971|mediastinum
null|Benign tumor of mediastinum|Disorder|false|false|C4299144;C0230147;C0025066;C4037971|mediastinumnull|Chest>Mediastinum|Anatomy|false|false|C0153956;C0496915|mediastinum
null|Mediastinum|Anatomy|false|false|C0153956;C0496915|mediastinumnull|Leftward|Modifier|false|false||leftwardnull|Protocol Deviation|Finding|false|false||deviationnull|Spatial Displacement|Modifier|false|false||deviation
null|Variant|Modifier|false|false||deviationnull|Carcinoma in situ of trachea|Disorder|false|false|C0040578;C4299086|trachea
null|Benign neoplasm of trachea|Disorder|false|false|C0040578;C4299086|trachea
null|Tracheal Diseases|Disorder|false|false|C0040578;C4299086|tracheanull|trachea findings|Finding|false|false|C0040578;C4299086|tracheanull|Procedure on trachea|Procedure|false|false|C0040578;C4299086|tracheanull|Neck+Chest>Trachea|Anatomy|false|false|C0040580;C0154070;C0153953;C0872391;C5848218;C1705923;C0947630;C2603343;C0008972|trachea
null|Trachea|Anatomy|false|false|C0040580;C0154070;C0153953;C0872391;C5848218;C1705923;C0947630;C2603343;C0008972|tracheanull|Trachea <Xyleninae>|Entity|false|false||tracheanull|Similarity|Modifier|false|false||similarnull|null|Time|false|false||priornull|Study Object|Finding|false|false|C0040578;C4299086|studynull|Scientific Study|Procedure|false|false|C0040578;C4299086|study
null|Study|Procedure|false|false|C0040578;C4299086|study
null|Clinical Research|Procedure|false|false|C0040578;C4299086|studynull|Room of building - Study|Device|false|false||studynull|findings aspects|Finding|false|false||Findingsnull|null|Attribute|false|false||Findingsnull|Present|Finding|false|false||presence ofnull|Providing presence (regime/therapy)|Procedure|false|false||presencenull|Presence (property)|Modifier|false|false||presencenull|Goiter|Disorder|false|false|C0040132|thyroid goiternull|THYROID DIAGNOSTIC RADIOPHARMACEUTICALS|Drug|false|false|C0040132|thyroid
null|THYROID|Drug|false|false|C0040132|thyroid
null|THYROID|Drug|false|false|C0040132|thyroid
null|thyroid (USP)|Drug|false|false|C0040132|thyroid
null|thyroid (USP)|Drug|false|false|C0040132|thyroid
null|thyroid (USP)|Drug|false|false|C0040132|thyroidnull|Thyroid Diseases|Disorder|false|false|C0040132|thyroidnull|examination of thyroid|Procedure|false|false|C0040132|thyroidnull|Thyroid Gland|Anatomy|false|false|C0018021;C0018021;C0040128;C2228489;C3540038;C0040134;C5781115|thyroidnull|Goiter|Disorder|false|false|C0040132|goiternull|Clinical NEC (not elsewhere classified in LNC)|Finding|false|false||clinicalnull|Clinical|Modifier|false|false||clinicalnull|Correlation|Modifier|false|false||correlationnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0741025|chest
null|Anterior thoracic region|Anatomy|false|false|C0741025|chestnull|Spine Problem|Finding|false|false|C2752558;C0037949|spinenull|Neuron spine|Anatomy|false|false|C4019020;C0150920|spine
null|Vertebral column|Anatomy|false|false|C4019020;C0150920|spinenull|Film Dosage Form|Drug|false|false||film
null|film - layer|Drug|false|false||filmnull|null|Finding|false|false|C2752558;C0037949|filmnull|film (photographic)|Device|false|false||film
null|Film Device|Device|false|false||film
null|Film Container Cap|Device|false|false||filmnull|Film (unit of presentation)|LabModifier|false|false||film
null|Film Dosing Unit|LabModifier|false|false||filmnull|Lumbar Region|Anatomy|false|false|C1420009;C1552651|lumbarnull|Type - ParameterizedDataType|Finding|false|false|C0024090;C0549207|type
null|SGCG gene|Finding|false|false|C0024090;C0549207|typenull|null|Modifier|false|false||typenull|Bone structure of spine|Anatomy|false|false|C1420009;C1552651|vertebralnull|Human body|Subject|false|false||bodiesnull|Present|Finding|false|false||present
null|Presentation|Finding|false|false||presentnull|Abnormal degeneration|Finding|false|false||degenerative changesnull|biologic degeneration|Finding|false|false||degenerative
null|Abnormal degeneration|Finding|false|false||degenerativenull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|Loss (adaptation)|Finding|false|false|C0442106;C0021815|lossnull|Loss (quantitative)|LabModifier|false|false||lossnull|Intervertebral disc structure|Anatomy|false|false|C1696131;C1444662;C5890125|intervertebral discnull|Intervertebral|Anatomy|false|false|C1696131;C1444662;C5890125|intervertebralnull|Disk Drug Form|Drug|false|false|C1621443;C1556138|discnull|Disc (List bullets)|Finding|false|false|C0442106;C0021815;C1621443;C1556138|disc
null|Discontinued|Finding|false|false|C0442106;C0021815;C1621443;C1556138|discnull|Disc - Body Part|Anatomy|false|false|C0993608;C1696131;C1444662|disc
null|death-inducing signaling complex location|Anatomy|false|false|C0993608;C1696131;C1444662|discnull|Disk Device|Device|false|false||discnull|Disk Shape|Modifier|false|false||discnull|Disk Dosing Unit|LabModifier|false|false||discnull|Height|LabModifier|false|false||heightnull|Numerous|LabModifier|false|false||multiplenull|Levels (qualifier value)|Modifier|false|false||levelsnull|Sclerotic (qualifier value)|Finding|false|false||sclerotic
null|Sclerosis|Finding|false|false||scleroticnull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|Adenohypophyseal Diseases|Disorder|false|false||anteriornull|Anterior|Modifier|false|false||anteriornull|Osteophyte formation|Finding|false|false||osteophyte formationnull|Osteophyte|Disorder|false|false||osteophyte
null|External hyperostosis|Disorder|false|false||osteophytenull|Formation|Finding|false|false||formationnull|Anabolism|Phenomenon|false|false||formationnull|Formations|Modifier|false|false||formationnull|Fracture|Disorder|true|false||fracturenull|Compression fracture of vertebral column|Finding|true|false|C0549207|vertebral compressionnull|Bone structure of spine|Anatomy|false|false|C0262431|vertebralnull|null|Finding|true|false||compression
null|Compressed structure|Finding|true|false||compressionnull|Compression Therapy|Procedure|true|false||compression
null|Data Compression|Procedure|true|false||compressionnull|Compression|Phenomenon|true|false||compressionnull|Deformity|Disorder|true|false||deformity
null|Congenital Abnormality|Disorder|true|false||deformitynull|null|Finding|true|false||deformitynull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Grade 1 (qualifier value)|Finding|false|false||grade 1
null|Tumor grade G1|Finding|false|false||grade 1
null|Simpson Grade 1|Finding|false|false||grade 1
null|First grade in elementary school|Finding|false|false||grade 1null|Histopathologic Grade|Finding|false|false||grade
null|Grade|Finding|false|false||grade
null|School Grade|Finding|false|false||gradenull|Anterolisthesis|Disorder|false|false||anterolisthesisnull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|biologic degeneration|Finding|false|false||degenerative
null|Abnormal degeneration|Finding|false|false||degenerativenull|Science of Etiology|Finding|false|false||etiology
null|Etiology aspects|Finding|false|false||etiology
null|Etiology|Finding|false|false||etiologynull|Structure of articular surface of bone|Anatomy|false|false||Facetnull|null|Disorder|false|false|C0024091;C3887615;C0024090;C2752558;C0037949|hypertrophicnull|Hypertrophic|Finding|false|false|C0024091;C3887615;C2752558;C0037949|hypertrophic
null|Hypertrophy|Finding|false|false|C0024091;C3887615;C2752558;C0037949|hypertrophicnull|Changing|Finding|false|false|C2752558;C0037949;C0024091;C3887615;C0024090|changesnull|Changed status|LabModifier|false|false||changesnull|Body Site Modifier - Lower|Anatomy|false|false|C2003888|lowernull|Lower (action)|Event|false|false|C1548802;C0024091;C3887615|lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Lumbar spine structure|Anatomy|false|false|C0263630;C2003888;C0333959;C0020564;C0150920;C0392747|lumbar spine
null|Bone structure of lumbar vertebra|Anatomy|false|false|C0263630;C2003888;C0333959;C0020564;C0150920;C0392747|lumbar spinenull|Lumbar Region|Anatomy|false|false|C0150920;C0263630;C0392747|lumbarnull|Spine Problem|Finding|false|false|C0024091;C3887615;C0024090;C2752558;C0037949|spinenull|Neuron spine|Anatomy|false|false|C0392747;C0333959;C0020564;C0263630;C0150920|spine
null|Vertebral column|Anatomy|false|false|C0392747;C0333959;C0020564;C0263630;C0150920|spinenull|Levels (qualifier value)|Modifier|false|false||levelsnull|Blood Vessel|Anatomy|false|false||Vascularnull|Vascular|Modifier|false|false||Vascularnull|Pathologic calcification, calcified structure|Finding|true|false||calcifications
null|Physiologic calcification|Finding|true|false||calcificationsnull|Calcified (qualifier value)|Modifier|false|false||calcificationsnull|Sacroiliac joint structure|Anatomy|false|false||sacroiliac jointsnull|sacroiliac|Anatomy|false|false||sacroiliacnull|Joints|Anatomy|false|false||joints
null|Articular system|Anatomy|false|false||jointsnull|impression (attitude)|Finding|false|false||IMPRESSION
null|EKG impression|Finding|false|false||IMPRESSIONnull|Fracture|Disorder|true|false||fracturenull|CAT scan of head|Procedure|false|false|C0018670;C0152336|CT headnull|null|Attribute|false|false|C0018670;C0152336|CT headnull|Problems with head|Disorder|false|false|C0018670;C0152336|headnull|Procedure on head|Procedure|false|false|C0018670;C0152336|headnull|Structure of head of caudate nucleus|Anatomy|false|false|C0876917;C0202691;C0881943;C0362076|head
null|Head|Anatomy|false|false|C0876917;C0202691;C0881943;C0362076|headnull|Head Device|Device|false|false||headnull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Intracranial Hemorrhage|Finding|true|false|C0524466|intracranial hemorrhagenull|Intracranial Route of Administration|Finding|false|false|C0524466|intracranialnull|Intracranial|Anatomy|false|false|C1522213;C0019080;C0151699|intracranialnull|Hemorrhage|Finding|true|false|C0524466|hemorrhagenull|Edema|Finding|true|false||edemanull|null|Attribute|true|false||edemanull|Admission Level of Care Code - Acute|Finding|true|false||acute
null|Acute - Triage Code|Finding|true|false||acutenull|acute|Time|false|false||acutenull|Blood Vessel|Anatomy|false|false||vascularnull|Vascular|Modifier|false|false||vascularnull|Infarction|Finding|false|false||infarctionnull|Areas <Spilosomini>|Entity|false|false||areasnull|Area|Modifier|false|false||areasnull|Encephalomalacia|Disorder|false|false|C0030560;C0796494|encephalomalacianull|Malignant neoplasm of parietal lobe|Disorder|false|false|C0030560;C0796494|parietal lobenull|Parietal Lobe|Anatomy|false|false|C0153637;C0014068;C3539671;C1428707|parietal lobenull|Parietal|Modifier|false|false||parietalnull|AKT1S1 wt Allele|Finding|false|false|C0796494;C0030560|lobe
null|AKT1S1 gene|Finding|false|false|C0796494;C0030560|lobenull|lobe|Anatomy|false|false|C3539671;C1428707;C0014068;C0153637|lobenull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|null|Finding|false|false||unchangednull|About The Same|Modifier|false|false||unchangednull|Academic Research Enhancement Awards|Event|false|false||areanull|Geographic Locations|Entity|false|false||areanull|Area|Modifier|false|false||areanull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Adjacent|Modifier|false|false||adjacent tonull|Adjacent|Modifier|false|false||adjacentnull|null|Finding|false|false||unchangednull|About The Same|Modifier|false|false||unchangednull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Coronal (qualifier value)|Modifier|false|false||frontalnull|Meningioma|Disorder|false|false||meningiomasnull|Greater|LabModifier|false|false||larger
null|Large|LabModifier|false|false||largernull|Calcified (qualifier value)|Modifier|false|false||calcifiednull|Observation Interpretation - better|Finding|false|false||betternull|Better|Modifier|false|false||betternull|null|Time|false|false||priornull|CYREN gene|Finding|false|false||MRInull|Magnetic resonance imaging service|Procedure|false|false||MRI
null|Magnetic Resonance Imaging|Procedure|false|false||MRInull|Maori Language|Entity|false|false||MRInull|Heart Ventricle|Anatomy|false|false||Ventriclesnull|Parenchymal volume loss|Finding|false|false||parenchymal volume lossnull|Volume (publication)|Finding|false|false||volumenull|Volume|LabModifier|false|false||volumenull|Loss (adaptation)|Finding|false|false||lossnull|Loss (quantitative)|LabModifier|false|false||lossnull|atherosclerotic|Finding|false|false||atheroscleroticnull|Physiologic calcification|Finding|false|false|C0007272|calcification
null|Calcification|Finding|false|false|C0007272|calcification
null|Calcinosis|Finding|false|false|C0007272|calcificationnull|Calcified (qualifier value)|Modifier|false|false||calcificationnull|Carotid Arteries|Anatomy|false|false|C1533591;C0006660;C0006663|carotidnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Fracture|Disorder|false|false||fracturenull|Pneumatic mastoid cell|Anatomy|false|false|C2681903;C1140091;C1866503;C2228459;C0001861;C3536832;C1550016|mastoid air cellsnull|examination of mastoid region|Procedure|false|false|C0229427;C0007634;C0446908;C4266570;C1521748|mastoidnull|Mastoid process|Anatomy|false|false|C1550016;C2681903;C1140091;C1866503;C2228459|mastoid
null|null|Anatomy|false|false|C1550016;C2681903;C1140091;C1866503;C2228459|mastoid
null|Head>Mastoid|Anatomy|false|false|C1550016;C2681903;C1140091;C1866503;C2228459|mastoidnull|Air (substance)|Drug|false|false|C0007634;C0229427|air
null|air|Drug|false|false|C0007634;C0229427|air
null|air|Drug|false|false|C0007634;C0229427|airnull|ACUTE INSULIN RESPONSE|Finding|false|false|C0229427;C0446908;C4266570;C1521748;C0007634|air
null|AIRN gene|Finding|false|false|C0229427;C0446908;C4266570;C1521748;C0007634|air
null|AI/RHEUM|Finding|false|false|C0229427;C0446908;C4266570;C1521748;C0007634|airnull|Cells|Anatomy|false|false|C0001861;C3536832;C2228459;C1550016;C2681903;C1140091;C1866503|cellsnull|Remote control command - Clear|Finding|false|false|C0446908;C4266570;C1521748;C0007634;C0229427|clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|impression (attitude)|Finding|false|false||IMPRESSION
null|EKG impression|Finding|false|false||IMPRESSIONnull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Intracranial Route of Administration|Finding|false|false|C0524466|intracranialnull|Intracranial|Anatomy|false|false|C1522213|intracranialnull|Congenital Abnormality|Disorder|false|false||abnormalitynull|Abnormality|Finding|false|false||abnormalitynull|null|Finding|false|false||unchangednull|About The Same|Modifier|false|false||unchangednull|Act Relationship Subset - previous|Time|false|false||previous
null|Previous|Time|false|false||previousnull|Infarction|Finding|false|false||infarctsnull|Meningioma|Disorder|false|false||meningiomasnull|Waveforms|Phenomenon|false|false|C0015809|Waveformsnull|Common Specifications in HL7 V3 Publishing|Finding|false|false|C0015809|common
null|shared attribute|Finding|false|false|C0015809|commonnull|Common (qualifier value)|LabModifier|false|false||commonnull|Femoral vein|Anatomy|false|false|C3245511;C1522138;C0450448;C0332516;C2699744;C0398102|femoral veinsnull|Femur|Anatomy|false|false|C0398102|femoralnull|Procedure on vein|Procedure|false|false|C0042449;C0015809;C0015811|veinsnull|Veins|Anatomy|false|false|C0398102;C0332516;C2699744|veinsnull|Symmetric Relationship|Finding|false|false|C0042449;C0015809|symmetric
null|Symmetrical|Finding|false|false|C0042449;C0015809|symmetricnull|Appropriate|Modifier|false|false||appropriatenull|Response process|Subject|false|false||responsesnull|Valsalva Maneuver|Procedure|false|false||Valsalva maneuversnull|valsalva|Procedure|false|false||Valsalvanull|Body Site Modifier - Lower|Anatomy|false|false|C2003888|lowernull|Lower (action)|Event|false|false|C1548802|lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|All extremities|Anatomy|false|false||extremities
null|Limb structure|Anatomy|false|false||extremitiesnull|Common Specifications in HL7 V3 Publishing|Finding|false|false||common
null|shared attribute|Finding|false|false||commonnull|Common (qualifier value)|LabModifier|false|false||commonnull|Femur|Anatomy|false|false||femoralnull|Proximal Resection Margin|Attribute|false|false||proximalnull|Proximal|Modifier|false|false||proximalnull|Greater|LabModifier|false|false||greaternull|Superficial|Modifier|false|false||superficialnull|Femur|Anatomy|false|false|C0398102|femoralnull|Structure of popliteal vein|Anatomy|false|false|C0398102|popliteal veinsnull|popliteal|Anatomy|false|false|C0398102|poplitealnull|Procedure on vein|Procedure|false|false|C0442037;C0015811;C0032652;C0042449|veinsnull|Veins|Anatomy|false|false|C0398102|veinsnull|Appropriate|Modifier|false|false||appropriatenull|Walls of a building|Device|false|false||wallnull|Walls of a building|Device|false|false||wallnull|Flow|Phenomenon|false|false||flownull|Color doppler ultrasound|Procedure|false|false||color Dopplernull|color additive|Drug|false|false||color
null|Coloring Excipient|Drug|false|false||colornull|color - solid dosage form|Modifier|false|false||color
null|Color|Modifier|false|false||colornull|Color quantity|LabModifier|false|false||colornull|Doppler studies|Procedure|false|false||Dopplernull|analysis aspect|Finding|false|false||analysisnull|Analysis of substances|Procedure|false|false||analysis
null|Analysis|Procedure|false|false||analysisnull|Communication Response|Finding|false|false||response
null|Disease Response|Finding|false|false||response
null|Answer (statement)|Finding|false|false||responsenull|Response process|Subject|false|false||responsenull|Waveforms|Phenomenon|false|false||waveformnull|Increased size (finding)|Finding|false|false||augmentationnull|Augmentation procedure|Procedure|false|false||augmentationnull|Walls of a building|Device|false|false||Wallnull|Walls of a building|Device|false|false||wallnull|Flow|Phenomenon|false|false||flownull|Posterior pituitary disease|Disorder|false|false||posteriornull|Dorsal|Modifier|false|false||posteriornull|Bone structure of tibia|Anatomy|false|false||tibialnull|Peroneal|Modifier|false|false||peronealnull|Procedure on vein|Procedure|false|false|C0042449|veinsnull|Veins|Anatomy|false|false|C0398102|veinsnull|impression (attitude)|Finding|false|false||IMPRESSION
null|EKG impression|Finding|false|false||IMPRESSIONnull|Deep Vein Thrombosis|Disorder|true|false|C0015385;C0023216;C0042449|deep venous thrombosisnull|Deep Resection Margin|Attribute|false|false||deepnull|Deep (qualifier value)|Modifier|false|false||deepnull|Venous thrombosis after immobility|Finding|true|false|C0023216;C0015385;C0042449|venous thrombosis
null|Venous Thrombosis|Finding|true|false|C0023216;C0015385;C0042449|venous thrombosisnull|Veins|Anatomy|false|false|C0149871;C0517555;C0042487|venousnull|Venous|Modifier|false|false||venousnull|Thrombosis|Finding|true|false|C0023216;C0015385|thrombosisnull|Lower Extremity|Anatomy|false|false|C2003888;C0517555;C0042487;C0149871;C0040053|lower extremitynull|Body Site Modifier - Lower|Anatomy|false|false|C2003888|lowernull|Lower (action)|Event|false|false|C0023216;C0015385;C1548802|lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Limb structure|Anatomy|false|false|C0149871;C2003888;C0517555;C0042487;C0040053|extremitynull|Microbiology Diagnostic Service Section ID|Finding|false|false||MICROBIOLOGY
null|Microbiological|Finding|false|false||MICROBIOLOGY
null|Microbiology - Laboratory Class|Finding|false|false||MICROBIOLOGYnull|Microbiology procedure|Procedure|false|false||MICROBIOLOGYnull|Science of Microbiology|Title|false|false||MICROBIOLOGYnull|Blood culture|Procedure|false|false||Blood culturenull|Blood and lymphatic system disorders|Disorder|false|false||Bloodnull|peripheral blood|Finding|false|false||Blood
null|Blood|Finding|false|false||Blood
null|In Blood|Finding|false|false||Bloodnull|Culture Dose Form|Drug|false|false||culturenull|Culture (Anthropological)|Finding|false|false||culture
null|Cultural aspects|Finding|false|false||culturenull|Microbial culture (procedure)|Procedure|false|false||culture
null|Laboratory culture|Procedure|false|false||culturenull|Growth & development aspects|Finding|true|false||growth
null|Tissue Growth|Finding|true|false||growth
null|Growth|Finding|true|false||growth
null|growth aspects|Finding|true|false||growthnull|Growth action|Phenomenon|true|false||growthnull|Atrial Fibrillation|Disorder|false|false||afibnull|Atrial Fibrillation by ECG Finding|Lab|false|false||afibnull|Congestive heart failure|Disorder|false|false|C0262212|CHFnull|Choroidal fissure|Anatomy|false|false|C0018802|CHFnull|Pulmonary Edema|Finding|false|false||pulm edemanull|Pulmonary ventilator management|Procedure|false|false||pulmnull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Congestive heart failure|Disorder|false|false|C0262212|CHFnull|Choroidal fissure|Anatomy|false|false|C0018802|CHFnull|Acute-on-chronic|Time|false|false||acute on chronicnull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Patient Outcome - Worsening|Finding|false|false||worseningnull|Worsening (qualifier value)|Modifier|false|false||worseningnull|Diastole|Attribute|false|false||diastolicnull|Congestive heart failure|Disorder|false|false|C4037974;C0018787|congestive heart failurenull|Congestive|Modifier|false|false||congestivenull|Congestive heart failure|Disorder|false|false|C4037974;C0018787|heart failure
null|Heart failure|Disorder|false|false|C4037974;C0018787|heart failurenull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787|heart
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787|heartnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|heartnull|Chest>Heart|Anatomy|false|false|C0680095;C0231174;C5200924;C0018801;C0018802;C0018802;C0153957;C0153500;C0795691|heart
null|Heart|Anatomy|false|false|C0680095;C0231174;C5200924;C0018801;C0018802;C0018802;C0153957;C0153500;C0795691|heartnull|Failure (biologic function)|Finding|false|false|C4037974;C0018787|failure
null|Failure|Finding|false|false|C4037974;C0018787|failure
null|Personal failure|Finding|false|false|C4037974;C0018787|failurenull|Most Recent|Time|false|false||most recentnull|Recent|Time|false|false||recentnull|LVEF (procedure)|Procedure|false|false||LVEFnull|Left ventricular ejection fraction|Attribute|false|false||LVEFnull|Recent|Time|false|false||recentnull|Reduced|Finding|false|false||decreasenull|Decrease|LabModifier|false|false||decreasenull|Mobility finding|Finding|false|false||mobilitynull|Range of Motion, Articular|Attribute|false|false||mobilitynull|Mobility (attribute)|Modifier|false|false||mobilitynull|Falls|Finding|false|false||fallnull|Autumn|Time|false|false||fallnull|Probable diagnosis|Finding|false|false||Likely
null|Probably|Finding|false|false||Likelynull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Medication Compliance|Finding|false|false||medication non-compliancenull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Patient Outcome - Worsening|Finding|false|false|C0003483|worseningnull|Worsening (qualifier value)|Modifier|false|false||worseningnull|Aortic Valve Stenosis|Finding|false|false|C0003483|aortic stenosisnull|Aorta|Anatomy|false|false|C0003507;C1546960;C1261287|aorticnull|Stenosis|Finding|false|false|C0003483|stenosisnull|Stenosis <Pimeliinae>|Entity|false|false||stenosisnull|Stenosis Morphology|Modifier|false|false||stenosisnull|Most Recent|Time|false|false||most recentnull|Recent|Time|false|false||recentnull|ECHO protocol|Procedure|false|false||echo
null|Extension for Community Healthcare Outcomes|Procedure|false|false||echonull|Echo <Calopterygidae>|Entity|false|false||echonull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|Never - AcknowledgementCondition|Time|false|false||never
null|Never (frequency)|Time|false|false||nevernull|Hypoxia|Finding|false|false||hypoxicnull|examination of lungs|Procedure|false|false|C4037972;C0024109|lung examnull|Lung diseases|Disorder|false|false|C4037972;C0024109|lungnull|Lung Problem|Finding|false|false|C4037972;C0024109|lungnull|Chest>Lung|Anatomy|false|false|C0582103;C0740941;C2228454;C4284036;C0024115|lung
null|Lung|Anatomy|false|false|C0582103;C0740941;C2228454;C4284036;C0024115|lungnull|Exam|Finding|false|false|C4037972;C0024109|examnull|Medical Examination|Procedure|false|false|C4037972;C0024109|examnull|Pulmonary ventilator management|Procedure|false|false||pulmnull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Leg|Anatomy|false|false|C0332459;C4551657;C0728907;C1257972;C0565514;C5781420|legsnull|null|Attribute|false|false|C1140621|legsnull|Compression Stockings|Device|false|false||compression stockings
null|Support stockings - garment|Device|false|false||compression stockingsnull|null|Finding|false|false|C1140621|compression
null|Compressed structure|Finding|false|false|C1140621|compressionnull|Compression Therapy|Procedure|false|false|C1140621|compression
null|Data Compression|Procedure|false|false|C1140621|compressionnull|Compression|Phenomenon|false|false|C1140621|compressionnull|Stocking (hosiery)|Device|false|false||stockings
null|Socks|Device|false|false||stockingsnull|torsemide|Drug|false|false||torsemide
null|torsemide|Drug|false|false||torsemidenull|Daily|Time|false|false||dailynull|Increase|Finding|false|false||increasenull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|wife|Subject|false|false||wifenull|Unable|Finding|false|false||unablenull|Clarify|Event|false|false||clarifynull|Intensity and Distress 1|Finding|false|false||slightnull|Slight (qualifier value)|Modifier|false|false||slight
null|Mild (qualifier value)|Modifier|false|false||slightnull|Improvement|Finding|false|false||improvementnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|On discharge|Time|false|false||on dischargenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Recent|Time|false|false||RECENTnull|Accidental Falls|Disorder|false|false||FALLSnull|Falls|Finding|false|false||FALLSnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Recent|Time|false|false||recentlynull|At home|Finding|false|false||at homenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|triptorelin|Drug|false|false||trip
null|triptorelin|Drug|false|false||trip
null|triptorelin|Drug|false|false||tripnull|TRAIP wt Allele|Finding|false|false||trip
null|TRAIP gene|Finding|false|false||trip
null|PIK3IP1 gene|Finding|false|false||trip
null|LRRFIP1 gene|Finding|false|false||tripnull|Tripping|Phenomenon|false|false||tripnull|Diagnostic Service Section ID - Physical Therapy|Finding|false|false||physical therapynull|Physical therapy|Procedure|false|false||physical therapynull|Physical therapy (field)|Title|false|false||physical therapynull|physical examination (physical finding)|Finding|false|false||physical
null|Physical|Finding|false|false||physicalnull|Physical Examination|Procedure|false|false||physicalnull|Therapy Object (animal model)|Finding|false|false||therapy
null|therapeutic aspects|Finding|false|false||therapynull|Therapeutic procedure|Procedure|false|false||therapynull|Unsteady|Modifier|false|false||unsteadynull|Foot|Anatomy|false|false||feetnull|Foot Unit of Length|LabModifier|false|false||feetnull|SAFE-Biopharma Standard|Finding|false|false||safenull|Discharge to home|Procedure|false|false||discharge homenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Walkers|Device|false|false||walkernull|Commodes|Device|false|false||commodenull|wife|Subject|false|false||wifenull|Hour|Time|false|false||hournull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Further|Modifier|false|false||furthernull|Accidental Falls|Disorder|false|false||fallsnull|Falls|Finding|false|false||fallsnull|On admission|Time|false|false||on admissionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|next - HtmlLinkType|Finding|false|false||nextnull|Following|Time|false|false||next
null|Then|Time|false|false||nextnull|Adjacent|Modifier|false|false||nextnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|BaseLine dental cement|Drug|false|false||baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|glipizide|Drug|false|false||Glipizide
null|glipizide|Drug|false|false||Glipizidenull|Actos|Drug|false|false||actos
null|Actos|Drug|false|false||actosnull|Hospitals|Device|false|false||in hospitalnull|Hospitals|Entity|false|false||in hospitalnull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|insulin, regular, human|Drug|false|false||insulin
null|Insulin [EPC]|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulinnull|INS gene|Finding|false|false||insulinnull|Insulin measurement|Procedure|false|false||insulinnull|Scale, LOINC Axis 5|Finding|false|false|C0222045|scale
null|Base Number|Finding|false|false|C0222045|scale
null|Scale - rank|Finding|false|false|C0222045|scalenull|Integumentary scale|Anatomy|false|false|C0349674;C2981742;C1522412;C1527415;C4521986;C1947916|scalenull|Weight measurement scales|Device|false|false||scalenull|Scaling|Event|false|false|C0222045|scalenull|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0222045;C0226896|oral
null|Oral (intended site)|Finding|false|false|C0222045;C0226896|oralnull|Oral cavity|Anatomy|false|false|C1272919;C4284232;C1527415;C4521986|oralnull|Oral|Modifier|false|false||oralnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false|C0226896|medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Hypertensive disease|Disorder|false|false||HTNnull|isosorbide|Drug|false|false||isosorbide
null|isosorbide|Drug|false|false||isosorbidenull|lisinopril|Drug|false|false||lisinopril
null|lisinopril|Drug|false|false||lisinoprilnull|One day|Time|false|false||one daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|null|Attribute|false|false||Metoprolol dosenull|metoprolol dose|LabModifier|false|false||Metoprolol dosenull|metoprolol|Drug|false|false||Metoprolol
null|metoprolol|Drug|false|false||Metoprololnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|Bradycardia by ECG Finding|Finding|false|false||bradycardia
null|Bradycardia|Finding|false|false||bradycardianull|Atrial Fibrillation|Disorder|false|false||Afibnull|Atrial Fibrillation by ECG Finding|Lab|false|false||Afibnull|Integrated Neuromusculoskeletal Release|Procedure|false|false||INR
null|International Normalized Ratio|Procedure|false|false||INRnull|Coagulation tissue factor induced.INR|Attribute|false|false||INRnull|On admission|Time|false|false||on admissionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Daily|Time|false|false||dailynull|Coumadin|Drug|false|false||coumadin
null|Coumadin|Drug|false|false||coumadinnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Daily|Time|false|false||dailynull|wife|Subject|false|false||wifenull|Home visit (procedure)|Procedure|false|false||home servicesnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Clinical Service|Procedure|false|false||servicesnull|Services|Event|false|false||servicesnull|Marketing basis - Transitional|Finding|false|false||TRANSITIONALnull|Transitional cell morphology|Modifier|false|false||TRANSITIONALnull|Blood culture|Procedure|false|false||Blood culturenull|Blood and lymphatic system disorders|Disorder|false|false||Bloodnull|peripheral blood|Finding|false|false||Blood
null|Blood|Finding|false|false||Blood
null|In Blood|Finding|false|false||Bloodnull|Culture Dose Form|Drug|false|false||culturenull|Culture (Anthropological)|Finding|false|false||culture
null|Cultural aspects|Finding|false|false||culturenull|Microbial culture (procedure)|Procedure|false|false||culture
null|Laboratory culture|Procedure|false|false||culturenull|Growth & development aspects|Finding|true|false||growth
null|Tissue Growth|Finding|true|false||growth
null|Growth|Finding|true|false||growth
null|growth aspects|Finding|true|false||growthnull|Growth action|Phenomenon|true|false||growthnull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|allopurinol|Drug|false|false||Allopurinol
null|allopurinol|Drug|false|false||Allopurinolnull|Tablet Dosage Form|Drug|false|false||TABLETnull|Tablet (unit of presentation)|LabModifier|false|false||TABLET
null|Tablet Dosing Unit|LabModifier|false|false||TABLETnull|Cyanocobalamin Drug Class|Drug|false|false||Cyanocobalamin
null|Cyanocobalamin Drug Class|Drug|false|false||Cyanocobalamin
null|vitamin B12|Drug|false|false||Cyanocobalamin
null|vitamin B12|Drug|false|false||Cyanocobalamin
null|vitamin B12|Drug|false|false||Cyanocobalaminnull|microgram|LabModifier|false|false||MCGnull|per milliliter|LabModifier|false|false||/MLnull|Vial device|Device|false|false||VIALnull|Vial (unit of presentation)|LabModifier|false|false||VIAL
null|Vial Dosing Unit|LabModifier|false|false||VIALnull|Take|Procedure|false|false||Takenull|dexamethasone|Drug|false|false||Dexamethasone
null|dexamethasone|Drug|false|false||Dexamethasonenull|Tablet Dosage Form|Drug|false|false||TABLETnull|Tablet (unit of presentation)|LabModifier|false|false||TABLET
null|Tablet Dosing Unit|LabModifier|false|false||TABLETnull|glipizide|Drug|false|false||Glipizide
null|glipizide|Drug|false|false||Glipizidenull|Tablet Dosage Form|Drug|false|false||TABLETnull|Tablet (unit of presentation)|LabModifier|false|false||TABLET
null|Tablet Dosing Unit|LabModifier|false|false||TABLETnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|goserelin acetate|Drug|false|false||Goserelin acetate
null|goserelin acetate|Drug|false|false||Goserelin acetate
null|goserelin acetate|Drug|false|false||Goserelin acetatenull|goserelin|Drug|false|false||Goserelin
null|goserelin|Drug|false|false||Goserelinnull|acetate|Drug|false|false||acetate
null|acetate|Drug|false|false||acetatenull|Drug Implant|Drug|false|false||IMPLANTnull|Traumatic implant|Disorder|false|false||IMPLANTnull|null|Finding|false|false||IMPLANT
null|Administration via Implantation|Finding|false|false||IMPLANTnull|Implantation procedure|Procedure|false|false||IMPLANTnull|null|Attribute|false|false||IMPLANTnull|Implants|Device|false|false||IMPLANTnull|Implant (unit of presentation)|LabModifier|false|false||IMPLANT
null|Implant Dosing Unit|LabModifier|false|false||IMPLANTnull|isosorbide dinitrate|Drug|false|false||Isosorbide dinitrate
null|isosorbide dinitrate|Drug|false|false||Isosorbide dinitratenull|isosorbide|Drug|false|false||Isosorbide
null|isosorbide|Drug|false|false||Isosorbidenull|Tablet Dosage Form|Drug|false|false||TABLETnull|Tablet (unit of presentation)|LabModifier|false|false||TABLET
null|Tablet Dosing Unit|LabModifier|false|false||TABLETnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|lisinopril|Drug|false|false||Lisinopril
null|lisinopril|Drug|false|false||Lisinoprilnull|Tablet Dosage Form|Drug|false|false||TABLETnull|Tablet (unit of presentation)|LabModifier|false|false||TABLET
null|Tablet Dosing Unit|LabModifier|false|false||TABLETnull|memantine|Drug|false|false||Memantine
null|memantine|Drug|false|false||Memantinenull|metoprolol tartrate|Drug|false|false||Metoprolol tartrate
null|metoprolol tartrate|Drug|false|false||Metoprolol tartratenull|metoprolol|Drug|false|false||Metoprolol
null|metoprolol|Drug|false|false||Metoprololnull|tartrate|Drug|false|false||tartrate
null|Tartrates|Drug|false|false||tartrate
null|tartrate|Drug|false|false||tartratenull|Tablet Dosage Form|Drug|false|false||TABLETnull|Tablet (unit of presentation)|LabModifier|false|false||TABLET
null|Tablet Dosing Unit|LabModifier|false|false||TABLETnull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|nilutamide|Drug|false|false||Nilutamide
null|nilutamide|Drug|false|false||Nilutamidenull|Tablet Dosage Form|Drug|false|false||TABLETnull|Tablet (unit of presentation)|LabModifier|false|false||TABLET
null|Tablet Dosing Unit|LabModifier|false|false||TABLETnull|nitroglycerin|Drug|false|false||Nitroglycerin
null|nitroglycerin|Drug|false|false||Nitroglycerinnull|oxycodone|Drug|false|false||Oxycodone
null|oxycodone|Drug|false|false||Oxycodonenull|Oxycodone measurement|Procedure|false|false||Oxycodonenull|Tablet Dosage Form|Drug|false|false||TABLETnull|Tablet (unit of presentation)|LabModifier|false|false||TABLET
null|Tablet Dosing Unit|LabModifier|false|false||TABLETnull|Take|Procedure|false|false||Takenull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|prednisone|Drug|false|false||Prednisone
null|prednisone|Drug|false|false||Prednisone
null|prednisone|Drug|false|false||Prednisonenull|null|Procedure|false|false||Tapernull|Tablet Dosage Form|Drug|false|false||TABLETnull|Tablet (unit of presentation)|LabModifier|false|false||TABLET
null|Tablet Dosing Unit|LabModifier|false|false||TABLETnull|day|Time|false|false||daysnull|simvastatin|Drug|false|false||Simvastatin
null|simvastatin|Drug|false|false||Simvastatinnull|Tablet Dosage Form|Drug|false|false||TABLETnull|Tablet (unit of presentation)|LabModifier|false|false||TABLET
null|Tablet Dosing Unit|LabModifier|false|false||TABLETnull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|torsemide|Drug|false|false||Torsemide
null|torsemide|Drug|false|false||Torsemidenull|Tablet Dosage Form|Drug|false|false||TABLETnull|Tablet (unit of presentation)|LabModifier|false|false||TABLET
null|Tablet Dosing Unit|LabModifier|false|false||TABLETnull|warfarin sodium|Drug|false|false||Warfarin sodium
null|warfarin sodium|Drug|false|false||Warfarin sodium
null|warfarin sodium|Drug|false|false||Warfarin sodiumnull|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarinnull|Sodium supplements|Drug|false|false||sodium
null|sodium|Drug|false|false||sodium
null|sodium|Drug|false|false||sodium
null|Sodium Drug Class|Drug|false|false||sodiumnull|Sodium metabolic function|Finding|false|false||sodiumnull|Sodium measurement|Procedure|false|false||sodiumnull|Tablet Dosage Form|Drug|false|false||TABLETnull|Tablet (unit of presentation)|LabModifier|false|false||TABLET
null|Tablet Dosing Unit|LabModifier|false|false||TABLETnull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|dexamethasone|Drug|false|false||dexamethasone
null|dexamethasone|Drug|false|false||dexamethasonenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|glipizide|Drug|false|false||glipizide
null|glipizide|Drug|false|false||glipizidenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Once A Day|Drug|false|false||once a daynull|Once daily|Time|false|false||once a daynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|goserelin|Drug|false|false||goserelin
null|goserelin|Drug|false|false||goserelinnull|Drug Implant|Drug|false|false||Implantnull|Traumatic implant|Disorder|false|false||Implantnull|null|Finding|false|false||Implant
null|Administration via Implantation|Finding|false|false||Implantnull|Implantation procedure|Procedure|false|false||Implantnull|null|Attribute|false|false||Implantnull|Implants|Device|false|false||Implantnull|Implant (unit of presentation)|LabModifier|false|false||Implant
null|Implant Dosing Unit|LabModifier|false|false||Implantnull|Drug Implant|Drug|false|false||implantnull|Traumatic implant|Disorder|false|false||implantnull|null|Finding|false|false||implant
null|Administration via Implantation|Finding|false|false||implantnull|Implantation procedure|Procedure|false|false||implantnull|null|Attribute|false|false||implantnull|Implants|Device|false|false||implantnull|Implant (unit of presentation)|LabModifier|false|false||implant
null|Implant Dosing Unit|LabModifier|false|false||implantnull|Subcutaneous Route of Administration|Finding|false|false||Subcutaneousnull|subcutaneous|Modifier|false|false||Subcutaneousnull|isosorbide dinitrate|Drug|false|false||isosorbide dinitrate
null|isosorbide dinitrate|Drug|false|false||isosorbide dinitratenull|isosorbide|Drug|false|false||isosorbide
null|isosorbide|Drug|false|false||isosorbidenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Twice a day|Time|false|false||twice a daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|lisinopril|Drug|false|false||lisinopril
null|lisinopril|Drug|false|false||lisinoprilnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Once A Day|Drug|false|false||once a daynull|Once daily|Time|false|false||once a daynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|metoprolol tartrate|Drug|false|false||metoprolol tartrate
null|metoprolol tartrate|Drug|false|false||metoprolol tartratenull|metoprolol|Drug|false|false||metoprolol
null|metoprolol|Drug|false|false||metoprololnull|tartrate|Drug|false|false||tartrate
null|Tartrates|Drug|false|false||tartrate
null|tartrate|Drug|false|false||tartratenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|nilutamide|Drug|false|false||nilutamide
null|nilutamide|Drug|false|false||nilutamidenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Once A Day|Drug|false|false||once a daynull|Once daily|Time|false|false||once a daynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|oxycodone|Drug|false|false||oxycodone
null|oxycodone|Drug|false|false||oxycodonenull|Oxycodone measurement|Procedure|false|false||oxycodonenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Hour|Time|false|false||hoursnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|simvastatin|Drug|false|false||simvastatin
null|simvastatin|Drug|false|false||simvastatinnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|torsemide|Drug|false|false||torsemide
null|torsemide|Drug|false|false||torsemidenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Once A Day|Drug|false|false||once a daynull|Once daily|Time|false|false||once a daynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|VITAMIN B12 MEASUREMENT|Procedure|false|false||cyanocobalamin (vitamin B-12)null|Cyanocobalamin Drug Class|Drug|false|false||cyanocobalamin
null|Cyanocobalamin Drug Class|Drug|false|false||cyanocobalamin
null|vitamin B12|Drug|false|false||cyanocobalamin
null|vitamin B12|Drug|false|false||cyanocobalamin
null|vitamin B12|Drug|false|false||cyanocobalaminnull|vitamin B12|Drug|false|false||vitamin B-12
null|cobalamins|Drug|false|false||vitamin B-12
null|cobalamins|Drug|false|false||vitamin B-12
null|vitamin B12|Drug|false|false||vitamin B-12
null|vitamin B12|Drug|false|false||vitamin B-12null|VITAMIN B12 MEASUREMENT|Procedure|false|false||vitamin B-12null|vitamin B complex|Drug|false|false||vitamin B
null|vitamin B complex|Drug|false|false||vitamin B
null|vitamin B complex|Drug|false|false||vitamin B
null|B Vitamin Family|Drug|false|false||vitamin B
null|B Vitamin Family|Drug|false|false||vitamin B
null|VITAMIN B|Drug|false|false||vitamin B
null|VITAMIN B|Drug|false|false||vitamin Bnull|Vitamins|Drug|false|false||vitamin
null|Vitamins|Drug|false|false||vitamin
null|Vitamins|Drug|false|false||vitaminnull|microgram|LabModifier|false|false||mcgnull|Liquid Dosage Form|Drug|false|false||Liquid
null|Liquid substance|Drug|false|false||Liquidnull|Liquid (finding)|Finding|false|false||Liquidnull|Liquid diet|Procedure|false|false||Liquidnull|Liquid (state of matter)|Modifier|false|false||Liquidnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Once a week|Time|false|false||once a weeknull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|memantine|Drug|false|false||memantine
null|memantine|Drug|false|false||memantinenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Twice a day|Time|false|false||twice a daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|allopurinol|Drug|false|false||allopurinol
null|allopurinol|Drug|false|false||allopurinolnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Once A Day|Drug|false|false||once a daynull|Once daily|Time|false|false||once a daynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarinnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||tabletsnull|Vitamin D Drug Class|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|D Vitamin|Drug|false|false||Vitamin D
null|Vitamin D [EPC]|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|Vitamin D Drug Class|Drug|false|false||Vitamin Dnull|Vitamin D measurement|Procedure|false|false||Vitamin Dnull|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitaminnull|Storage Unit|Device|false|false||unit
null|Unit device|Device|false|false||unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||unit
null|Unit of Measure|LabModifier|false|false||unit
null|Unit|LabModifier|false|false||unit
null|Enzyme Unit|LabModifier|false|false||unitnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|insulin glargine|Drug|false|false||insulin glargine
null|insulin glargine|Drug|false|false||insulin glargine
null|insulin glargine|Drug|false|false||insulin glarginenull|insulin, regular, human|Drug|false|false||insulin
null|Insulin [EPC]|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulinnull|INS gene|Finding|false|false||insulinnull|Insulin measurement|Procedure|false|false||insulinnull|insulin glargine|Drug|false|false||glargine
null|insulin glargine|Drug|false|false||glargine
null|insulin glargine|Drug|false|false||glarginenull|Unit per Milliliter|LabModifier|false|false||unit/mLnull|Storage Unit|Device|false|false||unit
null|Unit device|Device|false|false||unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||unit
null|Unit of Measure|LabModifier|false|false||unit
null|Unit|LabModifier|false|false||unit
null|Enzyme Unit|LabModifier|false|false||unitnull|per milliliter|LabModifier|false|false||/mLnull|Cartridge - package type|Finding|false|false||Cartridgenull|Cartridge device|Device|false|false||Cartridge
null|Cartridge|Device|false|false||Cartridgenull|Cartridge (unit of presentation)|LabModifier|false|false||Cartridge
null|Cartridge Dosing Unit|LabModifier|false|false||Cartridgenull|Unit - NCI Thesaurus Property|LabModifier|false|false||units
null|Unit of Measure|LabModifier|false|false||units
null|Unit|LabModifier|false|false||unitsnull|Subcutaneous Route of Administration|Finding|false|false||Subcutaneousnull|subcutaneous|Modifier|false|false||Subcutaneousnull|Once a day, at bedtime|Time|false|false||at bedtimenull|Once a day, at bedtime|Time|false|false||bedtime
null|Bedtime (qualifier value)|Time|false|false||bedtimenull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|ADMIN.FACILITY|Finding|false|false||Facilitynull|Facility (object)|Device|false|false||Facilitynull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|True primary (qualifier value)|Time|false|false||PRIMARYnull|Primary|Modifier|false|false||PRIMARYnull|Acute on chronic diastolic heart failure|Disorder|false|false|C4037974;C0018787|Acute on chronic diastolic congestive heart failurenull|Acute-on-chronic|Time|false|false||Acute on chronicnull|Admission Level of Care Code - Acute|Finding|false|false||Acute
null|Acute - Triage Code|Finding|false|false||Acutenull|acute|Time|false|false||Acutenull|Chronic diastolic heart failure|Disorder|false|false|C4037974;C0018787|chronic diastolic congestive heart failurenull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|diastolic congestive heart failure|Disorder|false|false|C4037974;C0018787|diastolic congestive heart failurenull|Diastole|Attribute|false|false||diastolicnull|Congestive heart failure|Disorder|false|false|C4037974;C0018787|congestive heart failurenull|Congestive|Modifier|false|false||congestivenull|Congestive heart failure|Disorder|false|false|C4037974;C0018787|heart failure
null|Heart failure|Disorder|false|false|C4037974;C0018787|heart failurenull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787|heart
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787|heartnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|heartnull|Chest>Heart|Anatomy|false|false|C2711480;C0795691;C0018801;C0018802;C2183328;C0018802;C0153957;C0153500;C2732749|heart
null|Heart|Anatomy|false|false|C2711480;C0795691;C0018801;C0018802;C2183328;C0018802;C0153957;C0153500;C2732749|heartnull|Failure (biologic function)|Finding|false|false||failure
null|Failure|Finding|false|false||failure
null|Personal failure|Finding|false|false||failurenull|Neoplasm Metastasis|Disorder|false|false||SECONDARYnull|metastatic qualifier|Finding|false|false||SECONDARYnull|Secondary to|Modifier|false|false||SECONDARYnull|second (number)|LabModifier|false|false||SECONDARYnull|Atrial Fibrillation|Disorder|false|false|C0018792|Atrial fibrillationnull|null|Attribute|false|false|C0018792|Atrial fibrillationnull|Atrial Fibrillation by ECG Finding|Lab|false|false|C0018792|Atrial fibrillationnull|Heart Atrium|Anatomy|false|false|C0232197;C0004238;C2926591;C0344434|Atrialnull|Fibrillation|Disorder|false|false|C0018792|fibrillationnull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||Diabetes
null|Diabetes|Disorder|false|false||Diabetes
null|Diabetes Mellitus|Disorder|false|false||Diabetesnull|Hypertensive disease|Disorder|false|false||Hypertensionnull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Helping Behavior|Finding|false|false||assistancenull|Assisted (qualifier value)|Modifier|false|false||assistancenull|AICDA protein, human|Drug|false|false||aid
null|AICDA protein, human|Drug|false|false||aidnull|AICDA wt Allele|Finding|false|false||aid
null|AICDA gene|Finding|false|false||aidnull|AID - Artificial insemination by donor|Procedure|false|false||aid
null|dacarbazine/doxorubicin/ifosfamide protocol|Procedure|false|false||aidnull|Aid (attribute)|Modifier|false|false||aid
null|Assisted (qualifier value)|Modifier|false|false||aidnull|Walkers|Device|false|false||walkernull|CANE, INCLUDES CANES OF ALL MATERIALS, ADJUSTABLE OR FIXED, WITH TIP|Device|false|false||canenull|Cane - plant part|Entity|false|false||canenull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Swelling|Finding|false|false|C1140621|swelling
null|Edema|Finding|false|false|C1140621|swellingnull|Leg|Anatomy|false|false|C5781420;C0013604;C0038999|legsnull|null|Attribute|false|false|C1140621|legsnull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Congestive heart failure|Disorder|false|false|C4037974;C0018787|heart failure
null|Heart failure|Disorder|false|false|C4037974;C0018787|heart failurenull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787|heart
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787|heartnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|heartnull|Chest>Heart|Anatomy|false|false|C0018801;C0018802;C0153957;C0153500;C0795691|heart
null|Heart|Anatomy|false|false|C0018801;C0018802;C0153957;C0153500;C0795691|heartnull|Failure (biologic function)|Finding|false|false||failure
null|Failure|Finding|false|false||failure
null|Personal failure|Finding|false|false||failurenull|Diuretic [APC]|Drug|false|false||diuretic
null|Diuretics|Drug|false|false||diureticnull|Diagnostic Service Section ID - Physical Therapy|Finding|false|false||physical therapynull|Physical therapy|Procedure|false|false||physical therapynull|Physical therapy (field)|Title|false|false||physical therapynull|physical examination (physical finding)|Finding|false|false||physical
null|Physical|Finding|false|false||physicalnull|Physical Examination|Procedure|false|false||physicalnull|Therapy Object (animal model)|Finding|false|false||therapy
null|therapeutic aspects|Finding|false|false||therapynull|Therapeutic procedure|Procedure|false|false||therapynull|Daily|Time|false|false||dailynull|Doctor - Title|Finding|false|false||doctornull|Physicians|Subject|false|false||doctornull|infant weight for previous delivery (history)|Finding|false|false||weight
null|Weight symptom (finding)|Finding|false|false||weightnull|Weighing patient|Procedure|false|false||weightnull|null|Attribute|false|false||weightnull|Body Weight|Subject|false|false||weightnull|Importance Weight|Modifier|false|false||weightnull|Weight|LabModifier|false|false||weightnull|Greater Than|LabModifier|false|false||more thannull|More|LabModifier|false|false||morenull|Pounds|LabModifier|false|false||poundsnull|Pharmaceutical Preparations|Drug|false|false||Medicationnull|medication - HL7 publishing domain|Finding|false|false||Medication
null|Medications|Finding|false|false||Medicationnull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|Continuous|Finding|false|false||CONTINUEnull|torsemide|Drug|false|false||torsemide
null|torsemide|Drug|false|false||torsemidenull|Daily|Time|false|false||dailynull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|metoprolol|Drug|false|false||metoprolol
null|metoprolol|Drug|false|false||metoprololnull|Daily|Time|false|false||dailynull|Blood pressure finding|Finding|false|false||blood pressure
null|Systemic arterial pressure|Finding|false|false||blood pressure
null|Blood Pressure|Finding|false|false||blood pressurenull|Blood pressure determination|Procedure|false|false||blood pressurenull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|IPSS-R Risk Category Low|Finding|false|false||low
null|IPSS Risk Category Low|Finding|false|false||low
null|low confidentiality|Finding|false|false||lownull|Low - MessageWaitingPriority|Modifier|false|false||low
null|low|Modifier|false|false||low
null|low exposure|Modifier|false|false||lownull|null|LabModifier|false|false||lownull|Doctor - Title|Finding|false|false||doctornull|Physicians|Subject|false|false||doctornull|Office Visits|Procedure|false|false||office visitnull|Address type - Office|Finding|false|false||officenull|Office|Device|false|false||officenull|Organization unit type - Office|Entity|false|false||officenull|Visit|Finding|false|false||visitnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions